module decoder_controller (

    
);


endmodule