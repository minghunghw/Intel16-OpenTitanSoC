// For DHM

`define DHM_STAGES_0       0
`define DHM_INCLUDE_RAM_0  0
`define DHM_STAGES_1       0
`define DHM_INCLUDE_RAM_1  0
`define DHM_STAGES_2       0
`define DHM_INCLUDE_RAM_2  0
`define DHM_LUT_WIDTH_IN   4
`define DHM_LUT_WIDTH_OUT  4

// For DHM_RAM

`define DHM_RAM_STAGES_0       0
`define DHM_RAM_INCLUDE_RAM_0  1
`define DHM_RAM_STAGES_1       0
`define DHM_RAM_INCLUDE_RAM_1  1
`define DHM_RAM_STAGES_2       0
`define DHM_RAM_INCLUDE_RAM_2  1
`define DHM_RAM_LUT_WIDTH_IN   4
`define DHM_RAM_LUT_WIDTH_OUT  4

// For DHM_UPF

`define DHM_UPF_STAGES_0       0
`define DHM_UPF_INCLUDE_RAM_0  0
`define DHM_UPF_STAGES_1       0
`define DHM_UPF_INCLUDE_RAM_1  0
`define DHM_UPF_STAGES_2       0
`define DHM_UPF_INCLUDE_RAM_2  0
`define DHM_UPF_LUT_WIDTH_IN   4
`define DHM_UPF_LUT_WIDTH_OUT  4

// For DSMA

`define DSMA_STAGES_0       0
`define DSMA_INCLUDE_RAM_0  0
`define DSMA_STAGES_1       0
`define DSMA_INCLUDE_RAM_1  0
`define DSMA_STAGES_2       0
`define DSMA_INCLUDE_RAM_2  0
`define DSMA_LUT_WIDTH_IN   4
`define DSMA_LUT_WIDTH_OUT  4

// For DSMB

`define DSMB_STAGES_0       0
`define DSMB_INCLUDE_RAM_0  0
`define DSMB_STAGES_1       0
`define DSMB_INCLUDE_RAM_1  0
`define DSMB_STAGES_2       0
`define DSMB_INCLUDE_RAM_2  0
`define DSMB_LUT_WIDTH_IN   4
`define DSMB_LUT_WIDTH_OUT  4

////////////////////////////////////////////////////////////////////////////////
// end of file
////////////////////////////////////////////////////////////////////////////////
