module spi_device_tlul (clk_i,
    rst_ni,
    spi_cs,
    spi_sclk,
    spi_sdi0,
    spi_sdi1,
    spi_sdi2,
    spi_sdi3,
    spi_sdo0,
    spi_sdo1,
    spi_sdo2,
    spi_sdo3,
    test_mode,
    spi_mode,
    tl_i,
    tl_o);
 input clk_i;
 input rst_ni;
 input spi_cs;
 input spi_sclk;
 input spi_sdi0;
 input spi_sdi1;
 input spi_sdi2;
 input spi_sdi3;
 output spi_sdo0;
 output spi_sdo1;
 output spi_sdo2;
 output spi_sdo3;
 input test_mode;
 output [1:0] spi_mode;
 input [65:0] tl_i;
 output [108:0] tl_o;

 wire ctrl_addr_valid;
 wire ctrl_data_tx_ready;
 wire ctrl_rd_wr;
 wire en_quad;
 wire n1455;
 wire n1456;
 wire n1691;
 wire n1694;
 wire n1697;
 wire n1700;
 wire n1703;
 wire n1706;
 wire n1709;
 wire n1712;
 wire n1715;
 wire n1718;
 wire n1721;
 wire n1724;
 wire n1727;
 wire n1730;
 wire n1733;
 wire n1736;
 wire n1739;
 wire n1742;
 wire n1745;
 wire n1748;
 wire n1751;
 wire n1754;
 wire n1757;
 wire n1760;
 wire n1763;
 wire n1766;
 wire n1769;
 wire n1772;
 wire n1775;
 wire n1778;
 wire n1781;
 wire n1784;
 wire n1787;
 wire n1790;
 wire n1793;
 wire n1796;
 wire n1799;
 wire n1802;
 wire n1869;
 wire n1878;
 wire n1881;
 wire n2656;
 wire n2723;
 wire n2726;
 wire n2727;
 wire n2728;
 wire n2729;
 wire n2730;
 wire n2731;
 wire n2732;
 wire n2733;
 wire n2734;
 wire n2735;
 wire n2736;
 wire n2737;
 wire n2738;
 wire n2739;
 wire n2740;
 wire n2741;
 wire n2742;
 wire n2743;
 wire n2744;
 wire n2745;
 wire n2746;
 wire n2747;
 wire n2748;
 wire n2749;
 wire n2750;
 wire n2751;
 wire n2763;
 wire n2764;
 wire n2765;
 wire n2766;
 wire n2767;
 wire n2768;
 wire n2769;
 wire n2770;
 wire n2771;
 wire n2772;
 wire n2773;
 wire n2774;
 wire n2775;
 wire n2776;
 wire n2777;
 wire n2778;
 wire n2779;
 wire n2780;
 wire n2781;
 wire n2782;
 wire n2783;
 wire n2784;
 wire n2787;
 wire n2788;
 wire n2789;
 wire n2790;
 wire n2791;
 wire n2792;
 wire n2793;
 wire n2794;
 wire n2795;
 wire n2796;
 wire n2797;
 wire n2798;
 wire n2799;
 wire n2802;
 wire n2803;
 wire n2804;
 wire n2805;
 wire n2806;
 wire n2807;
 wire n2808;
 wire n2809;
 wire n2810;
 wire n2811;
 wire n2812;
 wire n2813;
 wire n2814;
 wire n2815;
 wire n2816;
 wire n2819;
 wire n2820;
 wire n2822;
 wire n2823;
 wire n2824;
 wire n2825;
 wire n2826;
 wire n2827;
 wire n2828;
 wire n2829;
 wire n2830;
 wire n2831;
 wire n2832;
 wire n2833;
 wire n2834;
 wire n2835;
 wire n2836;
 wire n2837;
 wire n2838;
 wire n2839;
 wire n2840;
 wire n2841;
 wire n2842;
 wire n2843;
 wire n2844;
 wire n2845;
 wire n2846;
 wire n2847;
 wire n2848;
 wire n2849;
 wire n2850;
 wire n2851;
 wire n2852;
 wire n2853;
 wire n2854;
 wire n2855;
 wire n2856;
 wire n2857;
 wire n2858;
 wire n2859;
 wire n2860;
 wire n2861;
 wire n2862;
 wire n2863;
 wire n2864;
 wire n2865;
 wire n2866;
 wire n2867;
 wire n2868;
 wire n2870;
 wire n2871;
 wire n2872;
 wire n2873;
 wire n2874;
 wire n2875;
 wire n2876;
 wire n2877;
 wire n2878;
 wire n2879;
 wire n2880;
 wire n2881;
 wire n2882;
 wire n2883;
 wire n2884;
 wire n2885;
 wire n2886;
 wire n2887;
 wire n2888;
 wire n2889;
 wire n2890;
 wire n2891;
 wire n2892;
 wire n2893;
 wire n2894;
 wire n2895;
 wire n2896;
 wire n2897;
 wire n2898;
 wire n2899;
 wire n2900;
 wire n2901;
 wire n2902;
 wire n2903;
 wire n2904;
 wire n2905;
 wire n2906;
 wire n2907;
 wire n2908;
 wire n2917;
 wire n2919;
 wire n2920;
 wire n2921;
 wire n2922;
 wire n2923;
 wire n2925;
 wire n2927;
 wire n2928;
 wire n2929;
 wire n2930;
 wire n2931;
 wire n2932;
 wire n2933;
 wire n2934;
 wire n2935;
 wire n2936;
 wire n2937;
 wire n2938;
 wire n2939;
 wire n2940;
 wire n2941;
 wire n2942;
 wire n2943;
 wire n2945;
 wire n2946;
 wire n2948;
 wire n2951;
 wire n2953;
 wire n2954;
 wire n2955;
 wire n2956;
 wire n2957;
 wire n2958;
 wire n2959;
 wire n2960;
 wire n2961;
 wire n2962;
 wire n2963;
 wire n2964;
 wire n2965;
 wire n2966;
 wire n2967;
 wire n2968;
 wire n2969;
 wire n2970;
 wire n2971;
 wire n2972;
 wire n2973;
 wire n2974;
 wire n2975;
 wire n2976;
 wire n2977;
 wire n2978;
 wire n2979;
 wire n2980;
 wire n2981;
 wire n3001;
 wire n3002;
 wire n3003;
 wire n3004;
 wire n3005;
 wire n3006;
 wire n3007;
 wire n3008;
 wire n3009;
 wire n3010;
 wire n3011;
 wire n3012;
 wire n3013;
 wire n3014;
 wire n3015;
 wire n3016;
 wire n3017;
 wire n3018;
 wire n3019;
 wire n3020;
 wire n3021;
 wire n3022;
 wire n3023;
 wire n3024;
 wire n3025;
 wire n3026;
 wire n3027;
 wire n3028;
 wire n3029;
 wire n3031;
 wire n3035;
 wire n3036;
 wire n3037;
 wire n3038;
 wire n3039;
 wire n3041;
 wire n3042;
 wire n3043;
 wire n3044;
 wire n3045;
 wire n3047;
 wire n3048;
 wire n3049;
 wire n3050;
 wire n3051;
 wire n3052;
 wire n3053;
 wire n3054;
 wire n3055;
 wire n3056;
 wire n3058;
 wire n3059;
 wire n3060;
 wire n3061;
 wire n3062;
 wire n3063;
 wire n3064;
 wire n3065;
 wire n3066;
 wire n3067;
 wire n3068;
 wire n3069;
 wire n3070;
 wire n3071;
 wire n3072;
 wire n3073;
 wire n3074;
 wire n3075;
 wire n3076;
 wire n3077;
 wire n3078;
 wire n3079;
 wire n3080;
 wire n3081;
 wire n3082;
 wire n3083;
 wire n3084;
 wire n3085;
 wire n3086;
 wire n3087;
 wire n3088;
 wire n3089;
 wire n3090;
 wire n3091;
 wire n3092;
 wire n3093;
 wire n3094;
 wire n3095;
 wire n3096;
 wire n3097;
 wire n3098;
 wire n3099;
 wire n3100;
 wire n3101;
 wire n3102;
 wire n3103;
 wire n3104;
 wire n3105;
 wire n3106;
 wire n3107;
 wire n3108;
 wire n3109;
 wire n3110;
 wire n3111;
 wire n3112;
 wire n3114;
 wire n3115;
 wire n3116;
 wire n3117;
 wire n3118;
 wire n3119;
 wire n3120;
 wire n3121;
 wire n3122;
 wire n3123;
 wire n3124;
 wire n3125;
 wire n3126;
 wire n3127;
 wire n3128;
 wire n3131;
 wire n3132;
 wire n3133;
 wire n3134;
 wire n3135;
 wire n3136;
 wire n3137;
 wire n3138;
 wire n3139;
 wire n3140;
 wire n3143;
 wire n3144;
 wire n3145;
 wire n3146;
 wire n3148;
 wire n3150;
 wire n3151;
 wire n3152;
 wire n3153;
 wire n3155;
 wire n3157;
 wire n3158;
 wire n3159;
 wire n3160;
 wire n3161;
 wire n3162;
 wire n3163;
 wire n3164;
 wire n3169;
 wire n3170;
 wire n3171;
 wire n3172;
 wire n3173;
 wire n3174;
 wire n3176;
 wire n3177;
 wire n3178;
 wire n3179;
 wire n3180;
 wire n3181;
 wire n3182;
 wire n3183;
 wire n3184;
 wire n3185;
 wire n3186;
 wire n3187;
 wire n3188;
 wire n3189;
 wire n3190;
 wire n3191;
 wire n3192;
 wire n3193;
 wire n3194;
 wire n3196;
 wire n3197;
 wire n3198;
 wire n3199;
 wire n3200;
 wire n3201;
 wire n3202;
 wire n3203;
 wire n3204;
 wire n3205;
 wire n3206;
 wire n3209;
 wire n3210;
 wire n3211;
 wire n3212;
 wire n3213;
 wire n3214;
 wire n3215;
 wire n3216;
 wire n3222;
 wire n3223;
 wire n3224;
 wire n3225;
 wire n3226;
 wire n3227;
 wire n3228;
 wire n3229;
 wire n3230;
 wire n3233;
 wire n3234;
 wire n3235;
 wire n3236;
 wire n3237;
 wire n3238;
 wire n3239;
 wire n3240;
 wire n3241;
 wire n3242;
 wire n3243;
 wire n3244;
 wire n3245;
 wire n3246;
 wire n3247;
 wire n3248;
 wire n3249;
 wire n3250;
 wire n3251;
 wire n3252;
 wire n3253;
 wire n3254;
 wire n3255;
 wire n3256;
 wire n3257;
 wire n3258;
 wire n3259;
 wire n3260;
 wire n3261;
 wire n3262;
 wire n3263;
 wire n3264;
 wire n3265;
 wire n3266;
 wire n3267;
 wire n3268;
 wire n3269;
 wire n3270;
 wire n3271;
 wire n3272;
 wire n3273;
 wire n3274;
 wire n3275;
 wire n3276;
 wire n3277;
 wire n3278;
 wire n3279;
 wire n3280;
 wire n3281;
 wire n3282;
 wire n3283;
 wire n3284;
 wire n3285;
 wire n3286;
 wire n3287;
 wire n3288;
 wire n3289;
 wire n3290;
 wire n3291;
 wire n3292;
 wire n3293;
 wire n3294;
 wire n3295;
 wire n3296;
 wire n3297;
 wire n3298;
 wire n3299;
 wire n3300;
 wire n3301;
 wire n3302;
 wire n3303;
 wire n3304;
 wire n3305;
 wire n3306;
 wire n3307;
 wire n3308;
 wire n3309;
 wire n3310;
 wire n3311;
 wire n3312;
 wire n3313;
 wire n3314;
 wire n3315;
 wire n3316;
 wire n3317;
 wire n3318;
 wire n3319;
 wire n3320;
 wire n3321;
 wire n3322;
 wire n3323;
 wire n3324;
 wire n3325;
 wire n3326;
 wire n3327;
 wire n3328;
 wire n3329;
 wire n3330;
 wire n3331;
 wire n3332;
 wire n3333;
 wire n3334;
 wire n3335;
 wire n3336;
 wire n3337;
 wire n3338;
 wire n3339;
 wire n3340;
 wire n3341;
 wire n3342;
 wire n3343;
 wire n3344;
 wire n3345;
 wire n3346;
 wire n3347;
 wire n3348;
 wire n3349;
 wire n3350;
 wire n3351;
 wire n3352;
 wire n3353;
 wire n3354;
 wire n3355;
 wire n3356;
 wire n3357;
 wire n3358;
 wire n3359;
 wire n3360;
 wire n3361;
 wire n3362;
 wire n3363;
 wire n3364;
 wire n3365;
 wire n3366;
 wire n3367;
 wire n3368;
 wire n3369;
 wire n3370;
 wire n3372;
 wire n3373;
 wire n3374;
 wire n3375;
 wire n3376;
 wire n3380;
 wire n3381;
 wire n3382;
 wire n3383;
 wire n3384;
 wire n3385;
 wire n3386;
 wire n3387;
 wire n3388;
 wire n3389;
 wire n3390;
 wire n3391;
 wire n3392;
 wire n3393;
 wire n3394;
 wire n3398;
 wire n3399;
 wire n3400;
 wire n3401;
 wire n3402;
 wire n3404;
 wire n3405;
 wire n3406;
 wire n3407;
 wire n3408;
 wire n3409;
 wire n3410;
 wire n3411;
 wire n3412;
 wire n3413;
 wire n3415;
 wire n3416;
 wire n3417;
 wire n3418;
 wire n3419;
 wire n3420;
 wire n3421;
 wire n3422;
 wire n3423;
 wire n3424;
 wire n3425;
 wire n3426;
 wire n3427;
 wire n3428;
 wire n3429;
 wire n3430;
 wire n3431;
 wire n3432;
 wire n3433;
 wire n3434;
 wire n3435;
 wire n3436;
 wire n3437;
 wire n3438;
 wire n3439;
 wire n3440;
 wire n3441;
 wire n3442;
 wire n3443;
 wire n3444;
 wire n3445;
 wire n3446;
 wire n3447;
 wire n3448;
 wire n3449;
 wire n3450;
 wire n3451;
 wire n3452;
 wire n3453;
 wire n3454;
 wire n3455;
 wire n3456;
 wire n3457;
 wire n3458;
 wire n3459;
 wire n3460;
 wire n3461;
 wire n3462;
 wire n3463;
 wire n3464;
 wire n3465;
 wire n3466;
 wire n3467;
 wire n3468;
 wire n3469;
 wire n3471;
 wire n3472;
 wire n3473;
 wire n3474;
 wire n3475;
 wire n3477;
 wire n3478;
 wire n3479;
 wire n3480;
 wire n3481;
 wire n3482;
 wire n3483;
 wire n3484;
 wire n3485;
 wire n3486;
 wire n3487;
 wire n3488;
 wire n3489;
 wire n3490;
 wire n3491;
 wire n3492;
 wire n3493;
 wire n3494;
 wire n3495;
 wire n3496;
 wire n3497;
 wire n3498;
 wire n3499;
 wire n3500;
 wire n3501;
 wire n3503;
 wire n3504;
 wire n3505;
 wire n3506;
 wire n3507;
 wire n3510;
 wire n3511;
 wire n3512;
 wire n3513;
 wire n3514;
 wire n3517;
 wire n3518;
 wire n3519;
 wire n3520;
 wire n3521;
 wire n3525;
 wire n3526;
 wire n3527;
 wire n3528;
 wire n3529;
 wire n3532;
 wire n3533;
 wire n3534;
 wire n3535;
 wire n3536;
 wire n3542;
 wire n3543;
 wire n3544;
 wire n3545;
 wire n3546;
 wire n3556;
 wire n3557;
 wire n3558;
 wire n3559;
 wire n3560;
 wire n3561;
 wire n3562;
 wire n3563;
 wire n3564;
 wire n3565;
 wire n3566;
 wire n3567;
 wire n3568;
 wire n3569;
 wire n3570;
 wire n3571;
 wire n3572;
 wire n3573;
 wire n3574;
 wire n3575;
 wire n3576;
 wire n3577;
 wire n3578;
 wire n3579;
 wire n3580;
 wire n3581;
 wire n3582;
 wire n3583;
 wire n3584;
 wire n3585;
 wire n3586;
 wire n3587;
 wire n3588;
 wire n3589;
 wire n3590;
 wire n3591;
 wire n3592;
 wire n3593;
 wire n3594;
 wire n3595;
 wire n3596;
 wire n3597;
 wire n3598;
 wire n3599;
 wire n3600;
 wire n3601;
 wire n3602;
 wire n3603;
 wire n3604;
 wire n3605;
 wire n3606;
 wire n3607;
 wire n3608;
 wire n3609;
 wire n3610;
 wire n3611;
 wire n3612;
 wire n3613;
 wire n3614;
 wire n3615;
 wire n3616;
 wire n3617;
 wire n3618;
 wire n3619;
 wire n3620;
 wire n3621;
 wire n3622;
 wire n3623;
 wire n3625;
 wire n3626;
 wire n3627;
 wire n3628;
 wire n3629;
 wire n3631;
 wire n3632;
 wire n3633;
 wire n3634;
 wire n3635;
 wire n3636;
 wire n3637;
 wire n3638;
 wire n3639;
 wire n3640;
 wire n3641;
 wire n3642;
 wire n3643;
 wire n3644;
 wire n3645;
 wire n3646;
 wire n3647;
 wire n3648;
 wire n3649;
 wire n3650;
 wire n3651;
 wire n3652;
 wire n3653;
 wire n3654;
 wire n3655;
 wire n3656;
 wire n3657;
 wire n3658;
 wire n3659;
 wire n3660;
 wire n3661;
 wire n3662;
 wire n3663;
 wire n3664;
 wire n3665;
 wire n3666;
 wire n3675;
 wire n3676;
 wire n3677;
 wire n3678;
 wire n3679;
 wire n3680;
 wire n3681;
 wire n3682;
 wire n3683;
 wire n3685;
 wire n3688;
 wire n3769;
 wire n3770;
 wire n3771;
 wire n3772;
 wire n3773;
 wire n3774;
 wire n3776;
 wire n3777;
 wire n3778;
 wire net94;
 wire net93;
 wire net92;
 wire net91;
 wire net90;
 wire net89;
 wire net88;
 wire net87;
 wire net86;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net81;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire net75;
 wire net74;
 wire net73;
 wire net72;
 wire net71;
 wire net70;
 wire net69;
 wire net68;
 wire n3807;
 wire net67;
 wire n3809;
 wire n3811;
 wire net66;
 wire n3813;
 wire n3815;
 wire n3817;
 wire n3818;
 wire n3819;
 wire n3820;
 wire n3821;
 wire n3822;
 wire net63;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire net54;
 wire net53;
 wire net52;
 wire net51;
 wire net50;
 wire net49;
 wire net48;
 wire net47;
 wire net46;
 wire net45;
 wire net44;
 wire net43;
 wire net42;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire net36;
 wire net35;
 wire net34;
 wire net33;
 wire net32;
 wire net31;
 wire net30;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire net11;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire net65;
 wire net64;
 wire net1;
 wire n604;
 wire net1954;
 wire rd_wr_sync;
 wire tx_counter_upd;
 wire tx_data_valid;
 wire tx_done;
 wire u_dcfifo_rx_u_din_buffer_N26;
 wire u_dcfifo_rx_u_din_buffer_N27;
 wire u_dcfifo_rx_u_din_buffer_N28;
 wire u_dcfifo_rx_u_din_buffer_N29;
 wire u_dcfifo_rx_u_din_buffer_N30;
 wire u_dcfifo_rx_u_din_buffer_N31;
 wire u_dcfifo_rx_u_din_buffer_N32;
 wire u_dcfifo_rx_u_din_buffer_N33;
 wire u_dcfifo_rx_u_din_buffer_net670;
 wire u_dcfifo_rx_u_din_buffer_net676;
 wire u_dcfifo_rx_u_din_buffer_net681;
 wire u_dcfifo_rx_u_din_buffer_net686;
 wire u_dcfifo_rx_u_din_buffer_net691;
 wire u_dcfifo_rx_u_din_buffer_net696;
 wire u_dcfifo_rx_u_din_buffer_net701;
 wire u_dcfifo_rx_u_din_buffer_net706;
 wire u_dcfifo_rx_u_din_buffer_net711;
 wire u_dcfifo_rx_u_din_buffer_net716;
 wire u_dcfifo_rx_u_din_buffer_net721;
 wire u_dcfifo_rx_u_din_buffer_net726;
 wire u_dcfifo_rx_u_din_buffer_net731;
 wire u_dcfifo_rx_u_din_buffer_net736;
 wire u_dcfifo_rx_u_din_buffer_net741;
 wire u_dcfifo_rx_u_din_buffer_net746;
 wire u_dcfifo_rx_u_din_full_N0;
 wire u_dcfifo_rx_u_din_full_full_dn;
 wire u_dcfifo_rx_u_din_full_full_synch_d_middle_0_;
 wire u_dcfifo_rx_u_din_full_full_up;
 wire u_dcfifo_rx_u_din_full_latched_full_s;
 wire u_dcfifo_rx_u_din_write_enable;
 wire u_dcfifo_rx_u_din_write_tr_net652;
 wire u_dcfifo_rx_u_dout_read_tr_net634;
 wire u_dcfifo_tx_u_din_buffer_N26;
 wire u_dcfifo_tx_u_din_buffer_N27;
 wire u_dcfifo_tx_u_din_buffer_N28;
 wire u_dcfifo_tx_u_din_buffer_N29;
 wire u_dcfifo_tx_u_din_buffer_N30;
 wire u_dcfifo_tx_u_din_buffer_N31;
 wire u_dcfifo_tx_u_din_buffer_N32;
 wire u_dcfifo_tx_u_din_buffer_N33;
 wire u_dcfifo_tx_u_din_buffer_net670;
 wire u_dcfifo_tx_u_din_buffer_net676;
 wire u_dcfifo_tx_u_din_buffer_net681;
 wire u_dcfifo_tx_u_din_buffer_net686;
 wire u_dcfifo_tx_u_din_buffer_net691;
 wire u_dcfifo_tx_u_din_buffer_net696;
 wire u_dcfifo_tx_u_din_buffer_net701;
 wire u_dcfifo_tx_u_din_buffer_net706;
 wire u_dcfifo_tx_u_din_buffer_net711;
 wire u_dcfifo_tx_u_din_buffer_net716;
 wire u_dcfifo_tx_u_din_buffer_net721;
 wire u_dcfifo_tx_u_din_buffer_net726;
 wire u_dcfifo_tx_u_din_buffer_net731;
 wire u_dcfifo_tx_u_din_buffer_net736;
 wire u_dcfifo_tx_u_din_buffer_net741;
 wire u_dcfifo_tx_u_din_buffer_net746;
 wire u_dcfifo_tx_u_din_full_N0;
 wire u_dcfifo_tx_u_din_full_full_dn;
 wire u_dcfifo_tx_u_din_full_full_synch_d_middle_0_;
 wire u_dcfifo_tx_u_din_full_full_up;
 wire u_dcfifo_tx_u_din_full_latched_full_s;
 wire u_dcfifo_tx_u_din_write_enable;
 wire u_dcfifo_tx_u_din_write_tr_net652;
 wire u_dcfifo_tx_u_dout_read_enable;
 wire u_dcfifo_tx_u_dout_read_tr_net634;
 wire u_device_sm_N163;
 wire u_device_sm_N174;
 wire u_device_sm_N175;
 wire u_device_sm_N176;
 wire u_device_sm_N177;
 wire u_device_sm_N178;
 wire u_device_sm_N179;
 wire u_device_sm_N180;
 wire u_device_sm_N181;
 wire u_device_sm_N182;
 wire u_device_sm_N183;
 wire u_device_sm_N184;
 wire u_device_sm_N185;
 wire u_device_sm_N186;
 wire u_device_sm_N187;
 wire u_device_sm_N188;
 wire u_device_sm_N189;
 wire u_device_sm_N190;
 wire u_device_sm_N191;
 wire u_device_sm_N192;
 wire u_device_sm_N193;
 wire u_device_sm_N194;
 wire u_device_sm_N195;
 wire u_device_sm_N196;
 wire u_device_sm_N197;
 wire u_device_sm_N198;
 wire u_device_sm_N199;
 wire u_device_sm_N200;
 wire u_device_sm_N201;
 wire u_device_sm_N202;
 wire u_device_sm_N203;
 wire u_device_sm_N204;
 wire u_device_sm_N205;
 wire u_device_sm_ctrl_data_tx_ready_next;
 wire u_device_sm_net763;
 wire u_device_sm_net769;
 wire u_device_sm_net774;
 wire u_device_sm_sample_ADDR;
 wire u_device_sm_sample_CMD;
 wire u_device_sm_tx_counter_next_3_;
 wire u_device_sm_tx_counter_upd_next;
 wire u_device_sm_tx_data_valid_next;
 wire u_device_sm_tx_done_reg;
 wire u_device_sm_u_spiregs_N31;
 wire u_device_sm_u_spiregs_N32;
 wire u_device_sm_u_spiregs_N33;
 wire u_device_sm_u_spiregs_N34;
 wire u_device_sm_u_spiregs_net791;
 wire u_device_sm_u_spiregs_net797;
 wire u_device_sm_u_spiregs_net802;
 wire u_device_sm_u_spiregs_net807;
 wire u_rxreg_N22;
 wire u_rxreg_N23;
 wire u_rxreg_N24;
 wire u_rxreg_N25;
 wire u_rxreg_N26;
 wire u_rxreg_N27;
 wire u_rxreg_N28;
 wire u_rxreg_N29;
 wire u_rxreg_N30;
 wire u_rxreg_N31;
 wire u_rxreg_N32;
 wire u_rxreg_N33;
 wire u_rxreg_N34;
 wire u_rxreg_N35;
 wire u_rxreg_N36;
 wire u_rxreg_N37;
 wire u_rxreg_N38;
 wire u_rxreg_N39;
 wire u_rxreg_N40;
 wire u_rxreg_N41;
 wire u_rxreg_N42;
 wire u_rxreg_N43;
 wire u_rxreg_N44;
 wire u_rxreg_N45;
 wire u_rxreg_N46;
 wire u_rxreg_N47;
 wire u_rxreg_N48;
 wire u_rxreg_N49;
 wire u_rxreg_N50;
 wire u_rxreg_N51;
 wire u_rxreg_N52;
 wire u_rxreg_N53;
 wire u_rxreg_N54;
 wire u_rxreg_N55;
 wire u_rxreg_N56;
 wire u_rxreg_N57;
 wire u_rxreg_N58;
 wire u_rxreg_N59;
 wire u_rxreg_N60;
 wire u_rxreg_N7;
 wire u_rxreg_N9;
 wire u_rxreg_net857;
 wire u_rxreg_net863;
 wire u_rxreg_net868;
 wire u_rxreg_net873;
 wire u_spi_device_tlul_plug_N61;
 wire u_spi_device_tlul_plug_net611;
 wire u_spi_device_tlul_plug_net617;
 wire u_spi_device_tlul_plug_we;
 wire u_syncro_cs_reg_0_;
 wire u_syncro_rdwr_reg_0_;
 wire u_txreg_N10;
 wire u_txreg_N11;
 wire u_txreg_N24;
 wire u_txreg_N25;
 wire u_txreg_N26;
 wire u_txreg_N27;
 wire u_txreg_N28;
 wire u_txreg_N29;
 wire u_txreg_N30;
 wire u_txreg_N31;
 wire u_txreg_N34;
 wire u_txreg_N35;
 wire u_txreg_N36;
 wire u_txreg_N37;
 wire u_txreg_N38;
 wire u_txreg_N39;
 wire u_txreg_N40;
 wire u_txreg_N41;
 wire u_txreg_N42;
 wire u_txreg_N43;
 wire u_txreg_N44;
 wire u_txreg_N45;
 wire u_txreg_N46;
 wire u_txreg_N47;
 wire u_txreg_N48;
 wire u_txreg_N49;
 wire u_txreg_N50;
 wire u_txreg_N51;
 wire u_txreg_N52;
 wire u_txreg_N53;
 wire u_txreg_N54;
 wire u_txreg_N55;
 wire u_txreg_N56;
 wire u_txreg_N57;
 wire u_txreg_N58;
 wire u_txreg_N59;
 wire u_txreg_N60;
 wire u_txreg_N61;
 wire u_txreg_N62;
 wire u_txreg_N63;
 wire u_txreg_N64;
 wire u_txreg_N65;
 wire u_txreg_net824;
 wire u_txreg_net830;
 wire u_txreg_net835;
 wire u_txreg_net840;
 wire u_txreg_running;
 wire clknet_0_clk_i;
 wire u_txreg_sclk_test;
 wire net1450;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire clknet_2_0_0_clk_i;
 wire clknet_2_1_0_clk_i;
 wire clknet_2_2_0_clk_i;
 wire clknet_2_3_0_clk_i;
 wire clknet_0_u_spi_device_tlul_plug_net611;
 wire clknet_1_0__leaf_u_spi_device_tlul_plug_net611;
 wire clknet_1_1__leaf_u_spi_device_tlul_plug_net611;
 wire clknet_0_u_spi_device_tlul_plug_net617;
 wire clknet_1_0__leaf_u_spi_device_tlul_plug_net617;
 wire clknet_1_1__leaf_u_spi_device_tlul_plug_net617;
 wire clknet_0_u_dcfifo_tx_u_din_write_tr_net652;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_write_tr_net652;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_write_tr_net652;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net670;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net670;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net670;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net676;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net676;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net676;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net681;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net681;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net681;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net686;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net686;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net686;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net691;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net691;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net691;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net696;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net696;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net696;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net701;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net701;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net701;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net706;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net706;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net706;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net711;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net711;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net711;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net716;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net716;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net716;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net721;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net721;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net721;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net726;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net726;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net726;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net731;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net731;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net731;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net736;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net736;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net736;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net741;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net741;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net741;
 wire clknet_0_u_dcfifo_tx_u_din_buffer_net746;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net746;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net746;
 wire clknet_0_u_dcfifo_rx_u_dout_read_tr_net634;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_dout_read_tr_net634;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_dout_read_tr_net634;
 wire clknet_0_spi_sclk;
 wire clknet_2_0_0_spi_sclk;
 wire clknet_2_1_0_spi_sclk;
 wire clknet_2_2_0_spi_sclk;
 wire clknet_2_3_0_spi_sclk;
 wire clknet_3_0__leaf_spi_sclk;
 wire clknet_3_1__leaf_spi_sclk;
 wire clknet_3_2__leaf_spi_sclk;
 wire clknet_3_3__leaf_spi_sclk;
 wire clknet_3_4__leaf_spi_sclk;
 wire clknet_3_5__leaf_spi_sclk;
 wire clknet_3_6__leaf_spi_sclk;
 wire clknet_3_7__leaf_spi_sclk;
 wire clknet_0_u_txreg_sclk_test;
 wire clknet_1_0__leaf_u_txreg_sclk_test;
 wire clknet_1_1__leaf_u_txreg_sclk_test;
 wire clknet_0_u_txreg_net830;
 wire clknet_1_0__leaf_u_txreg_net830;
 wire clknet_1_1__leaf_u_txreg_net830;
 wire clknet_0_u_txreg_net835;
 wire clknet_1_0__leaf_u_txreg_net835;
 wire clknet_1_1__leaf_u_txreg_net835;
 wire clknet_0_u_txreg_net840;
 wire clknet_1_0__leaf_u_txreg_net840;
 wire clknet_1_1__leaf_u_txreg_net840;
 wire clknet_0_u_txreg_net824;
 wire clknet_1_0__leaf_u_txreg_net824;
 wire clknet_1_1__leaf_u_txreg_net824;
 wire clknet_0_u_rxreg_net863;
 wire clknet_1_0__leaf_u_rxreg_net863;
 wire clknet_1_1__leaf_u_rxreg_net863;
 wire clknet_0_u_rxreg_net868;
 wire clknet_1_0__leaf_u_rxreg_net868;
 wire clknet_1_1__leaf_u_rxreg_net868;
 wire clknet_0_u_rxreg_net873;
 wire clknet_1_0__leaf_u_rxreg_net873;
 wire clknet_1_1__leaf_u_rxreg_net873;
 wire clknet_0_u_rxreg_net857;
 wire clknet_1_0__leaf_u_rxreg_net857;
 wire clknet_1_1__leaf_u_rxreg_net857;
 wire clknet_0_u_device_sm_u_spiregs_net791;
 wire clknet_1_0__leaf_u_device_sm_u_spiregs_net791;
 wire clknet_1_1__leaf_u_device_sm_u_spiregs_net791;
 wire clknet_0_u_device_sm_u_spiregs_net807;
 wire clknet_1_0__leaf_u_device_sm_u_spiregs_net807;
 wire clknet_1_1__leaf_u_device_sm_u_spiregs_net807;
 wire clknet_0_u_device_sm_u_spiregs_net802;
 wire clknet_1_0__leaf_u_device_sm_u_spiregs_net802;
 wire clknet_1_1__leaf_u_device_sm_u_spiregs_net802;
 wire clknet_0_u_device_sm_u_spiregs_net797;
 wire clknet_1_0__leaf_u_device_sm_u_spiregs_net797;
 wire clknet_1_1__leaf_u_device_sm_u_spiregs_net797;
 wire clknet_0_u_device_sm_net774;
 wire clknet_1_0__leaf_u_device_sm_net774;
 wire clknet_1_1__leaf_u_device_sm_net774;
 wire clknet_0_u_device_sm_net763;
 wire clknet_1_0__leaf_u_device_sm_net763;
 wire clknet_1_1__leaf_u_device_sm_net763;
 wire clknet_0_u_device_sm_net769;
 wire clknet_1_0__leaf_u_device_sm_net769;
 wire clknet_1_1__leaf_u_device_sm_net769;
 wire clknet_0_u_dcfifo_tx_u_dout_read_tr_net634;
 wire clknet_1_0__leaf_u_dcfifo_tx_u_dout_read_tr_net634;
 wire clknet_1_1__leaf_u_dcfifo_tx_u_dout_read_tr_net634;
 wire clknet_0_u_dcfifo_rx_u_din_write_tr_net652;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_write_tr_net652;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_write_tr_net652;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net670;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net670;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net670;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net676;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net676;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net676;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net681;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net681;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net681;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net686;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net686;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net686;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net691;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net691;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net691;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net696;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net696;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net696;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net701;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net701;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net701;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net706;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net706;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net706;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net711;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net711;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net711;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net716;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net716;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net716;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net721;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net721;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net721;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net726;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net726;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net726;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net731;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net731;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net731;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net736;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net736;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net736;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net741;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net741;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net741;
 wire clknet_0_u_dcfifo_rx_u_din_buffer_net746;
 wire clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net746;
 wire clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net746;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire [31:0] addr_sync;
 wire [31:0] ctrl_data_rx;
 wire [7:0] tx_counter;
 wire [31:0] tx_data;
 wire [255:0] u_dcfifo_rx_u_din_buffer_data;
 wire [7:0] u_dcfifo_rx_u_dout_empty_synch_d_middle;
 wire [7:0] u_dcfifo_rx_u_dout_read_token;
 wire [7:0] u_dcfifo_rx_u_dout_write_token_dn;
 wire [7:0] u_dcfifo_rx_write_token;
 wire [255:0] u_dcfifo_tx_u_din_buffer_data;
 wire [7:0] u_dcfifo_tx_u_dout_empty_synch_d_middle;
 wire [7:0] u_dcfifo_tx_u_dout_read_token;
 wire [7:0] u_dcfifo_tx_u_dout_write_token_dn;
 wire [7:0] u_dcfifo_tx_write_token;
 wire [7:0] u_device_sm_cmd_reg;
 wire [7:0] u_device_sm_s_dummy_cycles;
 wire [2:0] u_device_sm_state;
 wire [2:0] u_device_sm_state_next;
 wire [16:0] u_device_sm_u_spiregs_n;
 wire [7:0] u_device_sm_u_spiregs_reg0;
 wire [7:0] u_rxreg_counter;
 wire [7:0] u_rxreg_counter_trgt;
 wire [7:0] u_rxreg_counter_trgt_next;
 wire [31:0] u_rxreg_data_int;
 wire [1:0] u_spi_device_tlul_plug_state;
 wire [1:0] u_spi_device_tlul_plug_state_next;
 wire [31:0] u_spi_device_tlul_plug_wdata_next;
 wire [2:0] u_syncro_valid_reg;
 wire [7:0] u_txreg_counter;
 wire [7:0] u_txreg_counter_trgt;
 wire [31:0] u_txreg_data_int;

 b15mbn022ar1n02x5 U2913 (.a(clknet_3_0__leaf_spi_sclk),
    .b(net1954),
    .o(u_txreg_sclk_test),
    .sa(net7));
 b15inv040as1n40x5 U2914 (.a(net2),
    .o1(n3769));
 b15inv000as1n28x5 U2915 (.a(net426),
    .o1(n3770));
 b15inv000as1n64x5 U2916 (.a(net426),
    .o1(n3771));
 b15inv020ah1n24x5 U2917 (.a(net2364),
    .o1(n2729));
 b15inv020as1n24x5 U2918 (.a(u_rxreg_data_int[4]),
    .o1(n2787));
 b15inv000as1n80x5 U2919 (.a(net2),
    .o1(n3772));
 b15aoi022ah1n32x5 U2920 (.a(net298),
    .b(n2729),
    .c(n2787),
    .d(net263),
    .o1(u_rxreg_N34));
 b15inv020ah1n80x5 U2921 (.a(net427),
    .o1(n3773));
 b15inv040aq1n05x5 U2922 (.a(u_rxreg_data_int[3]),
    .o1(n2726));
 b15inv040aq1n60x5 U2923 (.a(net426),
    .o1(n3774));
 b15inv000ar1n03x5 U2924 (.a(net466),
    .o1(tl_o[0]));
 b15inv000as1n80x5 U2925 (.a(net426),
    .o1(n3776));
 b15aoi022as1n08x5 U2926 (.a(net298),
    .b(net6),
    .c(u_rxreg_data_int[2]),
    .d(n3817),
    .o1(n2778));
 b15inv040as1n48x5 U2927 (.a(net2),
    .o1(n3777));
 b15inv000as1n48x5 U2928 (.a(net427),
    .o1(n3778));
 b15aoi022ah1n12x5 U2929 (.a(net346),
    .b(n2726),
    .c(n2778),
    .d(n3807),
    .o1(ctrl_data_rx[3]));
 b15inv000ar1n16x5 U2931 (.a(net2350),
    .o1(n2798));
 b15aoi022as1n08x5 U2932 (.a(net298),
    .b(n2726),
    .c(n2798),
    .d(n3817),
    .o1(u_rxreg_N36));
 b15ztpn00an1n08x5 PHY_95 ();
 b15oa0022aq1n06x5 U2934 (.a(n3809),
    .b(u_rxreg_data_int[7]),
    .c(u_rxreg_N36),
    .d(net349),
    .o(ctrl_data_rx[7]));
 b15ztpn00an1n08x5 PHY_94 ();
 b15oai022al1n08x5 U2936 (.a(n3817),
    .b(u_rxreg_data_int[2]),
    .c(net294),
    .d(net298),
    .o1(n2776));
 b15aoi022aq1n12x5 U2937 (.a(net346),
    .b(n2798),
    .c(n2776),
    .d(n3807),
    .o1(ctrl_data_rx[6]));
 b15nand02aq1n04x5 U2938 (.a(net296),
    .b(net4),
    .o1(n2727));
 b15aob012al1n12x5 U2939 (.a(n2727),
    .b(n3817),
    .c(u_rxreg_data_int[0]),
    .out0(u_rxreg_N30));
 b15ztpn00an1n08x5 PHY_93 ();
 b15aboi22as1n24x5 U2941 (.a(u_rxreg_N30),
    .b(n3807),
    .c(net346),
    .d(n2729),
    .out0(ctrl_data_rx[1]));
 b15nandp2ar1n05x5 U2942 (.a(net296),
    .b(net5),
    .o1(n2728));
 b15oai012aq1n16x5 U2943 (.a(n2728),
    .b(net296),
    .c(n2729),
    .o1(u_rxreg_N31));
 b15oa0022al1n32x5 U2944 (.a(n3809),
    .b(u_rxreg_data_int[2]),
    .c(u_rxreg_N31),
    .d(net346),
    .o(ctrl_data_rx[2]));
 b15oai022an1n24x5 U2945 (.a(n3817),
    .b(u_rxreg_data_int[0]),
    .c(u_rxreg_data_int[3]),
    .d(net298),
    .o1(n2777));
 b15aoi022as1n48x5 U2946 (.a(net346),
    .b(n2787),
    .c(n2777),
    .d(n3807),
    .o1(ctrl_data_rx[4]));
 b15inv040as1n06x5 U2947 (.a(u_rxreg_counter_trgt[4]),
    .o1(n2871));
 b15inv000ar1n05x5 U2948 (.a(u_rxreg_counter_trgt[6]),
    .o1(n2731));
 b15aoi022an1n06x5 U2949 (.a(n2871),
    .b(u_rxreg_counter[4]),
    .c(u_rxreg_counter[6]),
    .d(n2731),
    .o1(n2730));
 b15oai122ah1n12x5 U2950 (.a(n2730),
    .b(n2871),
    .c(u_rxreg_counter[4]),
    .d(n2731),
    .e(u_rxreg_counter[6]),
    .o1(n2742));
 b15inv020ah1n10x5 U2951 (.a(u_rxreg_counter_trgt[0]),
    .o1(n2874));
 b15inv000ah1n04x5 U2952 (.a(u_rxreg_counter_trgt[2]),
    .o1(n2733));
 b15aoi022ah1n06x5 U2953 (.a(n2874),
    .b(u_rxreg_counter[0]),
    .c(u_rxreg_counter[2]),
    .d(n2733),
    .o1(n2732));
 b15oai122as1n16x5 U2954 (.a(n2732),
    .b(n2874),
    .c(u_rxreg_counter[0]),
    .d(n2733),
    .e(u_rxreg_counter[2]),
    .o1(n2741));
 b15inv020an1n06x5 U2955 (.a(u_rxreg_counter_trgt[5]),
    .o1(n2736));
 b15inv000ah1n04x5 U2956 (.a(u_rxreg_counter_trgt[1]),
    .o1(n2735));
 b15aoi022an1n04x5 U2957 (.a(n2736),
    .b(u_rxreg_counter[5]),
    .c(u_rxreg_counter[1]),
    .d(n2735),
    .o1(n2734));
 b15oai122aq1n12x5 U2958 (.a(n2734),
    .b(n2736),
    .c(u_rxreg_counter[5]),
    .d(n2735),
    .e(u_rxreg_counter[1]),
    .o1(n2740));
 b15inv020as1n05x5 U2959 (.a(u_rxreg_counter_trgt[7]),
    .o1(n2738));
 b15inv040as1n06x5 U2960 (.a(u_rxreg_counter_trgt[3]),
    .o1(n2870));
 b15aoi022ah1n04x5 U2961 (.a(n2738),
    .b(u_rxreg_counter[7]),
    .c(u_rxreg_counter[3]),
    .d(n2870),
    .o1(n2737));
 b15oai122al1n16x5 U2962 (.a(n2737),
    .b(n2738),
    .c(u_rxreg_counter[7]),
    .d(n2870),
    .e(u_rxreg_counter[3]),
    .o1(n2739));
 b15nor004as1n12x5 U2963 (.a(n2742),
    .b(n2741),
    .c(n2740),
    .d(n2739),
    .o1(n2781));
 b15inv000as1n20x5 U2964 (.a(n2781),
    .o1(n2868));
 b15norp02ah1n48x5 U2965 (.a(n2868),
    .b(n1869),
    .o1(n2878));
 b15inv000ar1n24x5 U2966 (.a(net355),
    .o1(n2840));
 b15inv020aq1n16x5 U2967 (.a(net359),
    .o1(n2841));
 b15nandp2as1n24x5 U2968 (.a(n2840),
    .b(n2841),
    .o1(n2876));
 b15norp02aq1n48x5 U2969 (.a(n2876),
    .b(net358),
    .o1(n2750));
 b15ztpn00an1n08x5 PHY_92 ();
 b15oai022as1n48x5 U2971 (.a(n3811),
    .b(net293),
    .c(u_rxreg_N34),
    .d(net346),
    .o1(n2802));
 b15nand02ar1n12x5 U2972 (.a(n3819),
    .b(u_device_sm_cmd_reg[5]),
    .o1(n2743));
 b15oai012ah1n12x5 U2973 (.a(n2743),
    .b(n3819),
    .c(n2802),
    .o1(n2751));
 b15inv020as1n08x5 U2974 (.a(n2751),
    .o1(n2746));
 b15nandp2ah1n05x5 U2975 (.a(n3819),
    .b(u_device_sm_cmd_reg[3]),
    .o1(n2744));
 b15aob012as1n24x5 U2976 (.a(n2744),
    .b(n2750),
    .c(net246),
    .out0(n2832));
 b15norp02al1n32x5 U2977 (.a(n2746),
    .b(n2832),
    .o1(n2858));
 b15oai022an1n08x5 U2978 (.a(n3811),
    .b(u_rxreg_data_int[0]),
    .c(net3),
    .d(net346),
    .o1(n2783));
 b15nandp2as1n05x5 U2979 (.a(n3819),
    .b(u_device_sm_cmd_reg[0]),
    .o1(n2745));
 b15oai012ah1n24x5 U2980 (.a(n2745),
    .b(n3819),
    .c(net264),
    .o1(n2833));
 b15inv000ah1n03x5 U2981 (.a(n2833),
    .o1(n2748));
 b15qgbna2an1n10x5 U2982 (.a(n2833),
    .b(n2746),
    .o1(n2831));
 b15norp02ar1n16x5 U2983 (.a(n2832),
    .b(n2831),
    .o1(n2826));
 b15orn003ah1n02x5 U2984 (.a(n3819),
    .b(net243),
    .c(net240),
    .o(n2747));
 b15oai013as1n12x5 U2985 (.a(n2747),
    .b(n2750),
    .c(u_device_sm_cmd_reg[7]),
    .d(u_device_sm_cmd_reg[6]),
    .o1(n2825));
 b15aoi022ar1n24x5 U2986 (.a(n2750),
    .b(net238),
    .c(u_device_sm_cmd_reg[1]),
    .d(n3819),
    .o1(n2822));
 b15aoi022ah1n24x5 U2987 (.a(n2750),
    .b(net235),
    .c(u_device_sm_cmd_reg[2]),
    .d(n3819),
    .o1(n2837));
 b15nand02ar1n16x5 U2988 (.a(n2822),
    .b(n2837),
    .o1(n2828));
 b15nonb02as1n16x5 U2989 (.a(n2825),
    .b(n2828),
    .out0(n2859));
 b15aoai13as1n08x5 U2990 (.a(n2859),
    .b(n2826),
    .c(n2858),
    .d(n2748),
    .o1(n2839));
 b15inv040an1n08x5 U2991 (.a(n2839),
    .o1(n2853));
 b15nandp2ah1n05x5 U2992 (.a(n3819),
    .b(u_device_sm_cmd_reg[4]),
    .o1(n2749));
 b15aob012ah1n24x5 U2993 (.a(n2749),
    .b(n2750),
    .c(net234),
    .out0(n2836));
 b15nor002aq1n04x5 U2994 (.a(n2822),
    .b(n2836),
    .o1(n2824));
 b15nand03aq1n16x5 U2995 (.a(n2837),
    .b(n2824),
    .c(n2825),
    .o1(n2830));
 b15nor004as1n12x5 U2996 (.a(n2833),
    .b(n2832),
    .c(n2751),
    .d(n2830),
    .o1(n2880));
 b15nor002ar1n24x5 U2997 (.a(n2853),
    .b(n2880),
    .o1(n2847));
 b15inv000aq1n20x5 U2998 (.a(net356),
    .o1(n2852));
 b15norp03as1n24x5 U2999 (.a(net360),
    .b(n2840),
    .c(n2852),
    .o1(n2890));
 b15nand03as1n24x5 U3000 (.a(n2878),
    .b(n2847),
    .c(n2890),
    .o1(n2877));
 b15nor002an1n08x5 U3001 (.a(n3813),
    .b(n2877),
    .o1(u_device_sm_N163));
 b15cbf000an1n16x5 clkbuf_0_clk_i (.clk(clk_i),
    .clkout(clknet_0_clk_i));
 b15ztpn00an1n08x5 PHY_91 ();
 b15ztpn00an1n08x5 PHY_90 ();
 b15ztpn00an1n08x5 PHY_89 ();
 b15ztpn00an1n08x5 PHY_88 ();
 b15ztpn00an1n08x5 PHY_87 ();
 b15ztpn00an1n08x5 PHY_86 ();
 b15ztpn00an1n08x5 PHY_85 ();
 b15ztpn00an1n08x5 PHY_84 ();
 b15ztpn00an1n08x5 PHY_83 ();
 b15ztpn00an1n08x5 PHY_82 ();
 b15ztpn00an1n08x5 PHY_81 ();
 b15ztpn00an1n08x5 PHY_80 ();
 b15ztpn00an1n08x5 PHY_79 ();
 b15ztpn00an1n08x5 PHY_78 ();
 b15ztpn00an1n08x5 PHY_77 ();
 b15ztpn00an1n08x5 PHY_76 ();
 b15ztpn00an1n08x5 PHY_75 ();
 b15ztpn00an1n08x5 PHY_74 ();
 b15ztpn00an1n08x5 PHY_73 ();
 b15ztpn00an1n08x5 PHY_72 ();
 b15ztpn00an1n08x5 PHY_71 ();
 b15ztpn00an1n08x5 PHY_70 ();
 b15ztpn00an1n08x5 PHY_69 ();
 b15inv000as1n80x5 U3026 (.a(net345),
    .o1(n3807));
 b15ztpn00an1n08x5 PHY_68 ();
 b15inv000ah1n64x5 U3028 (.a(net350),
    .o1(n3809));
 b15inv000ar1n03x5 U3029 (.a(net1450),
    .o1(tl_o[1]));
 b15qgbin1an1n40x5 U3030 (.a(net346),
    .o1(n3811));
 b15ztpn00an1n08x5 PHY_67 ();
 b15inv000as1n56x5 U3032 (.a(net300),
    .o1(n3813));
 b15inv000ah1n32x5 U3034 (.a(net296),
    .o1(n3815));
 b15inv000ar1n03x5 U3035 (.a(net467),
    .o1(tl_o[2]));
 b15inv000aq1n80x5 U3036 (.a(net298),
    .o1(n3817));
 b15inv000as1n32x5 U3037 (.a(net264),
    .o1(n3818));
 b15inv040ah1n36x5 U3038 (.a(n2750),
    .o1(n3819));
 b15inv000as1n56x5 U3039 (.a(n2802),
    .o1(n3820));
 b15inv000al1n10x5 U3040 (.a(n3664),
    .o1(n3821));
 b15inv020aq1n10x5 U3041 (.a(n3681),
    .o1(n3822));
 b15inv000ar1n03x5 U3043 (.a(net1451),
    .o1(tl_o[3]));
 b15inv000ar1n03x5 U3045 (.a(net468),
    .o1(tl_o[4]));
 b15inv000ar1n03x5 U3047 (.a(net1452),
    .o1(tl_o[5]));
 b15nand02aq1n24x5 U3049 (.a(net307),
    .b(net306),
    .o1(n3645));
 b15nor002as1n03x5 U3050 (.a(u_dcfifo_tx_u_dout_write_token_dn[1]),
    .b(n3645),
    .o1(n2775));
 b15inv020ah1n03x5 U3051 (.a(u_dcfifo_tx_u_dout_write_token_dn[5]),
    .o1(n2765));
 b15nandp2ah1n08x5 U3052 (.a(u_dcfifo_tx_u_dout_read_token[4]),
    .b(u_dcfifo_tx_u_dout_read_token[5]),
    .o1(n3647));
 b15inv000ah1n08x5 U3053 (.a(n3647),
    .o1(n3001));
 b15and003al1n04x5 U3054 (.a(n2765),
    .b(n3001),
    .c(u_dcfifo_tx_u_dout_write_token_dn[6]),
    .o(n2774));
 b15nand02al1n12x5 U3055 (.a(net306),
    .b(u_dcfifo_tx_u_dout_read_token[2]),
    .o1(n3638));
 b15inv040aq1n05x5 U3056 (.a(n3638),
    .o1(n3635));
 b15inv000al1n02x5 U3057 (.a(u_dcfifo_tx_u_dout_write_token_dn[2]),
    .o1(n2764));
 b15nandp2an1n08x5 U3058 (.a(u_dcfifo_tx_u_dout_read_token[5]),
    .b(u_dcfifo_tx_u_dout_read_token[6]),
    .o1(n3653));
 b15nonb03al1n02x5 U3059 (.a(u_dcfifo_tx_u_dout_write_token_dn[7]),
    .b(u_dcfifo_tx_u_dout_write_token_dn[6]),
    .c(n3653),
    .out0(n2763));
 b15aoi013al1n03x5 U3060 (.a(n2763),
    .b(n3635),
    .c(u_dcfifo_tx_u_dout_write_token_dn[3]),
    .d(n2764),
    .o1(n2772));
 b15nandp2as1n05x5 U3061 (.a(u_dcfifo_tx_u_dout_read_token[2]),
    .b(net305),
    .o1(n3637));
 b15inv020ah1n04x5 U3062 (.a(n3637),
    .o1(n3650));
 b15inv000al1n02x5 U3063 (.a(u_dcfifo_tx_u_dout_write_token_dn[3]),
    .o1(n2767));
 b15nandp2as1n12x5 U3064 (.a(u_dcfifo_tx_u_dout_read_token[4]),
    .b(net305),
    .o1(n3640));
 b15norp03ar1n02x5 U3065 (.a(u_dcfifo_tx_u_dout_write_token_dn[4]),
    .b(n2765),
    .c(n3640),
    .o1(n2766));
 b15aoi013aq1n02x5 U3066 (.a(n2766),
    .b(n3650),
    .c(u_dcfifo_tx_u_dout_write_token_dn[4]),
    .d(n2767),
    .o1(n2771));
 b15nand02as1n48x5 U3067 (.a(net307),
    .b(net303),
    .o1(n3008));
 b15inv020aq1n16x5 U3068 (.a(n3008),
    .o1(n3633));
 b15inv000as1n02x5 U3069 (.a(net2351),
    .o1(n2769));
 b15nandp2ah1n05x5 U3070 (.a(net304),
    .b(u_dcfifo_tx_u_dout_read_token[6]),
    .o1(n3641));
 b15oai013aq1n02x5 U3071 (.a(ctrl_data_tx_ready),
    .b(u_dcfifo_tx_u_dout_write_token_dn[7]),
    .c(n3641),
    .d(n2769),
    .o1(n2768));
 b15aoi013ar1n03x5 U3072 (.a(n2768),
    .b(n3633),
    .c(u_dcfifo_tx_u_dout_write_token_dn[1]),
    .d(n2769),
    .o1(n2770));
 b15nand03ah1n06x5 U3073 (.a(n2772),
    .b(n2771),
    .c(n2770),
    .o1(n2773));
 b15aoi112ah1n08x5 U3074 (.a(n2774),
    .b(net2352),
    .c(n2775),
    .d(u_dcfifo_tx_u_dout_write_token_dn[2]),
    .o1(u_dcfifo_tx_u_dout_read_enable));
 b15nand02an1n32x5 U3075 (.a(n2840),
    .b(net2089),
    .o1(n2842));
 b15norp02an1n24x5 U3076 (.a(n2852),
    .b(net2090),
    .o1(n2860));
 b15nor002ah1n16x5 U3077 (.a(net2091),
    .b(n3813),
    .o1(net56));
 b15oai022as1n16x5 U3078 (.a(net263),
    .b(u_rxreg_data_int[25]),
    .c(u_rxreg_data_int[28]),
    .d(net297),
    .o1(n2784));
 b15inv020as1n06x5 U3079 (.a(n2784),
    .o1(u_rxreg_N58));
 b15inv000as1n02x5 U3080 (.a(n2776),
    .o1(u_rxreg_N35));
 b15inv040ar1n03x5 U3081 (.a(n2777),
    .o1(u_rxreg_N33));
 b15norp02ah1n04x5 U3082 (.a(u_rxreg_counter[0]),
    .b(n2781),
    .o1(u_rxreg_N22));
 b15oai022as1n06x5 U3083 (.a(n3817),
    .b(u_rxreg_data_int[20]),
    .c(u_rxreg_data_int[23]),
    .d(net297),
    .o1(n2811));
 b15inv020aq1n03x5 U3084 (.a(n2811),
    .o1(u_rxreg_N53));
 b15oai022an1n24x5 U3085 (.a(n3817),
    .b(u_rxreg_data_int[22]),
    .c(u_rxreg_data_int[25]),
    .d(net297),
    .o1(n2807));
 b15inv040aq1n04x5 U3086 (.a(n2807),
    .o1(u_rxreg_N55));
 b15oai022an1n24x5 U3087 (.a(n3817),
    .b(u_rxreg_data_int[17]),
    .c(u_rxreg_data_int[20]),
    .d(net296),
    .o1(n2813));
 b15inv020as1n03x5 U3088 (.a(n2813),
    .o1(u_rxreg_N50));
 b15oai022al1n32x5 U3089 (.a(net263),
    .b(net294),
    .c(net292),
    .d(net298),
    .o1(n2803));
 b15inv040ar1n02x5 U3090 (.a(n2803),
    .o1(u_rxreg_N38));
 b15oai022as1n24x5 U3091 (.a(n3817),
    .b(net295),
    .c(u_rxreg_data_int[17]),
    .d(net296),
    .o1(n2805));
 b15inv000al1n03x5 U3092 (.a(n2805),
    .o1(u_rxreg_N47));
 b15oai022ah1n12x5 U3093 (.a(net263),
    .b(u_rxreg_data_int[8]),
    .c(u_rxreg_data_int[11]),
    .d(net296),
    .o1(n2815));
 b15inv040ar1n03x5 U3094 (.a(n2815),
    .o1(u_rxreg_N41));
 b15oai022as1n16x5 U3095 (.a(net263),
    .b(u_rxreg_data_int[23]),
    .c(u_rxreg_data_int[26]),
    .d(net297),
    .o1(n2809));
 b15inv040as1n02x5 U3096 (.a(n2809),
    .o1(u_rxreg_N56));
 b15oai022an1n24x5 U3097 (.a(n3817),
    .b(u_rxreg_data_int[11]),
    .c(u_rxreg_data_int[14]),
    .d(net296),
    .o1(n2819));
 b15inv000aq1n04x5 U3098 (.a(n2819),
    .o1(u_rxreg_N44));
 b15inv000aq1n02x5 U3099 (.a(n2778),
    .o1(u_rxreg_N32));
 b15inv020an1n03x5 U3100 (.a(u_rxreg_counter[2]),
    .o1(n2779));
 b15nand02aq1n06x5 U3101 (.a(u_rxreg_counter[0]),
    .b(u_rxreg_counter[1]),
    .o1(n2788));
 b15and003al1n08x5 U3102 (.a(u_rxreg_counter[0]),
    .b(u_rxreg_counter[2]),
    .c(u_rxreg_counter[1]),
    .o(n2791));
 b15aoi112ah1n06x5 U3103 (.a(n2791),
    .b(n2781),
    .c(n2779),
    .d(n2788),
    .o1(u_rxreg_N24));
 b15inv040ar1n04x5 U3104 (.a(u_rxreg_counter[4]),
    .o1(n2780));
 b15nandp2an1n08x5 U3105 (.a(u_rxreg_counter[3]),
    .b(n2791),
    .o1(n2790));
 b15nor002ah1n06x5 U3106 (.a(n2780),
    .b(n2790),
    .o1(n2794));
 b15aoi112an1n06x5 U3107 (.a(n2794),
    .b(n2781),
    .c(n2780),
    .d(n2790),
    .o1(u_rxreg_N26));
 b15inv000ah1n02x5 U3108 (.a(u_rxreg_counter[6]),
    .o1(n2782));
 b15nand02an1n08x5 U3109 (.a(u_rxreg_counter[5]),
    .b(n2794),
    .o1(n2793));
 b15norp02ah1n04x5 U3110 (.a(n2782),
    .b(n2793),
    .o1(n2797));
 b15aoi112ah1n03x5 U3111 (.a(n2797),
    .b(n2781),
    .c(n2782),
    .d(n2793),
    .o1(u_rxreg_N28));
 b15nand02an1n16x5 U3112 (.a(net2078),
    .b(net301),
    .o1(n3619));
 b15norp02an1n32x5 U3113 (.a(n2842),
    .b(net2079),
    .o1(net55));
 b15inv000ar1n03x5 U3114 (.a(net469),
    .o1(tl_o[6]));
 b15inv020aq1n10x5 U3115 (.a(u_rxreg_data_int[29]),
    .o1(n2799));
 b15oai022ah1n32x5 U3116 (.a(n3811),
    .b(n2799),
    .c(n2784),
    .d(net345),
    .o1(ctrl_data_rx[29]));
 b15aboi22ah1n16x5 U3118 (.a(u_rxreg_data_int[7]),
    .b(net263),
    .c(net298),
    .d(n2787),
    .out0(u_rxreg_N37));
 b15oa0022as1n32x5 U3119 (.a(u_rxreg_N37),
    .b(net346),
    .c(net292),
    .d(n3807),
    .o(ctrl_data_rx[8]));
 b15inv000ah1n16x5 U3120 (.a(u_rxreg_data_int[27]),
    .o1(n2810));
 b15aboi22as1n08x5 U3121 (.a(net2342),
    .b(net263),
    .c(net297),
    .d(n2810),
    .out0(u_rxreg_N60));
 b15ao0022aq1n24x5 U3122 (.a(u_rxreg_data_int[31]),
    .b(net345),
    .c(u_rxreg_N60),
    .d(n3807),
    .o(ctrl_data_rx[31]));
 b15oai112an1n02x5 U3123 (.a(n2788),
    .b(n2868),
    .c(u_rxreg_counter[0]),
    .d(u_rxreg_counter[1]),
    .o1(n2789));
 b15inv040as1n02x5 U3124 (.a(n2789),
    .o1(u_rxreg_N23));
 b15oai112aq1n16x5 U3125 (.a(n2790),
    .b(n2868),
    .c(u_rxreg_counter[3]),
    .d(n2791),
    .o1(n2792));
 b15inv020an1n03x5 U3126 (.a(n2792),
    .o1(u_rxreg_N25));
 b15oai112aq1n16x5 U3127 (.a(n2793),
    .b(n2868),
    .c(u_rxreg_counter[5]),
    .d(n2794),
    .o1(n2795));
 b15inv020ar1n04x5 U3128 (.a(n2795),
    .o1(u_rxreg_N27));
 b15oa0022al1n12x5 U3129 (.a(net263),
    .b(u_rxreg_data_int[7]),
    .c(u_rxreg_data_int[10]),
    .d(net296),
    .o(u_rxreg_N40));
 b15oa0022aq1n24x5 U3130 (.a(u_rxreg_N40),
    .b(net346),
    .c(u_rxreg_data_int[11]),
    .d(n3807),
    .o(ctrl_data_rx[11]));
 b15oa0022ah1n06x5 U3131 (.a(n3815),
    .b(u_rxreg_data_int[16]),
    .c(u_rxreg_data_int[19]),
    .d(net297),
    .o(u_rxreg_N49));
 b15oa0022as1n16x5 U3132 (.a(n3809),
    .b(u_rxreg_data_int[20]),
    .c(u_rxreg_N49),
    .d(net346),
    .o(ctrl_data_rx[20]));
 b15oa0022al1n08x5 U3133 (.a(n3815),
    .b(u_rxreg_data_int[13]),
    .c(u_rxreg_data_int[16]),
    .d(net296),
    .o(u_rxreg_N46));
 b15oa0022ar1n08x5 U3134 (.a(n3809),
    .b(u_rxreg_data_int[17]),
    .c(u_rxreg_N46),
    .d(net345),
    .o(ctrl_data_rx[17]));
 b15oa0022as1n06x5 U3135 (.a(n3815),
    .b(u_rxreg_data_int[19]),
    .c(u_rxreg_data_int[22]),
    .d(net297),
    .o(u_rxreg_N52));
 b15oa0022al1n24x5 U3136 (.a(n3809),
    .b(u_rxreg_data_int[23]),
    .c(u_rxreg_N52),
    .d(net348),
    .o(ctrl_data_rx[23]));
 b15oa0022ar1n12x5 U3137 (.a(n3815),
    .b(u_rxreg_data_int[10]),
    .c(u_rxreg_data_int[13]),
    .d(net296),
    .o(u_rxreg_N43));
 b15oa0022al1n24x5 U3138 (.a(n3809),
    .b(net295),
    .c(u_rxreg_N43),
    .d(net345),
    .o(ctrl_data_rx[14]));
 b15oai012ar1n03x5 U3139 (.a(n2868),
    .b(u_rxreg_counter[7]),
    .c(n2797),
    .o1(n2796));
 b15aoi012as1n02x5 U3140 (.a(n2796),
    .b(net2370),
    .c(n2797),
    .o1(u_rxreg_N29));
 b15inv000an1n28x5 U3141 (.a(u_rxreg_data_int[18]),
    .o1(n2806));
 b15inv000ah1n16x5 U3142 (.a(u_rxreg_data_int[21]),
    .o1(n2814));
 b15aoi022an1n24x5 U3143 (.a(net296),
    .b(n2806),
    .c(n2814),
    .d(n3817),
    .o1(u_rxreg_N51));
 b15oa0022ar1n32x5 U3144 (.a(n3809),
    .b(u_rxreg_data_int[22]),
    .c(u_rxreg_N51),
    .d(net346),
    .o(ctrl_data_rx[22]));
 b15inv040as1n16x5 U3145 (.a(net2339),
    .o1(n2804));
 b15aoi022aq1n32x5 U3146 (.a(net298),
    .b(n2798),
    .c(n2804),
    .d(n3817),
    .o1(u_rxreg_N39));
 b15oa0022aq1n24x5 U3147 (.a(n3809),
    .b(u_rxreg_data_int[10]),
    .c(u_rxreg_N39),
    .d(net345),
    .o(ctrl_data_rx[10]));
 b15inv020aq1n28x5 U3148 (.a(u_rxreg_data_int[15]),
    .o1(n2820));
 b15aoi022al1n32x5 U3149 (.a(net296),
    .b(n2820),
    .c(n2806),
    .d(n3817),
    .o1(u_rxreg_N48));
 b15oa0022al1n24x5 U3150 (.a(n3809),
    .b(u_rxreg_data_int[19]),
    .c(u_rxreg_N48),
    .d(net345),
    .o(ctrl_data_rx[19]));
 b15inv040as1n08x5 U3151 (.a(net2333),
    .o1(n2816));
 b15aoi022aq1n12x5 U3152 (.a(net296),
    .b(n2804),
    .c(n2816),
    .d(net263),
    .o1(u_rxreg_N42));
 b15oa0022ah1n12x5 U3153 (.a(n3809),
    .b(u_rxreg_data_int[13]),
    .c(u_rxreg_N42),
    .d(net346),
    .o(ctrl_data_rx[13]));
 b15aoi022an1n16x5 U3154 (.a(net296),
    .b(n2816),
    .c(n2820),
    .d(net263),
    .o1(u_rxreg_N45));
 b15oa0022an1n24x5 U3155 (.a(n3809),
    .b(u_rxreg_data_int[16]),
    .c(u_rxreg_N45),
    .d(net345),
    .o(ctrl_data_rx[16]));
 b15inv000as1n10x5 U3156 (.a(net2354),
    .o1(n2812));
 b15aoi022an1n12x5 U3157 (.a(net297),
    .b(n2814),
    .c(n2812),
    .d(n3815),
    .o1(u_rxreg_N54));
 b15oa0022ar1n04x5 U3158 (.a(n3809),
    .b(u_rxreg_data_int[25]),
    .c(u_rxreg_N54),
    .d(net345),
    .o(ctrl_data_rx[25]));
 b15inv040ah1n08x5 U3159 (.a(u_rxreg_data_int[26]),
    .o1(n2808));
 b15aoi022aq1n12x5 U3160 (.a(net297),
    .b(n2808),
    .c(n2799),
    .d(net263),
    .o1(u_rxreg_N59));
 b15ao0022aq1n16x5 U3161 (.a(net345),
    .b(net2514),
    .c(u_rxreg_N59),
    .d(n3811),
    .o(ctrl_data_rx[30]));
 b15aoi022al1n32x5 U3162 (.a(net297),
    .b(n2812),
    .c(n2810),
    .d(n3815),
    .o1(u_rxreg_N57));
 b15ao0022aq1n16x5 U3163 (.a(net345),
    .b(u_rxreg_data_int[28]),
    .c(u_rxreg_N57),
    .d(n3811),
    .o(ctrl_data_rx[28]));
 b15inv000ar1n03x5 U3164 (.a(net1453),
    .o1(tl_o[7]));
 b15aoi022as1n48x5 U3165 (.a(net345),
    .b(n2804),
    .c(n2803),
    .d(n3807),
    .o1(ctrl_data_rx[9]));
 b15aoi022ah1n48x5 U3166 (.a(net345),
    .b(n2806),
    .c(n2805),
    .d(n3807),
    .o1(ctrl_data_rx[18]));
 b15aoi022an1n48x5 U3167 (.a(net345),
    .b(n2808),
    .c(n2807),
    .d(n3807),
    .o1(ctrl_data_rx[26]));
 b15aoi022an1n48x5 U3168 (.a(net346),
    .b(n2810),
    .c(n2809),
    .d(n3807),
    .o1(ctrl_data_rx[27]));
 b15aoi022as1n04x5 U3169 (.a(net346),
    .b(n2812),
    .c(n2811),
    .d(n3807),
    .o1(ctrl_data_rx[24]));
 b15aoi022ah1n48x5 U3170 (.a(net347),
    .b(n2814),
    .c(n2813),
    .d(n3807),
    .o1(ctrl_data_rx[21]));
 b15aoi022an1n32x5 U3171 (.a(net345),
    .b(n2816),
    .c(n2815),
    .d(n3811),
    .o1(ctrl_data_rx[12]));
 b15aoi022as1n48x5 U3172 (.a(net345),
    .b(n2820),
    .c(n2819),
    .d(n3807),
    .o1(ctrl_data_rx[15]));
 b15inv020aq1n32x5 U3173 (.a(n2878),
    .o1(n2862));
 b15nandp3as1n24x5 U3174 (.a(net355),
    .b(n2852),
    .c(n2841),
    .o1(n2889));
 b15norp02as1n32x5 U3175 (.a(n2862),
    .b(n2889),
    .o1(n2865));
 b15inv020ah1n16x5 U3176 (.a(n2865),
    .o1(n2898));
 b15inv020an1n16x5 U3177 (.a(n2836),
    .o1(n2829));
 b15nand04as1n16x5 U3178 (.a(n2826),
    .b(n2822),
    .c(n2829),
    .d(n2825),
    .o1(n3228));
 b15nor002ah1n04x5 U3179 (.a(n2898),
    .b(n3228),
    .o1(u_device_sm_u_spiregs_N32));
 b15nand02ar1n32x5 U3180 (.a(n2858),
    .b(n2859),
    .o1(n2823));
 b15nor002as1n24x5 U3181 (.a(n2829),
    .b(n2823),
    .o1(n3665));
 b15and002ar1n03x5 U3182 (.a(n3665),
    .b(n2865),
    .o(u_device_sm_u_spiregs_N31));
 b15nor002al1n32x5 U3183 (.a(n2836),
    .b(n2823),
    .o1(n3663));
 b15and002ar1n04x5 U3184 (.a(n3663),
    .b(n2865),
    .o(u_device_sm_u_spiregs_N34));
 b15nanb02as1n02x5 U3185 (.a(n2837),
    .b(n2824),
    .out0(n2827));
 b15nand02aq1n08x5 U3186 (.a(n2826),
    .b(n2825),
    .o1(n2835));
 b15oaoi13as1n08x5 U3187 (.a(n2835),
    .b(n2827),
    .c(n2829),
    .d(n2828),
    .o1(n3664));
 b15qgbno2an1n05x5 U3189 (.o1(u_device_sm_u_spiregs_N33),
    .a(n2898),
    .b(n3821));
 b15nanb02al1n24x5 U3190 (.a(n2876),
    .b(net357),
    .out0(n2879));
 b15inv000ah1n08x5 U3191 (.a(net2332),
    .o1(n3194));
 b15norp02an1n24x5 U3192 (.a(net356),
    .b(n2842),
    .o1(n2891));
 b15inv020ah1n16x5 U3193 (.a(n2891),
    .o1(n2851));
 b15nonb03as1n12x5 U3194 (.a(n2832),
    .b(n2831),
    .c(n2830),
    .out0(n2886));
 b15inv020aq1n10x5 U3195 (.a(n2886),
    .o1(n2846));
 b15norp02al1n24x5 U3196 (.a(n2862),
    .b(n2846),
    .o1(n3611));
 b15inv020ah1n16x5 U3197 (.a(n3611),
    .o1(n3613));
 b15oaoi13as1n08x5 U3198 (.a(n3613),
    .b(n2851),
    .c(n2879),
    .d(n3194),
    .o1(u_rxreg_counter_trgt_next[5]));
 b15aoi013ah1n04x5 U3199 (.a(n2886),
    .b(n2858),
    .c(n2833),
    .d(n2859),
    .o1(n2834));
 b15oai013as1n12x5 U3200 (.a(n2834),
    .b(n2837),
    .c(n2836),
    .d(n2835),
    .o1(ctrl_rd_wr));
 b15norp02al1n24x5 U3201 (.a(n2862),
    .b(n3819),
    .o1(u_device_sm_sample_CMD));
 b15inv000as1n08x5 U3202 (.a(ctrl_rd_wr),
    .o1(n2845));
 b15nandp2ar1n12x5 U3203 (.a(n2891),
    .b(n2878),
    .o1(n2856));
 b15norp02as1n03x5 U3204 (.a(n2878),
    .b(n2879),
    .o1(n2838));
 b15nor002ah1n16x5 U3205 (.a(n2880),
    .b(n2886),
    .o1(n3617));
 b15nandp2an1n05x5 U3206 (.a(n3617),
    .b(u_device_sm_tx_done_reg),
    .o1(n2861));
 b15and003ar1n08x5 U3207 (.a(net360),
    .b(net356),
    .c(n2861),
    .o(n2849));
 b15aoi112an1n06x5 U3208 (.a(n2838),
    .b(n2849),
    .c(u_device_sm_sample_CMD),
    .d(n2839),
    .o1(n2844));
 b15aoi012al1n12x5 U3209 (.a(n2840),
    .b(n2878),
    .c(n2841),
    .o1(n3618));
 b15oai112al1n12x5 U3210 (.a(net357),
    .b(n2842),
    .c(n2847),
    .d(n3618),
    .o1(n2843));
 b15oai112ah1n16x5 U3211 (.a(n2844),
    .b(n2843),
    .c(n2845),
    .d(n2856),
    .o1(u_device_sm_state_next[0]));
 b15norp02aq1n08x5 U3212 (.a(n2879),
    .b(n2862),
    .o1(u_device_sm_sample_ADDR));
 b15nandp2an1n24x5 U3213 (.a(n2846),
    .b(ctrl_rd_wr),
    .o1(n3627));
 b15inv040aq1n05x5 U3214 (.a(u_device_sm_sample_ADDR),
    .o1(n2857));
 b15inv020an1n16x5 U3215 (.a(n2847),
    .o1(n3620));
 b15norp02ah1n16x5 U3216 (.a(n2886),
    .b(n3620),
    .o1(n3632));
 b15aobi12aq1n08x5 U3217 (.a(n2877),
    .b(u_device_sm_sample_CMD),
    .c(n3632),
    .out0(n2855));
 b15oaoi13ar1n08x5 U3218 (.a(n2851),
    .b(n2878),
    .c(n2886),
    .d(n3620),
    .o1(n2848));
 b15aoi112ah1n06x5 U3219 (.a(n2849),
    .b(n2848),
    .c(net360),
    .d(net355),
    .o1(n2850));
 b15oai112as1n16x5 U3220 (.a(n2855),
    .b(n2850),
    .c(n3627),
    .d(n2857),
    .o1(u_device_sm_state_next[1]));
 b15oai012aq1n24x5 U3221 (.a(n2851),
    .b(n2876),
    .c(n2852),
    .o1(n3626));
 b15nano22as1n06x5 U3222 (.a(n3626),
    .b(n2878),
    .c(n3632),
    .out0(n2866));
 b15aoi112aq1n06x5 U3223 (.a(n2866),
    .b(n3618),
    .c(u_device_sm_sample_CMD),
    .d(n2853),
    .o1(n2854));
 b15nand02as1n08x5 U3224 (.a(n2890),
    .b(n3620),
    .o1(n2863));
 b15oai112as1n16x5 U3225 (.a(n2854),
    .b(n2863),
    .c(n3617),
    .d(n2889),
    .o1(u_device_sm_state_next[2]));
 b15nanb03ah1n16x5 U3226 (.a(n3617),
    .b(n2860),
    .c(u_device_sm_tx_done_reg),
    .out0(n2875));
 b15oai112as1n16x5 U3227 (.a(n2855),
    .b(n2875),
    .c(n3627),
    .d(n2856),
    .o1(u_device_sm_tx_data_valid_next));
 b15oabi12aq1n16x5 U3228 (.a(u_device_sm_tx_data_valid_next),
    .b(n3627),
    .c(n2857),
    .out0(u_device_sm_tx_counter_upd_next));
 b15aoi012aq1n32x5 U3229 (.a(n3664),
    .b(n2859),
    .c(n2858),
    .o1(n3666));
 b15inv020as1n04x5 U3230 (.a(n3666),
    .o1(n3174));
 b15inv040an1n04x5 U3231 (.a(n3228),
    .o1(n3176));
 b15nor002aq1n08x5 U3232 (.a(n3174),
    .b(n3176),
    .o1(n3681));
 b15ao0012an1n03x5 U3233 (.a(u_dcfifo_rx_u_din_full_full_up),
    .b(n3681),
    .c(n2865),
    .o(u_dcfifo_rx_u_din_full_N0));
 b15inv000al1n10x5 U3234 (.a(n2860),
    .o1(n3622));
 b15nor002ah1n04x5 U3235 (.a(n2861),
    .b(n3622),
    .o1(n2867));
 b15oaoi13ar1n08x5 U3236 (.a(n2862),
    .b(n2863),
    .c(n3632),
    .d(n3819),
    .o1(n2864));
 b15nor004as1n12x5 U3237 (.a(n2867),
    .b(n2866),
    .c(n2865),
    .d(n2864),
    .o1(n2656));
 b15nandp2al1n03x5 U3238 (.a(n2656),
    .b(n2868),
    .o1(u_rxreg_N9));
 b15nor004ah1n04x5 U3239 (.a(u_rxreg_counter_trgt[2]),
    .b(u_rxreg_counter_trgt[5]),
    .c(u_rxreg_counter_trgt[1]),
    .d(u_rxreg_counter_trgt[7]),
    .o1(n2872));
 b15nand04aq1n08x5 U3240 (.a(n2872),
    .b(n2871),
    .c(n2870),
    .d(n3813),
    .o1(n2873));
 b15oai013as1n12x5 U3241 (.a(n2656),
    .b(u_rxreg_counter_trgt[6]),
    .c(n2874),
    .d(n2873),
    .o1(u_rxreg_N7));
 b15inv000ar1n03x5 U3242 (.a(net470),
    .o1(tl_o[15]));
 b15oai112ah1n16x5 U3244 (.a(n2876),
    .b(n2875),
    .c(net138),
    .d(n2877),
    .o1(u_device_sm_ctrl_data_tx_ready_next));
 b15nand02an1n24x5 U3245 (.a(n2878),
    .b(net301),
    .o1(n3628));
 b15aoi022as1n08x5 U3246 (.a(n2886),
    .b(u_device_sm_s_dummy_cycles[4]),
    .c(n3613),
    .d(n3628),
    .o1(n2885));
 b15nor002an1n08x5 U3247 (.a(n2656),
    .b(n2879),
    .o1(n3612));
 b15inv020as1n10x5 U3248 (.a(n3612),
    .o1(n2896));
 b15nor003aq1n06x5 U3249 (.a(net302),
    .b(n3819),
    .c(net138),
    .o1(n2884));
 b15nor002as1n03x5 U3250 (.a(n2880),
    .b(n2886),
    .o1(n2882));
 b15aoi012ah1n02x5 U3251 (.a(n2890),
    .b(n2891),
    .c(n3613),
    .o1(n2881));
 b15inv040ah1n08x5 U3252 (.a(n3628),
    .o1(n3631));
 b15oaoi13an1n08x5 U3253 (.a(n3631),
    .b(n2881),
    .c(n2882),
    .d(n2889),
    .o1(n2883));
 b15oabi12al1n16x5 U3254 (.a(n2656),
    .b(n2884),
    .c(n2883),
    .out0(n2887));
 b15oai012ah1n12x5 U3255 (.a(n2887),
    .b(n2885),
    .c(n2896),
    .o1(u_rxreg_counter_trgt_next[4]));
 b15aoi022as1n08x5 U3256 (.a(n2886),
    .b(u_device_sm_s_dummy_cycles[3]),
    .c(n3613),
    .d(n3628),
    .o1(n2888));
 b15oai012ah1n12x5 U3257 (.a(n2887),
    .b(n2888),
    .c(n2896),
    .o1(u_rxreg_counter_trgt_next[3]));
 b15inv020as1n08x5 U3258 (.a(net2346),
    .o1(n3185));
 b15nor002aq1n04x5 U3259 (.a(n3617),
    .b(n2889),
    .o1(n2894));
 b15oai022as1n08x5 U3260 (.a(net301),
    .b(n3622),
    .c(n3631),
    .d(n2889),
    .o1(n2893));
 b15aoi112as1n08x5 U3261 (.a(n2890),
    .b(n2656),
    .c(n2891),
    .d(n3613),
    .o1(n3616));
 b15aoai13ah1n06x5 U3262 (.a(n3616),
    .b(n3819),
    .c(n3631),
    .d(net138),
    .o1(n2892));
 b15oai013as1n12x5 U3263 (.a(u_rxreg_N7),
    .b(n2894),
    .c(n2893),
    .d(n2892),
    .o1(n2895));
 b15aoai13as1n08x5 U3264 (.a(n2895),
    .b(n2896),
    .c(n3611),
    .d(n3185),
    .o1(u_rxreg_counter_trgt_next[2]));
 b15inv000ah1n03x5 U3265 (.a(u_device_sm_s_dummy_cycles[1]),
    .o1(n2897));
 b15aoai13as1n08x5 U3266 (.a(n2895),
    .b(n2896),
    .c(n3611),
    .d(n2897),
    .o1(u_rxreg_counter_trgt_next[1]));
 b15aoi112ah1n04x5 U3267 (.a(net139),
    .b(n2898),
    .c(u_dcfifo_rx_u_din_full_full_up),
    .d(u_dcfifo_rx_u_din_full_latched_full_s),
    .o1(u_dcfifo_rx_u_din_write_enable));
 b15nand02an1n12x5 U3268 (.a(net329),
    .b(net330),
    .o1(n3238));
 b15nand02as1n06x5 U3269 (.a(net331),
    .b(net333),
    .o1(n3248));
 b15nandp2ar1n08x5 U3270 (.a(u_dcfifo_rx_write_token[6]),
    .b(net327),
    .o1(n3246));
 b15nand02al1n12x5 U3271 (.a(u_dcfifo_rx_write_token[0]),
    .b(net336),
    .o1(n3242));
 b15nand04as1n16x5 U3272 (.a(n3238),
    .b(n3248),
    .c(n3246),
    .d(n3242),
    .o1(n2908));
 b15oa0012al1n32x5 U3273 (.a(u_dcfifo_rx_write_token[6]),
    .b(net329),
    .c(net327),
    .o(n3239));
 b15oaoi13as1n08x5 U3274 (.a(n3239),
    .b(u_dcfifo_rx_write_token[4]),
    .c(u_dcfifo_rx_write_token[5]),
    .d(u_dcfifo_rx_write_token[3]),
    .o1(n2903));
 b15oai012ah1n48x5 U3275 (.a(net334),
    .b(net332),
    .c(net335),
    .o1(n3235));
 b15nona23ah1n32x5 U3276 (.a(n3239),
    .b(n2903),
    .c(n3235),
    .d(net134),
    .out0(n2899));
 b15nor002ah1n16x5 U3277 (.a(n2908),
    .b(n2899),
    .o1(u_dcfifo_rx_u_din_buffer_N30));
 b15inv020aq1n32x5 U3278 (.a(n2908),
    .o1(n2906));
 b15nor002ah1n16x5 U3279 (.a(n2906),
    .b(n2899),
    .o1(u_dcfifo_rx_u_din_buffer_N31));
 b15inv040al1n12x5 U3280 (.a(n3235),
    .o1(n2905));
 b15and002ah1n08x5 U3281 (.a(net134),
    .b(n2903),
    .o(n2901));
 b15nand02as1n16x5 U3282 (.a(n2905),
    .b(n2901),
    .o1(n2900));
 b15norp02as1n12x5 U3283 (.a(n2906),
    .b(n2900),
    .o1(u_dcfifo_rx_u_din_buffer_N29));
 b15nor002aq1n02x5 U3284 (.a(n2908),
    .b(n2900),
    .o1(u_dcfifo_rx_u_din_buffer_N28));
 b15nand02ah1n32x5 U3285 (.a(n2901),
    .b(n3235),
    .o1(n2902));
 b15norp02ar1n48x5 U3286 (.a(n2906),
    .b(n2902),
    .o1(u_dcfifo_rx_u_din_buffer_N27));
 b15nor002aq1n16x5 U3287 (.a(n2908),
    .b(n2902),
    .o1(u_dcfifo_rx_u_din_buffer_N26));
 b15nonb02al1n12x5 U3288 (.a(net134),
    .b(n2903),
    .out0(n2904));
 b15oai012al1n48x5 U3289 (.a(n2904),
    .b(n2905),
    .c(n3239),
    .o1(n2907));
 b15norp02al1n32x5 U3290 (.a(n2906),
    .b(n2907),
    .o1(u_dcfifo_rx_u_din_buffer_N33));
 b15norp02ah1n16x5 U3291 (.a(n2908),
    .b(n2907),
    .o1(u_dcfifo_rx_u_din_buffer_N32));
 b15inv000ar1n03x5 U3292 (.a(net1454),
    .o1(tl_o[16]));
 b15inv000ar1n03x5 U3294 (.a(net1455),
    .o1(tl_o[17]));
 b15norp02al1n08x5 U3296 (.a(tx_counter_upd),
    .b(u_txreg_running),
    .o1(n2966));
 b15inv020as1n10x5 U3297 (.a(n2966),
    .o1(u_txreg_N11));
 b15inv000ar1n03x5 U3298 (.a(net471),
    .o1(tl_o[18]));
 b15inv000ar1n03x5 U3300 (.a(net1456),
    .o1(tl_o[19]));
 b15inv000ar1n03x5 U3302 (.a(net1457),
    .o1(tl_o[20]));
 b15inv000ar1n03x5 U3304 (.a(net1458),
    .o1(tl_o[21]));
 b15inv000ar1n03x5 U3306 (.a(net1459),
    .o1(tl_o[22]));
 b15ao0022an1n16x5 U3307 (.a(net296),
    .b(net255),
    .c(net250),
    .d(net262),
    .o(net57));
 b15nonb02al1n12x5 U3308 (.a(net251),
    .b(net262),
    .out0(net59));
 b15nonb02al1n08x5 U3309 (.a(net249),
    .b(net262),
    .out0(net60));
 b15nonb02as1n06x5 U3310 (.a(net253),
    .b(net262),
    .out0(net58));
 b15and002an1n08x5 U3312 (.a(net2298),
    .b(net2196),
    .o(u_txreg_N34));
 b15qgbno2an1n10x5 U3313 (.a(net298),
    .b(net354),
    .o1(n2917));
 b15inv000ar1n03x5 U3314 (.a(net1460),
    .o1(tl_o[23]));
 b15ao0022al1n04x5 U3316 (.a(net352),
    .b(net2214),
    .c(net260),
    .d(u_txreg_data_int[2]),
    .o(u_txreg_N37));
 b15ao0022ah1n02x5 U3317 (.a(net352),
    .b(net2315),
    .c(net260),
    .d(u_txreg_data_int[1]),
    .o(u_txreg_N36));
 b15ao0022ar1n02x5 U3318 (.a(net352),
    .b(net2312),
    .c(net261),
    .d(u_txreg_data_int[0]),
    .o(u_txreg_N35));
 b15norp02aq1n08x5 U3319 (.a(net353),
    .b(n3815),
    .o1(n2919));
 b15inv000ar1n03x5 U3320 (.a(net472),
    .o1(tl_o[56]));
 b15inv000ar1n03x5 U3322 (.a(net473),
    .o1(tl_o[57]));
 b15aoi022ar1n02x5 U3324 (.a(net353),
    .b(net2163),
    .c(net261),
    .d(u_txreg_data_int[24]),
    .o1(n2920));
 b15aob012al1n04x5 U3325 (.a(net2164),
    .b(net257),
    .c(u_txreg_data_int[21]),
    .out0(u_txreg_N59));
 b15aoi022ar1n04x5 U3326 (.a(net2299),
    .b(tx_data[29]),
    .c(net261),
    .d(u_txreg_data_int[28]),
    .o1(n2921));
 b15aob012ar1n08x5 U3327 (.a(net2300),
    .b(net257),
    .c(u_txreg_data_int[25]),
    .out0(u_txreg_N63));
 b15aoi022an1n02x5 U3328 (.a(net353),
    .b(net2166),
    .c(net261),
    .d(u_txreg_data_int[26]),
    .o1(n2922));
 b15aob012aq1n08x5 U3329 (.a(net2167),
    .b(net257),
    .c(u_txreg_data_int[23]),
    .out0(u_txreg_N61));
 b15aoi022ah1n08x5 U3330 (.a(net352),
    .b(net2231),
    .c(net260),
    .d(u_txreg_data_int[29]),
    .o1(n2923));
 b15aob012al1n06x5 U3331 (.a(net2232),
    .b(net257),
    .c(u_txreg_data_int[26]),
    .out0(u_txreg_N64));
 b15aoi022as1n04x5 U3332 (.a(net353),
    .b(net2179),
    .c(net261),
    .d(u_txreg_data_int[25]),
    .o1(n2925));
 b15aob012al1n08x5 U3333 (.a(net2180),
    .b(net257),
    .c(u_txreg_data_int[22]),
    .out0(u_txreg_N60));
 b15inv000ar1n03x5 U3334 (.a(net474),
    .o1(tl_o[58]));
 b15aoi022ar1n08x5 U3336 (.a(net353),
    .b(net2170),
    .c(net261),
    .d(u_txreg_data_int[19]),
    .o1(n2927));
 b15aob012as1n04x5 U3337 (.a(net2171),
    .b(net256),
    .c(u_txreg_data_int[16]),
    .out0(u_txreg_N54));
 b15aoi022an1n04x5 U3338 (.a(net352),
    .b(net2141),
    .c(net261),
    .d(u_txreg_data_int[18]),
    .o1(n2928));
 b15aob012al1n06x5 U3339 (.a(net2142),
    .b(net257),
    .c(u_txreg_data_int[15]),
    .out0(u_txreg_N53));
 b15inv000ar1n03x5 U3340 (.a(net475),
    .o1(tl_o[59]));
 b15aoi022an1n04x5 U3341 (.a(net353),
    .b(net2176),
    .c(net260),
    .d(u_txreg_data_int[11]),
    .o1(n2929));
 b15aob012ar1n04x5 U3342 (.a(net2177),
    .b(net256),
    .c(u_txreg_data_int[8]),
    .out0(u_txreg_N46));
 b15aoi022an1n06x5 U3343 (.a(net352),
    .b(net2288),
    .c(net260),
    .d(u_txreg_data_int[30]),
    .o1(n2930));
 b15aob012aq1n06x5 U3344 (.a(net2289),
    .b(net257),
    .c(u_txreg_data_int[27]),
    .out0(u_txreg_N65));
 b15aoi022aq1n04x5 U3345 (.a(net352),
    .b(net2189),
    .c(net261),
    .d(u_txreg_data_int[14]),
    .o1(n2931));
 b15aob012as1n04x5 U3346 (.a(net2190),
    .b(net256),
    .c(u_txreg_data_int[11]),
    .out0(u_txreg_N49));
 b15aoi022al1n06x5 U3347 (.a(net352),
    .b(net2204),
    .c(net260),
    .d(u_txreg_data_int[9]),
    .o1(n2932));
 b15aob012ar1n06x5 U3348 (.a(net2205),
    .b(net256),
    .c(u_txreg_data_int[6]),
    .out0(u_txreg_N44));
 b15aoi022as1n06x5 U3349 (.a(net353),
    .b(net2201),
    .c(net260),
    .d(u_txreg_data_int[13]),
    .o1(n2933));
 b15aob012ar1n02x5 U3350 (.a(net2202),
    .b(net256),
    .c(u_txreg_data_int[10]),
    .out0(u_txreg_N48));
 b15aoi022an1n04x5 U3351 (.a(net353),
    .b(net2209),
    .c(net261),
    .d(u_txreg_data_int[22]),
    .o1(n2934));
 b15aob012ah1n06x5 U3352 (.a(net2210),
    .b(net257),
    .c(u_txreg_data_int[19]),
    .out0(u_txreg_N57));
 b15aoi022al1n02x5 U3353 (.a(net353),
    .b(net2183),
    .c(net260),
    .d(u_txreg_data_int[12]),
    .o1(n2935));
 b15aob012ah1n03x5 U3354 (.a(net2184),
    .b(net256),
    .c(u_txreg_data_int[9]),
    .out0(u_txreg_N47));
 b15aoi022ar1n02x5 U3355 (.a(net352),
    .b(net2192),
    .c(net260),
    .d(u_txreg_data_int[8]),
    .o1(n2936));
 b15aob012ar1n02x5 U3356 (.a(net2193),
    .b(net256),
    .c(u_txreg_data_int[5]),
    .out0(u_txreg_N43));
 b15aoi022ar1n06x5 U3357 (.a(net352),
    .b(net2198),
    .c(net260),
    .d(u_txreg_data_int[16]),
    .o1(n2937));
 b15aob012ar1n08x5 U3358 (.a(net2199),
    .b(net256),
    .c(u_txreg_data_int[13]),
    .out0(u_txreg_N51));
 b15aoi022ar1n08x5 U3359 (.a(net353),
    .b(net2155),
    .c(net261),
    .d(u_txreg_data_int[17]),
    .o1(n2938));
 b15aob012ar1n06x5 U3360 (.a(net2156),
    .b(net256),
    .c(u_txreg_data_int[14]),
    .out0(u_txreg_N52));
 b15aoi022ar1n02x5 U3361 (.a(net352),
    .b(net2173),
    .c(net260),
    .d(u_txreg_data_int[10]),
    .o1(n2939));
 b15aob012al1n03x5 U3362 (.a(net2174),
    .b(net256),
    .c(u_txreg_data_int[7]),
    .out0(u_txreg_N45));
 b15aoi022an1n04x5 U3363 (.a(net353),
    .b(net2152),
    .c(net261),
    .d(u_txreg_data_int[15]),
    .o1(n2940));
 b15aob012al1n08x5 U3364 (.a(net2153),
    .b(net256),
    .c(u_txreg_data_int[12]),
    .out0(u_txreg_N50));
 b15aoi022al1n04x5 U3365 (.a(net353),
    .b(net2186),
    .c(net261),
    .d(u_txreg_data_int[20]),
    .o1(n2941));
 b15aob012al1n06x5 U3366 (.a(net2187),
    .b(net257),
    .c(u_txreg_data_int[17]),
    .out0(u_txreg_N55));
 b15aoi022ar1n08x5 U3367 (.a(net352),
    .b(net2238),
    .c(net260),
    .d(u_txreg_data_int[7]),
    .o1(n2942));
 b15aob012aq1n03x5 U3368 (.a(net2239),
    .b(net256),
    .c(u_txreg_data_int[4]),
    .out0(u_txreg_N42));
 b15aoi022an1n04x5 U3369 (.a(net353),
    .b(net2206),
    .c(net261),
    .d(u_txreg_data_int[21]),
    .o1(n2943));
 b15aob012al1n08x5 U3370 (.a(net2207),
    .b(net257),
    .c(u_txreg_data_int[18]),
    .out0(u_txreg_N56));
 b15aoi022an1n02x5 U3371 (.a(net353),
    .b(net2144),
    .c(net261),
    .d(u_txreg_data_int[23]),
    .o1(n2945));
 b15aob012an1n03x5 U3372 (.a(net2145),
    .b(net257),
    .c(u_txreg_data_int[20]),
    .out0(u_txreg_N58));
 b15aoi022an1n02x5 U3373 (.a(net352),
    .b(net2219),
    .c(net260),
    .d(u_txreg_data_int[5]),
    .o1(n2946));
 b15aob012ar1n06x5 U3374 (.a(net2220),
    .b(net256),
    .c(u_txreg_data_int[2]),
    .out0(u_txreg_N40));
 b15aoi022as1n06x5 U3375 (.a(net352),
    .b(net2225),
    .c(net260),
    .d(u_txreg_data_int[6]),
    .o1(n2948));
 b15aob012ah1n04x5 U3376 (.a(net2226),
    .b(net256),
    .c(u_txreg_data_int[3]),
    .out0(u_txreg_N41));
 b15aoi022ar1n12x5 U3377 (.a(net353),
    .b(net2234),
    .c(u_txreg_data_int[27]),
    .d(net261),
    .o1(n2951));
 b15aob012ah1n06x5 U3378 (.a(net2235),
    .b(net257),
    .c(u_txreg_data_int[24]),
    .out0(u_txreg_N62));
 b15inv020as1n10x5 U3379 (.a(u_txreg_counter[2]),
    .o1(n2980));
 b15inv040al1n03x5 U3380 (.a(u_txreg_counter[5]),
    .o1(n2962));
 b15xor002as1n03x5 U3381 (.a(u_txreg_counter_trgt[3]),
    .b(u_txreg_counter[3]),
    .out0(n2961));
 b15inv000al1n02x5 U3382 (.a(u_txreg_counter[0]),
    .o1(n2958));
 b15xor002al1n02x5 U3383 (.a(u_txreg_counter_trgt[7]),
    .b(u_txreg_counter[7]),
    .out0(n2957));
 b15nand02ar1n02x5 U3384 (.a(u_txreg_counter[4]),
    .b(u_txreg_counter_trgt[4]),
    .o1(n2954));
 b15xor002ar1n02x5 U3385 (.a(u_txreg_counter_trgt[6]),
    .b(u_txreg_counter[6]),
    .out0(n2953));
 b15oaoi13ar1n03x5 U3386 (.a(n2953),
    .b(n2954),
    .c(u_txreg_counter[4]),
    .d(u_txreg_counter_trgt[4]),
    .o1(n2955));
 b15oai012ar1n02x5 U3387 (.a(n2955),
    .b(u_txreg_counter_trgt[0]),
    .c(n2958),
    .o1(n2956));
 b15aoi112ar1n02x5 U3388 (.a(n2957),
    .b(n2956),
    .c(u_txreg_counter_trgt[0]),
    .d(n2958),
    .o1(n2959));
 b15oai012aq1n03x5 U3389 (.a(n2959),
    .b(n2962),
    .c(u_txreg_counter_trgt[5]),
    .o1(n2960));
 b15aoi112an1n06x5 U3390 (.a(n2961),
    .b(n2960),
    .c(n2962),
    .d(u_txreg_counter_trgt[5]),
    .o1(n2965));
 b15xor002al1n03x5 U3391 (.a(u_txreg_counter_trgt[1]),
    .b(u_txreg_counter[1]),
    .out0(n2963));
 b15aoi012ar1n06x5 U3392 (.a(n2963),
    .b(u_txreg_counter_trgt[2]),
    .c(n2980),
    .o1(n2964));
 b15oai112as1n16x5 U3393 (.a(n2965),
    .b(n2964),
    .c(u_txreg_counter_trgt[2]),
    .d(n2980),
    .o1(n2981));
 b15norp02as1n12x5 U3394 (.a(n2966),
    .b(n2981),
    .o1(tx_done));
 b15nandp2ar1n05x5 U3395 (.a(u_txreg_counter[1]),
    .b(u_txreg_counter[0]),
    .o1(n2979));
 b15oai112ar1n04x5 U3396 (.a(n2979),
    .b(n2981),
    .c(u_txreg_counter[1]),
    .d(u_txreg_counter[0]),
    .o1(n2967));
 b15inv020an1n04x5 U3397 (.a(n2967),
    .o1(u_txreg_N25));
 b15inv020al1n05x5 U3398 (.a(u_txreg_counter[4]),
    .o1(n2973));
 b15and003aq1n04x5 U3399 (.a(net2372),
    .b(u_txreg_counter[1]),
    .c(u_txreg_counter[0]),
    .o(n2978));
 b15nand02an1n08x5 U3400 (.a(u_txreg_counter[3]),
    .b(n2978),
    .o1(n2972));
 b15nor002as1n04x5 U3401 (.a(n2973),
    .b(n2972),
    .o1(n2971));
 b15nandp2al1n08x5 U3402 (.a(u_txreg_counter[5]),
    .b(n2971),
    .o1(n2975));
 b15oai112aq1n02x5 U3403 (.a(n2975),
    .b(n2981),
    .c(u_txreg_counter[5]),
    .d(n2971),
    .o1(n2968));
 b15inv000aq1n02x5 U3404 (.a(n2968),
    .o1(u_txreg_N29));
 b15oai112an1n02x5 U3405 (.a(n2972),
    .b(n2981),
    .c(u_txreg_counter[3]),
    .d(n2978),
    .o1(n2969));
 b15inv040as1n02x5 U3406 (.a(n2969),
    .o1(u_txreg_N27));
 b15inv020as1n08x5 U3407 (.a(n2981),
    .o1(n2977));
 b15norp02as1n03x5 U3408 (.a(u_txreg_counter[0]),
    .b(n2977),
    .o1(u_txreg_N24));
 b15inv000aq1n05x5 U3409 (.a(u_txreg_counter[6]),
    .o1(n2976));
 b15nor002al1n06x5 U3410 (.a(n2976),
    .b(n2975),
    .o1(n2974));
 b15oai012al1n02x5 U3411 (.a(n2981),
    .b(u_txreg_counter[7]),
    .c(n2974),
    .o1(n2970));
 b15aoi012an1n04x5 U3412 (.a(n2970),
    .b(u_txreg_counter[7]),
    .c(n2974),
    .o1(u_txreg_N31));
 b15aoi112al1n06x5 U3413 (.a(n2971),
    .b(n2977),
    .c(n2973),
    .d(n2972),
    .o1(u_txreg_N28));
 b15aoi112ar1n08x5 U3414 (.a(n2974),
    .b(n2977),
    .c(n2976),
    .d(n2975),
    .o1(u_txreg_N30));
 b15aoi112al1n06x5 U3415 (.a(n2978),
    .b(n2977),
    .c(n2980),
    .d(n2979),
    .o1(u_txreg_N26));
 b15nanb02ah1n08x5 U3416 (.a(tx_counter_upd),
    .b(n2981),
    .out0(u_txreg_N10));
 b15orn002ar1n02x5 U3417 (.a(u_dcfifo_tx_u_din_full_full_up),
    .b(net53),
    .o(u_dcfifo_tx_u_din_full_N0));
 b15inv000ar1n03x5 U3419 (.a(net1461),
    .o1(tl_o[60]));
 b15inv000ar1n03x5 U3421 (.a(net1462),
    .o1(tl_o[61]));
 b15inv000ar1n03x5 U3423 (.a(net1463),
    .o1(tl_o[93]));
 b15inv000ar1n03x5 U3425 (.a(net1464),
    .o1(tl_o[94]));
 b15inv000ar1n03x5 U3427 (.a(net1465),
    .o1(tl_o[95]));
 b15inv000ar1n03x5 U3429 (.a(net1466),
    .o1(tl_o[96]));
 b15inv000ar1n03x5 U3431 (.a(net1467),
    .o1(tl_o[97]));
 b15inv000ar1n03x5 U3433 (.a(net1468),
    .o1(tl_o[98]));
 b15inv000ar1n03x5 U3435 (.a(net1469),
    .o1(tl_o[99]));
 b15inv000ar1n03x5 U3437 (.a(net1470),
    .o1(tl_o[100]));
 b15inv000ar1n03x5 U3439 (.a(net476),
    .o1(tl_o[101]));
 b15inv000ar1n03x5 U3441 (.a(net1471),
    .o1(tl_o[102]));
 b15inv000ar1n03x5 U3443 (.a(net1472),
    .o1(tl_o[103]));
 b15inv000ar1n03x5 U3445 (.a(net1473),
    .o1(tl_o[104]));
 b15inv000ar1n03x5 U3447 (.a(net1474),
    .o1(tl_o[105]));
 b15inv000ar1n03x5 U3449 (.a(net1475),
    .o1(tl_o[106]));
 b15ztpn00an1n08x5 PHY_66 ();
 b15ztpn00an1n08x5 PHY_65 ();
 b15ztpn00an1n08x5 PHY_64 ();
 b15ztpn00an1n08x5 PHY_63 ();
 b15ztpn00an1n08x5 PHY_62 ();
 b15ztpn00an1n08x5 PHY_61 ();
 b15ztpn00an1n08x5 PHY_60 ();
 b15ztpn00an1n08x5 PHY_59 ();
 b15ztpn00an1n08x5 PHY_58 ();
 b15ztpn00an1n08x5 PHY_57 ();
 b15ztpn00an1n08x5 PHY_56 ();
 b15ztpn00an1n08x5 PHY_55 ();
 b15ztpn00an1n08x5 PHY_54 ();
 b15ztpn00an1n08x5 PHY_53 ();
 b15ztpn00an1n08x5 PHY_52 ();
 b15ztpn00an1n08x5 PHY_51 ();
 b15ztpn00an1n08x5 PHY_50 ();
 b15ztpn00an1n08x5 PHY_49 ();
 b15ztpn00an1n08x5 PHY_48 ();
 b15nandp2ar1n32x5 U3471 (.a(n3008),
    .b(n3645),
    .o1(n3634));
 b15oaoi13as1n08x5 U3472 (.a(n3634),
    .b(u_dcfifo_tx_u_dout_read_token[4]),
    .c(u_dcfifo_tx_u_dout_read_token[5]),
    .d(net305),
    .o1(n3014));
 b15nandp2al1n16x5 U3473 (.a(n3647),
    .b(n3640),
    .o1(n3649));
 b15oaoi13as1n08x5 U3474 (.a(n3649),
    .b(u_dcfifo_tx_u_dout_read_token[2]),
    .c(u_dcfifo_tx_u_dout_read_token[1]),
    .d(u_dcfifo_tx_u_dout_read_token[3]),
    .o1(n3012));
 b15aoi022aq1n32x5 U3475 (.a(u_dcfifo_tx_u_dout_read_token[0]),
    .b(net306),
    .c(net304),
    .d(u_dcfifo_tx_u_dout_read_token[6]),
    .o1(n3007));
 b15inv000as1n06x5 U3476 (.a(n3007),
    .o1(n3005));
 b15aoi112as1n08x5 U3477 (.a(n3001),
    .b(n3005),
    .c(u_dcfifo_tx_u_dout_read_token[2]),
    .d(u_dcfifo_tx_u_dout_read_token[3]),
    .o1(n3013));
 b15nanb02as1n24x5 U3478 (.a(n3012),
    .b(n3013),
    .out0(n3003));
 b15norp02as1n48x5 U3479 (.a(n3014),
    .b(n3003),
    .o1(n3002));
 b15ztpn00an1n08x5 PHY_47 ();
 b15ztpn00an1n08x5 PHY_46 ();
 b15inv020an1n16x5 U3482 (.a(n3014),
    .o1(n3017));
 b15norp02al1n24x5 U3483 (.a(n3017),
    .b(n3003),
    .o1(n3004));
 b15ztpn00an1n08x5 PHY_45 ();
 b15ztpn00an1n08x5 PHY_44 ();
 b15aoi022an1n08x5 U3486 (.a(net188),
    .b(u_dcfifo_tx_u_din_buffer_data[203]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[139]),
    .o1(n3024));
 b15nandp2ar1n24x5 U3487 (.a(n3012),
    .b(n3005),
    .o1(n3019));
 b15nor002aq1n04x5 U3488 (.a(n3634),
    .b(n3019),
    .o1(n3006));
 b15ztpn00an1n08x5 PHY_43 ();
 b15ztpn00an1n08x5 PHY_42 ();
 b15nand02ah1n48x5 U3491 (.a(n3012),
    .b(n3007),
    .o1(n3010));
 b15norp02aq1n48x5 U3492 (.a(n3008),
    .b(n3010),
    .o1(n3009));
 b15ztpn00an1n08x5 PHY_41 ();
 b15aoi022aq1n16x5 U3495 (.a(net182),
    .b(u_dcfifo_tx_u_din_buffer_data[43]),
    .c(net180),
    .d(u_dcfifo_tx_u_din_buffer_data[75]),
    .o1(n3023));
 b15qgbno2an1n05x5 U3496 (.o1(n3011),
    .a(n3633),
    .b(n3010));
 b15ztpn00an1n08x5 PHY_40 ();
 b15ztpn00an1n08x5 PHY_39 ();
 b15orn002al1n32x5 U3499 (.a(n3013),
    .b(n3012),
    .o(n3016));
 b15nor002an1n24x5 U3500 (.a(n3014),
    .b(n3016),
    .o1(n3015));
 b15ztpn00an1n08x5 PHY_38 ();
 b15ztpn00an1n08x5 PHY_37 ();
 b15aoi022ah1n16x5 U3503 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[11]),
    .c(net174),
    .d(u_dcfifo_tx_u_din_buffer_data[235]),
    .o1(n3022));
 b15norp02aq1n48x5 U3504 (.a(n3017),
    .b(n3016),
    .o1(n3018));
 b15ztpn00an1n08x5 PHY_36 ();
 b15ztpn00an1n08x5 PHY_35 ();
 b15nonb02ah1n03x5 U3507 (.a(n3634),
    .b(n3019),
    .out0(n3020));
 b15ztpn00an1n08x5 PHY_34 ();
 b15ztpn00an1n08x5 PHY_33 ();
 b15aoi022ah1n08x5 U3510 (.a(net172),
    .b(u_dcfifo_tx_u_din_buffer_data[171]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[107]),
    .o1(n3021));
 b15nand04as1n16x5 U3511 (.a(n3024),
    .b(n3023),
    .c(n3022),
    .d(n3021),
    .o1(n3025));
 b15ztpn00an1n08x5 PHY_32 ();
 b15nonb02ar1n02x3 U3513 (.a(n3025),
    .b(net135),
    .out0(u_device_sm_N185));
 b15ztpn00an1n08x5 PHY_31 ();
 b15ztpn00an1n08x5 PHY_30 ();
 b15aoi022as1n08x5 U3516 (.a(net183),
    .b(u_dcfifo_tx_u_din_buffer_data[59]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[123]),
    .o1(n3029));
 b15ztpn00an1n08x5 PHY_29 ();
 b15aoi022an1n08x5 U3519 (.a(net189),
    .b(u_dcfifo_tx_u_din_buffer_data[219]),
    .c(net175),
    .d(u_dcfifo_tx_u_din_buffer_data[251]),
    .o1(n3028));
 b15ztpn00an1n08x5 PHY_28 ();
 b15aoi022as1n06x5 U3522 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[27]),
    .c(net173),
    .d(u_dcfifo_tx_u_din_buffer_data[187]),
    .o1(n3027));
 b15ztpn00an1n08x5 PHY_27 ();
 b15ztpn00an1n08x5 PHY_26 ();
 b15aoi022ar1n32x5 U3525 (.a(net181),
    .b(u_dcfifo_tx_u_din_buffer_data[91]),
    .c(net186),
    .d(u_dcfifo_tx_u_din_buffer_data[155]),
    .o1(n3026));
 b15nand04as1n16x5 U3526 (.a(n3029),
    .b(n3028),
    .c(n3027),
    .d(n3026),
    .o1(n3031));
 b15ztpn00an1n08x5 PHY_25 ();
 b15nonb02aq1n16x5 U3528 (.a(n3031),
    .b(net137),
    .out0(u_device_sm_N201));
 b15aoi022as1n06x5 U3529 (.a(net188),
    .b(u_dcfifo_tx_u_din_buffer_data[204]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[140]),
    .o1(n3038));
 b15aoi022al1n08x5 U3530 (.a(net182),
    .b(u_dcfifo_tx_u_din_buffer_data[44]),
    .c(net180),
    .d(u_dcfifo_tx_u_din_buffer_data[76]),
    .o1(n3037));
 b15ztpn00an1n08x5 PHY_24 ();
 b15ztpn00an1n08x5 PHY_23 ();
 b15aoi022as1n08x5 U3533 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[12]),
    .c(net172),
    .d(u_dcfifo_tx_u_din_buffer_data[172]),
    .o1(n3036));
 b15ztpn00an1n08x5 PHY_22 ();
 b15aoi022ar1n32x5 U3535 (.a(net174),
    .b(u_dcfifo_tx_u_din_buffer_data[236]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[108]),
    .o1(n3035));
 b15nand04aq1n16x5 U3536 (.a(n3038),
    .b(n3037),
    .c(n3036),
    .d(n3035),
    .o1(n3039));
 b15nonb02ar1n08x5 U3537 (.a(n3039),
    .b(net135),
    .out0(u_device_sm_N186));
 b15aoi022ah1n08x5 U3538 (.a(net180),
    .b(u_dcfifo_tx_u_din_buffer_data[77]),
    .c(net172),
    .d(u_dcfifo_tx_u_din_buffer_data[173]),
    .o1(n3044));
 b15ztpn00an1n08x5 PHY_21 ();
 b15aoi022an1n12x5 U3540 (.a(net188),
    .b(u_dcfifo_tx_u_din_buffer_data[205]),
    .c(net174),
    .d(u_dcfifo_tx_u_din_buffer_data[237]),
    .o1(n3043));
 b15aoi022aq1n16x5 U3541 (.a(net182),
    .b(u_dcfifo_tx_u_din_buffer_data[45]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[109]),
    .o1(n3042));
 b15aoi022aq1n08x5 U3542 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[13]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[141]),
    .o1(n3041));
 b15nand04aq1n16x5 U3543 (.a(n3044),
    .b(n3043),
    .c(n3042),
    .d(n3041),
    .o1(n3045));
 b15nonb02ar1n08x5 U3544 (.a(n3045),
    .b(net136),
    .out0(u_device_sm_N187));
 b15aoi022ar1n12x5 U3545 (.a(net189),
    .b(u_dcfifo_tx_u_din_buffer_data[215]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[119]),
    .o1(n3050));
 b15aoi022ar1n16x5 U3546 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[23]),
    .c(net175),
    .d(u_dcfifo_tx_u_din_buffer_data[247]),
    .o1(n3049));
 b15ztpn00an1n08x5 PHY_20 ();
 b15aoi022as1n06x5 U3548 (.a(net181),
    .b(u_dcfifo_tx_u_din_buffer_data[87]),
    .c(net173),
    .d(u_dcfifo_tx_u_din_buffer_data[183]),
    .o1(n3048));
 b15aoi022an1n08x5 U3549 (.a(net183),
    .b(u_dcfifo_tx_u_din_buffer_data[55]),
    .c(net186),
    .d(u_dcfifo_tx_u_din_buffer_data[151]),
    .o1(n3047));
 b15nand04as1n16x5 U3550 (.a(n3050),
    .b(n3049),
    .c(n3048),
    .d(n3047),
    .o1(n3051));
 b15nonb02as1n16x5 U3551 (.a(n3051),
    .b(net137),
    .out0(u_device_sm_N197));
 b15aoi022ar1n16x5 U3552 (.a(net183),
    .b(u_dcfifo_tx_u_din_buffer_data[51]),
    .c(net175),
    .d(u_dcfifo_tx_u_din_buffer_data[243]),
    .o1(n3055));
 b15aoi022aq1n08x5 U3553 (.a(net189),
    .b(u_dcfifo_tx_u_din_buffer_data[211]),
    .c(net181),
    .d(u_dcfifo_tx_u_din_buffer_data[83]),
    .o1(n3054));
 b15aoi022as1n08x5 U3554 (.a(net173),
    .b(u_dcfifo_tx_u_din_buffer_data[179]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[115]),
    .o1(n3053));
 b15aoi022an1n08x5 U3555 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[19]),
    .c(net186),
    .d(u_dcfifo_tx_u_din_buffer_data[147]),
    .o1(n3052));
 b15nand04as1n16x5 U3556 (.a(n3055),
    .b(n3054),
    .c(n3053),
    .d(n3052),
    .o1(n3056));
 b15nonb02ah1n16x5 U3557 (.a(n3056),
    .b(net137),
    .out0(u_device_sm_N193));
 b15ztpn00an1n08x5 PHY_19 ();
 b15aoi022as1n08x5 U3559 (.a(net183),
    .b(u_dcfifo_tx_u_din_buffer_data[63]),
    .c(net189),
    .d(u_dcfifo_tx_u_din_buffer_data[223]),
    .o1(n3061));
 b15aoi022aq1n08x5 U3560 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[31]),
    .c(net181),
    .d(u_dcfifo_tx_u_din_buffer_data[95]),
    .o1(n3060));
 b15aoi022aq1n32x5 U3561 (.a(net186),
    .b(u_dcfifo_tx_u_din_buffer_data[159]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[127]),
    .o1(n3059));
 b15aoi022ar1n16x5 U3562 (.a(net173),
    .b(u_dcfifo_tx_u_din_buffer_data[191]),
    .c(net175),
    .d(u_dcfifo_tx_u_din_buffer_data[255]),
    .o1(n3058));
 b15nand04as1n16x5 U3563 (.a(n3061),
    .b(n3060),
    .c(n3059),
    .d(n3058),
    .o1(n3062));
 b15nonb02aq1n06x5 U3564 (.a(n3062),
    .b(net136),
    .out0(u_device_sm_N205));
 b15aoi022an1n16x5 U3565 (.a(net183),
    .b(u_dcfifo_tx_u_din_buffer_data[50]),
    .c(net175),
    .d(u_dcfifo_tx_u_din_buffer_data[242]),
    .o1(n3066));
 b15aoi022as1n08x5 U3566 (.a(net189),
    .b(u_dcfifo_tx_u_din_buffer_data[210]),
    .c(net173),
    .d(u_dcfifo_tx_u_din_buffer_data[178]),
    .o1(n3065));
 b15aoi022as1n12x5 U3567 (.a(net186),
    .b(u_dcfifo_tx_u_din_buffer_data[146]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[114]),
    .o1(n3064));
 b15aoi022aq1n12x5 U3568 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[18]),
    .c(net181),
    .d(u_dcfifo_tx_u_din_buffer_data[82]),
    .o1(n3063));
 b15nand04as1n16x5 U3569 (.a(n3066),
    .b(n3065),
    .c(n3064),
    .d(n3063),
    .o1(n3067));
 b15nonb02ah1n16x5 U3570 (.a(n3067),
    .b(net137),
    .out0(u_device_sm_N192));
 b15aoi022aq1n12x5 U3571 (.a(net183),
    .b(u_dcfifo_tx_u_din_buffer_data[48]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[112]),
    .o1(n3071));
 b15aoi022ah1n08x5 U3572 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[16]),
    .c(net173),
    .d(u_dcfifo_tx_u_din_buffer_data[176]),
    .o1(n3070));
 b15aoi022al1n12x5 U3573 (.a(net189),
    .b(u_dcfifo_tx_u_din_buffer_data[208]),
    .c(net175),
    .d(u_dcfifo_tx_u_din_buffer_data[240]),
    .o1(n3069));
 b15aoi022ar1n24x5 U3574 (.a(net181),
    .b(u_dcfifo_tx_u_din_buffer_data[80]),
    .c(net186),
    .d(u_dcfifo_tx_u_din_buffer_data[144]),
    .o1(n3068));
 b15nand04as1n16x5 U3575 (.a(n3071),
    .b(n3070),
    .c(n3069),
    .d(n3068),
    .o1(n3072));
 b15nonb02aq1n16x5 U3576 (.a(n3072),
    .b(net137),
    .out0(u_device_sm_N190));
 b15aoi022as1n06x5 U3577 (.a(net189),
    .b(u_dcfifo_tx_u_din_buffer_data[222]),
    .c(net175),
    .d(u_dcfifo_tx_u_din_buffer_data[254]),
    .o1(n3076));
 b15aoi022al1n16x5 U3578 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[30]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[126]),
    .o1(n3075));
 b15aoi022aq1n16x5 U3579 (.a(net173),
    .b(u_dcfifo_tx_u_din_buffer_data[190]),
    .c(net186),
    .d(u_dcfifo_tx_u_din_buffer_data[158]),
    .o1(n3074));
 b15aoi022as1n06x5 U3580 (.a(net183),
    .b(u_dcfifo_tx_u_din_buffer_data[62]),
    .c(net181),
    .d(u_dcfifo_tx_u_din_buffer_data[94]),
    .o1(n3073));
 b15nand04as1n16x5 U3581 (.a(n3076),
    .b(n3075),
    .c(n3074),
    .d(n3073),
    .o1(n3077));
 b15nonb02ah1n06x5 U3582 (.a(n3077),
    .b(net136),
    .out0(u_device_sm_N204));
 b15aoi022an1n16x5 U3583 (.a(net188),
    .b(u_dcfifo_tx_u_din_buffer_data[206]),
    .c(net174),
    .d(u_dcfifo_tx_u_din_buffer_data[238]),
    .o1(n3081));
 b15aoi022as1n04x5 U3584 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[14]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[110]),
    .o1(n3080));
 b15aoi022al1n24x5 U3585 (.a(net180),
    .b(u_dcfifo_tx_u_din_buffer_data[78]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[142]),
    .o1(n3079));
 b15aoi022ah1n08x5 U3586 (.a(net182),
    .b(u_dcfifo_tx_u_din_buffer_data[46]),
    .c(net172),
    .d(u_dcfifo_tx_u_din_buffer_data[174]),
    .o1(n3078));
 b15nand04aq1n16x5 U3587 (.a(n3081),
    .b(n3080),
    .c(n3079),
    .d(n3078),
    .o1(n3082));
 b15nonb02al1n04x5 U3588 (.a(n3082),
    .b(net135),
    .out0(u_device_sm_N188));
 b15aoi022as1n06x5 U3589 (.a(net173),
    .b(u_dcfifo_tx_u_din_buffer_data[185]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[121]),
    .o1(n3086));
 b15aoi022an1n08x5 U3590 (.a(net183),
    .b(u_dcfifo_tx_u_din_buffer_data[57]),
    .c(net181),
    .d(u_dcfifo_tx_u_din_buffer_data[89]),
    .o1(n3085));
 b15aoi022ar1n24x5 U3591 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[25]),
    .c(net189),
    .d(u_dcfifo_tx_u_din_buffer_data[217]),
    .o1(n3084));
 b15aoi022al1n12x5 U3592 (.a(net175),
    .b(u_dcfifo_tx_u_din_buffer_data[249]),
    .c(net186),
    .d(u_dcfifo_tx_u_din_buffer_data[153]),
    .o1(n3083));
 b15nand04as1n16x5 U3593 (.a(n3086),
    .b(n3085),
    .c(n3084),
    .d(n3083),
    .o1(n3087));
 b15nonb02as1n16x5 U3594 (.a(n3087),
    .b(net136),
    .out0(u_device_sm_N199));
 b15aoi022ah1n16x5 U3595 (.a(net181),
    .b(u_dcfifo_tx_u_din_buffer_data[85]),
    .c(net186),
    .d(u_dcfifo_tx_u_din_buffer_data[149]),
    .o1(n3091));
 b15aoi022ah1n12x5 U3596 (.a(net183),
    .b(u_dcfifo_tx_u_din_buffer_data[53]),
    .c(net175),
    .d(u_dcfifo_tx_u_din_buffer_data[245]),
    .o1(n3090));
 b15aoi022ar1n12x5 U3597 (.a(net173),
    .b(u_dcfifo_tx_u_din_buffer_data[181]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[117]),
    .o1(n3089));
 b15aoi022ar1n32x5 U3598 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[21]),
    .c(net189),
    .d(u_dcfifo_tx_u_din_buffer_data[213]),
    .o1(n3088));
 b15nand04as1n16x5 U3599 (.a(n3091),
    .b(n3090),
    .c(n3089),
    .d(n3088),
    .o1(n3092));
 b15nonb02as1n16x5 U3600 (.a(n3092),
    .b(net136),
    .out0(u_device_sm_N195));
 b15aoi022ah1n08x5 U3601 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[24]),
    .c(net173),
    .d(u_dcfifo_tx_u_din_buffer_data[184]),
    .o1(n3096));
 b15aoi022as1n16x5 U3602 (.a(net181),
    .b(u_dcfifo_tx_u_din_buffer_data[88]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[120]),
    .o1(n3095));
 b15aoi022an1n08x5 U3603 (.a(net183),
    .b(u_dcfifo_tx_u_din_buffer_data[56]),
    .c(net186),
    .d(u_dcfifo_tx_u_din_buffer_data[152]),
    .o1(n3094));
 b15aoi022an1n12x5 U3604 (.a(net189),
    .b(u_dcfifo_tx_u_din_buffer_data[216]),
    .c(net175),
    .d(u_dcfifo_tx_u_din_buffer_data[248]),
    .o1(n3093));
 b15nand04as1n16x5 U3605 (.a(n3096),
    .b(n3095),
    .c(n3094),
    .d(n3093),
    .o1(n3097));
 b15nonb02as1n16x5 U3606 (.a(n3097),
    .b(net137),
    .out0(u_device_sm_N198));
 b15aoi022ah1n06x5 U3607 (.a(net180),
    .b(u_dcfifo_tx_u_din_buffer_data[74]),
    .c(net172),
    .d(u_dcfifo_tx_u_din_buffer_data[170]),
    .o1(n3101));
 b15aoi022an1n12x5 U3608 (.a(net182),
    .b(u_dcfifo_tx_u_din_buffer_data[42]),
    .c(net188),
    .d(u_dcfifo_tx_u_din_buffer_data[202]),
    .o1(n3100));
 b15aoi022an1n24x5 U3609 (.a(net174),
    .b(u_dcfifo_tx_u_din_buffer_data[234]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[106]),
    .o1(n3099));
 b15aoi022aq1n16x5 U3610 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[10]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[138]),
    .o1(n3098));
 b15nand04as1n16x5 U3611 (.a(n3101),
    .b(n3100),
    .c(n3099),
    .d(n3098),
    .o1(n3102));
 b15nonb02an1n02x5 U3612 (.a(n3102),
    .b(net135),
    .out0(u_device_sm_N184));
 b15aoi022aq1n12x5 U3613 (.a(net183),
    .b(u_dcfifo_tx_u_din_buffer_data[54]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[118]),
    .o1(n3106));
 b15aoi022aq1n12x5 U3614 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[22]),
    .c(net181),
    .d(u_dcfifo_tx_u_din_buffer_data[86]),
    .o1(n3105));
 b15aoi022aq1n12x5 U3615 (.a(net189),
    .b(u_dcfifo_tx_u_din_buffer_data[214]),
    .c(net173),
    .d(u_dcfifo_tx_u_din_buffer_data[182]),
    .o1(n3104));
 b15aoi022ar1n24x5 U3616 (.a(net175),
    .b(u_dcfifo_tx_u_din_buffer_data[246]),
    .c(net186),
    .d(u_dcfifo_tx_u_din_buffer_data[150]),
    .o1(n3103));
 b15nand04as1n16x5 U3617 (.a(n3106),
    .b(n3105),
    .c(n3104),
    .d(n3103),
    .o1(n3107));
 b15nonb02ah1n16x5 U3618 (.a(n3107),
    .b(net137),
    .out0(u_device_sm_N196));
 b15aoi022ah1n12x5 U3619 (.a(net188),
    .b(u_dcfifo_tx_u_din_buffer_data[207]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[111]),
    .o1(n3111));
 b15aoi022an1n16x5 U3620 (.a(net180),
    .b(u_dcfifo_tx_u_din_buffer_data[79]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[143]),
    .o1(n3110));
 b15aoi022ah1n08x5 U3621 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[15]),
    .c(net174),
    .d(u_dcfifo_tx_u_din_buffer_data[239]),
    .o1(n3109));
 b15aoi022ah1n08x5 U3622 (.a(net182),
    .b(u_dcfifo_tx_u_din_buffer_data[47]),
    .c(net172),
    .d(u_dcfifo_tx_u_din_buffer_data[175]),
    .o1(n3108));
 b15nand04as1n16x5 U3623 (.a(n3111),
    .b(n3110),
    .c(n3109),
    .d(n3108),
    .o1(n3112));
 b15nonb02an1n02x5 U3624 (.a(n3112),
    .b(net135),
    .out0(u_device_sm_N189));
 b15ztpn00an1n08x5 PHY_18 ();
 b15aoi022aq1n12x5 U3626 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[20]),
    .c(net183),
    .d(u_dcfifo_tx_u_din_buffer_data[52]),
    .o1(n3117));
 b15aoi022ah1n06x5 U3627 (.a(net189),
    .b(u_dcfifo_tx_u_din_buffer_data[212]),
    .c(net175),
    .d(u_dcfifo_tx_u_din_buffer_data[244]),
    .o1(n3116));
 b15aoi022al1n24x5 U3628 (.a(net181),
    .b(u_dcfifo_tx_u_din_buffer_data[84]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[116]),
    .o1(n3115));
 b15aoi022ah1n16x5 U3629 (.a(net173),
    .b(u_dcfifo_tx_u_din_buffer_data[180]),
    .c(net186),
    .d(u_dcfifo_tx_u_din_buffer_data[148]),
    .o1(n3114));
 b15nand04as1n16x5 U3630 (.a(n3117),
    .b(n3116),
    .c(n3115),
    .d(n3114),
    .o1(n3118));
 b15nonb02as1n16x5 U3631 (.a(n3118),
    .b(net136),
    .out0(u_device_sm_N194));
 b15aoi022as1n08x5 U3632 (.a(net173),
    .b(u_dcfifo_tx_u_din_buffer_data[186]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[122]),
    .o1(n3122));
 b15aoi022as1n08x5 U3633 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[26]),
    .c(net183),
    .d(u_dcfifo_tx_u_din_buffer_data[58]),
    .o1(n3121));
 b15aoi022ah1n08x5 U3634 (.a(net189),
    .b(u_dcfifo_tx_u_din_buffer_data[218]),
    .c(net175),
    .d(u_dcfifo_tx_u_din_buffer_data[250]),
    .o1(n3120));
 b15aoi022ar1n32x5 U3635 (.a(net181),
    .b(u_dcfifo_tx_u_din_buffer_data[90]),
    .c(net186),
    .d(u_dcfifo_tx_u_din_buffer_data[154]),
    .o1(n3119));
 b15nand04as1n16x5 U3636 (.a(n3122),
    .b(n3121),
    .c(n3120),
    .d(n3119),
    .o1(n3123));
 b15nonb02al1n16x5 U3637 (.a(n3123),
    .b(net137),
    .out0(u_device_sm_N200));
 b15aoi022as1n06x5 U3638 (.a(net173),
    .b(u_dcfifo_tx_u_din_buffer_data[189]),
    .c(net175),
    .d(u_dcfifo_tx_u_din_buffer_data[253]),
    .o1(n3127));
 b15aoi022as1n16x5 U3639 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[29]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[125]),
    .o1(n3126));
 b15aoi022as1n08x5 U3640 (.a(net183),
    .b(u_dcfifo_tx_u_din_buffer_data[61]),
    .c(net189),
    .d(u_dcfifo_tx_u_din_buffer_data[221]),
    .o1(n3125));
 b15aoi022an1n24x5 U3641 (.a(net181),
    .b(u_dcfifo_tx_u_din_buffer_data[93]),
    .c(net186),
    .d(u_dcfifo_tx_u_din_buffer_data[157]),
    .o1(n3124));
 b15nand04as1n16x5 U3642 (.a(n3127),
    .b(n3126),
    .c(n3125),
    .d(n3124),
    .o1(n3128));
 b15nonb02as1n08x5 U3643 (.a(n3128),
    .b(net136),
    .out0(u_device_sm_N203));
 b15aoi022aq1n08x5 U3644 (.a(net183),
    .b(u_dcfifo_tx_u_din_buffer_data[49]),
    .c(net173),
    .d(u_dcfifo_tx_u_din_buffer_data[177]),
    .o1(n3134));
 b15aoi022an1n12x5 U3645 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[17]),
    .c(net189),
    .d(u_dcfifo_tx_u_din_buffer_data[209]),
    .o1(n3133));
 b15aoi022al1n32x5 U3646 (.a(net175),
    .b(u_dcfifo_tx_u_din_buffer_data[241]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[113]),
    .o1(n3132));
 b15aoi022al1n24x5 U3647 (.a(net181),
    .b(u_dcfifo_tx_u_din_buffer_data[81]),
    .c(net186),
    .d(u_dcfifo_tx_u_din_buffer_data[145]),
    .o1(n3131));
 b15nand04ah1n16x5 U3648 (.a(n3134),
    .b(n3133),
    .c(n3132),
    .d(n3131),
    .o1(n3135));
 b15nonb02as1n16x5 U3649 (.a(n3135),
    .b(net136),
    .out0(u_device_sm_N191));
 b15aoi022ah1n06x5 U3650 (.a(net188),
    .b(u_dcfifo_tx_u_din_buffer_data[201]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[137]),
    .o1(n3139));
 b15aoi022ah1n12x5 U3651 (.a(net174),
    .b(u_dcfifo_tx_u_din_buffer_data[233]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[105]),
    .o1(n3138));
 b15aoi022aq1n12x5 U3652 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[9]),
    .c(net182),
    .d(u_dcfifo_tx_u_din_buffer_data[41]),
    .o1(n3137));
 b15aoi022aq1n12x5 U3653 (.a(net180),
    .b(u_dcfifo_tx_u_din_buffer_data[73]),
    .c(net172),
    .d(u_dcfifo_tx_u_din_buffer_data[169]),
    .o1(n3136));
 b15nand04an1n16x5 U3654 (.a(n3139),
    .b(n3138),
    .c(n3137),
    .d(n3136),
    .o1(n3140));
 b15nonb02aq1n06x5 U3655 (.a(n3140),
    .b(net136),
    .out0(u_device_sm_N183));
 b15aoi022al1n12x5 U3656 (.a(net178),
    .b(u_dcfifo_tx_u_din_buffer_data[28]),
    .c(net181),
    .d(u_dcfifo_tx_u_din_buffer_data[92]),
    .o1(n3146));
 b15aoi022as1n24x5 U3657 (.a(net186),
    .b(u_dcfifo_tx_u_din_buffer_data[156]),
    .c(net170),
    .d(u_dcfifo_tx_u_din_buffer_data[124]),
    .o1(n3145));
 b15aoi022as1n08x5 U3658 (.a(net173),
    .b(u_dcfifo_tx_u_din_buffer_data[188]),
    .c(net175),
    .d(u_dcfifo_tx_u_din_buffer_data[252]),
    .o1(n3144));
 b15aoi022ah1n08x5 U3659 (.a(net183),
    .b(u_dcfifo_tx_u_din_buffer_data[60]),
    .c(net189),
    .d(u_dcfifo_tx_u_din_buffer_data[220]),
    .o1(n3143));
 b15nand04ah1n16x5 U3660 (.a(n3146),
    .b(n3145),
    .c(n3144),
    .d(n3143),
    .o1(n3148));
 b15nonb02ar1n16x5 U3661 (.a(n3148),
    .b(net136),
    .out0(u_device_sm_N202));
 b15aoi022an1n16x5 U3662 (.a(net182),
    .b(u_dcfifo_tx_u_din_buffer_data[40]),
    .c(net174),
    .d(u_dcfifo_tx_u_din_buffer_data[232]),
    .o1(n3153));
 b15aoi022an1n32x5 U3663 (.a(net172),
    .b(u_dcfifo_tx_u_din_buffer_data[168]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[136]),
    .o1(n3152));
 b15aoi022ar1n12x5 U3664 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[8]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[104]),
    .o1(n3151));
 b15aoi022al1n12x5 U3665 (.a(net188),
    .b(u_dcfifo_tx_u_din_buffer_data[200]),
    .c(net180),
    .d(u_dcfifo_tx_u_din_buffer_data[72]),
    .o1(n3150));
 b15nand04as1n16x5 U3666 (.a(n3153),
    .b(n3152),
    .c(n3151),
    .d(n3150),
    .o1(n3155));
 b15nonb02ah1n04x5 U3667 (.a(n3155),
    .b(net135),
    .out0(u_device_sm_N182));
 b15aoi022an1n16x5 U3668 (.a(net188),
    .b(u_dcfifo_tx_u_din_buffer_data[199]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[103]),
    .o1(n3160));
 b15aoi022al1n24x5 U3669 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[7]),
    .c(net182),
    .d(u_dcfifo_tx_u_din_buffer_data[39]),
    .o1(n3159));
 b15aoi022al1n16x5 U3671 (.a(net174),
    .b(u_dcfifo_tx_u_din_buffer_data[231]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[135]),
    .o1(n3158));
 b15aoi022ar1n16x5 U3672 (.a(net180),
    .b(u_dcfifo_tx_u_din_buffer_data[71]),
    .c(net172),
    .d(u_dcfifo_tx_u_din_buffer_data[167]),
    .o1(n3157));
 b15nand04as1n16x5 U3673 (.a(n3160),
    .b(n3159),
    .c(n3158),
    .d(n3157),
    .o1(n3164));
 b15aoi022an1n02x5 U3674 (.a(n3663),
    .b(u_device_sm_u_spiregs_n[9]),
    .c(n3665),
    .d(u_device_sm_u_spiregs_n[1]),
    .o1(n3161));
 b15aob012aq1n08x5 U3675 (.a(n3161),
    .b(n3664),
    .c(u_device_sm_s_dummy_cycles[7]),
    .out0(n3162));
 b15oaoi13as1n08x5 U3676 (.a(n3162),
    .b(n3666),
    .c(u_device_sm_u_spiregs_reg0[7]),
    .d(n3228),
    .o1(n3163));
 b15oab012al1n02x5 U3677 (.a(n3163),
    .b(n3164),
    .c(net139),
    .out0(u_device_sm_N181));
 b15aoi022aq1n32x5 U3678 (.a(net172),
    .b(u_dcfifo_tx_u_din_buffer_data[160]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[128]),
    .o1(n3172));
 b15aoi022ar1n24x5 U3679 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[0]),
    .c(net180),
    .d(u_dcfifo_tx_u_din_buffer_data[64]),
    .o1(n3171));
 b15aoi022as1n08x5 U3680 (.a(net182),
    .b(u_dcfifo_tx_u_din_buffer_data[32]),
    .c(net174),
    .d(u_dcfifo_tx_u_din_buffer_data[224]),
    .o1(n3170));
 b15aoi022ah1n16x5 U3681 (.a(net188),
    .b(u_dcfifo_tx_u_din_buffer_data[192]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[96]),
    .o1(n3169));
 b15nand04as1n16x5 U3682 (.a(n3172),
    .b(n3171),
    .c(n3170),
    .d(n3169),
    .o1(n3179));
 b15aoi022aq1n12x5 U3683 (.a(n3663),
    .b(u_device_sm_u_spiregs_n[16]),
    .c(n3665),
    .d(u_device_sm_u_spiregs_n[8]),
    .o1(n3173));
 b15aoai13ah1n03x5 U3684 (.a(n3173),
    .b(n3174),
    .c(n3176),
    .d(n3817),
    .o1(n3177));
 b15aoi012aq1n08x5 U3685 (.a(n3177),
    .b(u_device_sm_s_dummy_cycles[0]),
    .c(n3664),
    .o1(n3178));
 b15oab012as1n08x5 U3686 (.c(n3179),
    .a(n3178),
    .b(net139),
    .out0(u_device_sm_N174));
 b15aoi022ar1n16x5 U3687 (.a(net182),
    .b(u_dcfifo_tx_u_din_buffer_data[34]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[98]),
    .o1(n3183));
 b15aoi022an1n24x5 U3688 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[2]),
    .c(net174),
    .d(u_dcfifo_tx_u_din_buffer_data[226]),
    .o1(n3182));
 b15aoi022ar1n32x5 U3689 (.a(net172),
    .b(u_dcfifo_tx_u_din_buffer_data[162]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[130]),
    .o1(n3181));
 b15aoi022al1n12x5 U3690 (.a(net188),
    .b(u_dcfifo_tx_u_din_buffer_data[194]),
    .c(net180),
    .d(u_dcfifo_tx_u_din_buffer_data[66]),
    .o1(n3180));
 b15nand04as1n16x5 U3691 (.a(n3183),
    .b(n3182),
    .c(n3181),
    .d(n3180),
    .o1(n3188));
 b15aoi022as1n04x5 U3692 (.a(n3663),
    .b(u_device_sm_u_spiregs_n[14]),
    .c(n3665),
    .d(u_device_sm_u_spiregs_n[6]),
    .o1(n3184));
 b15oai012ah1n12x5 U3693 (.a(n3184),
    .b(n3821),
    .c(n3185),
    .o1(n3186));
 b15oaoi13as1n08x5 U3694 (.a(n3186),
    .b(n3666),
    .c(u_device_sm_u_spiregs_reg0[2]),
    .d(n3228),
    .o1(n3187));
 b15oab012ar1n04x5 U3695 (.a(n3187),
    .b(net138),
    .c(n3188),
    .out0(u_device_sm_N176));
 b15aoi022as1n06x5 U3696 (.a(net188),
    .b(u_dcfifo_tx_u_din_buffer_data[197]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[133]),
    .o1(n3192));
 b15aoi022an1n08x5 U3697 (.a(net182),
    .b(u_dcfifo_tx_u_din_buffer_data[37]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[101]),
    .o1(n3191));
 b15aoi022as1n08x5 U3698 (.a(net180),
    .b(u_dcfifo_tx_u_din_buffer_data[69]),
    .c(net172),
    .d(u_dcfifo_tx_u_din_buffer_data[165]),
    .o1(n3190));
 b15aoi022al1n32x5 U3699 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[5]),
    .c(net174),
    .d(u_dcfifo_tx_u_din_buffer_data[229]),
    .o1(n3189));
 b15nand04as1n16x5 U3700 (.a(n3192),
    .b(n3191),
    .c(n3190),
    .d(n3189),
    .o1(n3198));
 b15aoi022al1n08x5 U3701 (.a(n3663),
    .b(u_device_sm_u_spiregs_n[11]),
    .c(n3665),
    .d(u_device_sm_u_spiregs_n[3]),
    .o1(n3193));
 b15oai012as1n12x5 U3702 (.a(n3193),
    .b(n3821),
    .c(n3194),
    .o1(n3196));
 b15oaoi13as1n08x5 U3703 (.a(n3196),
    .b(n3666),
    .c(u_device_sm_u_spiregs_reg0[5]),
    .d(n3228),
    .o1(n3197));
 b15oab012aq1n03x5 U3704 (.a(n3197),
    .b(net138),
    .c(n3198),
    .out0(u_device_sm_N179));
 b15aoi022ah1n06x5 U3705 (.a(net188),
    .b(u_dcfifo_tx_u_din_buffer_data[198]),
    .c(net180),
    .d(u_dcfifo_tx_u_din_buffer_data[70]),
    .o1(n3202));
 b15aoi022aq1n12x5 U3706 (.a(net174),
    .b(u_dcfifo_tx_u_din_buffer_data[230]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[102]),
    .o1(n3201));
 b15aoi022aq1n12x5 U3707 (.a(net182),
    .b(u_dcfifo_tx_u_din_buffer_data[38]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[134]),
    .o1(n3200));
 b15aoi022aq1n08x5 U3708 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[6]),
    .c(net172),
    .d(u_dcfifo_tx_u_din_buffer_data[166]),
    .o1(n3199));
 b15nand04as1n16x5 U3709 (.a(n3202),
    .b(n3201),
    .c(n3200),
    .d(n3199),
    .o1(n3206));
 b15aoi022ah1n08x5 U3710 (.a(n3664),
    .b(u_device_sm_s_dummy_cycles[6]),
    .c(n3665),
    .d(u_device_sm_u_spiregs_n[2]),
    .o1(n3203));
 b15aob012aq1n12x5 U3711 (.a(n3203),
    .b(n3663),
    .c(u_device_sm_u_spiregs_n[10]),
    .out0(n3204));
 b15oaoi13as1n08x5 U3712 (.a(n3204),
    .b(n3666),
    .c(u_device_sm_u_spiregs_reg0[6]),
    .d(n3228),
    .o1(n3205));
 b15oab012ah1n03x5 U3713 (.a(n3205),
    .b(net138),
    .c(n3206),
    .out0(u_device_sm_N180));
 b15aoi022ar1n12x5 U3714 (.a(net182),
    .b(u_dcfifo_tx_u_din_buffer_data[35]),
    .c(net172),
    .d(u_dcfifo_tx_u_din_buffer_data[163]),
    .o1(n3212));
 b15aoi022an1n16x5 U3715 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[3]),
    .c(net180),
    .d(u_dcfifo_tx_u_din_buffer_data[67]),
    .o1(n3211));
 b15aoi022al1n16x5 U3716 (.a(net188),
    .b(u_dcfifo_tx_u_din_buffer_data[195]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[131]),
    .o1(n3210));
 b15aoi022as1n08x5 U3717 (.a(net174),
    .b(u_dcfifo_tx_u_din_buffer_data[227]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[99]),
    .o1(n3209));
 b15nand04as1n16x5 U3718 (.a(n3212),
    .b(n3211),
    .c(n3210),
    .d(n3209),
    .o1(n3216));
 b15aoi022an1n06x5 U3719 (.a(n3663),
    .b(u_device_sm_u_spiregs_n[13]),
    .c(n3665),
    .d(u_device_sm_u_spiregs_n[5]),
    .o1(n3213));
 b15aob012an1n12x5 U3720 (.a(n3213),
    .b(n3664),
    .c(u_device_sm_s_dummy_cycles[3]),
    .out0(n3214));
 b15oaoi13as1n08x5 U3721 (.a(n3214),
    .b(n3666),
    .c(u_device_sm_u_spiregs_reg0[3]),
    .d(n3228),
    .o1(n3215));
 b15oab012aq1n06x5 U3722 (.a(n3215),
    .b(net139),
    .c(n3216),
    .out0(u_device_sm_N177));
 b15aoi022aq1n16x5 U3723 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[4]),
    .c(net188),
    .d(u_dcfifo_tx_u_din_buffer_data[196]),
    .o1(n3225));
 b15aoi022ah1n08x5 U3724 (.a(net182),
    .b(u_dcfifo_tx_u_din_buffer_data[36]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[100]),
    .o1(n3224));
 b15aoi022aq1n16x5 U3725 (.a(net172),
    .b(u_dcfifo_tx_u_din_buffer_data[164]),
    .c(net174),
    .d(u_dcfifo_tx_u_din_buffer_data[228]),
    .o1(n3223));
 b15aoi022as1n08x5 U3726 (.a(net180),
    .b(u_dcfifo_tx_u_din_buffer_data[68]),
    .c(net185),
    .d(u_dcfifo_tx_u_din_buffer_data[132]),
    .o1(n3222));
 b15nand04as1n16x5 U3727 (.a(n3225),
    .b(n3224),
    .c(n3223),
    .d(n3222),
    .o1(n3230));
 b15aoi022ah1n06x5 U3728 (.a(n3663),
    .b(u_device_sm_u_spiregs_n[12]),
    .c(n3665),
    .d(u_device_sm_u_spiregs_n[4]),
    .o1(n3226));
 b15aob012al1n16x5 U3729 (.a(n3226),
    .b(n3664),
    .c(u_device_sm_s_dummy_cycles[4]),
    .out0(n3227));
 b15oaoi13as1n08x5 U3730 (.a(n3227),
    .b(n3666),
    .c(u_device_sm_u_spiregs_reg0[4]),
    .d(n3228),
    .o1(n3229));
 b15oab012al1n04x5 U3731 (.a(n3229),
    .b(net138),
    .c(n3230),
    .out0(u_device_sm_N178));
 b15ztpn00an1n08x5 PHY_17 ();
 b15inv000aq1n16x5 U3733 (.a(net2465),
    .o1(n3276));
 b15nor002ah1n12x5 U3734 (.a(net1975),
    .b(n3276),
    .o1(net62));
 b15inv000an1n03x5 U3735 (.a(net131),
    .o1(n3234));
 b15nandp3ar1n04x5 U3736 (.a(net62),
    .b(net8),
    .c(n3234),
    .o1(n3233));
 b15aoai13as1n08x5 U3737 (.a(n3233),
    .b(n3234),
    .c(net8),
    .d(net62),
    .o1(n604));
 b15nandp2ah1n04x5 U3738 (.a(u_dcfifo_rx_u_dout_read_token[7]),
    .b(u_dcfifo_rx_u_dout_read_token[6]),
    .o1(n3269));
 b15inv040as1n05x5 U3739 (.a(n3269),
    .o1(n3255));
 b15aoi012an1n12x5 U3740 (.a(n3255),
    .b(net325),
    .c(u_dcfifo_rx_u_dout_read_token[4]),
    .o1(n3346));
 b15oai012al1n06x5 U3741 (.a(n3239),
    .b(net328),
    .c(n3255),
    .o1(n3258));
 b15oai012al1n03x5 U3742 (.a(net330),
    .b(net328),
    .c(net331),
    .o1(n3237));
 b15oai012ar1n04x5 U3743 (.a(u_dcfifo_rx_u_dout_read_token[4]),
    .b(net326),
    .c(net325),
    .o1(n3236));
 b15qgbna2an1n10x5 U3744 (.a(u_dcfifo_rx_u_dout_read_token[1]),
    .b(u_dcfifo_rx_u_dout_read_token[2]),
    .o1(n3243));
 b15nandp2ah1n16x5 U3745 (.a(net326),
    .b(u_dcfifo_rx_u_dout_read_token[2]),
    .o1(n3344));
 b15nandp2ah1n16x5 U3746 (.a(n3243),
    .b(n3344),
    .o1(n3348));
 b15inv020as1n10x5 U3747 (.a(n3348),
    .o1(n3358));
 b15oai022an1n06x5 U3748 (.a(n3237),
    .b(n3236),
    .c(n3358),
    .d(n3235),
    .o1(n3254));
 b15nand02ah1n12x5 U3749 (.a(u_dcfifo_rx_u_dout_read_token[0]),
    .b(u_dcfifo_rx_u_dout_read_token[7]),
    .o1(n3245));
 b15nandp2ah1n16x5 U3750 (.a(u_dcfifo_rx_u_dout_read_token[0]),
    .b(u_dcfifo_rx_u_dout_read_token[1]),
    .o1(n3345));
 b15nand02as1n24x5 U3751 (.a(n3245),
    .b(n3345),
    .o1(n3354));
 b15inv020ar1n06x5 U3752 (.a(n3354),
    .o1(n3244));
 b15inv040al1n02x5 U3753 (.a(n3238),
    .o1(n3240));
 b15oai112as1n06x5 U3754 (.a(u_dcfifo_rx_u_dout_read_token[5]),
    .b(u_dcfifo_rx_u_dout_read_token[6]),
    .c(n3240),
    .d(n3239),
    .o1(n3241));
 b15aoai13ah1n03x5 U3755 (.a(n3241),
    .b(n3242),
    .c(n3244),
    .d(n3243),
    .o1(n3253));
 b15nandp2ar1n03x5 U3756 (.a(u_dcfifo_rx_u_dout_read_token[4]),
    .b(net326),
    .o1(n3247));
 b15oai022ar1n04x5 U3757 (.a(n3248),
    .b(n3247),
    .c(n3246),
    .d(n3245),
    .o1(n3252));
 b15nandp2ar1n02x5 U3758 (.a(net330),
    .b(net331),
    .o1(n3250));
 b15nand02al1n04x5 U3759 (.a(net333),
    .b(net336),
    .o1(n3249));
 b15oai022aq1n02x5 U3760 (.a(n3250),
    .b(n3344),
    .c(n3345),
    .d(n3249),
    .o1(n3251));
 b15nor004an1n06x5 U3761 (.a(n3254),
    .b(n3253),
    .c(n3252),
    .d(n3251),
    .o1(n3257));
 b15oai112ah1n06x5 U3762 (.a(u_dcfifo_rx_write_token[0]),
    .b(net327),
    .c(n3255),
    .d(n3354),
    .o1(n3256));
 b15oai112ah1n12x5 U3763 (.a(n3257),
    .b(n3256),
    .c(n3346),
    .d(n3258),
    .o1(u_dcfifo_rx_u_din_full_full_dn));
 b15aobi12as1n16x5 U3764 (.a(net53),
    .b(u_dcfifo_tx_u_din_full_full_up),
    .c(net2329),
    .out0(u_dcfifo_tx_u_din_write_enable));
 b15aoi022al1n16x5 U3765 (.a(u_dcfifo_tx_write_token[7]),
    .b(net312),
    .c(net314),
    .d(u_dcfifo_tx_write_token[4]),
    .o1(n3259));
 b15nand02ar1n24x5 U3766 (.a(net322),
    .b(net324),
    .o1(n3661));
 b15nand02as1n24x5 U3767 (.a(net318),
    .b(net320),
    .o1(n3639));
 b15nandp3as1n24x5 U3768 (.a(n3259),
    .b(n3661),
    .c(n3639),
    .o1(n3286));
 b15oai012al1n32x5 U3769 (.a(net311),
    .b(net309),
    .c(net314),
    .o1(n3643));
 b15oai012as1n16x5 U3770 (.a(net320),
    .b(net322),
    .c(net318),
    .o1(n3636));
 b15nandp2ah1n24x5 U3771 (.a(n3643),
    .b(n3636),
    .o1(n3282));
 b15inv040an1n08x5 U3772 (.a(n3282),
    .o1(n3280));
 b15and002an1n03x5 U3773 (.a(u_dcfifo_tx_write_token[7]),
    .b(net312),
    .o(n3260));
 b15oaoi13as1n08x5 U3774 (.a(n3260),
    .b(u_dcfifo_tx_write_token[5]),
    .c(net312),
    .d(net316),
    .o1(n3654));
 b15aob012as1n24x5 U3775 (.a(n3654),
    .b(u_dcfifo_tx_write_token[3]),
    .c(net316),
    .out0(n3279));
 b15nandp3as1n24x5 U3776 (.a(n3280),
    .b(u_dcfifo_tx_u_din_write_enable),
    .c(n3279),
    .o1(n3278));
 b15nor002ah1n32x5 U3777 (.a(n3286),
    .b(n3278),
    .o1(u_dcfifo_tx_u_din_buffer_N30));
 b15nandp3as1n24x5 U3778 (.a(u_dcfifo_tx_u_din_write_enable),
    .b(n3282),
    .c(n3279),
    .o1(n3277));
 b15norp02as1n32x5 U3779 (.a(n3286),
    .b(n3277),
    .o1(u_dcfifo_tx_u_din_buffer_N32));
 b15inv020ar1n06x5 U3780 (.a(u_dcfifo_rx_u_dout_read_token[3]),
    .o1(n3262));
 b15aoai13as1n03x5 U3781 (.a(u_dcfifo_rx_u_dout_read_token[4]),
    .b(u_dcfifo_rx_u_dout_write_token_dn[5]),
    .c(net325),
    .d(u_dcfifo_rx_u_dout_write_token_dn[6]),
    .o1(n3261));
 b15oaoi13as1n08x5 U3782 (.a(n3261),
    .b(u_dcfifo_rx_u_dout_write_token_dn[5]),
    .c(u_dcfifo_rx_u_dout_write_token_dn[4]),
    .d(n3262),
    .o1(n3274));
 b15inv000as1n05x5 U3783 (.a(u_dcfifo_rx_u_dout_write_token_dn[2]),
    .o1(n3264));
 b15inv040as1n04x5 U3784 (.a(u_dcfifo_rx_u_dout_write_token_dn[0]),
    .o1(n3270));
 b15nand04as1n02x5 U3785 (.a(u_dcfifo_rx_u_dout_read_token[7]),
    .b(u_dcfifo_rx_u_dout_read_token[0]),
    .c(u_dcfifo_rx_u_dout_write_token_dn[1]),
    .d(n3270),
    .o1(n3263));
 b15oai013as1n06x5 U3786 (.a(n3263),
    .b(net2366),
    .c(n3345),
    .d(n3264),
    .o1(n3273));
 b15inv040ar1n03x5 U3787 (.a(u_dcfifo_rx_u_dout_write_token_dn[4]),
    .o1(n3266));
 b15nand04ah1n04x5 U3788 (.a(u_dcfifo_rx_u_dout_read_token[1]),
    .b(u_dcfifo_rx_u_dout_read_token[2]),
    .c(u_dcfifo_rx_u_dout_write_token_dn[3]),
    .d(n3264),
    .o1(n3265));
 b15oai013an1n12x5 U3789 (.a(n3265),
    .b(u_dcfifo_rx_u_dout_write_token_dn[3]),
    .c(n3266),
    .d(n3344),
    .o1(n3272));
 b15inv000al1n02x5 U3790 (.a(u_dcfifo_rx_u_dout_write_token_dn[6]),
    .o1(n3267));
 b15nand04as1n03x5 U3791 (.a(u_dcfifo_rx_u_dout_read_token[5]),
    .b(u_dcfifo_rx_u_dout_read_token[6]),
    .c(u_dcfifo_rx_u_dout_write_token_dn[7]),
    .d(n3267),
    .o1(n3268));
 b15oai013al1n08x5 U3792 (.a(n3268),
    .b(u_dcfifo_rx_u_dout_write_token_dn[7]),
    .c(n3270),
    .d(n3269),
    .o1(n3271));
 b15nor004as1n12x5 U3793 (.a(n3274),
    .b(n3273),
    .c(n3272),
    .d(n3271),
    .o1(n2723));
 b15inv000ar1n12x5 U3794 (.a(n2723),
    .o1(n3308));
 b15nonb03as1n06x5 U3795 (.a(u_syncro_valid_reg[1]),
    .b(net344),
    .c(u_syncro_valid_reg[2]),
    .out0(n3307));
 b15aoi012aq1n04x5 U3796 (.a(net361),
    .b(rd_wr_sync),
    .c(n3307),
    .o1(n3275));
 b15aoi013as1n08x5 U3797 (.a(n3275),
    .b(net362),
    .c(n3276),
    .d(n3308),
    .o1(u_spi_device_tlul_plug_state_next[1]));
 b15inv020an1n64x5 U3798 (.a(n3286),
    .o1(n3284));
 b15norp02al1n48x5 U3799 (.a(n3284),
    .b(n3277),
    .o1(u_dcfifo_tx_u_din_buffer_N33));
 b15norp02al1n48x5 U3800 (.a(n3284),
    .b(n3278),
    .o1(u_dcfifo_tx_u_din_buffer_N31));
 b15nonb02al1n16x5 U3801 (.a(u_dcfifo_tx_u_din_write_enable),
    .b(n3279),
    .out0(n3283));
 b15nand02aq1n32x5 U3802 (.a(n3280),
    .b(n3283),
    .o1(n3281));
 b15norp02ar1n48x5 U3803 (.a(n3284),
    .b(n3281),
    .o1(u_dcfifo_tx_u_din_buffer_N27));
 b15norp02aq1n48x5 U3804 (.a(n3286),
    .b(n3281),
    .o1(u_dcfifo_tx_u_din_buffer_N26));
 b15nand02an1n48x5 U3805 (.a(n3283),
    .b(n3282),
    .o1(n3285));
 b15norp02as1n48x5 U3806 (.a(n3284),
    .b(n3285),
    .o1(u_dcfifo_tx_u_din_buffer_N29));
 b15nor002aq1n32x5 U3807 (.a(n3286),
    .b(n3285),
    .o1(u_dcfifo_tx_u_din_buffer_N28));
 b15inv020as1n05x5 U3808 (.a(net48),
    .o1(n3288));
 b15aboi22al1n12x5 U3809 (.a(net52),
    .b(n3288),
    .c(net48),
    .d(net52),
    .out0(n3305));
 b15inv000aq1n02x5 U3810 (.a(net49),
    .o1(n3302));
 b15xor002ar1n03x5 U3811 (.a(net10),
    .b(net52),
    .out0(n3294));
 b15xor002an1n04x5 U3812 (.a(net52),
    .b(net54),
    .out0(n3290));
 b15qgbin1an1n05x5 U3813 (.a(net51),
    .o1(n3298));
 b15aboi22an1n12x5 U3814 (.a(net50),
    .b(net51),
    .c(net50),
    .d(n3298),
    .out0(n3287));
 b15qgbxo2an1n05x5 U3815 (.a(net49),
    .b(n3287),
    .out0(n3289));
 b15xor002aq1n06x5 U3816 (.a(n3289),
    .b(n3288),
    .out0(n3291));
 b15xor002al1n02x5 U3817 (.a(n3290),
    .b(n3291),
    .out0(n3293));
 b15xnr002ar1n03x5 U3818 (.a(net9),
    .b(n3291),
    .out0(n3292));
 b15nor004aq1n02x5 U3819 (.a(net19),
    .b(n3294),
    .c(n3293),
    .d(n3292),
    .o1(n3296));
 b15nand04aq1n02x5 U3820 (.a(net19),
    .b(n3294),
    .c(n3293),
    .d(n3292),
    .o1(n3295));
 b15nanb02ah1n03x5 U3821 (.a(n3296),
    .b(n3295),
    .out0(n3300));
 b15oai022ar1n02x5 U3822 (.a(n3298),
    .b(net14),
    .c(net13),
    .d(net50),
    .o1(n3297));
 b15aoi122aq1n02x5 U3823 (.a(n3297),
    .b(n3298),
    .c(net14),
    .d(net50),
    .e(net13),
    .o1(n3299));
 b15oai112aq1n02x5 U3824 (.a(n3300),
    .b(n3299),
    .c(n3302),
    .d(net12),
    .o1(n3301));
 b15aoi012as1n02x5 U3825 (.a(n3301),
    .b(n3302),
    .c(net12),
    .o1(n3303));
 b15oai012as1n04x5 U3826 (.a(n3303),
    .b(n3305),
    .c(net11),
    .o1(n3304));
 b15aoai13as1n08x5 U3827 (.a(net53),
    .b(n3304),
    .c(net11),
    .d(n3305),
    .o1(n3306));
 b15nanb02an1n02x5 U3828 (.a(net2320),
    .b(n3306),
    .out0(n1456));
 b15inv000ah1n10x5 U3829 (.a(n3307),
    .o1(n3610));
 b15inv040aq1n05x5 U3830 (.a(net361),
    .o1(n3310));
 b15norp03aq1n24x5 U3831 (.a(net344),
    .b(n3310),
    .c(n3308),
    .o1(n3309));
 b15ztpn00an1n08x5 PHY_16 ();
 b15oaoi13as1n08x5 U3834 (.a(net167),
    .b(n3310),
    .c(rd_wr_sync),
    .d(n3610),
    .o1(u_spi_device_tlul_plug_state_next[0]));
 b15inv000aq1n10x5 U3835 (.a(net2013),
    .o1(net61));
 b15inv040as1n06x5 U3836 (.a(net2111),
    .o1(n3339));
 b15aboi22as1n24x5 U3837 (.a(net2098),
    .b(n3339),
    .c(net2111),
    .d(net2098),
    .out0(n3561));
 b15inv020ah1n05x5 U3838 (.a(net2118),
    .o1(n3317));
 b15inv000aq1n16x5 U3839 (.a(net2103),
    .o1(n3318));
 b15aoi022aq1n12x5 U3840 (.a(net2103),
    .b(net2498),
    .c(n3317),
    .d(n3318),
    .o1(n3312));
 b15inv020an1n32x5 U3841 (.a(net275),
    .o1(n3595));
 b15inv020as1n16x5 U3842 (.a(net271),
    .o1(n3580));
 b15aoi022an1n48x5 U3843 (.a(net271),
    .b(net274),
    .c(n3595),
    .d(n3580),
    .o1(n3326));
 b15qgbin1an1n15x5 U3844 (.a(net2122),
    .o1(n3334));
 b15aboi22aq1n16x5 U3845 (.a(n3326),
    .b(net2512),
    .c(n3326),
    .d(n3334),
    .out0(n3311));
 b15xor002an1n12x5 U3846 (.a(n3312),
    .b(n3311),
    .out0(n3315));
 b15inv000as1n06x5 U3847 (.a(net2128),
    .o1(n3340));
 b15aoi022ah1n24x5 U3848 (.a(net339),
    .b(net2084),
    .c(n3340),
    .d(net2014),
    .o1(n3314));
 b15inv020an1n32x5 U3849 (.a(net268),
    .o1(n3322));
 b15aboi22al1n16x5 U3850 (.a(net273),
    .b(n3322),
    .c(net273),
    .d(net103),
    .out0(n3313));
 b15xor002ah1n12x5 U3851 (.a(n3314),
    .b(n3313),
    .out0(n3585));
 b15xor002ah1n06x5 U3852 (.a(n3315),
    .b(n3585),
    .out0(n3316));
 b15xor002an1n12x5 U3853 (.a(n3561),
    .b(net2513),
    .out0(net128));
 b15inv000as1n05x5 U3854 (.a(net2132),
    .o1(n3564));
 b15aoi022aq1n16x5 U3855 (.a(net2504),
    .b(net2118),
    .c(n3317),
    .d(n3564),
    .o1(n3333));
 b15inv040al1n12x5 U3856 (.a(net117),
    .o1(n3572));
 b15aoi022ah1n24x5 U3857 (.a(net2104),
    .b(net2134),
    .c(n3572),
    .d(n3318),
    .o1(n3320));
 b15inv040aq1n05x5 U3858 (.a(net2055),
    .o1(n3581));
 b15inv020as1n10x5 U3859 (.a(net2125),
    .o1(n3330));
 b15aoi022ah1n16x5 U3860 (.a(net2125),
    .b(n3581),
    .c(net2055),
    .d(n3330),
    .o1(n3319));
 b15xor002as1n12x5 U3861 (.a(n3320),
    .b(n3319),
    .out0(n3599));
 b15inv020aq1n10x5 U3862 (.a(net2114),
    .o1(n3569));
 b15aboi22aq1n24x5 U3863 (.a(net113),
    .b(net2487),
    .c(net113),
    .d(n3569),
    .out0(n3321));
 b15xor002ah1n03x5 U3864 (.a(n3599),
    .b(n3321),
    .out0(n3324));
 b15aboi22as1n08x5 U3865 (.a(net277),
    .b(n3322),
    .c(net277),
    .d(net2149),
    .out0(n3323));
 b15xor002an1n08x5 U3866 (.a(n3324),
    .b(n3323),
    .out0(n3325));
 b15xor002as1n08x5 U3867 (.a(n3333),
    .b(n3325),
    .out0(n3328));
 b15xor002ah1n16x5 U3868 (.a(net2071),
    .b(n3326),
    .out0(n3562));
 b15inv040an1n08x5 U3869 (.a(net2120),
    .o1(n3331));
 b15inv040ah1n10x5 U3870 (.a(net2036),
    .o1(n3573));
 b15aoi022ah1n32x5 U3871 (.a(net2036),
    .b(net2502),
    .c(n3331),
    .d(n3573),
    .o1(n3593));
 b15xor002as1n04x5 U3872 (.a(net2072),
    .b(n3593),
    .out0(n3327));
 b15xor002as1n06x5 U3873 (.a(n3328),
    .b(net2073),
    .out0(net66));
 b15inv020as1n32x5 U3874 (.a(net278),
    .o1(n3583));
 b15inv000aq1n32x5 U3875 (.a(net284),
    .o1(n3596));
 b15aoi022ah1n32x5 U3876 (.a(net283),
    .b(n3583),
    .c(net279),
    .d(n3596),
    .o1(n3329));
 b15xor002ah1n08x5 U3877 (.a(net277),
    .b(n3329),
    .out0(n3578));
 b15aoi022an1n12x5 U3878 (.a(net2125),
    .b(net2120),
    .c(n3331),
    .d(n3330),
    .o1(n3332));
 b15xor002aq1n02x5 U3879 (.a(n3333),
    .b(n3332),
    .out0(n3336));
 b15inv020aq1n16x5 U3880 (.a(net2159),
    .o1(n3582));
 b15aoi022as1n48x5 U3881 (.a(net2069),
    .b(net2123),
    .c(n3334),
    .d(n3582),
    .o1(n3608));
 b15xor002as1n08x5 U3882 (.a(net2106),
    .b(n3608),
    .out0(n3335));
 b15xor002aq1n03x5 U3883 (.a(n3336),
    .b(n3335),
    .out0(n3338));
 b15inv000aq1n20x5 U3884 (.a(net2048),
    .o1(n3566));
 b15aboi22as1n24x5 U3885 (.a(net290),
    .b(net288),
    .c(net290),
    .d(n3566),
    .out0(n3337));
 b15xor002an1n06x5 U3886 (.a(n3338),
    .b(n3337),
    .out0(n3342));
 b15aoi022aq1n12x5 U3887 (.a(net2111),
    .b(net2128),
    .c(n3340),
    .d(n3339),
    .o1(n3341));
 b15xor002an1n08x5 U3888 (.a(n3342),
    .b(n3341),
    .out0(n3343));
 b15xor002ar1n12x5 U3889 (.a(n3578),
    .b(net2129),
    .out0(net67));
 b15ztpn00an1n08x5 PHY_15 ();
 b15nandp3as1n24x5 U3891 (.a(n3346),
    .b(n3345),
    .c(n3344),
    .o1(n3360));
 b15inv000ah1n32x5 U3892 (.a(n3360),
    .o1(n3364));
 b15oaoi13as1n08x5 U3893 (.a(n3348),
    .b(u_dcfifo_rx_u_dout_read_token[4]),
    .c(net326),
    .d(net325),
    .o1(n3355));
 b15oaoi13as1n08x5 U3894 (.a(n3354),
    .b(u_dcfifo_rx_u_dout_read_token[4]),
    .c(net326),
    .d(net325),
    .o1(n3357));
 b15orn002ah1n24x5 U3895 (.a(n3355),
    .b(n3357),
    .o(n3350));
 b15nor002an1n32x5 U3896 (.a(n3364),
    .b(n3350),
    .o1(n3347));
 b15ztpn00an1n08x5 PHY_14 ();
 b15nandp2al1n48x5 U3899 (.a(n3357),
    .b(n3348),
    .o1(n3352));
 b15nor002aq1n32x5 U3900 (.a(n3360),
    .b(n3352),
    .o1(n3349));
 b15ztpn00an1n08x5 PHY_13 ();
 b15aoi022ah1n06x5 U3903 (.a(net155),
    .b(u_dcfifo_rx_u_din_buffer_data[232]),
    .c(net164),
    .d(u_dcfifo_rx_u_din_buffer_data[136]),
    .o1(n3369));
 b15norp02ah1n32x5 U3904 (.a(n3360),
    .b(n3350),
    .o1(n3351));
 b15norp02ar1n48x5 U3907 (.a(n3364),
    .b(n3352),
    .o1(n3353));
 b15ztpn00an1n08x5 PHY_12 ();
 b15ztpn00an1n08x5 PHY_11 ();
 b15aoi022as1n08x5 U3910 (.a(net162),
    .b(u_dcfifo_rx_u_din_buffer_data[200]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[168]),
    .o1(n3368));
 b15nandp2ah1n32x5 U3911 (.a(n3355),
    .b(n3354),
    .o1(n3361));
 b15norp02ah1n32x5 U3912 (.a(n3364),
    .b(n3361),
    .o1(n3356));
 b15ztpn00an1n08x5 PHY_10 ();
 b15nandp2an1n48x5 U3915 (.a(n3358),
    .b(n3357),
    .o1(n3363));
 b15norp02al1n48x5 U3916 (.a(n3360),
    .b(n3363),
    .o1(n3359));
 b15ztpn00an1n08x5 PHY_9 ();
 b15ztpn00an1n08x5 PHY_8 ();
 b15aoi022as1n16x5 U3919 (.a(net151),
    .b(u_dcfifo_rx_u_din_buffer_data[104]),
    .c(net160),
    .d(u_dcfifo_rx_u_din_buffer_data[8]),
    .o1(n3367));
 b15norp02aq1n48x5 U3920 (.a(n3361),
    .b(n3360),
    .o1(n3362));
 b15ztpn00an1n08x5 PHY_7 ();
 b15norp02ah1n48x5 U3923 (.a(n3364),
    .b(n3363),
    .o1(n3365));
 b15ztpn00an1n08x5 PHY_6 ();
 b15ztpn00an1n08x5 PHY_5 ();
 b15aoi022as1n16x5 U3926 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[72]),
    .c(net149),
    .d(u_dcfifo_rx_u_din_buffer_data[40]),
    .o1(n3366));
 b15nand04as1n16x5 U3927 (.a(n3369),
    .b(n3368),
    .c(n3367),
    .d(n3366),
    .o1(n3370));
 b15and002ar1n08x5 U3928 (.a(net168),
    .b(n3370),
    .o(u_spi_device_tlul_plug_wdata_next[8]));
 b15ztpn00an1n08x5 PHY_4 ();
 b15ztpn00an1n08x5 PHY_3 ();
 b15ztpn00an1n08x5 PHY_2 ();
 b15aoi022ah1n08x5 U3932 (.a(net156),
    .b(u_dcfifo_rx_u_din_buffer_data[250]),
    .c(net152),
    .d(u_dcfifo_rx_u_din_buffer_data[122]),
    .o1(n3375));
 b15ztpn00an1n08x5 PHY_1 ();
 b15ztpn00an1n08x5 PHY_0 ();
 b15aoi022ah1n06x5 U3935 (.a(net163),
    .b(u_dcfifo_rx_u_din_buffer_data[218]),
    .c(net166),
    .d(u_dcfifo_rx_u_din_buffer_data[154]),
    .o1(n3374));
 b15aoi022ah1n08x5 U3938 (.a(net161),
    .b(u_dcfifo_rx_u_din_buffer_data[26]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[186]),
    .o1(n3373));
 b15aoi022an1n24x5 U3940 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[90]),
    .c(net150),
    .d(u_dcfifo_rx_u_din_buffer_data[58]),
    .o1(n3372));
 b15nand04an1n16x5 U3941 (.a(n3375),
    .b(n3374),
    .c(n3373),
    .d(n3372),
    .o1(n3376));
 b15and002as1n16x5 U3942 (.a(net167),
    .b(net146),
    .o(u_spi_device_tlul_plug_wdata_next[26]));
 b15aoi022ah1n06x5 U3944 (.a(net160),
    .b(u_dcfifo_rx_u_din_buffer_data[4]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[164]),
    .o1(n3383));
 b15aoi022as1n16x5 U3945 (.a(net162),
    .b(u_dcfifo_rx_u_din_buffer_data[196]),
    .c(net164),
    .d(u_dcfifo_rx_u_din_buffer_data[132]),
    .o1(n3382));
 b15aoi022aq1n08x5 U3947 (.a(net155),
    .b(u_dcfifo_rx_u_din_buffer_data[228]),
    .c(net151),
    .d(u_dcfifo_rx_u_din_buffer_data[100]),
    .o1(n3381));
 b15aoi022aq1n32x5 U3949 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[68]),
    .c(net149),
    .d(u_dcfifo_rx_u_din_buffer_data[36]),
    .o1(n3380));
 b15nand04an1n16x5 U3950 (.a(n3383),
    .b(n3382),
    .c(n3381),
    .d(n3380),
    .o1(n3384));
 b15and002al1n04x5 U3951 (.a(net168),
    .b(n3384),
    .o(u_spi_device_tlul_plug_wdata_next[4]));
 b15aoi022ah1n06x5 U3952 (.a(net156),
    .b(u_dcfifo_rx_u_din_buffer_data[240]),
    .c(net164),
    .d(u_dcfifo_rx_u_din_buffer_data[144]),
    .o1(n3388));
 b15aoi022al1n32x5 U3953 (.a(net152),
    .b(u_dcfifo_rx_u_din_buffer_data[112]),
    .c(net161),
    .d(u_dcfifo_rx_u_din_buffer_data[16]),
    .o1(n3387));
 b15aoi022aq1n12x5 U3954 (.a(net163),
    .b(u_dcfifo_rx_u_din_buffer_data[208]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[176]),
    .o1(n3386));
 b15aoi022aq1n24x5 U3955 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[80]),
    .c(net149),
    .d(u_dcfifo_rx_u_din_buffer_data[48]),
    .o1(n3385));
 b15nand04as1n16x5 U3956 (.a(n3388),
    .b(n3387),
    .c(n3386),
    .d(n3385),
    .o1(n3389));
 b15and002al1n02x5 U3957 (.a(n3309),
    .b(n3389),
    .o(u_spi_device_tlul_plug_wdata_next[16]));
 b15aoi022ah1n06x5 U3959 (.a(net150),
    .b(u_dcfifo_rx_u_din_buffer_data[62]),
    .c(net152),
    .d(u_dcfifo_rx_u_din_buffer_data[126]),
    .o1(n3393));
 b15aoi022an1n08x5 U3960 (.a(net163),
    .b(u_dcfifo_rx_u_din_buffer_data[222]),
    .c(net161),
    .d(u_dcfifo_rx_u_din_buffer_data[30]),
    .o1(n3392));
 b15aoi022aq1n12x5 U3961 (.a(net156),
    .b(u_dcfifo_rx_u_din_buffer_data[254]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[190]),
    .o1(n3391));
 b15aoi022as1n08x5 U3962 (.a(net159),
    .b(net337),
    .c(net166),
    .d(u_dcfifo_rx_u_din_buffer_data[158]),
    .o1(n3390));
 b15nand04as1n16x5 U3963 (.a(n3393),
    .b(n3392),
    .c(n3391),
    .d(n3390),
    .o1(n3394));
 b15and002ar1n02x5 U3964 (.a(net167),
    .b(n3394),
    .o(u_spi_device_tlul_plug_wdata_next[30]));
 b15aoi022al1n12x5 U3966 (.a(n3349),
    .b(u_dcfifo_rx_u_din_buffer_data[157]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[189]),
    .o1(n3401));
 b15aoi022ar1n32x5 U3968 (.a(net150),
    .b(u_dcfifo_rx_u_din_buffer_data[61]),
    .c(net163),
    .d(u_dcfifo_rx_u_din_buffer_data[221]),
    .o1(n3400));
 b15aoi022aq1n08x5 U3969 (.a(net156),
    .b(u_dcfifo_rx_u_din_buffer_data[253]),
    .c(net152),
    .d(u_dcfifo_rx_u_din_buffer_data[125]),
    .o1(n3399));
 b15aoi022as1n06x5 U3971 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[93]),
    .c(net161),
    .d(u_dcfifo_rx_u_din_buffer_data[29]),
    .o1(n3398));
 b15nand04as1n16x5 U3972 (.a(n3401),
    .b(n3400),
    .c(n3399),
    .d(n3398),
    .o1(n3402));
 b15and002ar1n02x5 U3973 (.a(net167),
    .b(n3402),
    .o(u_spi_device_tlul_plug_wdata_next[29]));
 b15aoi022ar1n32x5 U3974 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[95]),
    .c(n3365),
    .d(u_dcfifo_rx_u_din_buffer_data[63]),
    .o1(n3407));
 b15aoi022ar1n16x5 U3976 (.a(net163),
    .b(u_dcfifo_rx_u_din_buffer_data[223]),
    .c(net156),
    .d(u_dcfifo_rx_u_din_buffer_data[255]),
    .o1(n3406));
 b15aoi022aq1n32x5 U3977 (.a(net152),
    .b(u_dcfifo_rx_u_din_buffer_data[127]),
    .c(net165),
    .d(u_dcfifo_rx_u_din_buffer_data[159]),
    .o1(n3405));
 b15aoi022aq1n12x5 U3978 (.a(net161),
    .b(u_dcfifo_rx_u_din_buffer_data[31]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[191]),
    .o1(n3404));
 b15nand04as1n16x5 U3979 (.a(n3407),
    .b(n3406),
    .c(n3405),
    .d(n3404),
    .o1(n3408));
 b15and002al1n02x5 U3980 (.a(net168),
    .b(n3408),
    .o(u_spi_device_tlul_plug_wdata_next[31]));
 b15aoi022ah1n08x5 U3981 (.a(net161),
    .b(u_dcfifo_rx_u_din_buffer_data[17]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[177]),
    .o1(n3412));
 b15aoi022an1n32x5 U3982 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[81]),
    .c(net150),
    .d(u_dcfifo_rx_u_din_buffer_data[49]),
    .o1(n3411));
 b15aoi022ah1n08x5 U3983 (.a(net163),
    .b(u_dcfifo_rx_u_din_buffer_data[209]),
    .c(net165),
    .d(u_dcfifo_rx_u_din_buffer_data[145]),
    .o1(n3410));
 b15aoi022ah1n08x5 U3984 (.a(net156),
    .b(u_dcfifo_rx_u_din_buffer_data[241]),
    .c(net152),
    .d(u_dcfifo_rx_u_din_buffer_data[113]),
    .o1(n3409));
 b15nand04as1n16x5 U3985 (.a(n3412),
    .b(n3411),
    .c(n3410),
    .d(n3409),
    .o1(n3413));
 b15and002an1n03x5 U3986 (.a(n3309),
    .b(n3413),
    .o(u_spi_device_tlul_plug_wdata_next[17]));
 b15aoi022ah1n06x5 U3987 (.a(net156),
    .b(u_dcfifo_rx_u_din_buffer_data[242]),
    .c(net161),
    .d(u_dcfifo_rx_u_din_buffer_data[18]),
    .o1(n3418));
 b15aoi022ar1n16x5 U3988 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[82]),
    .c(net166),
    .d(u_dcfifo_rx_u_din_buffer_data[146]),
    .o1(n3417));
 b15aoi022al1n16x5 U3989 (.a(net163),
    .b(u_dcfifo_rx_u_din_buffer_data[210]),
    .c(net152),
    .d(u_dcfifo_rx_u_din_buffer_data[114]),
    .o1(n3416));
 b15aoi022an1n08x5 U3991 (.a(net150),
    .b(u_dcfifo_rx_u_din_buffer_data[50]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[178]),
    .o1(n3415));
 b15nand04as1n16x5 U3992 (.a(n3418),
    .b(n3417),
    .c(n3416),
    .d(n3415),
    .o1(n3419));
 b15and002ar1n02x5 U3993 (.a(net168),
    .b(n3419),
    .o(u_spi_device_tlul_plug_wdata_next[18]));
 b15aoi022ah1n12x5 U3994 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[86]),
    .c(net163),
    .d(u_dcfifo_rx_u_din_buffer_data[214]),
    .o1(n3423));
 b15aoi022an1n08x5 U3995 (.a(net150),
    .b(u_dcfifo_rx_u_din_buffer_data[54]),
    .c(net166),
    .d(u_dcfifo_rx_u_din_buffer_data[150]),
    .o1(n3422));
 b15aoi022an1n48x5 U3996 (.a(net152),
    .b(u_dcfifo_rx_u_din_buffer_data[118]),
    .c(net161),
    .d(u_dcfifo_rx_u_din_buffer_data[22]),
    .o1(n3421));
 b15aoi022an1n08x5 U3997 (.a(net156),
    .b(u_dcfifo_rx_u_din_buffer_data[246]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[182]),
    .o1(n3420));
 b15nand04as1n16x5 U3998 (.a(n3423),
    .b(n3422),
    .c(n3421),
    .d(n3420),
    .o1(n3424));
 b15and002al1n02x5 U3999 (.a(net168),
    .b(n3424),
    .o(u_spi_device_tlul_plug_wdata_next[22]));
 b15aoi022ar1n32x5 U4000 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[76]),
    .c(net162),
    .d(u_dcfifo_rx_u_din_buffer_data[204]),
    .o1(n3428));
 b15aoi022al1n32x5 U4001 (.a(net164),
    .b(u_dcfifo_rx_u_din_buffer_data[140]),
    .c(net160),
    .d(u_dcfifo_rx_u_din_buffer_data[12]),
    .o1(n3427));
 b15aoi022as1n06x5 U4002 (.a(net155),
    .b(u_dcfifo_rx_u_din_buffer_data[236]),
    .c(net151),
    .d(u_dcfifo_rx_u_din_buffer_data[108]),
    .o1(n3426));
 b15aoi022ar1n12x5 U4003 (.a(net149),
    .b(net338),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[172]),
    .o1(n3425));
 b15nand04as1n16x5 U4004 (.a(n3428),
    .b(n3427),
    .c(n3426),
    .d(n3425),
    .o1(n3429));
 b15and002al1n04x5 U4005 (.a(net167),
    .b(n3429),
    .o(u_spi_device_tlul_plug_wdata_next[12]));
 b15aoi022ar1n32x5 U4006 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[84]),
    .c(net150),
    .d(u_dcfifo_rx_u_din_buffer_data[52]),
    .o1(n3433));
 b15aoi022an1n02x5 U4007 (.a(net156),
    .b(u_dcfifo_rx_u_din_buffer_data[244]),
    .c(net166),
    .d(u_dcfifo_rx_u_din_buffer_data[148]),
    .o1(n3432));
 b15aoi022as1n12x5 U4008 (.a(net163),
    .b(u_dcfifo_rx_u_din_buffer_data[212]),
    .c(net161),
    .d(u_dcfifo_rx_u_din_buffer_data[20]),
    .o1(n3431));
 b15aoi022ah1n08x5 U4009 (.a(net152),
    .b(u_dcfifo_rx_u_din_buffer_data[116]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[180]),
    .o1(n3430));
 b15nand04as1n08x5 U4010 (.a(n3433),
    .b(n3432),
    .c(n3431),
    .d(n3430),
    .o1(n3434));
 b15and002ar1n02x5 U4011 (.a(net167),
    .b(net145),
    .o(u_spi_device_tlul_plug_wdata_next[20]));
 b15aoi022aq1n12x5 U4012 (.a(net151),
    .b(u_dcfifo_rx_u_din_buffer_data[97]),
    .c(net164),
    .d(u_dcfifo_rx_u_din_buffer_data[129]),
    .o1(n3438));
 b15aoi022al1n16x5 U4013 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[65]),
    .c(net162),
    .d(u_dcfifo_rx_u_din_buffer_data[193]),
    .o1(n3437));
 b15aoi022ah1n08x5 U4014 (.a(net155),
    .b(u_dcfifo_rx_u_din_buffer_data[225]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[161]),
    .o1(n3436));
 b15aoi022aq1n12x5 U4015 (.a(net149),
    .b(u_dcfifo_rx_u_din_buffer_data[33]),
    .c(net160),
    .d(u_dcfifo_rx_u_din_buffer_data[1]),
    .o1(n3435));
 b15nand04as1n16x5 U4016 (.a(n3438),
    .b(n3437),
    .c(n3436),
    .d(n3435),
    .o1(n3439));
 b15and002as1n02x5 U4017 (.a(net167),
    .b(n3439),
    .o(u_spi_device_tlul_plug_wdata_next[1]));
 b15aoi022as1n08x5 U4018 (.a(net165),
    .b(u_dcfifo_rx_u_din_buffer_data[137]),
    .c(net160),
    .d(u_dcfifo_rx_u_din_buffer_data[9]),
    .o1(n3443));
 b15aoi022ar1n24x5 U4019 (.a(net150),
    .b(u_dcfifo_rx_u_din_buffer_data[41]),
    .c(net155),
    .d(u_dcfifo_rx_u_din_buffer_data[233]),
    .o1(n3442));
 b15aoi022as1n06x5 U4020 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[73]),
    .c(net151),
    .d(u_dcfifo_rx_u_din_buffer_data[105]),
    .o1(n3441));
 b15aoi022an1n12x5 U4021 (.a(net162),
    .b(u_dcfifo_rx_u_din_buffer_data[201]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[169]),
    .o1(n3440));
 b15nand04as1n16x5 U4022 (.a(n3443),
    .b(n3442),
    .c(n3441),
    .d(n3440),
    .o1(n3444));
 b15and002al1n02x5 U4023 (.a(net167),
    .b(n3444),
    .o(u_spi_device_tlul_plug_wdata_next[9]));
 b15aoi022aq1n12x5 U4024 (.a(net149),
    .b(u_dcfifo_rx_u_din_buffer_data[38]),
    .c(net160),
    .d(u_dcfifo_rx_u_din_buffer_data[6]),
    .o1(n3448));
 b15aoi022ah1n08x5 U4025 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[70]),
    .c(net164),
    .d(u_dcfifo_rx_u_din_buffer_data[134]),
    .o1(n3447));
 b15aoi022ah1n12x5 U4026 (.a(net162),
    .b(u_dcfifo_rx_u_din_buffer_data[198]),
    .c(net155),
    .d(u_dcfifo_rx_u_din_buffer_data[230]),
    .o1(n3446));
 b15aoi022ah1n08x5 U4027 (.a(net151),
    .b(u_dcfifo_rx_u_din_buffer_data[102]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[166]),
    .o1(n3445));
 b15nand04as1n16x5 U4028 (.a(n3448),
    .b(n3447),
    .c(n3446),
    .d(n3445),
    .o1(n3449));
 b15and002an1n24x5 U4029 (.a(net168),
    .b(n3449),
    .o(u_spi_device_tlul_plug_wdata_next[6]));
 b15aoi022ah1n12x5 U4030 (.a(net162),
    .b(u_dcfifo_rx_u_din_buffer_data[197]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[165]),
    .o1(n3453));
 b15aoi022ar1n16x5 U4031 (.a(net149),
    .b(u_dcfifo_rx_u_din_buffer_data[37]),
    .c(net151),
    .d(u_dcfifo_rx_u_din_buffer_data[101]),
    .o1(n3452));
 b15aoi022aq1n16x5 U4032 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[69]),
    .c(net155),
    .d(u_dcfifo_rx_u_din_buffer_data[229]),
    .o1(n3451));
 b15aoi022an1n04x5 U4033 (.a(net164),
    .b(u_dcfifo_rx_u_din_buffer_data[133]),
    .c(net160),
    .d(u_dcfifo_rx_u_din_buffer_data[5]),
    .o1(n3450));
 b15nand04as1n06x5 U4034 (.a(n3453),
    .b(n3452),
    .c(n3451),
    .d(n3450),
    .o1(n3454));
 b15and002ar1n04x5 U4035 (.a(net168),
    .b(n3454),
    .o(u_spi_device_tlul_plug_wdata_next[5]));
 b15aoi022ah1n08x5 U4036 (.a(net150),
    .b(u_dcfifo_rx_u_din_buffer_data[55]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[183]),
    .o1(n3458));
 b15aoi022aq1n16x5 U4037 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[87]),
    .c(net156),
    .d(u_dcfifo_rx_u_din_buffer_data[247]),
    .o1(n3457));
 b15aoi022an1n16x5 U4038 (.a(net163),
    .b(u_dcfifo_rx_u_din_buffer_data[215]),
    .c(net161),
    .d(u_dcfifo_rx_u_din_buffer_data[23]),
    .o1(n3456));
 b15aoi022aq1n16x5 U4039 (.a(net152),
    .b(u_dcfifo_rx_u_din_buffer_data[119]),
    .c(net166),
    .d(u_dcfifo_rx_u_din_buffer_data[151]),
    .o1(n3455));
 b15nand04as1n16x5 U4040 (.a(n3458),
    .b(n3457),
    .c(n3456),
    .d(n3455),
    .o1(n3459));
 b15and002an1n03x5 U4041 (.a(net168),
    .b(n3459),
    .o(u_spi_device_tlul_plug_wdata_next[23]));
 b15aoi022al1n24x5 U4042 (.a(net166),
    .b(u_dcfifo_rx_u_din_buffer_data[153]),
    .c(net161),
    .d(u_dcfifo_rx_u_din_buffer_data[25]),
    .o1(n3463));
 b15aoi022an1n16x5 U4043 (.a(net163),
    .b(u_dcfifo_rx_u_din_buffer_data[217]),
    .c(net156),
    .d(u_dcfifo_rx_u_din_buffer_data[249]),
    .o1(n3462));
 b15aoi022an1n16x5 U4044 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[89]),
    .c(net152),
    .d(u_dcfifo_rx_u_din_buffer_data[121]),
    .o1(n3461));
 b15aoi022al1n12x5 U4045 (.a(net150),
    .b(u_dcfifo_rx_u_din_buffer_data[57]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[185]),
    .o1(n3460));
 b15nand04as1n16x5 U4046 (.a(n3463),
    .b(n3462),
    .c(n3461),
    .d(n3460),
    .o1(n3464));
 b15and002aq1n16x5 U4047 (.a(net167),
    .b(net144),
    .o(u_spi_device_tlul_plug_wdata_next[25]));
 b15aoi022aq1n08x5 U4048 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[71]),
    .c(net164),
    .d(u_dcfifo_rx_u_din_buffer_data[135]),
    .o1(n3468));
 b15aoi022al1n12x5 U4049 (.a(net155),
    .b(u_dcfifo_rx_u_din_buffer_data[231]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[167]),
    .o1(n3467));
 b15aoi022ah1n24x5 U4050 (.a(net149),
    .b(u_dcfifo_rx_u_din_buffer_data[39]),
    .c(net162),
    .d(u_dcfifo_rx_u_din_buffer_data[199]),
    .o1(n3466));
 b15aoi022ah1n24x5 U4051 (.a(net151),
    .b(u_dcfifo_rx_u_din_buffer_data[103]),
    .c(net160),
    .d(u_dcfifo_rx_u_din_buffer_data[7]),
    .o1(n3465));
 b15nand04as1n16x5 U4052 (.a(n3468),
    .b(n3467),
    .c(n3466),
    .d(n3465),
    .o1(n3469));
 b15and002ah1n04x5 U4053 (.a(net168),
    .b(n3469),
    .o(u_spi_device_tlul_plug_wdata_next[7]));
 b15aoi022as1n06x5 U4054 (.a(net151),
    .b(u_dcfifo_rx_u_din_buffer_data[111]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[175]),
    .o1(n3474));
 b15aoi022aq1n16x5 U4055 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[79]),
    .c(net149),
    .d(u_dcfifo_rx_u_din_buffer_data[47]),
    .o1(n3473));
 b15aoi022as1n06x5 U4056 (.a(net155),
    .b(u_dcfifo_rx_u_din_buffer_data[239]),
    .c(net160),
    .d(u_dcfifo_rx_u_din_buffer_data[15]),
    .o1(n3472));
 b15aoi022ar1n12x5 U4057 (.a(net162),
    .b(u_dcfifo_rx_u_din_buffer_data[207]),
    .c(net164),
    .d(u_dcfifo_rx_u_din_buffer_data[143]),
    .o1(n3471));
 b15nand04as1n16x5 U4058 (.a(n3474),
    .b(n3473),
    .c(n3472),
    .d(n3471),
    .o1(n3475));
 b15and002al1n02x5 U4059 (.a(net167),
    .b(n3475),
    .o(u_spi_device_tlul_plug_wdata_next[15]));
 b15aoi022as1n08x5 U4060 (.a(net150),
    .b(u_dcfifo_rx_u_din_buffer_data[53]),
    .c(net161),
    .d(u_dcfifo_rx_u_din_buffer_data[21]),
    .o1(n3480));
 b15aoi022aq1n12x5 U4061 (.a(net156),
    .b(u_dcfifo_rx_u_din_buffer_data[245]),
    .c(net166),
    .d(u_dcfifo_rx_u_din_buffer_data[149]),
    .o1(n3479));
 b15aoi022al1n32x5 U4062 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[85]),
    .c(net163),
    .d(u_dcfifo_rx_u_din_buffer_data[213]),
    .o1(n3478));
 b15aoi022aq1n08x5 U4063 (.a(net152),
    .b(u_dcfifo_rx_u_din_buffer_data[117]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[181]),
    .o1(n3477));
 b15nand04as1n16x5 U4064 (.a(n3480),
    .b(n3479),
    .c(n3478),
    .d(n3477),
    .o1(n3481));
 b15and002ar1n02x5 U4065 (.a(net168),
    .b(n3481),
    .o(u_spi_device_tlul_plug_wdata_next[21]));
 b15aoi022ah1n12x5 U4066 (.a(net151),
    .b(u_dcfifo_rx_u_din_buffer_data[110]),
    .c(net164),
    .d(u_dcfifo_rx_u_din_buffer_data[142]),
    .o1(n3485));
 b15aoi022ar1n16x5 U4067 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[78]),
    .c(net162),
    .d(u_dcfifo_rx_u_din_buffer_data[206]),
    .o1(n3484));
 b15aoi022aq1n12x5 U4068 (.a(net149),
    .b(u_dcfifo_rx_u_din_buffer_data[46]),
    .c(net160),
    .d(u_dcfifo_rx_u_din_buffer_data[14]),
    .o1(n3483));
 b15aoi022al1n12x5 U4069 (.a(net155),
    .b(u_dcfifo_rx_u_din_buffer_data[238]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[174]),
    .o1(n3482));
 b15nand04as1n16x5 U4070 (.a(n3485),
    .b(n3484),
    .c(n3483),
    .d(n3482),
    .o1(n3486));
 b15and002ah1n03x5 U4071 (.a(net168),
    .b(n3486),
    .o(u_spi_device_tlul_plug_wdata_next[14]));
 b15aoi022al1n16x5 U4072 (.a(net151),
    .b(u_dcfifo_rx_u_din_buffer_data[109]),
    .c(net160),
    .d(u_dcfifo_rx_u_din_buffer_data[13]),
    .o1(n3490));
 b15aoi022ah1n12x5 U4073 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[77]),
    .c(net162),
    .d(u_dcfifo_rx_u_din_buffer_data[205]),
    .o1(n3489));
 b15aoi022ar1n24x5 U4074 (.a(net149),
    .b(u_dcfifo_rx_u_din_buffer_data[45]),
    .c(net164),
    .d(u_dcfifo_rx_u_din_buffer_data[141]),
    .o1(n3488));
 b15aoi022aq1n08x5 U4075 (.a(net155),
    .b(u_dcfifo_rx_u_din_buffer_data[237]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[173]),
    .o1(n3487));
 b15nand04as1n16x5 U4076 (.a(n3490),
    .b(n3489),
    .c(n3488),
    .d(n3487),
    .o1(n3491));
 b15and002an1n04x5 U4077 (.a(net168),
    .b(n3491),
    .o(u_spi_device_tlul_plug_wdata_next[13]));
 b15aoi022as1n04x5 U4078 (.a(net160),
    .b(u_dcfifo_rx_u_din_buffer_data[2]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[162]),
    .o1(n3495));
 b15aoi022al1n16x5 U4079 (.a(net149),
    .b(u_dcfifo_rx_u_din_buffer_data[34]),
    .c(net162),
    .d(u_dcfifo_rx_u_din_buffer_data[194]),
    .o1(n3494));
 b15aoi022an1n08x5 U4080 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[66]),
    .c(net151),
    .d(u_dcfifo_rx_u_din_buffer_data[98]),
    .o1(n3493));
 b15aoi022ar1n16x5 U4081 (.a(net155),
    .b(u_dcfifo_rx_u_din_buffer_data[226]),
    .c(net164),
    .d(u_dcfifo_rx_u_din_buffer_data[130]),
    .o1(n3492));
 b15nand04as1n16x5 U4082 (.a(n3495),
    .b(n3494),
    .c(n3493),
    .d(n3492),
    .o1(n3496));
 b15and002an1n02x5 U4083 (.a(net167),
    .b(n3496),
    .o(u_spi_device_tlul_plug_wdata_next[2]));
 b15aoi022ar1n24x5 U4084 (.a(net152),
    .b(u_dcfifo_rx_u_din_buffer_data[124]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[188]),
    .o1(n3500));
 b15aoi022al1n24x5 U4085 (.a(net166),
    .b(u_dcfifo_rx_u_din_buffer_data[156]),
    .c(net161),
    .d(u_dcfifo_rx_u_din_buffer_data[28]),
    .o1(n3499));
 b15aoi022al1n16x5 U4086 (.a(net150),
    .b(u_dcfifo_rx_u_din_buffer_data[60]),
    .c(net163),
    .d(u_dcfifo_rx_u_din_buffer_data[220]),
    .o1(n3498));
 b15aoi022ar1n24x5 U4087 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[92]),
    .c(net156),
    .d(u_dcfifo_rx_u_din_buffer_data[252]),
    .o1(n3497));
 b15nand04as1n16x5 U4088 (.a(n3500),
    .b(n3499),
    .c(n3498),
    .d(n3497),
    .o1(n3501));
 b15and002ar1n02x5 U4089 (.a(net168),
    .b(n3501),
    .o(u_spi_device_tlul_plug_wdata_next[28]));
 b15aoi022ar1n16x5 U4090 (.a(net149),
    .b(u_dcfifo_rx_u_din_buffer_data[35]),
    .c(net151),
    .d(u_dcfifo_rx_u_din_buffer_data[99]),
    .o1(n3506));
 b15aoi022an1n08x5 U4091 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[67]),
    .c(net160),
    .d(u_dcfifo_rx_u_din_buffer_data[3]),
    .o1(n3505));
 b15aoi022ar1n12x5 U4092 (.a(net164),
    .b(u_dcfifo_rx_u_din_buffer_data[131]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[163]),
    .o1(n3504));
 b15aoi022al1n16x5 U4093 (.a(net162),
    .b(u_dcfifo_rx_u_din_buffer_data[195]),
    .c(net155),
    .d(u_dcfifo_rx_u_din_buffer_data[227]),
    .o1(n3503));
 b15nand04as1n16x5 U4094 (.a(n3506),
    .b(n3505),
    .c(n3504),
    .d(n3503),
    .o1(n3507));
 b15and002ar1n02x5 U4095 (.a(net167),
    .b(n3507),
    .o(u_spi_device_tlul_plug_wdata_next[3]));
 b15aoi022an1n32x5 U4096 (.a(net166),
    .b(u_dcfifo_rx_u_din_buffer_data[155]),
    .c(net161),
    .d(u_dcfifo_rx_u_din_buffer_data[27]),
    .o1(n3513));
 b15aoi022as1n06x5 U4097 (.a(net156),
    .b(u_dcfifo_rx_u_din_buffer_data[251]),
    .c(net152),
    .d(u_dcfifo_rx_u_din_buffer_data[123]),
    .o1(n3512));
 b15aoi022as1n08x5 U4098 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[91]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[187]),
    .o1(n3511));
 b15aoi022as1n06x5 U4099 (.a(net150),
    .b(u_dcfifo_rx_u_din_buffer_data[59]),
    .c(net163),
    .d(u_dcfifo_rx_u_din_buffer_data[219]),
    .o1(n3510));
 b15nand04as1n16x5 U4100 (.a(n3513),
    .b(n3512),
    .c(n3511),
    .d(n3510),
    .o1(n3514));
 b15and002ar1n02x5 U4101 (.a(net168),
    .b(n3514),
    .o(u_spi_device_tlul_plug_wdata_next[27]));
 b15aoi022an1n12x5 U4102 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[75]),
    .c(net164),
    .d(u_dcfifo_rx_u_din_buffer_data[139]),
    .o1(n3520));
 b15aoi022an1n08x5 U4103 (.a(net160),
    .b(u_dcfifo_rx_u_din_buffer_data[11]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[171]),
    .o1(n3519));
 b15aoi022aq1n32x5 U4104 (.a(net149),
    .b(u_dcfifo_rx_u_din_buffer_data[43]),
    .c(net162),
    .d(u_dcfifo_rx_u_din_buffer_data[203]),
    .o1(n3518));
 b15aoi022aq1n08x5 U4105 (.a(net155),
    .b(u_dcfifo_rx_u_din_buffer_data[235]),
    .c(net151),
    .d(u_dcfifo_rx_u_din_buffer_data[107]),
    .o1(n3517));
 b15nand04as1n16x5 U4106 (.a(n3520),
    .b(n3519),
    .c(n3518),
    .d(n3517),
    .o1(n3521));
 b15and002an1n03x5 U4107 (.a(net167),
    .b(n3521),
    .o(u_spi_device_tlul_plug_wdata_next[11]));
 b15aoi022al1n24x5 U4108 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[64]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[160]),
    .o1(n3528));
 b15aoi022aq1n24x5 U4109 (.a(net151),
    .b(u_dcfifo_rx_u_din_buffer_data[96]),
    .c(net160),
    .d(u_dcfifo_rx_u_din_buffer_data[0]),
    .o1(n3527));
 b15aoi022as1n08x5 U4110 (.a(net155),
    .b(u_dcfifo_rx_u_din_buffer_data[224]),
    .c(net164),
    .d(u_dcfifo_rx_u_din_buffer_data[128]),
    .o1(n3526));
 b15aoi022aq1n12x5 U4111 (.a(net149),
    .b(u_dcfifo_rx_u_din_buffer_data[32]),
    .c(net162),
    .d(u_dcfifo_rx_u_din_buffer_data[192]),
    .o1(n3525));
 b15nand04as1n16x5 U4112 (.a(n3528),
    .b(n3527),
    .c(n3526),
    .d(n3525),
    .o1(n3529));
 b15and002ar1n12x5 U4113 (.a(n3309),
    .b(n3529),
    .o(u_spi_device_tlul_plug_wdata_next[0]));
 b15aoi022ar1n16x5 U4114 (.a(net152),
    .b(u_dcfifo_rx_u_din_buffer_data[115]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[179]),
    .o1(n3535));
 b15aoi022as1n08x5 U4115 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[83]),
    .c(net156),
    .d(u_dcfifo_rx_u_din_buffer_data[243]),
    .o1(n3534));
 b15aoi022ar1n32x5 U4116 (.a(net166),
    .b(u_dcfifo_rx_u_din_buffer_data[147]),
    .c(net161),
    .d(u_dcfifo_rx_u_din_buffer_data[19]),
    .o1(n3533));
 b15aoi022ar1n16x5 U4117 (.a(net150),
    .b(u_dcfifo_rx_u_din_buffer_data[51]),
    .c(net163),
    .d(u_dcfifo_rx_u_din_buffer_data[211]),
    .o1(n3532));
 b15nand04an1n12x5 U4118 (.a(n3535),
    .b(n3534),
    .c(n3533),
    .d(n3532),
    .o1(n3536));
 b15and002ar1n02x5 U4119 (.a(net167),
    .b(net143),
    .o(u_spi_device_tlul_plug_wdata_next[19]));
 b15aoi022aq1n16x5 U4120 (.a(net150),
    .b(u_dcfifo_rx_u_din_buffer_data[56]),
    .c(net152),
    .d(u_dcfifo_rx_u_din_buffer_data[120]),
    .o1(n3545));
 b15aoi022as1n06x5 U4121 (.a(net156),
    .b(u_dcfifo_rx_u_din_buffer_data[248]),
    .c(net154),
    .d(u_dcfifo_rx_u_din_buffer_data[184]),
    .o1(n3544));
 b15aoi022ar1n48x5 U4122 (.a(net166),
    .b(u_dcfifo_rx_u_din_buffer_data[152]),
    .c(net161),
    .d(u_dcfifo_rx_u_din_buffer_data[24]),
    .o1(n3543));
 b15aoi022al1n16x5 U4123 (.a(net159),
    .b(u_dcfifo_rx_u_din_buffer_data[88]),
    .c(net163),
    .d(u_dcfifo_rx_u_din_buffer_data[216]),
    .o1(n3542));
 b15nand04as1n16x5 U4124 (.a(n3545),
    .b(n3544),
    .c(n3543),
    .d(n3542),
    .o1(n3546));
 b15and002an1n24x5 U4125 (.a(net167),
    .b(n3546),
    .o(u_spi_device_tlul_plug_wdata_next[24]));
 b15aoi022as1n08x5 U4126 (.a(net149),
    .b(u_dcfifo_rx_u_din_buffer_data[42]),
    .c(net153),
    .d(u_dcfifo_rx_u_din_buffer_data[170]),
    .o1(n3559));
 b15aoi022as1n16x5 U4127 (.a(net164),
    .b(u_dcfifo_rx_u_din_buffer_data[138]),
    .c(net160),
    .d(u_dcfifo_rx_u_din_buffer_data[10]),
    .o1(n3558));
 b15aoi022as1n06x5 U4128 (.a(net155),
    .b(u_dcfifo_rx_u_din_buffer_data[234]),
    .c(net151),
    .d(u_dcfifo_rx_u_din_buffer_data[106]),
    .o1(n3557));
 b15aoi022ar1n24x5 U4129 (.a(net158),
    .b(u_dcfifo_rx_u_din_buffer_data[74]),
    .c(net162),
    .d(u_dcfifo_rx_u_din_buffer_data[202]),
    .o1(n3556));
 b15nand04as1n16x5 U4130 (.a(n3559),
    .b(n3558),
    .c(n3557),
    .d(n3556),
    .o1(n3560));
 b15and002aq1n02x5 U4131 (.a(net167),
    .b(n3560),
    .o(u_spi_device_tlul_plug_wdata_next[10]));
 b15xor002ah1n16x5 U4132 (.a(n3561),
    .b(net267),
    .out0(n3601));
 b15xor002as1n08x5 U4133 (.a(net291),
    .b(n3601),
    .out0(n3563));
 b15xor002an1n12x5 U4134 (.a(n3563),
    .b(net2072),
    .out0(n3575));
 b15inv020ar1n32x5 U4135 (.a(net265),
    .o1(n3571));
 b15aoi022an1n12x5 U4136 (.a(net2132),
    .b(net265),
    .c(n3571),
    .d(n3564),
    .o1(n3565));
 b15xor002as1n06x5 U4137 (.a(n3575),
    .b(n3565),
    .out0(n3568));
 b15inv040as1n08x5 U4138 (.a(net110),
    .o1(n3597));
 b15aoi022ar1n24x5 U4139 (.a(net2049),
    .b(net110),
    .c(n3597),
    .d(n3566),
    .o1(n3567));
 b15xor002as1n16x5 U4140 (.a(net2116),
    .b(n3567),
    .out0(n3586));
 b15xor002aq1n06x5 U4141 (.a(n3568),
    .b(n3586),
    .out0(n3570));
 b15aboi22as1n24x5 U4142 (.a(net2137),
    .b(net2114),
    .c(net2137),
    .d(n3569),
    .out0(n3605));
 b15xor002as1n08x5 U4143 (.a(n3570),
    .b(net2138),
    .out0(net132));
 b15inv040as1n12x5 U4144 (.a(net2059),
    .o1(n3598));
 b15aoi022an1n48x5 U4145 (.a(net2044),
    .b(net2060),
    .c(n3598),
    .d(n3571),
    .o1(n3590));
 b15xor002as1n04x5 U4146 (.a(net2061),
    .b(net339),
    .out0(n3577));
 b15aoi022al1n32x5 U4147 (.a(net117),
    .b(net2037),
    .c(n3573),
    .d(n3572),
    .o1(n3574));
 b15xor002as1n03x5 U4148 (.a(n3575),
    .b(n3574),
    .out0(n3576));
 b15xor002as1n06x5 U4149 (.a(net2062),
    .b(n3576),
    .out0(n3579));
 b15xor002an1n08x5 U4150 (.a(net2063),
    .b(n3578),
    .out0(net63));
 b15aoi022an1n16x5 U4151 (.a(net2029),
    .b(net2055),
    .c(n3581),
    .d(n3580),
    .o1(n3589));
 b15aoi022ar1n24x5 U4152 (.a(net2068),
    .b(net2021),
    .c(n3583),
    .d(n3582),
    .o1(n3584));
 b15xor002as1n02x5 U4153 (.a(n3585),
    .b(n3584),
    .out0(n3587));
 b15xor002al1n04x5 U4154 (.a(n3587),
    .b(n3586),
    .out0(n3588));
 b15xor002aq1n04x5 U4155 (.a(n3589),
    .b(n3588),
    .out0(n3591));
 b15xor002as1n06x5 U4156 (.a(n3591),
    .b(net2061),
    .out0(n3592));
 b15xor002an1n16x5 U4157 (.a(n3593),
    .b(n3592),
    .out0(n3594));
 b15xor002an1n06x5 U4158 (.a(n3594),
    .b(net2094),
    .out0(net65));
 b15aoi022aq1n16x5 U4159 (.a(net275),
    .b(n3596),
    .c(net284),
    .d(n3595),
    .o1(n3604));
 b15aoi022ar1n48x5 U4160 (.a(net2147),
    .b(net286),
    .c(n3598),
    .d(n3597),
    .o1(n3600));
 b15xor002an1n12x5 U4161 (.a(n3600),
    .b(n3599),
    .out0(n3602));
 b15xor002ar1n12x5 U4162 (.a(n3602),
    .b(n3601),
    .out0(n3603));
 b15xor002ar1n08x5 U4163 (.a(n3604),
    .b(n3603),
    .out0(n3606));
 b15xor002an1n08x5 U4164 (.a(n3606),
    .b(net2138),
    .out0(n3607));
 b15xor002as1n06x5 U4165 (.a(net273),
    .b(n3607),
    .out0(n3609));
 b15xor002as1n16x5 U4166 (.a(n3609),
    .b(net2160),
    .out0(net64));
 b15nor002al1n32x5 U4167 (.a(net361),
    .b(n3610),
    .o1(u_spi_device_tlul_plug_N61));
 b15and003ar1n08x5 U4168 (.a(n3612),
    .b(n3611),
    .c(u_device_sm_s_dummy_cycles[6]),
    .o(u_rxreg_counter_trgt_next[6]));
 b15and003an1n08x5 U4169 (.a(n3612),
    .b(n3611),
    .c(u_device_sm_s_dummy_cycles[7]),
    .o(u_rxreg_counter_trgt_next[7]));
 b15inv000al1n03x5 U4170 (.a(u_rxreg_N7),
    .o1(n3615));
 b15oai012ar1n06x5 U4171 (.a(n3612),
    .b(u_device_sm_s_dummy_cycles[0]),
    .c(n3613),
    .o1(n3614));
 b15aoai13as1n08x5 U4172 (.a(n3614),
    .b(n3615),
    .c(n3616),
    .d(n3626),
    .o1(u_rxreg_counter_trgt_next[0]));
 b15nonb02al1n03x5 U4174 (.a(u_device_sm_tx_done_reg),
    .b(n3617),
    .out0(n3623));
 b15oaoi13an1n04x5 U4175 (.a(n3618),
    .b(u_device_sm_state[2]),
    .c(n3620),
    .d(n3619),
    .o1(n3621));
 b15aoai13al1n02x5 U4176 (.a(n3621),
    .b(n3622),
    .c(net301),
    .d(n3623),
    .o1(n3625));
 b15oaoi13aq1n03x5 U4177 (.a(n3625),
    .b(n3626),
    .c(n3628),
    .d(n3627),
    .o1(n3629));
 b15aoai13as1n08x5 U4178 (.a(n3629),
    .b(n3819),
    .c(n3632),
    .d(n3631),
    .o1(u_device_sm_tx_counter_next_3_));
 b15aoai13as1n04x5 U4179 (.a(net309),
    .b(net324),
    .c(n3633),
    .d(net311),
    .o1(n3662));
 b15aoi012as1n12x5 U4180 (.a(n3634),
    .b(net321),
    .c(n3635),
    .o1(n3660));
 b15inv000an1n08x5 U4181 (.a(n3636),
    .o1(n3658));
 b15oai112al1n16x5 U4182 (.a(n3638),
    .b(n3637),
    .c(n3640),
    .d(n3639),
    .o1(n3657));
 b15nandp2an1n02x5 U4183 (.a(net323),
    .b(net308),
    .o1(n3642));
 b15aoi012aq1n04x5 U4184 (.a(n3641),
    .b(n3643),
    .c(n3642),
    .o1(n3656));
 b15nand02an1n02x5 U4185 (.a(net310),
    .b(net313),
    .o1(n3646));
 b15nand02ar1n02x5 U4186 (.a(net321),
    .b(net319),
    .o1(n3644));
 b15oai022al1n04x5 U4187 (.a(n3647),
    .b(n3646),
    .c(n3645),
    .d(n3644),
    .o1(n3648));
 b15aoi013ar1n04x5 U4188 (.a(n3648),
    .b(net313),
    .c(net315),
    .d(n3649),
    .o1(n3652));
 b15oai112al1n08x5 U4189 (.a(net317),
    .b(net315),
    .c(n3650),
    .d(n3649),
    .o1(n3651));
 b15oai112al1n12x5 U4190 (.a(n3652),
    .b(n3651),
    .c(n3654),
    .d(n3653),
    .o1(n3655));
 b15aoi112as1n08x5 U4191 (.a(n3656),
    .b(n3655),
    .c(n3658),
    .d(n3657),
    .o1(n3659));
 b15aoai13as1n08x5 U4192 (.a(n3659),
    .b(n3660),
    .c(n3662),
    .d(n3661),
    .o1(u_dcfifo_tx_u_din_full_full_dn));
 b15aoi022ar1n32x5 U4193 (.a(n3664),
    .b(u_device_sm_s_dummy_cycles[1]),
    .c(n3663),
    .d(u_device_sm_u_spiregs_n[15]),
    .o1(n3683));
 b15aoi022aq1n12x5 U4194 (.a(n3666),
    .b(u_device_sm_u_spiregs_reg0[1]),
    .c(n3665),
    .d(u_device_sm_u_spiregs_n[7]),
    .o1(n3682));
 b15aoi022aq1n16x5 U4195 (.a(net177),
    .b(u_dcfifo_tx_u_din_buffer_data[1]),
    .c(net182),
    .d(u_dcfifo_tx_u_din_buffer_data[33]),
    .o1(n3678));
 b15aoi022ar1n16x5 U4196 (.a(net188),
    .b(u_dcfifo_tx_u_din_buffer_data[193]),
    .c(net180),
    .d(u_dcfifo_tx_u_din_buffer_data[65]),
    .o1(n3677));
 b15aoi022ah1n12x5 U4197 (.a(net172),
    .b(u_dcfifo_tx_u_din_buffer_data[161]),
    .c(net174),
    .d(u_dcfifo_tx_u_din_buffer_data[225]),
    .o1(n3676));
 b15aoi022an1n16x5 U4198 (.a(net185),
    .b(u_dcfifo_tx_u_din_buffer_data[129]),
    .c(net169),
    .d(u_dcfifo_tx_u_din_buffer_data[97]),
    .o1(n3675));
 b15nand04as1n16x5 U4199 (.a(n3678),
    .b(n3677),
    .c(n3676),
    .d(n3675),
    .o1(n3679));
 b15nand02aq1n02x5 U4200 (.a(n3681),
    .b(n3679),
    .o1(n3680));
 b15aoai13aq1n08x5 U4201 (.a(n3680),
    .b(n3681),
    .c(n3683),
    .d(n3682),
    .o1(u_device_sm_N175));
 b15aoi022ar1n02x5 U4204 (.a(net352),
    .b(net2222),
    .c(net260),
    .d(u_txreg_data_int[4]),
    .o1(n3685));
 b15aob012an1n04x5 U4205 (.a(net2223),
    .b(net256),
    .c(u_txreg_data_int[1]),
    .out0(u_txreg_N39));
 b15aoi022al1n04x5 U4206 (.a(net352),
    .b(net2217),
    .c(net260),
    .d(u_txreg_data_int[3]),
    .o1(n3688));
 b15aob012al1n04x5 U4207 (.a(net2218),
    .b(net256),
    .c(u_txreg_data_int[0]),
    .out0(u_txreg_N38));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_0__0_latch (.clk(clknet_3_6__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net746),
    .en(u_dcfifo_rx_u_din_buffer_N26),
    .te(net477));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_0__latch (.clk(clknet_3_6__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net741),
    .en(u_dcfifo_rx_u_din_buffer_N26),
    .te(net478));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_1__0_latch (.clk(clknet_3_7__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net736),
    .en(u_dcfifo_rx_u_din_buffer_N27),
    .te(net479));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_1__latch (.clk(clknet_3_7__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net731),
    .en(u_dcfifo_rx_u_din_buffer_N27),
    .te(net480));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_2__0_latch (.clk(clknet_3_7__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net726),
    .en(net133),
    .te(net481));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_2__latch (.clk(clknet_3_5__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net721),
    .en(net133),
    .te(net482));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_3__0_latch (.clk(clknet_3_6__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net716),
    .en(u_dcfifo_rx_u_din_buffer_N29),
    .te(net483));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_3__latch (.clk(clknet_3_4__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net711),
    .en(u_dcfifo_rx_u_din_buffer_N29),
    .te(net484));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_4__0_latch (.clk(clknet_3_7__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net706),
    .en(u_dcfifo_rx_u_din_buffer_N30),
    .te(net485));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_4__latch (.clk(clknet_3_4__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net701),
    .en(u_dcfifo_rx_u_din_buffer_N30),
    .te(net486));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_5__0_latch (.clk(clknet_3_7__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net696),
    .en(u_dcfifo_rx_u_din_buffer_N31),
    .te(net487));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_5__latch (.clk(clknet_3_5__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net691),
    .en(u_dcfifo_rx_u_din_buffer_N31),
    .te(net488));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_6__0_latch (.clk(clknet_3_7__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net686),
    .en(u_dcfifo_rx_u_din_buffer_N32),
    .te(net489));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_6__latch (.clk(clknet_3_7__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net681),
    .en(u_dcfifo_rx_u_din_buffer_N32),
    .te(net490));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_7__0_latch (.clk(clknet_3_7__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net676),
    .en(u_dcfifo_rx_u_din_buffer_N33),
    .te(net491));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_7__latch (.clk(clknet_3_5__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_buffer_net670),
    .en(u_dcfifo_rx_u_din_buffer_N33),
    .te(net492));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__0__u_dcfifo_rx_u_din_buffer_data_reg_0__1_ (.rb(net445),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net741),
    .d1(n3818),
    .d2(ctrl_data_rx[1]),
    .o1(u_dcfifo_rx_u_din_buffer_data[0]),
    .o2(u_dcfifo_rx_u_din_buffer_data[1]),
    .si1(net493),
    .si2(net494),
    .ssb(net1476));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__10__u_dcfifo_rx_u_din_buffer_data_reg_0__11_ (.rb(net445),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net741),
    .d1(ctrl_data_rx[10]),
    .d2(ctrl_data_rx[11]),
    .o1(u_dcfifo_rx_u_din_buffer_data[10]),
    .o2(u_dcfifo_rx_u_din_buffer_data[11]),
    .si1(net495),
    .si2(net496),
    .ssb(net1477));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__12__u_dcfifo_rx_u_din_buffer_data_reg_0__13_ (.rb(net445),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net741),
    .d1(net194),
    .d2(net214),
    .o1(u_dcfifo_rx_u_din_buffer_data[12]),
    .o2(u_dcfifo_rx_u_din_buffer_data[13]),
    .si1(net497),
    .si2(net498),
    .ssb(net1478));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__14__u_dcfifo_rx_u_din_buffer_data_reg_0__15_ (.rb(net445),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net741),
    .d1(ctrl_data_rx[14]),
    .d2(net192),
    .o1(u_dcfifo_rx_u_din_buffer_data[14]),
    .o2(u_dcfifo_rx_u_din_buffer_data[15]),
    .si1(net499),
    .si2(net500),
    .ssb(net1479));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__16__u_dcfifo_rx_u_din_buffer_data_reg_0__17_ (.rb(net443),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net746),
    .d1(ctrl_data_rx[16]),
    .d2(net226),
    .o1(u_dcfifo_rx_u_din_buffer_data[16]),
    .o2(u_dcfifo_rx_u_din_buffer_data[17]),
    .si1(net501),
    .si2(net502),
    .ssb(net1480));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__18__u_dcfifo_rx_u_din_buffer_data_reg_0__19_ (.rb(net443),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net746),
    .d1(net204),
    .d2(net216),
    .o1(u_dcfifo_rx_u_din_buffer_data[18]),
    .o2(u_dcfifo_rx_u_din_buffer_data[19]),
    .si1(net503),
    .si2(net504),
    .ssb(net1481));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__20__u_dcfifo_rx_u_din_buffer_data_reg_0__21_ (.rb(net443),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net746),
    .d1(net228),
    .d2(net196),
    .o1(u_dcfifo_rx_u_din_buffer_data[20]),
    .o2(u_dcfifo_rx_u_din_buffer_data[21]),
    .si1(net505),
    .si2(net506),
    .ssb(net1482));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__22__u_dcfifo_rx_u_din_buffer_data_reg_0__23_ (.rb(net444),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net746),
    .d1(net219),
    .d2(net223),
    .o1(u_dcfifo_rx_u_din_buffer_data[22]),
    .o2(u_dcfifo_rx_u_din_buffer_data[23]),
    .si1(net507),
    .si2(net508),
    .ssb(net1483));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__24__u_dcfifo_rx_u_din_buffer_data_reg_0__25_ (.rb(net444),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net746),
    .d1(net198),
    .d2(net210),
    .o1(u_dcfifo_rx_u_din_buffer_data[24]),
    .o2(u_dcfifo_rx_u_din_buffer_data[25]),
    .si1(net509),
    .si2(net510),
    .ssb(net1484));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__26__u_dcfifo_rx_u_din_buffer_data_reg_0__27_ (.rb(net443),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net746),
    .d1(net202),
    .d2(net200),
    .o1(u_dcfifo_rx_u_din_buffer_data[26]),
    .o2(u_dcfifo_rx_u_din_buffer_data[27]),
    .si1(net511),
    .si2(net512),
    .ssb(net1485));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__28__u_dcfifo_rx_u_din_buffer_data_reg_0__29_ (.rb(net444),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net746),
    .d1(net206),
    .d2(net232),
    .o1(u_dcfifo_rx_u_din_buffer_data[28]),
    .o2(u_dcfifo_rx_u_din_buffer_data[29]),
    .si1(net513),
    .si2(net514),
    .ssb(net1486));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__2__u_dcfifo_rx_u_din_buffer_data_reg_0__3_ (.rb(net445),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net741),
    .d1(net237),
    .d2(net247),
    .o1(u_dcfifo_rx_u_din_buffer_data[2]),
    .o2(u_dcfifo_rx_u_din_buffer_data[3]),
    .si1(net515),
    .si2(net516),
    .ssb(net1487));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__30__u_dcfifo_rx_u_din_buffer_data_reg_0__31_ (.rb(net443),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net746),
    .d1(net208),
    .d2(ctrl_data_rx[31]),
    .o1(u_dcfifo_rx_u_din_buffer_data[30]),
    .o2(u_dcfifo_rx_u_din_buffer_data[31]),
    .si1(net517),
    .si2(net518),
    .ssb(net1488));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__4__u_dcfifo_rx_u_din_buffer_data_reg_0__5_ (.rb(net445),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net741),
    .d1(ctrl_data_rx[4]),
    .d2(n3820),
    .o1(u_dcfifo_rx_u_din_buffer_data[4]),
    .o2(u_dcfifo_rx_u_din_buffer_data[5]),
    .si1(net519),
    .si2(net520),
    .ssb(net1489));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__6__u_dcfifo_rx_u_din_buffer_data_reg_0__7_ (.rb(net445),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net741),
    .d1(net242),
    .d2(net245),
    .o1(u_dcfifo_rx_u_din_buffer_data[6]),
    .o2(u_dcfifo_rx_u_din_buffer_data[7]),
    .si1(net521),
    .si2(net522),
    .ssb(net1490));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_0__8__u_dcfifo_rx_u_din_buffer_data_reg_0__9_ (.rb(net445),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net741),
    .d1(ctrl_data_rx[8]),
    .d2(ctrl_data_rx[9]),
    .o1(u_dcfifo_rx_u_din_buffer_data[8]),
    .o2(u_dcfifo_rx_u_din_buffer_data[9]),
    .si1(net523),
    .si2(net524),
    .ssb(net1491));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__0__u_dcfifo_rx_u_din_buffer_data_reg_1__1_ (.rb(net461),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net731),
    .d1(net259),
    .d2(net239),
    .o1(u_dcfifo_rx_u_din_buffer_data[32]),
    .o2(u_dcfifo_rx_u_din_buffer_data[33]),
    .si1(net525),
    .si2(net526),
    .ssb(net1492));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__10__u_dcfifo_rx_u_din_buffer_data_reg_1__11_ (.rb(net462),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net731),
    .d1(net217),
    .d2(net229),
    .o1(u_dcfifo_rx_u_din_buffer_data[42]),
    .o2(u_dcfifo_rx_u_din_buffer_data[43]),
    .si1(net527),
    .si2(net528),
    .ssb(net1493));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__12__u_dcfifo_rx_u_din_buffer_data_reg_1__13_ (.rb(net462),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net731),
    .d1(net193),
    .d2(net213),
    .o1(u_dcfifo_rx_u_din_buffer_data[44]),
    .o2(u_dcfifo_rx_u_din_buffer_data[45]),
    .si1(net529),
    .si2(net530),
    .ssb(net1494));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__14__u_dcfifo_rx_u_din_buffer_data_reg_1__15_ (.rb(net461),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net731),
    .d1(net220),
    .d2(net192),
    .o1(u_dcfifo_rx_u_din_buffer_data[46]),
    .o2(u_dcfifo_rx_u_din_buffer_data[47]),
    .si1(net531),
    .si2(net532),
    .ssb(net1495));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__16__u_dcfifo_rx_u_din_buffer_data_reg_1__17_ (.rb(net462),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net736),
    .d1(net211),
    .d2(net224),
    .o1(u_dcfifo_rx_u_din_buffer_data[48]),
    .o2(u_dcfifo_rx_u_din_buffer_data[49]),
    .si1(net533),
    .si2(net534),
    .ssb(net1496));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__18__u_dcfifo_rx_u_din_buffer_data_reg_1__19_ (.rb(net462),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net736),
    .d1(net203),
    .d2(net215),
    .o1(u_dcfifo_rx_u_din_buffer_data[50]),
    .o2(u_dcfifo_rx_u_din_buffer_data[51]),
    .si1(net535),
    .si2(net536),
    .ssb(net1497));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__20__u_dcfifo_rx_u_din_buffer_data_reg_1__21_ (.rb(net462),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net736),
    .d1(net228),
    .d2(net196),
    .o1(u_dcfifo_rx_u_din_buffer_data[52]),
    .o2(u_dcfifo_rx_u_din_buffer_data[53]),
    .si1(net537),
    .si2(net538),
    .ssb(net1498));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__22__u_dcfifo_rx_u_din_buffer_data_reg_1__23_ (.rb(net462),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net736),
    .d1(net218),
    .d2(net222),
    .o1(u_dcfifo_rx_u_din_buffer_data[54]),
    .o2(u_dcfifo_rx_u_din_buffer_data[55]),
    .si1(net539),
    .si2(net540),
    .ssb(net1499));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__24__u_dcfifo_rx_u_din_buffer_data_reg_1__25_ (.rb(net462),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net736),
    .d1(net197),
    .d2(net209),
    .o1(u_dcfifo_rx_u_din_buffer_data[56]),
    .o2(u_dcfifo_rx_u_din_buffer_data[57]),
    .si1(net541),
    .si2(net542),
    .ssb(net1500));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__26__u_dcfifo_rx_u_din_buffer_data_reg_1__27_ (.rb(net462),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net736),
    .d1(net201),
    .d2(net199),
    .o1(u_dcfifo_rx_u_din_buffer_data[58]),
    .o2(u_dcfifo_rx_u_din_buffer_data[59]),
    .si1(net543),
    .si2(net544),
    .ssb(net1501));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__28__u_dcfifo_rx_u_din_buffer_data_reg_1__29_ (.rb(net463),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net736),
    .d1(net205),
    .d2(net231),
    .o1(u_dcfifo_rx_u_din_buffer_data[60]),
    .o2(u_dcfifo_rx_u_din_buffer_data[61]),
    .si1(net545),
    .si2(net546),
    .ssb(net1502));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__2__u_dcfifo_rx_u_din_buffer_data_reg_1__3_ (.rb(net461),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net731),
    .d1(net236),
    .d2(net248),
    .o1(u_dcfifo_rx_u_din_buffer_data[34]),
    .o2(u_dcfifo_rx_u_din_buffer_data[35]),
    .si1(net547),
    .si2(net548),
    .ssb(net1503));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__30__u_dcfifo_rx_u_din_buffer_data_reg_1__31_ (.rb(net463),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net736),
    .d1(net207),
    .d2(net230),
    .o1(u_dcfifo_rx_u_din_buffer_data[62]),
    .o2(u_dcfifo_rx_u_din_buffer_data[63]),
    .si1(net549),
    .si2(net550),
    .ssb(net1504));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__4__u_dcfifo_rx_u_din_buffer_data_reg_1__5_ (.rb(net461),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net731),
    .d1(net233),
    .d2(net190),
    .o1(u_dcfifo_rx_u_din_buffer_data[36]),
    .o2(u_dcfifo_rx_u_din_buffer_data[37]),
    .si1(net551),
    .si2(net552),
    .ssb(net1505));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__6__u_dcfifo_rx_u_din_buffer_data_reg_1__7_ (.rb(net462),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net731),
    .d1(net242),
    .d2(net245),
    .o1(u_dcfifo_rx_u_din_buffer_data[38]),
    .o2(u_dcfifo_rx_u_din_buffer_data[39]),
    .si1(net553),
    .si2(net554),
    .ssb(net1506));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_1__8__u_dcfifo_rx_u_din_buffer_data_reg_1__9_ (.rb(net461),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net731),
    .d1(ctrl_data_rx[8]),
    .d2(ctrl_data_rx[9]),
    .o1(u_dcfifo_rx_u_din_buffer_data[40]),
    .o2(u_dcfifo_rx_u_din_buffer_data[41]),
    .si1(net555),
    .si2(net556),
    .ssb(net1507));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__0__u_dcfifo_rx_u_din_buffer_data_reg_2__1_ (.rb(net451),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net721),
    .d1(net259),
    .d2(net239),
    .o1(u_dcfifo_rx_u_din_buffer_data[64]),
    .o2(u_dcfifo_rx_u_din_buffer_data[65]),
    .si1(net557),
    .si2(net558),
    .ssb(net1508));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__10__u_dcfifo_rx_u_din_buffer_data_reg_2__11_ (.rb(net451),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net721),
    .d1(net217),
    .d2(net229),
    .o1(u_dcfifo_rx_u_din_buffer_data[74]),
    .o2(u_dcfifo_rx_u_din_buffer_data[75]),
    .si1(net559),
    .si2(net560),
    .ssb(net1509));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__12__u_dcfifo_rx_u_din_buffer_data_reg_2__13_ (.rb(net451),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net721),
    .d1(net193),
    .d2(net213),
    .o1(u_dcfifo_rx_u_din_buffer_data[76]),
    .o2(u_dcfifo_rx_u_din_buffer_data[77]),
    .si1(net561),
    .si2(net562),
    .ssb(net1510));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__14__u_dcfifo_rx_u_din_buffer_data_reg_2__15_ (.rb(net451),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net721),
    .d1(net221),
    .d2(ctrl_data_rx[15]),
    .o1(u_dcfifo_rx_u_din_buffer_data[78]),
    .o2(u_dcfifo_rx_u_din_buffer_data[79]),
    .si1(net563),
    .si2(net564),
    .ssb(net1511));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__16__u_dcfifo_rx_u_din_buffer_data_reg_2__17_ (.rb(net462),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net726),
    .d1(net211),
    .d2(net224),
    .o1(u_dcfifo_rx_u_din_buffer_data[80]),
    .o2(u_dcfifo_rx_u_din_buffer_data[81]),
    .si1(net565),
    .si2(net566),
    .ssb(net1512));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__18__u_dcfifo_rx_u_din_buffer_data_reg_2__19_ (.rb(net462),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net726),
    .d1(net203),
    .d2(net215),
    .o1(u_dcfifo_rx_u_din_buffer_data[82]),
    .o2(u_dcfifo_rx_u_din_buffer_data[83]),
    .si1(net567),
    .si2(net568),
    .ssb(net1513));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__20__u_dcfifo_rx_u_din_buffer_data_reg_2__21_ (.rb(net462),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net726),
    .d1(net227),
    .d2(net195),
    .o1(u_dcfifo_rx_u_din_buffer_data[84]),
    .o2(u_dcfifo_rx_u_din_buffer_data[85]),
    .si1(net569),
    .si2(net570),
    .ssb(net1514));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__22__u_dcfifo_rx_u_din_buffer_data_reg_2__23_ (.rb(net463),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net726),
    .d1(net218),
    .d2(net222),
    .o1(u_dcfifo_rx_u_din_buffer_data[86]),
    .o2(u_dcfifo_rx_u_din_buffer_data[87]),
    .si1(net571),
    .si2(net572),
    .ssb(net1515));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__24__u_dcfifo_rx_u_din_buffer_data_reg_2__25_ (.rb(net462),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net726),
    .d1(net197),
    .d2(net209),
    .o1(u_dcfifo_rx_u_din_buffer_data[88]),
    .o2(u_dcfifo_rx_u_din_buffer_data[89]),
    .si1(net573),
    .si2(net574),
    .ssb(net1516));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__26__u_dcfifo_rx_u_din_buffer_data_reg_2__27_ (.rb(net462),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net726),
    .d1(net201),
    .d2(net199),
    .o1(u_dcfifo_rx_u_din_buffer_data[90]),
    .o2(u_dcfifo_rx_u_din_buffer_data[91]),
    .si1(net575),
    .si2(net576),
    .ssb(net1517));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__28__u_dcfifo_rx_u_din_buffer_data_reg_2__29_ (.rb(net462),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net726),
    .d1(net205),
    .d2(net231),
    .o1(u_dcfifo_rx_u_din_buffer_data[92]),
    .o2(u_dcfifo_rx_u_din_buffer_data[93]),
    .si1(net577),
    .si2(net578),
    .ssb(net1518));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__2__u_dcfifo_rx_u_din_buffer_data_reg_2__3_ (.rb(net451),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net721),
    .d1(ctrl_data_rx[2]),
    .d2(net248),
    .o1(u_dcfifo_rx_u_din_buffer_data[66]),
    .o2(u_dcfifo_rx_u_din_buffer_data[67]),
    .si1(net579),
    .si2(net580),
    .ssb(net1519));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__30__u_dcfifo_rx_u_din_buffer_data_reg_2__31_ (.rb(net462),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net726),
    .d1(net207),
    .d2(net230),
    .o1(u_dcfifo_rx_u_din_buffer_data[94]),
    .o2(u_dcfifo_rx_u_din_buffer_data[95]),
    .si1(net581),
    .si2(net582),
    .ssb(net1520));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__4__u_dcfifo_rx_u_din_buffer_data_reg_2__5_ (.rb(net451),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net721),
    .d1(net233),
    .d2(net190),
    .o1(u_dcfifo_rx_u_din_buffer_data[68]),
    .o2(u_dcfifo_rx_u_din_buffer_data[69]),
    .si1(net583),
    .si2(net584),
    .ssb(net1521));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__6__u_dcfifo_rx_u_din_buffer_data_reg_2__7_ (.rb(net451),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net721),
    .d1(net241),
    .d2(net244),
    .o1(u_dcfifo_rx_u_din_buffer_data[70]),
    .o2(u_dcfifo_rx_u_din_buffer_data[71]),
    .si1(net585),
    .si2(net586),
    .ssb(net1522));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_2__8__u_dcfifo_rx_u_din_buffer_data_reg_2__9_ (.rb(net451),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net721),
    .d1(ctrl_data_rx[8]),
    .d2(ctrl_data_rx[9]),
    .o1(u_dcfifo_rx_u_din_buffer_data[72]),
    .o2(u_dcfifo_rx_u_din_buffer_data[73]),
    .si1(net587),
    .si2(net588),
    .ssb(net1523));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__0__u_dcfifo_rx_u_din_buffer_data_reg_3__1_ (.rb(net445),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net711),
    .d1(n3818),
    .d2(ctrl_data_rx[1]),
    .o1(u_dcfifo_rx_u_din_buffer_data[96]),
    .o2(u_dcfifo_rx_u_din_buffer_data[97]),
    .si1(net589),
    .si2(net590),
    .ssb(net1524));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__10__u_dcfifo_rx_u_din_buffer_data_reg_3__11_ (.rb(net445),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net711),
    .d1(ctrl_data_rx[10]),
    .d2(ctrl_data_rx[11]),
    .o1(u_dcfifo_rx_u_din_buffer_data[106]),
    .o2(u_dcfifo_rx_u_din_buffer_data[107]),
    .si1(net591),
    .si2(net592),
    .ssb(net1525));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__12__u_dcfifo_rx_u_din_buffer_data_reg_3__13_ (.rb(net445),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net711),
    .d1(net194),
    .d2(net214),
    .o1(u_dcfifo_rx_u_din_buffer_data[108]),
    .o2(u_dcfifo_rx_u_din_buffer_data[109]),
    .si1(net593),
    .si2(net594),
    .ssb(net1526));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__14__u_dcfifo_rx_u_din_buffer_data_reg_3__15_ (.rb(net445),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net711),
    .d1(ctrl_data_rx[14]),
    .d2(net192),
    .o1(u_dcfifo_rx_u_din_buffer_data[110]),
    .o2(u_dcfifo_rx_u_din_buffer_data[111]),
    .si1(net595),
    .si2(net596),
    .ssb(net1527));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__16__u_dcfifo_rx_u_din_buffer_data_reg_3__17_ (.rb(net443),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net716),
    .d1(ctrl_data_rx[16]),
    .d2(net226),
    .o1(u_dcfifo_rx_u_din_buffer_data[112]),
    .o2(u_dcfifo_rx_u_din_buffer_data[113]),
    .si1(net597),
    .si2(net598),
    .ssb(net1528));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__18__u_dcfifo_rx_u_din_buffer_data_reg_3__19_ (.rb(net443),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net716),
    .d1(net203),
    .d2(net215),
    .o1(u_dcfifo_rx_u_din_buffer_data[114]),
    .o2(u_dcfifo_rx_u_din_buffer_data[115]),
    .si1(net599),
    .si2(net600),
    .ssb(net1529));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__20__u_dcfifo_rx_u_din_buffer_data_reg_3__21_ (.rb(net459),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net716),
    .d1(net227),
    .d2(net195),
    .o1(u_dcfifo_rx_u_din_buffer_data[116]),
    .o2(u_dcfifo_rx_u_din_buffer_data[117]),
    .si1(net601),
    .si2(net602),
    .ssb(net1530));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__22__u_dcfifo_rx_u_din_buffer_data_reg_3__23_ (.rb(net443),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net716),
    .d1(net219),
    .d2(net223),
    .o1(u_dcfifo_rx_u_din_buffer_data[118]),
    .o2(u_dcfifo_rx_u_din_buffer_data[119]),
    .si1(net603),
    .si2(net604),
    .ssb(net1531));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__24__u_dcfifo_rx_u_din_buffer_data_reg_3__25_ (.rb(net443),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net716),
    .d1(net198),
    .d2(net210),
    .o1(u_dcfifo_rx_u_din_buffer_data[120]),
    .o2(u_dcfifo_rx_u_din_buffer_data[121]),
    .si1(net605),
    .si2(net606),
    .ssb(net1532));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__26__u_dcfifo_rx_u_din_buffer_data_reg_3__27_ (.rb(net459),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net716),
    .d1(net202),
    .d2(net200),
    .o1(u_dcfifo_rx_u_din_buffer_data[122]),
    .o2(u_dcfifo_rx_u_din_buffer_data[123]),
    .si1(net607),
    .si2(net608),
    .ssb(net1533));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__28__u_dcfifo_rx_u_din_buffer_data_reg_3__29_ (.rb(net443),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net716),
    .d1(net205),
    .d2(net231),
    .o1(u_dcfifo_rx_u_din_buffer_data[124]),
    .o2(u_dcfifo_rx_u_din_buffer_data[125]),
    .si1(net609),
    .si2(net610),
    .ssb(net1534));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__2__u_dcfifo_rx_u_din_buffer_data_reg_3__3_ (.rb(net458),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net711),
    .d1(net237),
    .d2(net247),
    .o1(u_dcfifo_rx_u_din_buffer_data[98]),
    .o2(u_dcfifo_rx_u_din_buffer_data[99]),
    .si1(net611),
    .si2(net612),
    .ssb(net1535));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__30__u_dcfifo_rx_u_din_buffer_data_reg_3__31_ (.rb(net459),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net716),
    .d1(net208),
    .d2(ctrl_data_rx[31]),
    .o1(u_dcfifo_rx_u_din_buffer_data[126]),
    .o2(u_dcfifo_rx_u_din_buffer_data[127]),
    .si1(net613),
    .si2(net614),
    .ssb(net1536));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__4__u_dcfifo_rx_u_din_buffer_data_reg_3__5_ (.rb(net445),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net711),
    .d1(ctrl_data_rx[4]),
    .d2(n3820),
    .o1(u_dcfifo_rx_u_din_buffer_data[100]),
    .o2(u_dcfifo_rx_u_din_buffer_data[101]),
    .si1(net615),
    .si2(net616),
    .ssb(net1537));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__6__u_dcfifo_rx_u_din_buffer_data_reg_3__7_ (.rb(net445),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net711),
    .d1(net242),
    .d2(net245),
    .o1(u_dcfifo_rx_u_din_buffer_data[102]),
    .o2(u_dcfifo_rx_u_din_buffer_data[103]),
    .si1(net617),
    .si2(net618),
    .ssb(net1538));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_3__8__u_dcfifo_rx_u_din_buffer_data_reg_3__9_ (.rb(net445),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net711),
    .d1(ctrl_data_rx[8]),
    .d2(ctrl_data_rx[9]),
    .o1(u_dcfifo_rx_u_din_buffer_data[104]),
    .o2(u_dcfifo_rx_u_din_buffer_data[105]),
    .si1(net619),
    .si2(net620),
    .ssb(net1539));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__0__u_dcfifo_rx_u_din_buffer_data_reg_4__1_ (.rb(net459),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net701),
    .d1(n3818),
    .d2(ctrl_data_rx[1]),
    .o1(u_dcfifo_rx_u_din_buffer_data[128]),
    .o2(u_dcfifo_rx_u_din_buffer_data[129]),
    .si1(net621),
    .si2(net622),
    .ssb(net1540));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__10__u_dcfifo_rx_u_din_buffer_data_reg_4__11_ (.rb(net458),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net701),
    .d1(ctrl_data_rx[10]),
    .d2(ctrl_data_rx[11]),
    .o1(u_dcfifo_rx_u_din_buffer_data[138]),
    .o2(u_dcfifo_rx_u_din_buffer_data[139]),
    .si1(net623),
    .si2(net624),
    .ssb(net1541));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__12__u_dcfifo_rx_u_din_buffer_data_reg_4__13_ (.rb(net458),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net701),
    .d1(net194),
    .d2(net214),
    .o1(u_dcfifo_rx_u_din_buffer_data[140]),
    .o2(u_dcfifo_rx_u_din_buffer_data[141]),
    .si1(net625),
    .si2(net626),
    .ssb(net1542));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__14__u_dcfifo_rx_u_din_buffer_data_reg_4__15_ (.rb(net458),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net701),
    .d1(net220),
    .d2(net192),
    .o1(u_dcfifo_rx_u_din_buffer_data[142]),
    .o2(u_dcfifo_rx_u_din_buffer_data[143]),
    .si1(net627),
    .si2(net628),
    .ssb(net1543));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__16__u_dcfifo_rx_u_din_buffer_data_reg_4__17_ (.rb(net443),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net706),
    .d1(ctrl_data_rx[16]),
    .d2(net226),
    .o1(u_dcfifo_rx_u_din_buffer_data[144]),
    .o2(u_dcfifo_rx_u_din_buffer_data[145]),
    .si1(net629),
    .si2(net630),
    .ssb(net1544));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__18__u_dcfifo_rx_u_din_buffer_data_reg_4__19_ (.rb(net443),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net706),
    .d1(net204),
    .d2(net216),
    .o1(u_dcfifo_rx_u_din_buffer_data[146]),
    .o2(u_dcfifo_rx_u_din_buffer_data[147]),
    .si1(net631),
    .si2(net632),
    .ssb(net1545));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__20__u_dcfifo_rx_u_din_buffer_data_reg_4__21_ (.rb(net443),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net706),
    .d1(net227),
    .d2(net195),
    .o1(u_dcfifo_rx_u_din_buffer_data[148]),
    .o2(u_dcfifo_rx_u_din_buffer_data[149]),
    .si1(net633),
    .si2(net634),
    .ssb(net1546));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__22__u_dcfifo_rx_u_din_buffer_data_reg_4__23_ (.rb(net443),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net706),
    .d1(net219),
    .d2(net223),
    .o1(u_dcfifo_rx_u_din_buffer_data[150]),
    .o2(u_dcfifo_rx_u_din_buffer_data[151]),
    .si1(net635),
    .si2(net636),
    .ssb(net1547));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__24__u_dcfifo_rx_u_din_buffer_data_reg_4__25_ (.rb(net443),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net706),
    .d1(net198),
    .d2(net210),
    .o1(u_dcfifo_rx_u_din_buffer_data[152]),
    .o2(u_dcfifo_rx_u_din_buffer_data[153]),
    .si1(net637),
    .si2(net638),
    .ssb(net1548));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__26__u_dcfifo_rx_u_din_buffer_data_reg_4__27_ (.rb(net443),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net706),
    .d1(net202),
    .d2(net200),
    .o1(u_dcfifo_rx_u_din_buffer_data[154]),
    .o2(u_dcfifo_rx_u_din_buffer_data[155]),
    .si1(net639),
    .si2(net640),
    .ssb(net1549));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__28__u_dcfifo_rx_u_din_buffer_data_reg_4__29_ (.rb(net444),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net706),
    .d1(net206),
    .d2(net232),
    .o1(u_dcfifo_rx_u_din_buffer_data[156]),
    .o2(u_dcfifo_rx_u_din_buffer_data[157]),
    .si1(net641),
    .si2(net642),
    .ssb(net1550));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__2__u_dcfifo_rx_u_din_buffer_data_reg_4__3_ (.rb(net459),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net701),
    .d1(net237),
    .d2(net247),
    .o1(u_dcfifo_rx_u_din_buffer_data[130]),
    .o2(u_dcfifo_rx_u_din_buffer_data[131]),
    .si1(net643),
    .si2(net644),
    .ssb(net1551));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__30__u_dcfifo_rx_u_din_buffer_data_reg_4__31_ (.rb(net444),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net706),
    .d1(net208),
    .d2(ctrl_data_rx[31]),
    .o1(u_dcfifo_rx_u_din_buffer_data[158]),
    .o2(u_dcfifo_rx_u_din_buffer_data[159]),
    .si1(net645),
    .si2(net646),
    .ssb(net1552));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__4__u_dcfifo_rx_u_din_buffer_data_reg_4__5_ (.rb(net459),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net701),
    .d1(ctrl_data_rx[4]),
    .d2(n3820),
    .o1(u_dcfifo_rx_u_din_buffer_data[132]),
    .o2(u_dcfifo_rx_u_din_buffer_data[133]),
    .si1(net647),
    .si2(net648),
    .ssb(net1553));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__6__u_dcfifo_rx_u_din_buffer_data_reg_4__7_ (.rb(net459),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net701),
    .d1(net242),
    .d2(net245),
    .o1(u_dcfifo_rx_u_din_buffer_data[134]),
    .o2(u_dcfifo_rx_u_din_buffer_data[135]),
    .si1(net649),
    .si2(net650),
    .ssb(net1554));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_4__8__u_dcfifo_rx_u_din_buffer_data_reg_4__9_ (.rb(net458),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net701),
    .d1(ctrl_data_rx[8]),
    .d2(ctrl_data_rx[9]),
    .o1(u_dcfifo_rx_u_din_buffer_data[136]),
    .o2(u_dcfifo_rx_u_din_buffer_data[137]),
    .si1(net651),
    .si2(net652),
    .ssb(net1555));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__0__u_dcfifo_rx_u_din_buffer_data_reg_5__1_ (.rb(net452),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net691),
    .d1(net259),
    .d2(net239),
    .o1(u_dcfifo_rx_u_din_buffer_data[160]),
    .o2(u_dcfifo_rx_u_din_buffer_data[161]),
    .si1(net653),
    .si2(net654),
    .ssb(net1556));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__10__u_dcfifo_rx_u_din_buffer_data_reg_5__11_ (.rb(net452),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net691),
    .d1(net217),
    .d2(net229),
    .o1(u_dcfifo_rx_u_din_buffer_data[170]),
    .o2(u_dcfifo_rx_u_din_buffer_data[171]),
    .si1(net655),
    .si2(net656),
    .ssb(net1557));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__12__u_dcfifo_rx_u_din_buffer_data_reg_5__13_ (.rb(net452),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net691),
    .d1(ctrl_data_rx[12]),
    .d2(ctrl_data_rx[13]),
    .o1(u_dcfifo_rx_u_din_buffer_data[172]),
    .o2(u_dcfifo_rx_u_din_buffer_data[173]),
    .si1(net657),
    .si2(net658),
    .ssb(net1558));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__14__u_dcfifo_rx_u_din_buffer_data_reg_5__15_ (.rb(net452),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net691),
    .d1(net221),
    .d2(ctrl_data_rx[15]),
    .o1(u_dcfifo_rx_u_din_buffer_data[174]),
    .o2(u_dcfifo_rx_u_din_buffer_data[175]),
    .si1(net659),
    .si2(net660),
    .ssb(net1559));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__16__u_dcfifo_rx_u_din_buffer_data_reg_5__17_ (.rb(net459),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net696),
    .d1(net211),
    .d2(net224),
    .o1(u_dcfifo_rx_u_din_buffer_data[176]),
    .o2(u_dcfifo_rx_u_din_buffer_data[177]),
    .si1(net661),
    .si2(net662),
    .ssb(net1560));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__18__u_dcfifo_rx_u_din_buffer_data_reg_5__19_ (.rb(net459),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net696),
    .d1(net204),
    .d2(net216),
    .o1(u_dcfifo_rx_u_din_buffer_data[178]),
    .o2(u_dcfifo_rx_u_din_buffer_data[179]),
    .si1(net663),
    .si2(net664),
    .ssb(net1561));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__20__u_dcfifo_rx_u_din_buffer_data_reg_5__21_ (.rb(net459),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net696),
    .d1(net228),
    .d2(net196),
    .o1(u_dcfifo_rx_u_din_buffer_data[180]),
    .o2(u_dcfifo_rx_u_din_buffer_data[181]),
    .si1(net665),
    .si2(net666),
    .ssb(net1562));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__22__u_dcfifo_rx_u_din_buffer_data_reg_5__23_ (.rb(net459),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net696),
    .d1(net218),
    .d2(net222),
    .o1(u_dcfifo_rx_u_din_buffer_data[182]),
    .o2(u_dcfifo_rx_u_din_buffer_data[183]),
    .si1(net667),
    .si2(net668),
    .ssb(net1563));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__24__u_dcfifo_rx_u_din_buffer_data_reg_5__25_ (.rb(net459),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net696),
    .d1(net198),
    .d2(net210),
    .o1(u_dcfifo_rx_u_din_buffer_data[184]),
    .o2(u_dcfifo_rx_u_din_buffer_data[185]),
    .si1(net669),
    .si2(net670),
    .ssb(net1564));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__26__u_dcfifo_rx_u_din_buffer_data_reg_5__27_ (.rb(net459),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net696),
    .d1(net201),
    .d2(net199),
    .o1(u_dcfifo_rx_u_din_buffer_data[186]),
    .o2(u_dcfifo_rx_u_din_buffer_data[187]),
    .si1(net671),
    .si2(net672),
    .ssb(net1565));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__28__u_dcfifo_rx_u_din_buffer_data_reg_5__29_ (.rb(net459),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net696),
    .d1(net205),
    .d2(net231),
    .o1(u_dcfifo_rx_u_din_buffer_data[188]),
    .o2(u_dcfifo_rx_u_din_buffer_data[189]),
    .si1(net673),
    .si2(net674),
    .ssb(net1566));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__2__u_dcfifo_rx_u_din_buffer_data_reg_5__3_ (.rb(net458),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net691),
    .d1(ctrl_data_rx[2]),
    .d2(net247),
    .o1(u_dcfifo_rx_u_din_buffer_data[162]),
    .o2(u_dcfifo_rx_u_din_buffer_data[163]),
    .si1(net675),
    .si2(net676),
    .ssb(net1567));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__30__u_dcfifo_rx_u_din_buffer_data_reg_5__31_ (.rb(net459),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net696),
    .d1(net207),
    .d2(net230),
    .o1(u_dcfifo_rx_u_din_buffer_data[190]),
    .o2(u_dcfifo_rx_u_din_buffer_data[191]),
    .si1(net677),
    .si2(net678),
    .ssb(net1568));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__4__u_dcfifo_rx_u_din_buffer_data_reg_5__5_ (.rb(net458),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net691),
    .d1(net233),
    .d2(net190),
    .o1(u_dcfifo_rx_u_din_buffer_data[164]),
    .o2(u_dcfifo_rx_u_din_buffer_data[165]),
    .si1(net679),
    .si2(net680),
    .ssb(net1569));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__6__u_dcfifo_rx_u_din_buffer_data_reg_5__7_ (.rb(net457),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net691),
    .d1(net241),
    .d2(net244),
    .o1(u_dcfifo_rx_u_din_buffer_data[166]),
    .o2(u_dcfifo_rx_u_din_buffer_data[167]),
    .si1(net681),
    .si2(net682),
    .ssb(net1570));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_5__8__u_dcfifo_rx_u_din_buffer_data_reg_5__9_ (.rb(net457),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net691),
    .d1(ctrl_data_rx[8]),
    .d2(ctrl_data_rx[9]),
    .o1(u_dcfifo_rx_u_din_buffer_data[168]),
    .o2(u_dcfifo_rx_u_din_buffer_data[169]),
    .si1(net683),
    .si2(net684),
    .ssb(net1571));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__0__u_dcfifo_rx_u_din_buffer_data_reg_6__1_ (.rb(net457),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net681),
    .d1(net259),
    .d2(net239),
    .o1(u_dcfifo_rx_u_din_buffer_data[192]),
    .o2(u_dcfifo_rx_u_din_buffer_data[193]),
    .si1(net685),
    .si2(net686),
    .ssb(net1572));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__10__u_dcfifo_rx_u_din_buffer_data_reg_6__11_ (.rb(net457),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net681),
    .d1(net217),
    .d2(net229),
    .o1(u_dcfifo_rx_u_din_buffer_data[202]),
    .o2(u_dcfifo_rx_u_din_buffer_data[203]),
    .si1(net687),
    .si2(net688),
    .ssb(net1573));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__12__u_dcfifo_rx_u_din_buffer_data_reg_6__13_ (.rb(net457),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net681),
    .d1(net193),
    .d2(net213),
    .o1(u_dcfifo_rx_u_din_buffer_data[204]),
    .o2(u_dcfifo_rx_u_din_buffer_data[205]),
    .si1(net689),
    .si2(net690),
    .ssb(net1574));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__14__u_dcfifo_rx_u_din_buffer_data_reg_6__15_ (.rb(net457),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net681),
    .d1(net220),
    .d2(net192),
    .o1(u_dcfifo_rx_u_din_buffer_data[206]),
    .o2(u_dcfifo_rx_u_din_buffer_data[207]),
    .si1(net691),
    .si2(net692),
    .ssb(net1575));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__16__u_dcfifo_rx_u_din_buffer_data_reg_6__17_ (.rb(net459),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net686),
    .d1(net211),
    .d2(net224),
    .o1(u_dcfifo_rx_u_din_buffer_data[208]),
    .o2(u_dcfifo_rx_u_din_buffer_data[209]),
    .si1(net693),
    .si2(net694),
    .ssb(net1576));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__18__u_dcfifo_rx_u_din_buffer_data_reg_6__19_ (.rb(net460),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net686),
    .d1(net203),
    .d2(net215),
    .o1(u_dcfifo_rx_u_din_buffer_data[210]),
    .o2(u_dcfifo_rx_u_din_buffer_data[211]),
    .si1(net695),
    .si2(net696),
    .ssb(net1577));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__20__u_dcfifo_rx_u_din_buffer_data_reg_6__21_ (.rb(net460),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net686),
    .d1(net227),
    .d2(net195),
    .o1(u_dcfifo_rx_u_din_buffer_data[212]),
    .o2(u_dcfifo_rx_u_din_buffer_data[213]),
    .si1(net697),
    .si2(net698),
    .ssb(net1578));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__22__u_dcfifo_rx_u_din_buffer_data_reg_6__23_ (.rb(net460),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net686),
    .d1(net218),
    .d2(net222),
    .o1(u_dcfifo_rx_u_din_buffer_data[214]),
    .o2(u_dcfifo_rx_u_din_buffer_data[215]),
    .si1(net699),
    .si2(net700),
    .ssb(net1579));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__24__u_dcfifo_rx_u_din_buffer_data_reg_6__25_ (.rb(net460),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net686),
    .d1(net197),
    .d2(net209),
    .o1(u_dcfifo_rx_u_din_buffer_data[216]),
    .o2(u_dcfifo_rx_u_din_buffer_data[217]),
    .si1(net701),
    .si2(net702),
    .ssb(net1580));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__26__u_dcfifo_rx_u_din_buffer_data_reg_6__27_ (.rb(net460),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net686),
    .d1(net201),
    .d2(net199),
    .o1(u_dcfifo_rx_u_din_buffer_data[218]),
    .o2(u_dcfifo_rx_u_din_buffer_data[219]),
    .si1(net703),
    .si2(net704),
    .ssb(net1581));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__28__u_dcfifo_rx_u_din_buffer_data_reg_6__29_ (.rb(net460),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net686),
    .d1(net205),
    .d2(net231),
    .o1(u_dcfifo_rx_u_din_buffer_data[220]),
    .o2(u_dcfifo_rx_u_din_buffer_data[221]),
    .si1(net705),
    .si2(net706),
    .ssb(net1582));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__2__u_dcfifo_rx_u_din_buffer_data_reg_6__3_ (.rb(net457),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net681),
    .d1(net237),
    .d2(net247),
    .o1(u_dcfifo_rx_u_din_buffer_data[194]),
    .o2(u_dcfifo_rx_u_din_buffer_data[195]),
    .si1(net707),
    .si2(net708),
    .ssb(net1583));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__30__u_dcfifo_rx_u_din_buffer_data_reg_6__31_ (.rb(net460),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net686),
    .d1(net207),
    .d2(net230),
    .o1(u_dcfifo_rx_u_din_buffer_data[222]),
    .o2(u_dcfifo_rx_u_din_buffer_data[223]),
    .si1(net709),
    .si2(net710),
    .ssb(net1584));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__4__u_dcfifo_rx_u_din_buffer_data_reg_6__5_ (.rb(net457),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net681),
    .d1(net233),
    .d2(net190),
    .o1(u_dcfifo_rx_u_din_buffer_data[196]),
    .o2(u_dcfifo_rx_u_din_buffer_data[197]),
    .si1(net711),
    .si2(net712),
    .ssb(net1585));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__6__u_dcfifo_rx_u_din_buffer_data_reg_6__7_ (.rb(net457),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net681),
    .d1(net242),
    .d2(net245),
    .o1(u_dcfifo_rx_u_din_buffer_data[198]),
    .o2(u_dcfifo_rx_u_din_buffer_data[199]),
    .si1(net713),
    .si2(net714),
    .ssb(net1586));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_6__8__u_dcfifo_rx_u_din_buffer_data_reg_6__9_ (.rb(net457),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net681),
    .d1(ctrl_data_rx[8]),
    .d2(ctrl_data_rx[9]),
    .o1(u_dcfifo_rx_u_din_buffer_data[200]),
    .o2(u_dcfifo_rx_u_din_buffer_data[201]),
    .si1(net715),
    .si2(net716),
    .ssb(net1587));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__0__u_dcfifo_rx_u_din_buffer_data_reg_7__1_ (.rb(net457),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net670),
    .d1(net259),
    .d2(net239),
    .o1(u_dcfifo_rx_u_din_buffer_data[224]),
    .o2(u_dcfifo_rx_u_din_buffer_data[225]),
    .si1(net717),
    .si2(net718),
    .ssb(net1588));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__10__u_dcfifo_rx_u_din_buffer_data_reg_7__11_ (.rb(net457),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net670),
    .d1(net217),
    .d2(net229),
    .o1(u_dcfifo_rx_u_din_buffer_data[234]),
    .o2(u_dcfifo_rx_u_din_buffer_data[235]),
    .si1(net719),
    .si2(net720),
    .ssb(net1589));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__12__u_dcfifo_rx_u_din_buffer_data_reg_7__13_ (.rb(net457),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net670),
    .d1(net193),
    .d2(net213),
    .o1(u_dcfifo_rx_u_din_buffer_data[236]),
    .o2(u_dcfifo_rx_u_din_buffer_data[237]),
    .si1(net721),
    .si2(net722),
    .ssb(net1590));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__14__u_dcfifo_rx_u_din_buffer_data_reg_7__15_ (.rb(net457),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net670),
    .d1(net220),
    .d2(net192),
    .o1(u_dcfifo_rx_u_din_buffer_data[238]),
    .o2(u_dcfifo_rx_u_din_buffer_data[239]),
    .si1(net723),
    .si2(net724),
    .ssb(net1591));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__16__u_dcfifo_rx_u_din_buffer_data_reg_7__17_ (.rb(net460),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net676),
    .d1(net211),
    .d2(net224),
    .o1(u_dcfifo_rx_u_din_buffer_data[240]),
    .o2(u_dcfifo_rx_u_din_buffer_data[241]),
    .si1(net725),
    .si2(net726),
    .ssb(net1592));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__18__u_dcfifo_rx_u_din_buffer_data_reg_7__19_ (.rb(net460),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net676),
    .d1(net203),
    .d2(net215),
    .o1(u_dcfifo_rx_u_din_buffer_data[242]),
    .o2(u_dcfifo_rx_u_din_buffer_data[243]),
    .si1(net727),
    .si2(net728),
    .ssb(net1593));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__20__u_dcfifo_rx_u_din_buffer_data_reg_7__21_ (.rb(net460),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net676),
    .d1(net228),
    .d2(net196),
    .o1(u_dcfifo_rx_u_din_buffer_data[244]),
    .o2(u_dcfifo_rx_u_din_buffer_data[245]),
    .si1(net729),
    .si2(net730),
    .ssb(net1594));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__22__u_dcfifo_rx_u_din_buffer_data_reg_7__23_ (.rb(net460),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net676),
    .d1(net218),
    .d2(net222),
    .o1(u_dcfifo_rx_u_din_buffer_data[246]),
    .o2(u_dcfifo_rx_u_din_buffer_data[247]),
    .si1(net731),
    .si2(net732),
    .ssb(net1595));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__24__u_dcfifo_rx_u_din_buffer_data_reg_7__25_ (.rb(net460),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net676),
    .d1(net197),
    .d2(net209),
    .o1(u_dcfifo_rx_u_din_buffer_data[248]),
    .o2(u_dcfifo_rx_u_din_buffer_data[249]),
    .si1(net733),
    .si2(net734),
    .ssb(net1596));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__26__u_dcfifo_rx_u_din_buffer_data_reg_7__27_ (.rb(net460),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net676),
    .d1(net201),
    .d2(net199),
    .o1(u_dcfifo_rx_u_din_buffer_data[250]),
    .o2(u_dcfifo_rx_u_din_buffer_data[251]),
    .si1(net735),
    .si2(net736),
    .ssb(net1597));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__28__u_dcfifo_rx_u_din_buffer_data_reg_7__29_ (.rb(net460),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net676),
    .d1(net205),
    .d2(net231),
    .o1(u_dcfifo_rx_u_din_buffer_data[252]),
    .o2(u_dcfifo_rx_u_din_buffer_data[253]),
    .si1(net737),
    .si2(net738),
    .ssb(net1598));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__2__u_dcfifo_rx_u_din_buffer_data_reg_7__3_ (.rb(net458),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net670),
    .d1(net236),
    .d2(net248),
    .o1(u_dcfifo_rx_u_din_buffer_data[226]),
    .o2(u_dcfifo_rx_u_din_buffer_data[227]),
    .si1(net739),
    .si2(net740),
    .ssb(net1599));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__30__u_dcfifo_rx_u_din_buffer_data_reg_7__31_ (.rb(net460),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net676),
    .d1(net207),
    .d2(net230),
    .o1(u_dcfifo_rx_u_din_buffer_data[254]),
    .o2(u_dcfifo_rx_u_din_buffer_data[255]),
    .si1(net741),
    .si2(net742),
    .ssb(net1600));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__4__u_dcfifo_rx_u_din_buffer_data_reg_7__5_ (.rb(net457),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net670),
    .d1(net233),
    .d2(net190),
    .o1(u_dcfifo_rx_u_din_buffer_data[228]),
    .o2(u_dcfifo_rx_u_din_buffer_data[229]),
    .si1(net743),
    .si2(net744),
    .ssb(net1601));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__6__u_dcfifo_rx_u_din_buffer_data_reg_7__7_ (.rb(net457),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net670),
    .d1(net241),
    .d2(net244),
    .o1(u_dcfifo_rx_u_din_buffer_data[230]),
    .o2(u_dcfifo_rx_u_din_buffer_data[231]),
    .si1(net745),
    .si2(net746),
    .ssb(net1602));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_buffer_data_reg_7__8__u_dcfifo_rx_u_din_buffer_data_reg_7__9_ (.rb(net461),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net670),
    .d1(ctrl_data_rx[8]),
    .d2(ctrl_data_rx[9]),
    .o1(u_dcfifo_rx_u_din_buffer_data[232]),
    .o2(u_dcfifo_rx_u_din_buffer_data[233]),
    .si1(net747),
    .si2(net748),
    .ssb(net1603));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_full_full_synch_d_middle_reg_0__u_dcfifo_rx_u_din_full_full_synch_d_out_reg_0_ (.rb(net445),
    .clk(clknet_3_4__leaf_spi_sclk),
    .d1(net157),
    .d2(net2285),
    .o1(u_dcfifo_rx_u_din_full_full_synch_d_middle_0_),
    .o2(u_dcfifo_rx_u_din_full_full_up),
    .si1(net749),
    .si2(net750),
    .ssb(net1604));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_full_latched_full_s_reg_u_dcfifo_tx_u_dout_empty_synch_d_out_reg_1_ (.rb(net442),
    .clk(clknet_3_3__leaf_spi_sclk),
    .d1(u_dcfifo_rx_u_din_full_N0),
    .d2(net2293),
    .o1(u_dcfifo_rx_u_din_full_latched_full_s),
    .o2(u_dcfifo_tx_u_dout_write_token_dn[1]),
    .si1(net751),
    .si2(net752),
    .ssb(net1605));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_din_write_tr_clk_gate_state_reg_latch (.clk(clknet_3_4__leaf_spi_sclk),
    .clkout(u_dcfifo_rx_u_din_write_tr_net652),
    .en(net134),
    .te(net753));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_write_tr_state_reg_0__u_dcfifo_rx_u_din_write_tr_state_reg_1_ (.rb(net452),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_write_tr_net652),
    .d1(net2360),
    .d2(u_dcfifo_rx_write_token[0]),
    .o1(u_dcfifo_rx_write_token[0]),
    .o2(u_dcfifo_rx_write_token[1]),
    .si1(net754),
    .si2(net755),
    .ssb(net1606));
 b15fqy00car1n02x5 u_dcfifo_rx_u_din_write_tr_state_reg_2_ (.clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_write_tr_net652),
    .d(net2290),
    .o(u_dcfifo_rx_write_token[2]),
    .psb(net452),
    .si(net756),
    .ssb(net1607));
 b15fqy00car1n02x5 u_dcfifo_rx_u_din_write_tr_state_reg_3_ (.clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_write_tr_net652),
    .d(net2307),
    .o(u_dcfifo_rx_write_token[3]),
    .psb(net452),
    .si(net757),
    .ssb(net1608));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_write_tr_state_reg_4__u_dcfifo_rx_u_din_write_tr_state_reg_5_ (.rb(net452),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_din_write_tr_net652),
    .d1(net2371),
    .d2(net2330),
    .o1(u_dcfifo_rx_write_token[4]),
    .o2(u_dcfifo_rx_write_token[5]),
    .si1(net758),
    .si2(net759),
    .ssb(net1609));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_din_write_tr_state_reg_6__u_dcfifo_rx_u_din_write_tr_state_reg_7_ (.rb(net452),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_din_write_tr_net652),
    .d1(net2355),
    .d2(u_dcfifo_rx_write_token[6]),
    .o1(u_dcfifo_rx_write_token[6]),
    .o2(u_dcfifo_rx_write_token[7]),
    .si1(net760),
    .si2(net761),
    .ssb(net1610));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_0__u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_1_ (.rb(net439),
    .clk(clknet_2_2_0_clk_i),
    .d1(u_dcfifo_rx_write_token[0]),
    .d2(net336),
    .o1(u_dcfifo_rx_u_dout_empty_synch_d_middle[0]),
    .o2(u_dcfifo_rx_u_dout_empty_synch_d_middle[1]),
    .si1(net762),
    .si2(net763),
    .ssb(net1611));
 b15fqy00car1n02x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_2_ (.clk(clknet_2_2_0_clk_i),
    .d(net333),
    .o(u_dcfifo_rx_u_dout_empty_synch_d_middle[2]),
    .psb(net449),
    .si(net764),
    .ssb(net1612));
 b15fqy00car1n02x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_3_ (.clk(clknet_2_2_0_clk_i),
    .d(net331),
    .o(u_dcfifo_rx_u_dout_empty_synch_d_middle[3]),
    .psb(net449),
    .si(net765),
    .ssb(net1613));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_4__u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_5_ (.rb(net449),
    .clk(clknet_2_2_0_clk_i),
    .d1(net330),
    .d2(net328),
    .o1(u_dcfifo_rx_u_dout_empty_synch_d_middle[4]),
    .o2(u_dcfifo_rx_u_dout_empty_synch_d_middle[5]),
    .si1(net766),
    .si2(net767),
    .ssb(net1614));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_6__u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_7_ (.rb(net449),
    .clk(clknet_2_3_0_clk_i),
    .d1(u_dcfifo_rx_write_token[6]),
    .d2(u_dcfifo_rx_write_token[7]),
    .o1(u_dcfifo_rx_u_dout_empty_synch_d_middle[6]),
    .o2(u_dcfifo_rx_u_dout_empty_synch_d_middle[7]),
    .si1(net768),
    .si2(net769),
    .ssb(net1615));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_0__u_dcfifo_rx_u_dout_empty_synch_d_out_reg_1_ (.rb(net439),
    .clk(clknet_2_2_0_clk_i),
    .d1(net2309),
    .d2(net2314),
    .o1(u_dcfifo_rx_u_dout_write_token_dn[0]),
    .o2(u_dcfifo_rx_u_dout_write_token_dn[1]),
    .si1(net770),
    .si2(net771),
    .ssb(net1616));
 b15fqy00car1n02x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_2_ (.clk(clknet_2_2_0_clk_i),
    .d(net2295),
    .o(u_dcfifo_rx_u_dout_write_token_dn[2]),
    .psb(net449),
    .si(net772),
    .ssb(net1617));
 b15fqy00car1n02x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_3_ (.clk(clknet_2_2_0_clk_i),
    .d(net2297),
    .o(u_dcfifo_rx_u_dout_write_token_dn[3]),
    .psb(net449),
    .si(net773),
    .ssb(net1618));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_4__u_dcfifo_rx_u_dout_empty_synch_d_out_reg_5_ (.rb(net449),
    .clk(clknet_2_2_0_clk_i),
    .d1(net2303),
    .d2(net2310),
    .o1(u_dcfifo_rx_u_dout_write_token_dn[4]),
    .o2(u_dcfifo_rx_u_dout_write_token_dn[5]),
    .si1(net774),
    .si2(net775),
    .ssb(net1619));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_6__u_dcfifo_rx_u_dout_empty_synch_d_out_reg_7_ (.rb(net449),
    .clk(clknet_2_3_0_clk_i),
    .d1(net2291),
    .d2(net2245),
    .o1(u_dcfifo_rx_u_dout_write_token_dn[6]),
    .o2(u_dcfifo_rx_u_dout_write_token_dn[7]),
    .si1(net776),
    .si2(net777),
    .ssb(net1620));
 b15cilb05ah1n02x3 u_dcfifo_rx_u_dout_read_tr_clk_gate_state_reg_latch (.clk(clknet_2_0_0_clk_i),
    .clkout(u_dcfifo_rx_u_dout_read_tr_net634),
    .en(n2723),
    .te(net778));
 b15fqy00car1n02x5 u_dcfifo_rx_u_dout_read_tr_state_reg_0_ (.clk(clknet_1_0__leaf_u_dcfifo_rx_u_dout_read_tr_net634),
    .d(net2327),
    .o(u_dcfifo_rx_u_dout_read_token[0]),
    .psb(net439),
    .si(net779),
    .ssb(net1621));
 b15fqy00car1n02x5 u_dcfifo_rx_u_dout_read_tr_state_reg_1_ (.clk(clknet_1_0__leaf_u_dcfifo_rx_u_dout_read_tr_net634),
    .d(u_dcfifo_rx_u_dout_read_token[0]),
    .o(u_dcfifo_rx_u_dout_read_token[1]),
    .psb(net439),
    .si(net780),
    .ssb(net1622));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_dout_read_tr_state_reg_2__u_dcfifo_rx_u_dout_read_tr_state_reg_3_ (.rb(net439),
    .clk(clknet_1_0__leaf_u_dcfifo_rx_u_dout_read_tr_net634),
    .d1(u_dcfifo_rx_u_dout_read_token[1]),
    .d2(u_dcfifo_rx_u_dout_read_token[2]),
    .o1(u_dcfifo_rx_u_dout_read_token[2]),
    .o2(u_dcfifo_rx_u_dout_read_token[3]),
    .si1(net781),
    .si2(net782),
    .ssb(net1623));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_dout_read_tr_state_reg_4__u_dcfifo_rx_u_dout_read_tr_state_reg_5_ (.rb(net439),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_dout_read_tr_net634),
    .d1(net2338),
    .d2(u_dcfifo_rx_u_dout_read_token[4]),
    .o1(u_dcfifo_rx_u_dout_read_token[4]),
    .o2(u_dcfifo_rx_u_dout_read_token[5]),
    .si1(net783),
    .si2(net784),
    .ssb(net1624));
 b15fqy203ar1n02x5 u_dcfifo_rx_u_dout_read_tr_state_reg_6__u_dcfifo_rx_u_dout_read_tr_state_reg_7_ (.rb(net439),
    .clk(clknet_1_1__leaf_u_dcfifo_rx_u_dout_read_tr_net634),
    .d1(net2362),
    .d2(net2345),
    .o1(u_dcfifo_rx_u_dout_read_token[6]),
    .o2(u_dcfifo_rx_u_dout_read_token[7]),
    .si1(net785),
    .si2(net786),
    .ssb(net1625));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_0__0_latch (.clk(clknet_2_3_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net746),
    .en(u_dcfifo_tx_u_din_buffer_N26),
    .te(net787));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_0__latch (.clk(clknet_2_1_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net741),
    .en(u_dcfifo_tx_u_din_buffer_N26),
    .te(net788));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_1__0_latch (.clk(clknet_2_3_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net736),
    .en(u_dcfifo_tx_u_din_buffer_N27),
    .te(net789));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_1__latch (.clk(clknet_2_0_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net731),
    .en(u_dcfifo_tx_u_din_buffer_N27),
    .te(net790));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_2__0_latch (.clk(clknet_2_2_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net726),
    .en(u_dcfifo_tx_u_din_buffer_N28),
    .te(net791));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_2__latch (.clk(clknet_2_0_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net721),
    .en(u_dcfifo_tx_u_din_buffer_N28),
    .te(net792));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_3__0_latch (.clk(clknet_2_2_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net716),
    .en(u_dcfifo_tx_u_din_buffer_N29),
    .te(net793));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_3__latch (.clk(clknet_2_0_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net711),
    .en(u_dcfifo_tx_u_din_buffer_N29),
    .te(net794));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_4__0_latch (.clk(clknet_2_2_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net706),
    .en(u_dcfifo_tx_u_din_buffer_N30),
    .te(net795));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_4__latch (.clk(clknet_2_0_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net701),
    .en(u_dcfifo_tx_u_din_buffer_N30),
    .te(net796));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_5__0_latch (.clk(clknet_2_3_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net696),
    .en(u_dcfifo_tx_u_din_buffer_N31),
    .te(net797));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_5__latch (.clk(clknet_2_0_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net691),
    .en(u_dcfifo_tx_u_din_buffer_N31),
    .te(net798));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_6__0_latch (.clk(clknet_2_3_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net686),
    .en(u_dcfifo_tx_u_din_buffer_N32),
    .te(net799));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_6__latch (.clk(clknet_2_0_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net681),
    .en(u_dcfifo_tx_u_din_buffer_N32),
    .te(net800));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_7__0_latch (.clk(clknet_2_2_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net676),
    .en(u_dcfifo_tx_u_din_buffer_N33),
    .te(net801));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_7__latch (.clk(clknet_2_0_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_buffer_net670),
    .en(u_dcfifo_tx_u_din_buffer_N33),
    .te(net802));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__0__u_dcfifo_tx_u_din_buffer_data_reg_0__1_ (.rb(net441),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net741),
    .d1(net435),
    .d2(net433),
    .o1(u_dcfifo_tx_u_din_buffer_data[0]),
    .o2(u_dcfifo_tx_u_din_buffer_data[1]),
    .si1(net803),
    .si2(net804),
    .ssb(net1626));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__10__u_dcfifo_tx_u_din_buffer_data_reg_0__11_ (.rb(net441),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net741),
    .d1(net413),
    .d2(net411),
    .o1(u_dcfifo_tx_u_din_buffer_data[10]),
    .o2(u_dcfifo_tx_u_din_buffer_data[11]),
    .si1(net805),
    .si2(net806),
    .ssb(net1627));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__12__u_dcfifo_tx_u_din_buffer_data_reg_0__13_ (.rb(net441),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net741),
    .d1(net409),
    .d2(net407),
    .o1(u_dcfifo_tx_u_din_buffer_data[12]),
    .o2(u_dcfifo_tx_u_din_buffer_data[13]),
    .si1(net807),
    .si2(net808),
    .ssb(net1628));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__14__u_dcfifo_tx_u_din_buffer_data_reg_0__15_ (.rb(net439),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net741),
    .d1(net405),
    .d2(net403),
    .o1(u_dcfifo_tx_u_din_buffer_data[14]),
    .o2(u_dcfifo_tx_u_din_buffer_data[15]),
    .si1(net809),
    .si2(net810),
    .ssb(net1629));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__16__u_dcfifo_tx_u_din_buffer_data_reg_0__17_ (.rb(net454),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net746),
    .d1(net401),
    .d2(net399),
    .o1(u_dcfifo_tx_u_din_buffer_data[16]),
    .o2(u_dcfifo_tx_u_din_buffer_data[17]),
    .si1(net811),
    .si2(net812),
    .ssb(net1630));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__18__u_dcfifo_tx_u_din_buffer_data_reg_0__19_ (.rb(net454),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net746),
    .d1(net397),
    .d2(net395),
    .o1(u_dcfifo_tx_u_din_buffer_data[18]),
    .o2(u_dcfifo_tx_u_din_buffer_data[19]),
    .si1(net813),
    .si2(net814),
    .ssb(net1631));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__20__u_dcfifo_tx_u_din_buffer_data_reg_0__21_ (.rb(net454),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net746),
    .d1(net392),
    .d2(net390),
    .o1(u_dcfifo_tx_u_din_buffer_data[20]),
    .o2(u_dcfifo_tx_u_din_buffer_data[21]),
    .si1(net815),
    .si2(net816),
    .ssb(net1632));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__22__u_dcfifo_tx_u_din_buffer_data_reg_0__23_ (.rb(net454),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net746),
    .d1(net389),
    .d2(net387),
    .o1(u_dcfifo_tx_u_din_buffer_data[22]),
    .o2(u_dcfifo_tx_u_din_buffer_data[23]),
    .si1(net817),
    .si2(net818),
    .ssb(net1633));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__24__u_dcfifo_tx_u_din_buffer_data_reg_0__25_ (.rb(net454),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net746),
    .d1(net385),
    .d2(net383),
    .o1(u_dcfifo_tx_u_din_buffer_data[24]),
    .o2(u_dcfifo_tx_u_din_buffer_data[25]),
    .si1(net819),
    .si2(net820),
    .ssb(net1634));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__26__u_dcfifo_tx_u_din_buffer_data_reg_0__27_ (.rb(net454),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net746),
    .d1(net381),
    .d2(net379),
    .o1(u_dcfifo_tx_u_din_buffer_data[26]),
    .o2(u_dcfifo_tx_u_din_buffer_data[27]),
    .si1(net821),
    .si2(net822),
    .ssb(net1635));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__28__u_dcfifo_tx_u_din_buffer_data_reg_0__29_ (.rb(net454),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net746),
    .d1(net377),
    .d2(net375),
    .o1(u_dcfifo_tx_u_din_buffer_data[28]),
    .o2(u_dcfifo_tx_u_din_buffer_data[29]),
    .si1(net823),
    .si2(net824),
    .ssb(net1636));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__2__u_dcfifo_tx_u_din_buffer_data_reg_0__3_ (.rb(net441),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net741),
    .d1(net431),
    .d2(net429),
    .o1(u_dcfifo_tx_u_din_buffer_data[2]),
    .o2(u_dcfifo_tx_u_din_buffer_data[3]),
    .si1(net825),
    .si2(net826),
    .ssb(net1637));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__30__u_dcfifo_tx_u_din_buffer_data_reg_0__31_ (.rb(net455),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net746),
    .d1(net373),
    .d2(net371),
    .o1(u_dcfifo_tx_u_din_buffer_data[30]),
    .o2(u_dcfifo_tx_u_din_buffer_data[31]),
    .si1(net827),
    .si2(net828),
    .ssb(net1638));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__4__u_dcfifo_tx_u_din_buffer_data_reg_0__5_ (.rb(net441),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net741),
    .d1(net425),
    .d2(net423),
    .o1(u_dcfifo_tx_u_din_buffer_data[4]),
    .o2(u_dcfifo_tx_u_din_buffer_data[5]),
    .si1(net829),
    .si2(net830),
    .ssb(net1639));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__6__u_dcfifo_tx_u_din_buffer_data_reg_0__7_ (.rb(net440),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net741),
    .d1(net420),
    .d2(net418),
    .o1(u_dcfifo_tx_u_din_buffer_data[6]),
    .o2(u_dcfifo_tx_u_din_buffer_data[7]),
    .si1(net831),
    .si2(net832),
    .ssb(net1640));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_0__8__u_dcfifo_tx_u_din_buffer_data_reg_0__9_ (.rb(net440),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net741),
    .d1(net417),
    .d2(net415),
    .o1(u_dcfifo_tx_u_din_buffer_data[8]),
    .o2(u_dcfifo_tx_u_din_buffer_data[9]),
    .si1(net833),
    .si2(net834),
    .ssb(net1641));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__0__u_dcfifo_tx_u_din_buffer_data_reg_1__1_ (.rb(net440),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net731),
    .d1(net435),
    .d2(net433),
    .o1(u_dcfifo_tx_u_din_buffer_data[32]),
    .o2(u_dcfifo_tx_u_din_buffer_data[33]),
    .si1(net835),
    .si2(net836),
    .ssb(net1642));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__10__u_dcfifo_tx_u_din_buffer_data_reg_1__11_ (.rb(net440),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net731),
    .d1(net413),
    .d2(net411),
    .o1(u_dcfifo_tx_u_din_buffer_data[42]),
    .o2(u_dcfifo_tx_u_din_buffer_data[43]),
    .si1(net837),
    .si2(net838),
    .ssb(net1643));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__12__u_dcfifo_tx_u_din_buffer_data_reg_1__13_ (.rb(net439),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net731),
    .d1(net408),
    .d2(net406),
    .o1(u_dcfifo_tx_u_din_buffer_data[44]),
    .o2(u_dcfifo_tx_u_din_buffer_data[45]),
    .si1(net839),
    .si2(net840),
    .ssb(net1644));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__14__u_dcfifo_tx_u_din_buffer_data_reg_1__15_ (.rb(net439),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net731),
    .d1(net405),
    .d2(net403),
    .o1(u_dcfifo_tx_u_din_buffer_data[46]),
    .o2(u_dcfifo_tx_u_din_buffer_data[47]),
    .si1(net841),
    .si2(net842),
    .ssb(net1645));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__16__u_dcfifo_tx_u_din_buffer_data_reg_1__17_ (.rb(net454),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net736),
    .d1(net401),
    .d2(net399),
    .o1(u_dcfifo_tx_u_din_buffer_data[48]),
    .o2(u_dcfifo_tx_u_din_buffer_data[49]),
    .si1(net843),
    .si2(net844),
    .ssb(net1646));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__18__u_dcfifo_tx_u_din_buffer_data_reg_1__19_ (.rb(net455),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net736),
    .d1(net397),
    .d2(net395),
    .o1(u_dcfifo_tx_u_din_buffer_data[50]),
    .o2(u_dcfifo_tx_u_din_buffer_data[51]),
    .si1(net845),
    .si2(net846),
    .ssb(net1647));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__20__u_dcfifo_tx_u_din_buffer_data_reg_1__21_ (.rb(net454),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net736),
    .d1(net392),
    .d2(net390),
    .o1(u_dcfifo_tx_u_din_buffer_data[52]),
    .o2(u_dcfifo_tx_u_din_buffer_data[53]),
    .si1(net847),
    .si2(net848),
    .ssb(net1648));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__22__u_dcfifo_tx_u_din_buffer_data_reg_1__23_ (.rb(net454),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net736),
    .d1(net389),
    .d2(net387),
    .o1(u_dcfifo_tx_u_din_buffer_data[54]),
    .o2(u_dcfifo_tx_u_din_buffer_data[55]),
    .si1(net849),
    .si2(net850),
    .ssb(net1649));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__24__u_dcfifo_tx_u_din_buffer_data_reg_1__25_ (.rb(net454),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net736),
    .d1(net384),
    .d2(net382),
    .o1(u_dcfifo_tx_u_din_buffer_data[56]),
    .o2(u_dcfifo_tx_u_din_buffer_data[57]),
    .si1(net851),
    .si2(net852),
    .ssb(net1650));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__26__u_dcfifo_tx_u_din_buffer_data_reg_1__27_ (.rb(net455),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net736),
    .d1(net381),
    .d2(net379),
    .o1(u_dcfifo_tx_u_din_buffer_data[58]),
    .o2(u_dcfifo_tx_u_din_buffer_data[59]),
    .si1(net853),
    .si2(net854),
    .ssb(net1651));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__28__u_dcfifo_tx_u_din_buffer_data_reg_1__29_ (.rb(net455),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net736),
    .d1(net377),
    .d2(net375),
    .o1(u_dcfifo_tx_u_din_buffer_data[60]),
    .o2(u_dcfifo_tx_u_din_buffer_data[61]),
    .si1(net855),
    .si2(net856),
    .ssb(net1652));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__2__u_dcfifo_tx_u_din_buffer_data_reg_1__3_ (.rb(net439),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net731),
    .d1(net430),
    .d2(net428),
    .o1(u_dcfifo_tx_u_din_buffer_data[34]),
    .o2(u_dcfifo_tx_u_din_buffer_data[35]),
    .si1(net857),
    .si2(net858),
    .ssb(net1653));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__30__u_dcfifo_tx_u_din_buffer_data_reg_1__31_ (.rb(net455),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net736),
    .d1(net373),
    .d2(net371),
    .o1(u_dcfifo_tx_u_din_buffer_data[62]),
    .o2(u_dcfifo_tx_u_din_buffer_data[63]),
    .si1(net859),
    .si2(net860),
    .ssb(net1654));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__4__u_dcfifo_tx_u_din_buffer_data_reg_1__5_ (.rb(net439),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net731),
    .d1(net425),
    .d2(net423),
    .o1(u_dcfifo_tx_u_din_buffer_data[36]),
    .o2(u_dcfifo_tx_u_din_buffer_data[37]),
    .si1(net861),
    .si2(net862),
    .ssb(net1655));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__6__u_dcfifo_tx_u_din_buffer_data_reg_1__7_ (.rb(net439),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net731),
    .d1(net421),
    .d2(net419),
    .o1(u_dcfifo_tx_u_din_buffer_data[38]),
    .o2(u_dcfifo_tx_u_din_buffer_data[39]),
    .si1(net863),
    .si2(net864),
    .ssb(net1656));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_1__8__u_dcfifo_tx_u_din_buffer_data_reg_1__9_ (.rb(net440),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net731),
    .d1(net417),
    .d2(net415),
    .o1(u_dcfifo_tx_u_din_buffer_data[40]),
    .o2(u_dcfifo_tx_u_din_buffer_data[41]),
    .si1(net865),
    .si2(net866),
    .ssb(net1657));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__0__u_dcfifo_tx_u_din_buffer_data_reg_2__1_ (.rb(net438),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net721),
    .d1(net434),
    .d2(net432),
    .o1(u_dcfifo_tx_u_din_buffer_data[64]),
    .o2(u_dcfifo_tx_u_din_buffer_data[65]),
    .si1(net867),
    .si2(net868),
    .ssb(net1658));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__10__u_dcfifo_tx_u_din_buffer_data_reg_2__11_ (.rb(net437),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net721),
    .d1(net412),
    .d2(net410),
    .o1(u_dcfifo_tx_u_din_buffer_data[74]),
    .o2(u_dcfifo_tx_u_din_buffer_data[75]),
    .si1(net869),
    .si2(net870),
    .ssb(net1659));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__12__u_dcfifo_tx_u_din_buffer_data_reg_2__13_ (.rb(net437),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net721),
    .d1(net409),
    .d2(net407),
    .o1(u_dcfifo_tx_u_din_buffer_data[76]),
    .o2(u_dcfifo_tx_u_din_buffer_data[77]),
    .si1(net871),
    .si2(net872),
    .ssb(net1660));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__14__u_dcfifo_tx_u_din_buffer_data_reg_2__15_ (.rb(net438),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net721),
    .d1(net405),
    .d2(net403),
    .o1(u_dcfifo_tx_u_din_buffer_data[78]),
    .o2(u_dcfifo_tx_u_din_buffer_data[79]),
    .si1(net873),
    .si2(net874),
    .ssb(net1661));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__16__u_dcfifo_tx_u_din_buffer_data_reg_2__17_ (.rb(net449),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net726),
    .d1(net400),
    .d2(net398),
    .o1(u_dcfifo_tx_u_din_buffer_data[80]),
    .o2(u_dcfifo_tx_u_din_buffer_data[81]),
    .si1(net875),
    .si2(net876),
    .ssb(net1662));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__18__u_dcfifo_tx_u_din_buffer_data_reg_2__19_ (.rb(net453),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net726),
    .d1(net396),
    .d2(net394),
    .o1(u_dcfifo_tx_u_din_buffer_data[82]),
    .o2(u_dcfifo_tx_u_din_buffer_data[83]),
    .si1(net877),
    .si2(net878),
    .ssb(net1663));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__20__u_dcfifo_tx_u_din_buffer_data_reg_2__21_ (.rb(net453),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net726),
    .d1(net392),
    .d2(net390),
    .o1(u_dcfifo_tx_u_din_buffer_data[84]),
    .o2(u_dcfifo_tx_u_din_buffer_data[85]),
    .si1(net879),
    .si2(net880),
    .ssb(net1664));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__22__u_dcfifo_tx_u_din_buffer_data_reg_2__23_ (.rb(net453),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net726),
    .d1(net388),
    .d2(net386),
    .o1(u_dcfifo_tx_u_din_buffer_data[86]),
    .o2(u_dcfifo_tx_u_din_buffer_data[87]),
    .si1(net881),
    .si2(net882),
    .ssb(net1665));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__24__u_dcfifo_tx_u_din_buffer_data_reg_2__25_ (.rb(net453),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net726),
    .d1(net384),
    .d2(net382),
    .o1(u_dcfifo_tx_u_din_buffer_data[88]),
    .o2(u_dcfifo_tx_u_din_buffer_data[89]),
    .si1(net883),
    .si2(net884),
    .ssb(net1666));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__26__u_dcfifo_tx_u_din_buffer_data_reg_2__27_ (.rb(net449),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net726),
    .d1(net380),
    .d2(net378),
    .o1(u_dcfifo_tx_u_din_buffer_data[90]),
    .o2(u_dcfifo_tx_u_din_buffer_data[91]),
    .si1(net885),
    .si2(net886),
    .ssb(net1667));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__28__u_dcfifo_tx_u_din_buffer_data_reg_2__29_ (.rb(net449),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net726),
    .d1(net376),
    .d2(net374),
    .o1(u_dcfifo_tx_u_din_buffer_data[92]),
    .o2(u_dcfifo_tx_u_din_buffer_data[93]),
    .si1(net887),
    .si2(net888),
    .ssb(net1668));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__2__u_dcfifo_tx_u_din_buffer_data_reg_2__3_ (.rb(net438),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net721),
    .d1(net431),
    .d2(net429),
    .o1(u_dcfifo_tx_u_din_buffer_data[66]),
    .o2(u_dcfifo_tx_u_din_buffer_data[67]),
    .si1(net889),
    .si2(net890),
    .ssb(net1669));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__30__u_dcfifo_tx_u_din_buffer_data_reg_2__31_ (.rb(net453),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net726),
    .d1(net373),
    .d2(net371),
    .o1(u_dcfifo_tx_u_din_buffer_data[94]),
    .o2(u_dcfifo_tx_u_din_buffer_data[95]),
    .si1(net891),
    .si2(net892),
    .ssb(net1670));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__4__u_dcfifo_tx_u_din_buffer_data_reg_2__5_ (.rb(net438),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net721),
    .d1(net424),
    .d2(net422),
    .o1(u_dcfifo_tx_u_din_buffer_data[68]),
    .o2(u_dcfifo_tx_u_din_buffer_data[69]),
    .si1(net893),
    .si2(net894),
    .ssb(net1671));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__6__u_dcfifo_tx_u_din_buffer_data_reg_2__7_ (.rb(net437),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net721),
    .d1(net420),
    .d2(net418),
    .o1(u_dcfifo_tx_u_din_buffer_data[70]),
    .o2(u_dcfifo_tx_u_din_buffer_data[71]),
    .si1(net895),
    .si2(net896),
    .ssb(net1672));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_2__8__u_dcfifo_tx_u_din_buffer_data_reg_2__9_ (.rb(net437),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net721),
    .d1(net416),
    .d2(net414),
    .o1(u_dcfifo_tx_u_din_buffer_data[72]),
    .o2(u_dcfifo_tx_u_din_buffer_data[73]),
    .si1(net897),
    .si2(net898),
    .ssb(net1673));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__0__u_dcfifo_tx_u_din_buffer_data_reg_3__1_ (.rb(net436),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net711),
    .d1(net434),
    .d2(net432),
    .o1(u_dcfifo_tx_u_din_buffer_data[96]),
    .o2(u_dcfifo_tx_u_din_buffer_data[97]),
    .si1(net899),
    .si2(net900),
    .ssb(net1674));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__10__u_dcfifo_tx_u_din_buffer_data_reg_3__11_ (.rb(net436),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net711),
    .d1(net412),
    .d2(net410),
    .o1(u_dcfifo_tx_u_din_buffer_data[106]),
    .o2(u_dcfifo_tx_u_din_buffer_data[107]),
    .si1(net901),
    .si2(net902),
    .ssb(net1675));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__12__u_dcfifo_tx_u_din_buffer_data_reg_3__13_ (.rb(net437),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net711),
    .d1(net408),
    .d2(net406),
    .o1(u_dcfifo_tx_u_din_buffer_data[108]),
    .o2(u_dcfifo_tx_u_din_buffer_data[109]),
    .si1(net903),
    .si2(net904),
    .ssb(net1676));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__14__u_dcfifo_tx_u_din_buffer_data_reg_3__15_ (.rb(net437),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net711),
    .d1(net404),
    .d2(net402),
    .o1(u_dcfifo_tx_u_din_buffer_data[110]),
    .o2(u_dcfifo_tx_u_din_buffer_data[111]),
    .si1(net905),
    .si2(net906),
    .ssb(net1677));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__16__u_dcfifo_tx_u_din_buffer_data_reg_3__17_ (.rb(net453),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net716),
    .d1(net401),
    .d2(net399),
    .o1(u_dcfifo_tx_u_din_buffer_data[112]),
    .o2(u_dcfifo_tx_u_din_buffer_data[113]),
    .si1(net907),
    .si2(net908),
    .ssb(net1678));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__18__u_dcfifo_tx_u_din_buffer_data_reg_3__19_ (.rb(net453),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net716),
    .d1(net396),
    .d2(net394),
    .o1(u_dcfifo_tx_u_din_buffer_data[114]),
    .o2(u_dcfifo_tx_u_din_buffer_data[115]),
    .si1(net909),
    .si2(net910),
    .ssb(net1679));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__20__u_dcfifo_tx_u_din_buffer_data_reg_3__21_ (.rb(net453),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net716),
    .d1(net392),
    .d2(net390),
    .o1(u_dcfifo_tx_u_din_buffer_data[116]),
    .o2(u_dcfifo_tx_u_din_buffer_data[117]),
    .si1(net911),
    .si2(net912),
    .ssb(net1680));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__22__u_dcfifo_tx_u_din_buffer_data_reg_3__23_ (.rb(net453),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net716),
    .d1(net388),
    .d2(net386),
    .o1(u_dcfifo_tx_u_din_buffer_data[118]),
    .o2(u_dcfifo_tx_u_din_buffer_data[119]),
    .si1(net913),
    .si2(net914),
    .ssb(net1681));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__24__u_dcfifo_tx_u_din_buffer_data_reg_3__25_ (.rb(net453),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net716),
    .d1(net384),
    .d2(net382),
    .o1(u_dcfifo_tx_u_din_buffer_data[120]),
    .o2(u_dcfifo_tx_u_din_buffer_data[121]),
    .si1(net915),
    .si2(net916),
    .ssb(net1682));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__26__u_dcfifo_tx_u_din_buffer_data_reg_3__27_ (.rb(net453),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net716),
    .d1(net381),
    .d2(net379),
    .o1(u_dcfifo_tx_u_din_buffer_data[122]),
    .o2(u_dcfifo_tx_u_din_buffer_data[123]),
    .si1(net917),
    .si2(net918),
    .ssb(net1683));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__28__u_dcfifo_tx_u_din_buffer_data_reg_3__29_ (.rb(net453),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net716),
    .d1(net377),
    .d2(net375),
    .o1(u_dcfifo_tx_u_din_buffer_data[124]),
    .o2(u_dcfifo_tx_u_din_buffer_data[125]),
    .si1(net919),
    .si2(net920),
    .ssb(net1684));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__2__u_dcfifo_tx_u_din_buffer_data_reg_3__3_ (.rb(net436),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net711),
    .d1(net430),
    .d2(net428),
    .o1(u_dcfifo_tx_u_din_buffer_data[98]),
    .o2(u_dcfifo_tx_u_din_buffer_data[99]),
    .si1(net921),
    .si2(net922),
    .ssb(net1685));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__30__u_dcfifo_tx_u_din_buffer_data_reg_3__31_ (.rb(net453),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net716),
    .d1(net373),
    .d2(net371),
    .o1(u_dcfifo_tx_u_din_buffer_data[126]),
    .o2(u_dcfifo_tx_u_din_buffer_data[127]),
    .si1(net923),
    .si2(net924),
    .ssb(net1686));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__4__u_dcfifo_tx_u_din_buffer_data_reg_3__5_ (.rb(net436),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net711),
    .d1(net424),
    .d2(net422),
    .o1(u_dcfifo_tx_u_din_buffer_data[100]),
    .o2(u_dcfifo_tx_u_din_buffer_data[101]),
    .si1(net925),
    .si2(net926),
    .ssb(net1687));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__6__u_dcfifo_tx_u_din_buffer_data_reg_3__7_ (.rb(net437),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net711),
    .d1(net421),
    .d2(net419),
    .o1(u_dcfifo_tx_u_din_buffer_data[102]),
    .o2(u_dcfifo_tx_u_din_buffer_data[103]),
    .si1(net927),
    .si2(net928),
    .ssb(net1688));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_3__8__u_dcfifo_tx_u_din_buffer_data_reg_3__9_ (.rb(net437),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net711),
    .d1(net416),
    .d2(net414),
    .o1(u_dcfifo_tx_u_din_buffer_data[104]),
    .o2(u_dcfifo_tx_u_din_buffer_data[105]),
    .si1(net929),
    .si2(net930),
    .ssb(net1689));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__0__u_dcfifo_tx_u_din_buffer_data_reg_4__1_ (.rb(net436),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net701),
    .d1(net434),
    .d2(net432),
    .o1(u_dcfifo_tx_u_din_buffer_data[128]),
    .o2(u_dcfifo_tx_u_din_buffer_data[129]),
    .si1(net931),
    .si2(net932),
    .ssb(net1690));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__10__u_dcfifo_tx_u_din_buffer_data_reg_4__11_ (.rb(net438),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net701),
    .d1(net412),
    .d2(net410),
    .o1(u_dcfifo_tx_u_din_buffer_data[138]),
    .o2(u_dcfifo_tx_u_din_buffer_data[139]),
    .si1(net933),
    .si2(net934),
    .ssb(net1691));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__12__u_dcfifo_tx_u_din_buffer_data_reg_4__13_ (.rb(net436),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net701),
    .d1(net409),
    .d2(net407),
    .o1(u_dcfifo_tx_u_din_buffer_data[140]),
    .o2(u_dcfifo_tx_u_din_buffer_data[141]),
    .si1(net935),
    .si2(net936),
    .ssb(net1692));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__14__u_dcfifo_tx_u_din_buffer_data_reg_4__15_ (.rb(net438),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net701),
    .d1(net405),
    .d2(net403),
    .o1(u_dcfifo_tx_u_din_buffer_data[142]),
    .o2(u_dcfifo_tx_u_din_buffer_data[143]),
    .si1(net937),
    .si2(net938),
    .ssb(net1693));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__16__u_dcfifo_tx_u_din_buffer_data_reg_4__17_ (.rb(net449),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net706),
    .d1(net400),
    .d2(net398),
    .o1(u_dcfifo_tx_u_din_buffer_data[144]),
    .o2(u_dcfifo_tx_u_din_buffer_data[145]),
    .si1(net939),
    .si2(net940),
    .ssb(net1694));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__18__u_dcfifo_tx_u_din_buffer_data_reg_4__19_ (.rb(net449),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net706),
    .d1(net396),
    .d2(net394),
    .o1(u_dcfifo_tx_u_din_buffer_data[146]),
    .o2(u_dcfifo_tx_u_din_buffer_data[147]),
    .si1(net941),
    .si2(net942),
    .ssb(net1695));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__20__u_dcfifo_tx_u_din_buffer_data_reg_4__21_ (.rb(net450),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net706),
    .d1(net393),
    .d2(net391),
    .o1(u_dcfifo_tx_u_din_buffer_data[148]),
    .o2(u_dcfifo_tx_u_din_buffer_data[149]),
    .si1(net943),
    .si2(net944),
    .ssb(net1696));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__22__u_dcfifo_tx_u_din_buffer_data_reg_4__23_ (.rb(net450),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net706),
    .d1(net388),
    .d2(net386),
    .o1(u_dcfifo_tx_u_din_buffer_data[150]),
    .o2(u_dcfifo_tx_u_din_buffer_data[151]),
    .si1(net945),
    .si2(net946),
    .ssb(net1697));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__24__u_dcfifo_tx_u_din_buffer_data_reg_4__25_ (.rb(net450),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net706),
    .d1(net384),
    .d2(net382),
    .o1(u_dcfifo_tx_u_din_buffer_data[152]),
    .o2(u_dcfifo_tx_u_din_buffer_data[153]),
    .si1(net947),
    .si2(net948),
    .ssb(net1698));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__26__u_dcfifo_tx_u_din_buffer_data_reg_4__27_ (.rb(net450),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net706),
    .d1(net380),
    .d2(net378),
    .o1(u_dcfifo_tx_u_din_buffer_data[154]),
    .o2(u_dcfifo_tx_u_din_buffer_data[155]),
    .si1(net949),
    .si2(net950),
    .ssb(net1699));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__28__u_dcfifo_tx_u_din_buffer_data_reg_4__29_ (.rb(net450),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net706),
    .d1(net376),
    .d2(net374),
    .o1(u_dcfifo_tx_u_din_buffer_data[156]),
    .o2(u_dcfifo_tx_u_din_buffer_data[157]),
    .si1(net951),
    .si2(net952),
    .ssb(net1700));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__2__u_dcfifo_tx_u_din_buffer_data_reg_4__3_ (.rb(net436),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net701),
    .d1(net431),
    .d2(net429),
    .o1(u_dcfifo_tx_u_din_buffer_data[130]),
    .o2(u_dcfifo_tx_u_din_buffer_data[131]),
    .si1(net953),
    .si2(net954),
    .ssb(net1701));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__30__u_dcfifo_tx_u_din_buffer_data_reg_4__31_ (.rb(net450),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net706),
    .d1(net372),
    .d2(net370),
    .o1(u_dcfifo_tx_u_din_buffer_data[158]),
    .o2(u_dcfifo_tx_u_din_buffer_data[159]),
    .si1(net955),
    .si2(net956),
    .ssb(net1702));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__4__u_dcfifo_tx_u_din_buffer_data_reg_4__5_ (.rb(net438),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net701),
    .d1(net424),
    .d2(net422),
    .o1(u_dcfifo_tx_u_din_buffer_data[132]),
    .o2(u_dcfifo_tx_u_din_buffer_data[133]),
    .si1(net957),
    .si2(net958),
    .ssb(net1703));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__6__u_dcfifo_tx_u_din_buffer_data_reg_4__7_ (.rb(net436),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net701),
    .d1(net420),
    .d2(net418),
    .o1(u_dcfifo_tx_u_din_buffer_data[134]),
    .o2(u_dcfifo_tx_u_din_buffer_data[135]),
    .si1(net959),
    .si2(net960),
    .ssb(net1704));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_4__8__u_dcfifo_tx_u_din_buffer_data_reg_4__9_ (.rb(net438),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net701),
    .d1(net416),
    .d2(net414),
    .o1(u_dcfifo_tx_u_din_buffer_data[136]),
    .o2(u_dcfifo_tx_u_din_buffer_data[137]),
    .si1(net961),
    .si2(net962),
    .ssb(net1705));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__0__u_dcfifo_tx_u_din_buffer_data_reg_5__1_ (.rb(net436),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net691),
    .d1(net434),
    .d2(net432),
    .o1(u_dcfifo_tx_u_din_buffer_data[160]),
    .o2(u_dcfifo_tx_u_din_buffer_data[161]),
    .si1(net963),
    .si2(net964),
    .ssb(net1706));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__10__u_dcfifo_tx_u_din_buffer_data_reg_5__11_ (.rb(net436),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net691),
    .d1(net412),
    .d2(net410),
    .o1(u_dcfifo_tx_u_din_buffer_data[170]),
    .o2(u_dcfifo_tx_u_din_buffer_data[171]),
    .si1(net965),
    .si2(net966),
    .ssb(net1707));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__12__u_dcfifo_tx_u_din_buffer_data_reg_5__13_ (.rb(net436),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net691),
    .d1(net409),
    .d2(net407),
    .o1(u_dcfifo_tx_u_din_buffer_data[172]),
    .o2(u_dcfifo_tx_u_din_buffer_data[173]),
    .si1(net967),
    .si2(net968),
    .ssb(net1708));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__14__u_dcfifo_tx_u_din_buffer_data_reg_5__15_ (.rb(net436),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net691),
    .d1(net404),
    .d2(net402),
    .o1(u_dcfifo_tx_u_din_buffer_data[174]),
    .o2(u_dcfifo_tx_u_din_buffer_data[175]),
    .si1(net969),
    .si2(net970),
    .ssb(net1709));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__16__u_dcfifo_tx_u_din_buffer_data_reg_5__17_ (.rb(net451),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net696),
    .d1(net400),
    .d2(net398),
    .o1(u_dcfifo_tx_u_din_buffer_data[176]),
    .o2(u_dcfifo_tx_u_din_buffer_data[177]),
    .si1(net971),
    .si2(net972),
    .ssb(net1710));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__18__u_dcfifo_tx_u_din_buffer_data_reg_5__19_ (.rb(net451),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net696),
    .d1(net396),
    .d2(net394),
    .o1(u_dcfifo_tx_u_din_buffer_data[178]),
    .o2(u_dcfifo_tx_u_din_buffer_data[179]),
    .si1(net973),
    .si2(net974),
    .ssb(net1711));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__20__u_dcfifo_tx_u_din_buffer_data_reg_5__21_ (.rb(net450),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net696),
    .d1(net393),
    .d2(net391),
    .o1(u_dcfifo_tx_u_din_buffer_data[180]),
    .o2(u_dcfifo_tx_u_din_buffer_data[181]),
    .si1(net975),
    .si2(net976),
    .ssb(net1712));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__22__u_dcfifo_tx_u_din_buffer_data_reg_5__23_ (.rb(net451),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net696),
    .d1(net389),
    .d2(net387),
    .o1(u_dcfifo_tx_u_din_buffer_data[182]),
    .o2(u_dcfifo_tx_u_din_buffer_data[183]),
    .si1(net977),
    .si2(net978),
    .ssb(net1713));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__24__u_dcfifo_tx_u_din_buffer_data_reg_5__25_ (.rb(net450),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net696),
    .d1(net385),
    .d2(net383),
    .o1(u_dcfifo_tx_u_din_buffer_data[184]),
    .o2(u_dcfifo_tx_u_din_buffer_data[185]),
    .si1(net979),
    .si2(net980),
    .ssb(net1714));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__26__u_dcfifo_tx_u_din_buffer_data_reg_5__27_ (.rb(net450),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net696),
    .d1(net380),
    .d2(net378),
    .o1(u_dcfifo_tx_u_din_buffer_data[186]),
    .o2(u_dcfifo_tx_u_din_buffer_data[187]),
    .si1(net981),
    .si2(net982),
    .ssb(net1715));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__28__u_dcfifo_tx_u_din_buffer_data_reg_5__29_ (.rb(net450),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net696),
    .d1(net376),
    .d2(net374),
    .o1(u_dcfifo_tx_u_din_buffer_data[188]),
    .o2(u_dcfifo_tx_u_din_buffer_data[189]),
    .si1(net983),
    .si2(net984),
    .ssb(net1716));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__2__u_dcfifo_tx_u_din_buffer_data_reg_5__3_ (.rb(net436),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net691),
    .d1(net431),
    .d2(net429),
    .o1(u_dcfifo_tx_u_din_buffer_data[162]),
    .o2(u_dcfifo_tx_u_din_buffer_data[163]),
    .si1(net985),
    .si2(net986),
    .ssb(net1717));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__30__u_dcfifo_tx_u_din_buffer_data_reg_5__31_ (.rb(net450),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net696),
    .d1(net372),
    .d2(net370),
    .o1(u_dcfifo_tx_u_din_buffer_data[190]),
    .o2(u_dcfifo_tx_u_din_buffer_data[191]),
    .si1(net987),
    .si2(net988),
    .ssb(net1718));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__4__u_dcfifo_tx_u_din_buffer_data_reg_5__5_ (.rb(net436),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net691),
    .d1(net424),
    .d2(net422),
    .o1(u_dcfifo_tx_u_din_buffer_data[164]),
    .o2(u_dcfifo_tx_u_din_buffer_data[165]),
    .si1(net989),
    .si2(net990),
    .ssb(net1719));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__6__u_dcfifo_tx_u_din_buffer_data_reg_5__7_ (.rb(net436),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net691),
    .d1(net420),
    .d2(net418),
    .o1(u_dcfifo_tx_u_din_buffer_data[166]),
    .o2(u_dcfifo_tx_u_din_buffer_data[167]),
    .si1(net991),
    .si2(net992),
    .ssb(net1720));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_5__8__u_dcfifo_tx_u_din_buffer_data_reg_5__9_ (.rb(net436),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net691),
    .d1(net416),
    .d2(net414),
    .o1(u_dcfifo_tx_u_din_buffer_data[168]),
    .o2(u_dcfifo_tx_u_din_buffer_data[169]),
    .si1(net993),
    .si2(net994),
    .ssb(net1721));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__0__u_dcfifo_tx_u_din_buffer_data_reg_6__1_ (.rb(net440),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net681),
    .d1(net435),
    .d2(net433),
    .o1(u_dcfifo_tx_u_din_buffer_data[192]),
    .o2(u_dcfifo_tx_u_din_buffer_data[193]),
    .si1(net995),
    .si2(net996),
    .ssb(net1722));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__10__u_dcfifo_tx_u_din_buffer_data_reg_6__11_ (.rb(net440),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net681),
    .d1(net413),
    .d2(net411),
    .o1(u_dcfifo_tx_u_din_buffer_data[202]),
    .o2(u_dcfifo_tx_u_din_buffer_data[203]),
    .si1(net997),
    .si2(net998),
    .ssb(net1723));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__12__u_dcfifo_tx_u_din_buffer_data_reg_6__13_ (.rb(net440),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net681),
    .d1(net408),
    .d2(net406),
    .o1(u_dcfifo_tx_u_din_buffer_data[204]),
    .o2(u_dcfifo_tx_u_din_buffer_data[205]),
    .si1(net999),
    .si2(net1000),
    .ssb(net1724));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__14__u_dcfifo_tx_u_din_buffer_data_reg_6__15_ (.rb(net440),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net681),
    .d1(net404),
    .d2(net402),
    .o1(u_dcfifo_tx_u_din_buffer_data[206]),
    .o2(u_dcfifo_tx_u_din_buffer_data[207]),
    .si1(net1001),
    .si2(net1002),
    .ssb(net1725));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__16__u_dcfifo_tx_u_din_buffer_data_reg_6__17_ (.rb(net454),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net686),
    .d1(net401),
    .d2(net399),
    .o1(u_dcfifo_tx_u_din_buffer_data[208]),
    .o2(u_dcfifo_tx_u_din_buffer_data[209]),
    .si1(net1003),
    .si2(net1004),
    .ssb(net1726));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__18__u_dcfifo_tx_u_din_buffer_data_reg_6__19_ (.rb(net451),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net686),
    .d1(net397),
    .d2(net395),
    .o1(u_dcfifo_tx_u_din_buffer_data[210]),
    .o2(u_dcfifo_tx_u_din_buffer_data[211]),
    .si1(net1005),
    .si2(net1006),
    .ssb(net1727));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__20__u_dcfifo_tx_u_din_buffer_data_reg_6__21_ (.rb(net454),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net686),
    .d1(net393),
    .d2(net391),
    .o1(u_dcfifo_tx_u_din_buffer_data[212]),
    .o2(u_dcfifo_tx_u_din_buffer_data[213]),
    .si1(net1007),
    .si2(net1008),
    .ssb(net1728));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__22__u_dcfifo_tx_u_din_buffer_data_reg_6__23_ (.rb(net451),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net686),
    .d1(net389),
    .d2(net387),
    .o1(u_dcfifo_tx_u_din_buffer_data[214]),
    .o2(u_dcfifo_tx_u_din_buffer_data[215]),
    .si1(net1009),
    .si2(net1010),
    .ssb(net1729));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__24__u_dcfifo_tx_u_din_buffer_data_reg_6__25_ (.rb(net454),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net686),
    .d1(net385),
    .d2(net383),
    .o1(u_dcfifo_tx_u_din_buffer_data[216]),
    .o2(u_dcfifo_tx_u_din_buffer_data[217]),
    .si1(net1011),
    .si2(net1012),
    .ssb(net1730));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__26__u_dcfifo_tx_u_din_buffer_data_reg_6__27_ (.rb(net454),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net686),
    .d1(net380),
    .d2(net378),
    .o1(u_dcfifo_tx_u_din_buffer_data[218]),
    .o2(u_dcfifo_tx_u_din_buffer_data[219]),
    .si1(net1013),
    .si2(net1014),
    .ssb(net1731));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__28__u_dcfifo_tx_u_din_buffer_data_reg_6__29_ (.rb(net451),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net686),
    .d1(net376),
    .d2(net374),
    .o1(u_dcfifo_tx_u_din_buffer_data[220]),
    .o2(u_dcfifo_tx_u_din_buffer_data[221]),
    .si1(net1015),
    .si2(net1016),
    .ssb(net1732));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__2__u_dcfifo_tx_u_din_buffer_data_reg_6__3_ (.rb(net437),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net681),
    .d1(net430),
    .d2(net428),
    .o1(u_dcfifo_tx_u_din_buffer_data[194]),
    .o2(u_dcfifo_tx_u_din_buffer_data[195]),
    .si1(net1017),
    .si2(net1018),
    .ssb(net1733));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__30__u_dcfifo_tx_u_din_buffer_data_reg_6__31_ (.rb(net454),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net686),
    .d1(net372),
    .d2(net370),
    .o1(u_dcfifo_tx_u_din_buffer_data[222]),
    .o2(u_dcfifo_tx_u_din_buffer_data[223]),
    .si1(net1019),
    .si2(net1020),
    .ssb(net1734));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__4__u_dcfifo_tx_u_din_buffer_data_reg_6__5_ (.rb(net437),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net681),
    .d1(net425),
    .d2(net423),
    .o1(u_dcfifo_tx_u_din_buffer_data[196]),
    .o2(u_dcfifo_tx_u_din_buffer_data[197]),
    .si1(net1021),
    .si2(net1022),
    .ssb(net1735));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__6__u_dcfifo_tx_u_din_buffer_data_reg_6__7_ (.rb(net437),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net681),
    .d1(net421),
    .d2(net419),
    .o1(u_dcfifo_tx_u_din_buffer_data[198]),
    .o2(u_dcfifo_tx_u_din_buffer_data[199]),
    .si1(net1023),
    .si2(net1024),
    .ssb(net1736));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_6__8__u_dcfifo_tx_u_din_buffer_data_reg_6__9_ (.rb(net437),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net681),
    .d1(net416),
    .d2(net414),
    .o1(u_dcfifo_tx_u_din_buffer_data[200]),
    .o2(u_dcfifo_tx_u_din_buffer_data[201]),
    .si1(net1025),
    .si2(net1026),
    .ssb(net1737));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__0__u_dcfifo_tx_u_din_buffer_data_reg_7__1_ (.rb(net440),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net670),
    .d1(net435),
    .d2(net433),
    .o1(u_dcfifo_tx_u_din_buffer_data[224]),
    .o2(u_dcfifo_tx_u_din_buffer_data[225]),
    .si1(net1027),
    .si2(net1028),
    .ssb(net1738));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__10__u_dcfifo_tx_u_din_buffer_data_reg_7__11_ (.rb(net440),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net670),
    .d1(net413),
    .d2(net411),
    .o1(u_dcfifo_tx_u_din_buffer_data[234]),
    .o2(u_dcfifo_tx_u_din_buffer_data[235]),
    .si1(net1029),
    .si2(net1030),
    .ssb(net1739));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__12__u_dcfifo_tx_u_din_buffer_data_reg_7__13_ (.rb(net440),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net670),
    .d1(net408),
    .d2(net406),
    .o1(u_dcfifo_tx_u_din_buffer_data[236]),
    .o2(u_dcfifo_tx_u_din_buffer_data[237]),
    .si1(net1031),
    .si2(net1032),
    .ssb(net1740));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__14__u_dcfifo_tx_u_din_buffer_data_reg_7__15_ (.rb(net439),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net670),
    .d1(net404),
    .d2(net402),
    .o1(u_dcfifo_tx_u_din_buffer_data[238]),
    .o2(u_dcfifo_tx_u_din_buffer_data[239]),
    .si1(net1033),
    .si2(net1034),
    .ssb(net1741));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__16__u_dcfifo_tx_u_din_buffer_data_reg_7__17_ (.rb(net453),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net676),
    .d1(net401),
    .d2(net399),
    .o1(u_dcfifo_tx_u_din_buffer_data[240]),
    .o2(u_dcfifo_tx_u_din_buffer_data[241]),
    .si1(net1035),
    .si2(net1036),
    .ssb(net1742));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__18__u_dcfifo_tx_u_din_buffer_data_reg_7__19_ (.rb(net453),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net676),
    .d1(net397),
    .d2(net395),
    .o1(u_dcfifo_tx_u_din_buffer_data[242]),
    .o2(u_dcfifo_tx_u_din_buffer_data[243]),
    .si1(net1037),
    .si2(net1038),
    .ssb(net1743));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__20__u_dcfifo_tx_u_din_buffer_data_reg_7__21_ (.rb(net453),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net676),
    .d1(net392),
    .d2(net390),
    .o1(u_dcfifo_tx_u_din_buffer_data[244]),
    .o2(u_dcfifo_tx_u_din_buffer_data[245]),
    .si1(net1039),
    .si2(net1040),
    .ssb(net1744));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__22__u_dcfifo_tx_u_din_buffer_data_reg_7__23_ (.rb(net456),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net676),
    .d1(net388),
    .d2(net386),
    .o1(u_dcfifo_tx_u_din_buffer_data[246]),
    .o2(u_dcfifo_tx_u_din_buffer_data[247]),
    .si1(net1041),
    .si2(net1042),
    .ssb(net1745));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__24__u_dcfifo_tx_u_din_buffer_data_reg_7__25_ (.rb(net456),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net676),
    .d1(net384),
    .d2(net382),
    .o1(u_dcfifo_tx_u_din_buffer_data[248]),
    .o2(u_dcfifo_tx_u_din_buffer_data[249]),
    .si1(net1043),
    .si2(net1044),
    .ssb(net1746));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__26__u_dcfifo_tx_u_din_buffer_data_reg_7__27_ (.rb(net456),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net676),
    .d1(net381),
    .d2(net379),
    .o1(u_dcfifo_tx_u_din_buffer_data[250]),
    .o2(u_dcfifo_tx_u_din_buffer_data[251]),
    .si1(net1045),
    .si2(net1046),
    .ssb(net1747));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__28__u_dcfifo_tx_u_din_buffer_data_reg_7__29_ (.rb(net456),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net676),
    .d1(net377),
    .d2(net375),
    .o1(u_dcfifo_tx_u_din_buffer_data[252]),
    .o2(u_dcfifo_tx_u_din_buffer_data[253]),
    .si1(net1047),
    .si2(net1048),
    .ssb(net1748));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__2__u_dcfifo_tx_u_din_buffer_data_reg_7__3_ (.rb(net440),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net670),
    .d1(net430),
    .d2(net428),
    .o1(u_dcfifo_tx_u_din_buffer_data[226]),
    .o2(u_dcfifo_tx_u_din_buffer_data[227]),
    .si1(net1049),
    .si2(net1050),
    .ssb(net1749));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__30__u_dcfifo_tx_u_din_buffer_data_reg_7__31_ (.rb(net456),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net676),
    .d1(net373),
    .d2(net371),
    .o1(u_dcfifo_tx_u_din_buffer_data[254]),
    .o2(u_dcfifo_tx_u_din_buffer_data[255]),
    .si1(net1051),
    .si2(net1052),
    .ssb(net1750));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__4__u_dcfifo_tx_u_din_buffer_data_reg_7__5_ (.rb(net439),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net670),
    .d1(net425),
    .d2(net423),
    .o1(u_dcfifo_tx_u_din_buffer_data[228]),
    .o2(u_dcfifo_tx_u_din_buffer_data[229]),
    .si1(net1053),
    .si2(net1054),
    .ssb(net1751));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__6__u_dcfifo_tx_u_din_buffer_data_reg_7__7_ (.rb(net440),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net670),
    .d1(net421),
    .d2(net419),
    .o1(u_dcfifo_tx_u_din_buffer_data[230]),
    .o2(u_dcfifo_tx_u_din_buffer_data[231]),
    .si1(net1055),
    .si2(net1056),
    .ssb(net1752));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_buffer_data_reg_7__8__u_dcfifo_tx_u_din_buffer_data_reg_7__9_ (.rb(net439),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net670),
    .d1(net417),
    .d2(net415),
    .o1(u_dcfifo_tx_u_din_buffer_data[232]),
    .o2(u_dcfifo_tx_u_din_buffer_data[233]),
    .si1(net1057),
    .si2(net1058),
    .ssb(net1753));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_full_full_synch_d_middle_reg_0__u_dcfifo_tx_u_din_full_full_synch_d_out_reg_0_ (.rb(net441),
    .clk(clknet_2_1_0_clk_i),
    .d1(u_dcfifo_tx_u_din_full_full_dn),
    .d2(net2284),
    .o1(u_dcfifo_tx_u_din_full_full_synch_d_middle_0_),
    .o2(u_dcfifo_tx_u_din_full_full_up),
    .si1(net1059),
    .si2(net1060),
    .ssb(net1754));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_full_latched_full_s_reg_u_spi_device_tlul_plug_state_reg_0_ (.rb(net438),
    .clk(clknet_2_1_0_clk_i),
    .d1(u_dcfifo_tx_u_din_full_N0),
    .d2(u_spi_device_tlul_plug_state_next[0]),
    .o1(u_dcfifo_tx_u_din_full_latched_full_s),
    .o2(u_spi_device_tlul_plug_state[0]),
    .si1(net1061),
    .si2(net1062),
    .ssb(net1755));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_din_write_tr_clk_gate_state_reg_latch (.clk(clknet_2_1_0_clk_i),
    .clkout(u_dcfifo_tx_u_din_write_tr_net652),
    .en(u_dcfifo_tx_u_din_write_enable),
    .te(net1063));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_write_tr_state_reg_0__u_dcfifo_tx_u_din_write_tr_state_reg_1_ (.rb(net438),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_write_tr_net652),
    .d1(u_dcfifo_tx_write_token[7]),
    .d2(net2308),
    .o1(u_dcfifo_tx_write_token[0]),
    .o2(u_dcfifo_tx_write_token[1]),
    .si1(net1064),
    .si2(net1065),
    .ssb(net1756));
 b15fqy00car1n02x5 u_dcfifo_tx_u_din_write_tr_state_reg_2_ (.clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_write_tr_net652),
    .d(net2304),
    .o(u_dcfifo_tx_write_token[2]),
    .psb(net438),
    .si(net1066),
    .ssb(net1757));
 b15fqy00car1n02x5 u_dcfifo_tx_u_din_write_tr_state_reg_3_ (.clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_write_tr_net652),
    .d(net2306),
    .o(u_dcfifo_tx_write_token[3]),
    .psb(net438),
    .si(net1067),
    .ssb(net1758));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_write_tr_state_reg_4__u_dcfifo_tx_u_din_write_tr_state_reg_5_ (.rb(net438),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_din_write_tr_net652),
    .d1(u_dcfifo_tx_write_token[3]),
    .d2(u_dcfifo_tx_write_token[4]),
    .o1(u_dcfifo_tx_write_token[4]),
    .o2(u_dcfifo_tx_write_token[5]),
    .si1(net1068),
    .si2(net1069),
    .ssb(net1759));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_din_write_tr_state_reg_6__u_dcfifo_tx_u_din_write_tr_state_reg_7_ (.rb(net438),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_din_write_tr_net652),
    .d1(net2356),
    .d2(net2311),
    .o1(u_dcfifo_tx_write_token[6]),
    .o2(u_dcfifo_tx_write_token[7]),
    .si1(net1070),
    .si2(net1071),
    .ssb(net1760));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_0__u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_1_ (.rb(net442),
    .clk(clknet_3_0__leaf_spi_sclk),
    .d1(net323),
    .d2(net321),
    .o1(u_dcfifo_tx_u_dout_empty_synch_d_middle[0]),
    .o2(u_dcfifo_tx_u_dout_empty_synch_d_middle[1]),
    .si1(net1072),
    .si2(net1073),
    .ssb(net1761));
 b15fqy00car1n02x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_2_ (.clk(clknet_3_2__leaf_spi_sclk),
    .d(net319),
    .o(u_dcfifo_tx_u_dout_empty_synch_d_middle[2]),
    .psb(net442),
    .si(net1074),
    .ssb(net1762));
 b15fqy00car1n02x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_3_ (.clk(clknet_3_0__leaf_spi_sclk),
    .d(net317),
    .o(u_dcfifo_tx_u_dout_empty_synch_d_middle[3]),
    .psb(net442),
    .si(net1075),
    .ssb(net1763));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_4__u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_5_ (.rb(net442),
    .clk(clknet_3_3__leaf_spi_sclk),
    .d1(net315),
    .d2(net313),
    .o1(u_dcfifo_tx_u_dout_empty_synch_d_middle[4]),
    .o2(u_dcfifo_tx_u_dout_empty_synch_d_middle[5]),
    .si1(net1076),
    .si2(net1077),
    .ssb(net1764));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_6__u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_7_ (.rb(net442),
    .clk(clknet_3_2__leaf_spi_sclk),
    .d1(net310),
    .d2(net308),
    .o1(u_dcfifo_tx_u_dout_empty_synch_d_middle[6]),
    .o2(u_dcfifo_tx_u_dout_empty_synch_d_middle[7]),
    .si1(net1078),
    .si2(net1079),
    .ssb(net1765));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_0__u_dcfifo_tx_u_dout_empty_synch_d_out_reg_5_ (.rb(net442),
    .clk(clknet_3_0__leaf_spi_sclk),
    .d1(net2294),
    .d2(net2326),
    .o1(u_dcfifo_tx_u_dout_write_token_dn[0]),
    .o2(u_dcfifo_tx_u_dout_write_token_dn[5]),
    .si1(net1080),
    .si2(net1081),
    .ssb(net1766));
 b15fqy00car1n02x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_2_ (.clk(clknet_3_6__leaf_spi_sclk),
    .d(u_dcfifo_tx_u_dout_empty_synch_d_middle[2]),
    .o(u_dcfifo_tx_u_dout_write_token_dn[2]),
    .psb(net444),
    .si(net1082),
    .ssb(net1767));
 b15fqy00car1n02x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_3_ (.clk(clknet_3_0__leaf_spi_sclk),
    .d(net2237),
    .o(u_dcfifo_tx_u_dout_write_token_dn[3]),
    .psb(net442),
    .si(net1083),
    .ssb(net1768));
 b15fqy003ar1n02x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_4_ (.rb(net442),
    .clk(clknet_3_2__leaf_spi_sclk),
    .d(net2322),
    .o(u_dcfifo_tx_u_dout_write_token_dn[4]),
    .si(net1084),
    .ssb(net1769));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_6__u_dcfifo_tx_u_dout_empty_synch_d_out_reg_7_ (.rb(net442),
    .clk(clknet_3_2__leaf_spi_sclk),
    .d1(net2305),
    .d2(net2292),
    .o1(u_dcfifo_tx_u_dout_write_token_dn[6]),
    .o2(u_dcfifo_tx_u_dout_write_token_dn[7]),
    .si1(net1085),
    .si2(net1086),
    .ssb(net1770));
 b15cilb05ah1n02x3 u_dcfifo_tx_u_dout_read_tr_clk_gate_state_reg_latch (.clk(clknet_3_2__leaf_spi_sclk),
    .clkout(u_dcfifo_tx_u_dout_read_tr_net634),
    .en(net2353),
    .te(net1087));
 b15fqy00car1n02x5 u_dcfifo_tx_u_dout_read_tr_state_reg_0_ (.clk(clknet_1_1__leaf_u_dcfifo_tx_u_dout_read_tr_net634),
    .d(net2302),
    .o(u_dcfifo_tx_u_dout_read_token[0]),
    .psb(net442),
    .si(net1088),
    .ssb(net1771));
 b15fqy00car1n02x5 u_dcfifo_tx_u_dout_read_tr_state_reg_1_ (.clk(clknet_1_0__leaf_u_dcfifo_tx_u_dout_read_tr_net634),
    .d(u_dcfifo_tx_u_dout_read_token[0]),
    .o(u_dcfifo_tx_u_dout_read_token[1]),
    .psb(net442),
    .si(net1089),
    .ssb(net1772));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_dout_read_tr_state_reg_2__u_dcfifo_tx_u_dout_read_tr_state_reg_3_ (.rb(net442),
    .clk(clknet_1_0__leaf_u_dcfifo_tx_u_dout_read_tr_net634),
    .d1(net2365),
    .d2(u_dcfifo_tx_u_dout_read_token[2]),
    .o1(u_dcfifo_tx_u_dout_read_token[2]),
    .o2(u_dcfifo_tx_u_dout_read_token[3]),
    .si1(net1090),
    .si2(net1091),
    .ssb(net1773));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_dout_read_tr_state_reg_4__u_dcfifo_tx_u_dout_read_tr_state_reg_5_ (.rb(net442),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_dout_read_tr_net634),
    .d1(net305),
    .d2(u_dcfifo_tx_u_dout_read_token[4]),
    .o1(u_dcfifo_tx_u_dout_read_token[4]),
    .o2(u_dcfifo_tx_u_dout_read_token[5]),
    .si1(net1092),
    .si2(net1093),
    .ssb(net1774));
 b15fqy203ar1n02x5 u_dcfifo_tx_u_dout_read_tr_state_reg_6__u_dcfifo_tx_u_dout_read_tr_state_reg_7_ (.rb(net442),
    .clk(clknet_1_1__leaf_u_dcfifo_tx_u_dout_read_tr_net634),
    .d1(u_dcfifo_tx_u_dout_read_token[5]),
    .d2(u_dcfifo_tx_u_dout_read_token[6]),
    .o1(u_dcfifo_tx_u_dout_read_token[6]),
    .o2(u_dcfifo_tx_u_dout_read_token[7]),
    .si1(net1094),
    .si2(net1095),
    .ssb(net1775));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_0__u_device_sm_addr_reg_reg_1_ (.rb(net366),
    .clk(clknet_1_0__leaf_u_device_sm_net763),
    .d1(net259),
    .d2(net239),
    .o1(addr_sync[0]),
    .o2(addr_sync[1]),
    .si1(net1096),
    .si2(net1097),
    .ssb(net1776));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_10__u_device_sm_addr_reg_reg_11_ (.rb(net366),
    .clk(clknet_1_0__leaf_u_device_sm_net763),
    .d1(net217),
    .d2(net229),
    .o1(addr_sync[10]),
    .o2(addr_sync[11]),
    .si1(net1098),
    .si2(net1099),
    .ssb(net1777));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_12__u_device_sm_addr_reg_reg_13_ (.rb(net366),
    .clk(clknet_1_1__leaf_u_device_sm_net763),
    .d1(net193),
    .d2(net213),
    .o1(addr_sync[12]),
    .o2(addr_sync[13]),
    .si1(net1100),
    .si2(net1101),
    .ssb(net1778));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_14__u_device_sm_addr_reg_reg_15_ (.rb(net366),
    .clk(clknet_1_1__leaf_u_device_sm_net763),
    .d1(net221),
    .d2(ctrl_data_rx[15]),
    .o1(addr_sync[14]),
    .o2(addr_sync[15]),
    .si1(net1102),
    .si2(net1103),
    .ssb(net1779));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_16__u_device_sm_addr_reg_reg_17_ (.rb(n3770),
    .clk(clknet_1_0__leaf_u_device_sm_net769),
    .d1(net212),
    .d2(net225),
    .o1(addr_sync[16]),
    .o2(addr_sync[17]),
    .si1(net1104),
    .si2(net1105),
    .ssb(net1780));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_18__u_device_sm_addr_reg_reg_19_ (.rb(n3770),
    .clk(clknet_1_0__leaf_u_device_sm_net769),
    .d1(ctrl_data_rx[18]),
    .d2(ctrl_data_rx[19]),
    .o1(addr_sync[18]),
    .o2(addr_sync[19]),
    .si1(net1106),
    .si2(net1107),
    .ssb(net1781));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_20__u_device_sm_addr_reg_reg_21_ (.rb(n3770),
    .clk(clknet_1_0__leaf_u_device_sm_net769),
    .d1(ctrl_data_rx[20]),
    .d2(ctrl_data_rx[21]),
    .o1(addr_sync[20]),
    .o2(addr_sync[21]),
    .si1(net1108),
    .si2(net1109),
    .ssb(net1782));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_22__u_device_sm_addr_reg_reg_23_ (.rb(n3770),
    .clk(clknet_1_0__leaf_u_device_sm_net769),
    .d1(ctrl_data_rx[22]),
    .d2(ctrl_data_rx[23]),
    .o1(addr_sync[22]),
    .o2(addr_sync[23]),
    .si1(net1110),
    .si2(net1111),
    .ssb(net1783));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_24__u_device_sm_addr_reg_reg_25_ (.rb(n3770),
    .clk(clknet_1_1__leaf_u_device_sm_net769),
    .d1(net197),
    .d2(net209),
    .o1(addr_sync[24]),
    .o2(addr_sync[25]),
    .si1(net1112),
    .si2(net1113),
    .ssb(net1784));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_26__u_device_sm_addr_reg_reg_27_ (.rb(n3770),
    .clk(clknet_1_1__leaf_u_device_sm_net769),
    .d1(ctrl_data_rx[26]),
    .d2(ctrl_data_rx[27]),
    .o1(addr_sync[26]),
    .o2(addr_sync[27]),
    .si1(net1114),
    .si2(net1115),
    .ssb(net1785));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_28__u_device_sm_addr_reg_reg_29_ (.rb(n3770),
    .clk(clknet_1_1__leaf_u_device_sm_net769),
    .d1(ctrl_data_rx[28]),
    .d2(ctrl_data_rx[29]),
    .o1(addr_sync[28]),
    .o2(addr_sync[29]),
    .si1(net1116),
    .si2(net1117),
    .ssb(net1786));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_2__u_device_sm_addr_reg_reg_3_ (.rb(n3774),
    .clk(clknet_1_0__leaf_u_device_sm_net763),
    .d1(net236),
    .d2(net248),
    .o1(addr_sync[2]),
    .o2(addr_sync[3]),
    .si1(net1118),
    .si2(net1119),
    .ssb(net1787));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_30__u_device_sm_addr_reg_reg_31_ (.rb(n3770),
    .clk(clknet_1_1__leaf_u_device_sm_net769),
    .d1(ctrl_data_rx[30]),
    .d2(net230),
    .o1(addr_sync[30]),
    .o2(addr_sync[31]),
    .si1(net1120),
    .si2(net1121),
    .ssb(net1788));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_4__u_device_sm_addr_reg_reg_5_ (.rb(net366),
    .clk(clknet_1_1__leaf_u_device_sm_net763),
    .d1(net233),
    .d2(net190),
    .o1(addr_sync[4]),
    .o2(addr_sync[5]),
    .si1(net1122),
    .si2(net1123),
    .ssb(net1789));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_6__u_device_sm_addr_reg_reg_7_ (.rb(net366),
    .clk(clknet_1_0__leaf_u_device_sm_net763),
    .d1(net241),
    .d2(net244),
    .o1(addr_sync[6]),
    .o2(addr_sync[7]),
    .si1(net1124),
    .si2(net1125),
    .ssb(net1790));
 b15fqy203ar1n02x5 u_device_sm_addr_reg_reg_8__u_device_sm_addr_reg_reg_9_ (.rb(net366),
    .clk(clknet_1_1__leaf_u_device_sm_net763),
    .d1(ctrl_data_rx[8]),
    .d2(ctrl_data_rx[9]),
    .o1(addr_sync[8]),
    .o2(addr_sync[9]),
    .si1(net1126),
    .si2(net1127),
    .ssb(net1791));
 b15cilb05ah1n02x3 u_device_sm_clk_gate_addr_reg_reg_0_latch (.clk(clknet_3_5__leaf_spi_sclk),
    .clkout(u_device_sm_net769),
    .en(net147),
    .te(net1128));
 b15cilb05ah1n02x3 u_device_sm_clk_gate_addr_reg_reg_latch (.clk(clknet_3_5__leaf_spi_sclk),
    .clkout(u_device_sm_net763),
    .en(net147),
    .te(net1129));
 b15cilb05ah1n02x3 u_device_sm_clk_gate_cmd_reg_reg_latch (.clk(clknet_3_2__leaf_spi_sclk),
    .clkout(u_device_sm_net774),
    .en(u_device_sm_sample_CMD),
    .te(net1130));
 b15fqy203ar1n02x5 u_device_sm_cmd_reg_reg_0__u_device_sm_cmd_reg_reg_1_ (.rb(net367),
    .clk(clknet_1_1__leaf_u_device_sm_net774),
    .d1(net258),
    .d2(net238),
    .o1(u_device_sm_cmd_reg[0]),
    .o2(u_device_sm_cmd_reg[1]),
    .si1(net1131),
    .si2(net1132),
    .ssb(net1792));
 b15fqy203ar1n02x5 u_device_sm_cmd_reg_reg_2__u_device_sm_cmd_reg_reg_3_ (.rb(n3774),
    .clk(clknet_1_0__leaf_u_device_sm_net774),
    .d1(net235),
    .d2(net246),
    .o1(u_device_sm_cmd_reg[2]),
    .o2(u_device_sm_cmd_reg[3]),
    .si1(net1133),
    .si2(net1134),
    .ssb(net1793));
 b15fqy203ar1n02x5 u_device_sm_cmd_reg_reg_4__u_device_sm_cmd_reg_reg_5_ (.rb(n3774),
    .clk(clknet_1_0__leaf_u_device_sm_net774),
    .d1(net234),
    .d2(net191),
    .o1(u_device_sm_cmd_reg[4]),
    .o2(u_device_sm_cmd_reg[5]),
    .si1(net1135),
    .si2(net1136),
    .ssb(net1794));
 b15fqy203ar1n02x5 u_device_sm_cmd_reg_reg_6__u_device_sm_cmd_reg_reg_7_ (.rb(n3774),
    .clk(clknet_1_1__leaf_u_device_sm_net774),
    .d1(net240),
    .d2(net243),
    .o1(u_device_sm_cmd_reg[6]),
    .o2(u_device_sm_cmd_reg[7]),
    .si1(net1137),
    .si2(net1138),
    .ssb(net1795));
 b15fqy203ar1n02x5 u_device_sm_ctrl_addr_valid_reg_u_device_sm_data_reg_reg_0_ (.rb(n3776),
    .clk(clknet_3_6__leaf_spi_sclk),
    .d1(net148),
    .d2(net2253),
    .o1(ctrl_addr_valid),
    .o2(n1712),
    .si1(net1139),
    .si2(net1140),
    .ssb(net1796));
 b15fqy203ar1n02x5 u_device_sm_ctrl_data_tx_ready_reg_u_device_sm_state_reg_1_ (.rb(net367),
    .clk(clknet_3_2__leaf_spi_sclk),
    .d1(u_device_sm_ctrl_data_tx_ready_next),
    .d2(u_device_sm_state_next[1]),
    .o1(ctrl_data_tx_ready),
    .o2(u_device_sm_state[1]),
    .si1(net1141),
    .si2(net1142),
    .ssb(net1797));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_10__u_device_sm_data_reg_reg_11_ (.rb(net368),
    .clk(clknet_3_6__leaf_spi_sclk),
    .d1(net2272),
    .d2(net2252),
    .o1(n1796),
    .o2(n1793),
    .si1(net1143),
    .si2(net1144),
    .ssb(net1798));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_12__u_device_sm_data_reg_reg_13_ (.rb(net364),
    .clk(clknet_3_3__leaf_spi_sclk),
    .d1(net2280),
    .d2(net2257),
    .o1(n1790),
    .o2(n1787),
    .si1(net1145),
    .si2(net1146),
    .ssb(net1799));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_14__u_device_sm_data_reg_reg_15_ (.rb(net368),
    .clk(clknet_3_3__leaf_spi_sclk),
    .d1(net2277),
    .d2(net2259),
    .o1(n1784),
    .o2(n1781),
    .si1(net1147),
    .si2(net1148),
    .ssb(net1800));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_16__u_device_sm_data_reg_reg_17_ (.rb(net365),
    .clk(clknet_3_4__leaf_spi_sclk),
    .d1(net2274),
    .d2(net2255),
    .o1(n1778),
    .o2(n1775),
    .si1(net1149),
    .si2(net1150),
    .ssb(net1801));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_18__u_device_sm_data_reg_reg_19_ (.rb(net364),
    .clk(clknet_3_6__leaf_spi_sclk),
    .d1(net2267),
    .d2(net2247),
    .o1(n1772),
    .o2(n1769),
    .si1(net1151),
    .si2(net1152),
    .ssb(net1802));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_1__u_device_sm_data_reg_reg_2_ (.rb(net364),
    .clk(clknet_3_3__leaf_spi_sclk),
    .d1(net2282),
    .d2(net2263),
    .o1(n1718),
    .o2(n1700),
    .si1(net1153),
    .si2(net1154),
    .ssb(net1803));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_20__u_device_sm_data_reg_reg_21_ (.rb(net369),
    .clk(clknet_3_3__leaf_spi_sclk),
    .d1(net2281),
    .d2(net2260),
    .o1(n1766),
    .o2(n1763),
    .si1(net1155),
    .si2(net1156),
    .ssb(net1804));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_22__u_device_sm_data_reg_reg_23_ (.rb(n3769),
    .clk(clknet_3_1__leaf_spi_sclk),
    .d1(net2265),
    .d2(net2244),
    .o1(n1760),
    .o2(n1757),
    .si1(net1157),
    .si2(net1158),
    .ssb(net1805));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_24__u_device_sm_data_reg_reg_25_ (.rb(net368),
    .clk(clknet_3_6__leaf_spi_sclk),
    .d1(net2268),
    .d2(net2248),
    .o1(n1754),
    .o2(n1751),
    .si1(net1159),
    .si2(net1160),
    .ssb(net1806));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_26__u_device_sm_data_reg_reg_27_ (.rb(n3769),
    .clk(clknet_3_6__leaf_spi_sclk),
    .d1(net2273),
    .d2(net2254),
    .o1(n1748),
    .o2(n1745),
    .si1(net1161),
    .si2(net1162),
    .ssb(net1807));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_28__u_device_sm_data_reg_reg_29_ (.rb(n3769),
    .clk(clknet_3_0__leaf_spi_sclk),
    .d1(net2264),
    .d2(net2243),
    .o1(n1742),
    .o2(n1739),
    .si1(net1163),
    .si2(net1164),
    .ssb(net1808));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_30__u_device_sm_data_reg_reg_31_ (.rb(net368),
    .clk(clknet_3_6__leaf_spi_sclk),
    .d1(net2266),
    .d2(net2246),
    .o1(n1736),
    .o2(n1733),
    .si1(net1165),
    .si2(net1166),
    .ssb(net1809));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_3__u_device_sm_data_reg_reg_4_ (.rb(net364),
    .clk(clknet_3_3__leaf_spi_sclk),
    .d1(net2276),
    .d2(net2258),
    .o1(n1694),
    .o2(n1706),
    .si1(net1167),
    .si2(net1168),
    .ssb(net1810));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_5__u_device_sm_state_reg_0_ (.rb(net369),
    .clk(clknet_3_2__leaf_spi_sclk),
    .d1(net2286),
    .d2(u_device_sm_state_next[0]),
    .o1(n1881),
    .o2(u_device_sm_state[0]),
    .si1(net1169),
    .si2(net1170),
    .ssb(net1811));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_6__u_device_sm_data_reg_reg_7_ (.rb(net364),
    .clk(clknet_3_6__leaf_spi_sclk),
    .d1(net2271),
    .d2(net2251),
    .o1(n1724),
    .o2(n1730),
    .si1(net1171),
    .si2(net1172),
    .ssb(net1812));
 b15fqy203ar1n02x5 u_device_sm_data_reg_reg_8__u_device_sm_data_reg_reg_9_ (.rb(net364),
    .clk(clknet_3_3__leaf_spi_sclk),
    .d1(net2278),
    .d2(net2261),
    .o1(n1802),
    .o2(n1799),
    .si1(net1173),
    .si2(net1174),
    .ssb(net1813));
 b15fqy203ar1n02x5 u_device_sm_mode_reg_reg_0__u_device_sm_mode_reg_reg_1_ (.rb(net368),
    .clk(clknet_3_3__leaf_spi_sclk),
    .d1(net2275),
    .d2(net2256),
    .o1(n1709),
    .o2(n1715),
    .si1(net1175),
    .si2(net1176),
    .ssb(net1814));
 b15fqy203ar1n02x5 u_device_sm_mode_reg_reg_2__u_device_sm_mode_reg_reg_3_ (.rb(net364),
    .clk(clknet_3_3__leaf_spi_sclk),
    .d1(net2279),
    .d2(net2262),
    .o1(n1697),
    .o2(n1691),
    .si1(net1177),
    .si2(net1178),
    .ssb(net1815));
 b15fqy203ar1n02x5 u_device_sm_mode_reg_reg_4__u_device_sm_mode_reg_reg_5_ (.rb(net364),
    .clk(clknet_3_6__leaf_spi_sclk),
    .d1(net2269),
    .d2(net2249),
    .o1(n1703),
    .o2(n1878),
    .si1(net1179),
    .si2(net1180),
    .ssb(net1816));
 b15fqy203ar1n02x5 u_device_sm_mode_reg_reg_6__u_device_sm_mode_reg_reg_7_ (.rb(net368),
    .clk(clknet_3_6__leaf_spi_sclk),
    .d1(net2270),
    .d2(net2250),
    .o1(n1721),
    .o2(n1727),
    .si1(net1181),
    .si2(net1182),
    .ssb(net1817));
 b15lsn000ar1n02x5 u_device_sm_pad_mode_next_reg_0_ (.clk(u_device_sm_N163),
    .d(net1818));
 b15lsn000ar1n02x5 u_device_sm_pad_mode_next_reg_1_ (.clk(u_device_sm_N163),
    .d(net1183));
 b15fqy203ar1n02x5 u_device_sm_state_reg_2__u_device_sm_tx_counter_reg_0_ (.rb(n3777),
    .clk(clknet_3_2__leaf_spi_sclk),
    .d1(u_device_sm_state_next[2]),
    .d2(net1819),
    .o1(u_device_sm_state[2]),
    .o2(tx_counter[0]),
    .si1(net1184),
    .si2(net1185),
    .ssb(net1820));
 b15fqy203ar1n02x5 u_device_sm_tx_counter_reg_1__u_device_sm_tx_data_reg_0_ (.rb(n3769),
    .clk(clknet_3_2__leaf_spi_sclk),
    .d1(net1821),
    .d2(u_device_sm_N174),
    .o1(tx_counter[1]),
    .o2(tx_data[0]),
    .si1(net1186),
    .si2(net1187),
    .ssb(net1822));
 b15fqy203ar1n02x5 u_device_sm_tx_counter_reg_2__u_device_sm_tx_counter_reg_3_ (.rb(net367),
    .clk(clknet_3_2__leaf_spi_sclk),
    .d1(net1823),
    .d2(u_device_sm_tx_counter_next_3_),
    .o1(tx_counter[2]),
    .o2(tx_counter[3]),
    .si1(net1188),
    .si2(net1189),
    .ssb(net1824));
 b15fqy203ar1n02x5 u_device_sm_tx_counter_reg_4__u_device_sm_tx_counter_upd_reg (.rb(net367),
    .clk(clknet_3_2__leaf_spi_sclk),
    .d1(u_device_sm_tx_counter_next_3_),
    .d2(u_device_sm_tx_counter_upd_next),
    .o1(tx_counter[4]),
    .o2(tx_counter_upd),
    .si1(net1190),
    .si2(net1191),
    .ssb(net1825));
 b15fqy203ar1n02x5 u_device_sm_tx_counter_reg_5__u_device_sm_tx_counter_reg_6_ (.rb(n3769),
    .clk(clknet_3_2__leaf_spi_sclk),
    .d1(net1192),
    .d2(net1193),
    .o1(tx_counter[5]),
    .o2(tx_counter[6]),
    .si1(net1194),
    .si2(net1195),
    .ssb(net1826));
 b15fqy003ar1n02x5 u_device_sm_tx_counter_reg_7_ (.rb(net365),
    .clk(clknet_3_0__leaf_spi_sclk),
    .d(net1196),
    .o(tx_counter[7]),
    .si(net1197),
    .ssb(net1827));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_11__u_device_sm_tx_data_reg_12_ (.rb(n3776),
    .clk(clknet_3_1__leaf_spi_sclk),
    .d1(u_device_sm_N185),
    .d2(u_device_sm_N186),
    .o1(tx_data[11]),
    .o2(tx_data[12]),
    .si1(net1198),
    .si2(net1199),
    .ssb(net1828));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_13__u_device_sm_tx_data_reg_14_ (.rb(n3776),
    .clk(clknet_3_1__leaf_spi_sclk),
    .d1(u_device_sm_N187),
    .d2(u_device_sm_N188),
    .o1(tx_data[13]),
    .o2(tx_data[14]),
    .si1(net1200),
    .si2(net1201),
    .ssb(net1829));
 b15fqy003ar1n02x5 u_device_sm_tx_data_reg_15_ (.rb(n3773),
    .clk(clknet_3_1__leaf_spi_sclk),
    .d(u_device_sm_N189),
    .o(tx_data[15]),
    .si(net1202),
    .ssb(net1830));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_16__u_device_sm_tx_data_reg_17_ (.rb(n3771),
    .clk(clknet_3_1__leaf_spi_sclk),
    .d1(u_device_sm_N190),
    .d2(u_device_sm_N191),
    .o1(tx_data[16]),
    .o2(tx_data[17]),
    .si1(net1203),
    .si2(net1204),
    .ssb(net1831));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_18__u_device_sm_tx_data_reg_19_ (.rb(n3771),
    .clk(clknet_3_1__leaf_spi_sclk),
    .d1(u_device_sm_N192),
    .d2(u_device_sm_N193),
    .o1(tx_data[18]),
    .o2(tx_data[19]),
    .si1(net1205),
    .si2(net1206),
    .ssb(net1832));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_1__u_device_sm_tx_data_reg_2_ (.rb(net363),
    .clk(clknet_3_2__leaf_spi_sclk),
    .d1(u_device_sm_N175),
    .d2(u_device_sm_N176),
    .o1(tx_data[1]),
    .o2(tx_data[2]),
    .si1(net1207),
    .si2(net1208),
    .ssb(net1833));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_20__u_device_sm_tx_data_reg_21_ (.rb(n3771),
    .clk(clknet_3_1__leaf_spi_sclk),
    .d1(u_device_sm_N194),
    .d2(u_device_sm_N195),
    .o1(tx_data[20]),
    .o2(tx_data[21]),
    .si1(net1209),
    .si2(net1210),
    .ssb(net1834));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_22__u_device_sm_tx_data_reg_23_ (.rb(n3771),
    .clk(clknet_3_4__leaf_spi_sclk),
    .d1(u_device_sm_N196),
    .d2(u_device_sm_N197),
    .o1(tx_data[22]),
    .o2(tx_data[23]),
    .si1(net1211),
    .si2(net1212),
    .ssb(net1835));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_24__u_device_sm_tx_data_reg_25_ (.rb(n3771),
    .clk(clknet_3_1__leaf_spi_sclk),
    .d1(u_device_sm_N198),
    .d2(u_device_sm_N199),
    .o1(tx_data[24]),
    .o2(tx_data[25]),
    .si1(net1213),
    .si2(net1214),
    .ssb(net1836));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_26__u_device_sm_tx_data_reg_27_ (.rb(n3771),
    .clk(clknet_3_1__leaf_spi_sclk),
    .d1(u_device_sm_N200),
    .d2(u_device_sm_N201),
    .o1(tx_data[26]),
    .o2(tx_data[27]),
    .si1(net1215),
    .si2(net1216),
    .ssb(net1837));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_28__u_device_sm_tx_data_reg_29_ (.rb(n3771),
    .clk(clknet_3_5__leaf_spi_sclk),
    .d1(u_device_sm_N202),
    .d2(u_device_sm_N203),
    .o1(tx_data[28]),
    .o2(tx_data[29]),
    .si1(net1217),
    .si2(net1218),
    .ssb(net1838));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_30__u_device_sm_tx_data_reg_31_ (.rb(n3771),
    .clk(clknet_3_4__leaf_spi_sclk),
    .d1(u_device_sm_N204),
    .d2(u_device_sm_N205),
    .o1(tx_data[30]),
    .o2(tx_data[31]),
    .si1(net1219),
    .si2(net1220),
    .ssb(net1839));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_3__u_device_sm_tx_data_reg_4_ (.rb(net363),
    .clk(clknet_3_0__leaf_spi_sclk),
    .d1(u_device_sm_N177),
    .d2(u_device_sm_N178),
    .o1(tx_data[3]),
    .o2(tx_data[4]),
    .si1(net1221),
    .si2(net1222),
    .ssb(net1840));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_5__u_device_sm_tx_data_reg_6_ (.rb(net363),
    .clk(clknet_3_0__leaf_spi_sclk),
    .d1(u_device_sm_N179),
    .d2(u_device_sm_N180),
    .o1(tx_data[5]),
    .o2(tx_data[6]),
    .si1(net1223),
    .si2(net1224),
    .ssb(net1841));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_7__u_device_sm_tx_data_reg_8_ (.rb(net368),
    .clk(clknet_3_1__leaf_spi_sclk),
    .d1(u_device_sm_N181),
    .d2(u_device_sm_N182),
    .o1(tx_data[7]),
    .o2(tx_data[8]),
    .si1(net1225),
    .si2(net1226),
    .ssb(net1842));
 b15fqy203ar1n02x5 u_device_sm_tx_data_reg_9__u_device_sm_tx_data_reg_10_ (.rb(n3778),
    .clk(clknet_3_1__leaf_spi_sclk),
    .d1(u_device_sm_N183),
    .d2(u_device_sm_N184),
    .o1(tx_data[9]),
    .o2(tx_data[10]),
    .si1(net1227),
    .si2(net1228),
    .ssb(net1843));
 b15fqy203ar1n03x5 u_device_sm_tx_data_valid_reg_u_device_sm_tx_done_reg_reg (.rb(net367),
    .clk(clknet_3_2__leaf_spi_sclk),
    .d1(u_device_sm_tx_data_valid_next),
    .d2(tx_done),
    .o1(tx_data_valid),
    .o2(u_device_sm_tx_done_reg),
    .si1(net1229),
    .si2(net1230),
    .ssb(net1844));
 b15cilb05ah1n02x3 u_device_sm_u_spiregs_clk_gate_reg0_reg_latch (.clk(clknet_3_3__leaf_spi_sclk),
    .clkout(u_device_sm_u_spiregs_net797),
    .en(u_device_sm_u_spiregs_N32),
    .te(net1231));
 b15cilb05ah1n02x3 u_device_sm_u_spiregs_clk_gate_reg1_reg_latch (.clk(clknet_3_3__leaf_spi_sclk),
    .clkout(u_device_sm_u_spiregs_net802),
    .en(u_device_sm_u_spiregs_N33),
    .te(net1232));
 b15cilb05ah1n02x3 u_device_sm_u_spiregs_clk_gate_reg2_reg_latch (.clk(clknet_3_3__leaf_spi_sclk),
    .clkout(u_device_sm_u_spiregs_net807),
    .en(u_device_sm_u_spiregs_N34),
    .te(net1233));
 b15cilb05ah1n02x3 u_device_sm_u_spiregs_clk_gate_reg3_reg_latch (.clk(clknet_3_3__leaf_spi_sclk),
    .clkout(u_device_sm_u_spiregs_net791),
    .en(u_device_sm_u_spiregs_N31),
    .te(net1234));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg0_reg_0__u_device_sm_u_spiregs_reg0_reg_1_ (.rb(net442),
    .clk(clknet_1_1__leaf_u_device_sm_u_spiregs_net797),
    .d1(net258),
    .d2(net238),
    .o1(en_quad),
    .o2(u_device_sm_u_spiregs_reg0[1]),
    .si1(net1235),
    .si2(net1236),
    .ssb(net1845));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg0_reg_2__u_device_sm_u_spiregs_reg0_reg_3_ (.rb(net446),
    .clk(clknet_1_1__leaf_u_device_sm_u_spiregs_net797),
    .d1(net235),
    .d2(net246),
    .o1(u_device_sm_u_spiregs_reg0[2]),
    .o2(u_device_sm_u_spiregs_reg0[3]),
    .si1(net1237),
    .si2(net1238),
    .ssb(net1846));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg0_reg_4__u_device_sm_u_spiregs_reg0_reg_5_ (.rb(net446),
    .clk(clknet_1_0__leaf_u_device_sm_u_spiregs_net797),
    .d1(net234),
    .d2(net191),
    .o1(u_device_sm_u_spiregs_reg0[4]),
    .o2(u_device_sm_u_spiregs_reg0[5]),
    .si1(net1239),
    .si2(net1240),
    .ssb(net1847));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg0_reg_6__u_device_sm_u_spiregs_reg0_reg_7_ (.rb(net446),
    .clk(clknet_1_0__leaf_u_device_sm_u_spiregs_net797),
    .d1(net240),
    .d2(net243),
    .o1(u_device_sm_u_spiregs_reg0[6]),
    .o2(u_device_sm_u_spiregs_reg0[7]),
    .si1(net1241),
    .si2(net1242),
    .ssb(net1848));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg1_reg_0__u_device_sm_u_spiregs_reg1_reg_1_ (.rb(net444),
    .clk(clknet_1_0__leaf_u_device_sm_u_spiregs_net802),
    .d1(net258),
    .d2(net238),
    .o1(u_device_sm_s_dummy_cycles[0]),
    .o2(u_device_sm_s_dummy_cycles[1]),
    .si1(net1243),
    .si2(net1244),
    .ssb(net1849));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg1_reg_2__u_device_sm_u_spiregs_reg1_reg_3_ (.rb(net444),
    .clk(clknet_1_1__leaf_u_device_sm_u_spiregs_net802),
    .d1(net235),
    .d2(net246),
    .o1(u_device_sm_s_dummy_cycles[2]),
    .o2(u_device_sm_s_dummy_cycles[3]),
    .si1(net1245),
    .si2(net1246),
    .ssb(net1850));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg1_reg_4__u_device_sm_u_spiregs_reg1_reg_6_ (.rb(net444),
    .clk(clknet_1_1__leaf_u_device_sm_u_spiregs_net802),
    .d1(net234),
    .d2(net240),
    .o1(u_device_sm_s_dummy_cycles[4]),
    .o2(u_device_sm_s_dummy_cycles[6]),
    .si1(net1247),
    .si2(net1248),
    .ssb(net1851));
 b15fqy00car1n02x5 u_device_sm_u_spiregs_reg1_reg_5_ (.clk(clknet_1_0__leaf_u_device_sm_u_spiregs_net802),
    .d(net191),
    .o(u_device_sm_s_dummy_cycles[5]),
    .psb(net444),
    .si(net1249),
    .ssb(net1852));
 b15fqy003ar1n02x5 u_device_sm_u_spiregs_reg1_reg_7_ (.rb(net444),
    .clk(clknet_1_0__leaf_u_device_sm_u_spiregs_net802),
    .d(net243),
    .o(u_device_sm_s_dummy_cycles[7]),
    .si(net1250),
    .ssb(net1853));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg2_reg_0__u_device_sm_u_spiregs_reg2_reg_1_ (.rb(net446),
    .clk(clknet_1_0__leaf_u_device_sm_u_spiregs_net807),
    .d1(net258),
    .d2(net238),
    .o1(u_device_sm_u_spiregs_n[16]),
    .o2(u_device_sm_u_spiregs_n[15]),
    .si1(net1251),
    .si2(net1252),
    .ssb(net1854));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg2_reg_2__u_device_sm_u_spiregs_reg2_reg_3_ (.rb(net446),
    .clk(clknet_1_0__leaf_u_device_sm_u_spiregs_net807),
    .d1(net235),
    .d2(net246),
    .o1(u_device_sm_u_spiregs_n[14]),
    .o2(u_device_sm_u_spiregs_n[13]),
    .si1(net1253),
    .si2(net1254),
    .ssb(net1855));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg2_reg_4__u_device_sm_u_spiregs_reg2_reg_5_ (.rb(net446),
    .clk(clknet_1_1__leaf_u_device_sm_u_spiregs_net807),
    .d1(net234),
    .d2(net191),
    .o1(u_device_sm_u_spiregs_n[12]),
    .o2(u_device_sm_u_spiregs_n[11]),
    .si1(net1255),
    .si2(net1256),
    .ssb(net1856));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg2_reg_6__u_device_sm_u_spiregs_reg2_reg_7_ (.rb(net446),
    .clk(clknet_1_1__leaf_u_device_sm_u_spiregs_net807),
    .d1(net240),
    .d2(net243),
    .o1(u_device_sm_u_spiregs_n[10]),
    .o2(u_device_sm_u_spiregs_n[9]),
    .si1(net1257),
    .si2(net1258),
    .ssb(net1857));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg3_reg_0__u_device_sm_u_spiregs_reg3_reg_1_ (.rb(net444),
    .clk(clknet_1_0__leaf_u_device_sm_u_spiregs_net791),
    .d1(net258),
    .d2(net238),
    .o1(u_device_sm_u_spiregs_n[8]),
    .o2(u_device_sm_u_spiregs_n[7]),
    .si1(net1259),
    .si2(net1260),
    .ssb(net1858));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg3_reg_2__u_device_sm_u_spiregs_reg3_reg_3_ (.rb(net444),
    .clk(clknet_1_1__leaf_u_device_sm_u_spiregs_net791),
    .d1(net235),
    .d2(net246),
    .o1(u_device_sm_u_spiregs_n[6]),
    .o2(u_device_sm_u_spiregs_n[5]),
    .si1(net1261),
    .si2(net1262),
    .ssb(net1859));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg3_reg_4__u_device_sm_u_spiregs_reg3_reg_5_ (.rb(net444),
    .clk(clknet_1_1__leaf_u_device_sm_u_spiregs_net791),
    .d1(net234),
    .d2(net191),
    .o1(u_device_sm_u_spiregs_n[4]),
    .o2(u_device_sm_u_spiregs_n[3]),
    .si1(net1263),
    .si2(net1264),
    .ssb(net1860));
 b15fqy203ar1n02x5 u_device_sm_u_spiregs_reg3_reg_6__u_device_sm_u_spiregs_reg3_reg_7_ (.rb(net444),
    .clk(clknet_1_0__leaf_u_device_sm_u_spiregs_net791),
    .d1(net240),
    .d2(net243),
    .o1(u_device_sm_u_spiregs_n[2]),
    .o2(u_device_sm_u_spiregs_n[1]),
    .si1(net1265),
    .si2(net1266),
    .ssb(net1861));
 b15cilb05ah1n02x3 u_rxreg_clk_gate_counter_reg_latch (.clk(clknet_3_2__leaf_spi_sclk),
    .clkout(u_rxreg_net857),
    .en(n3809),
    .te(net1267));
 b15cilb05ah1n02x3 u_rxreg_clk_gate_counter_trgt_reg_latch (.clk(clknet_3_2__leaf_spi_sclk),
    .clkout(u_rxreg_net873),
    .en(u_rxreg_N7),
    .te(net1268));
 b15cilb05ah1n02x3 u_rxreg_clk_gate_data_int_reg_0_latch (.clk(clknet_3_4__leaf_spi_sclk),
    .clkout(u_rxreg_net868),
    .en(n3809),
    .te(net1269));
 b15cilb05ah1n02x3 u_rxreg_clk_gate_data_int_reg_latch (.clk(clknet_3_1__leaf_spi_sclk),
    .clkout(u_rxreg_net863),
    .en(n3809),
    .te(net1270));
 b15fqy203ar1n02x5 u_rxreg_counter_reg_0__u_rxreg_counter_reg_1_ (.rb(net369),
    .clk(clknet_1_1__leaf_u_rxreg_net857),
    .d1(u_rxreg_N22),
    .d2(u_rxreg_N23),
    .o1(u_rxreg_counter[0]),
    .o2(u_rxreg_counter[1]),
    .si1(net1271),
    .si2(net1272),
    .ssb(net1862));
 b15fqy203ar1n02x5 u_rxreg_counter_reg_2__u_rxreg_counter_reg_3_ (.rb(net363),
    .clk(clknet_1_0__leaf_u_rxreg_net857),
    .d1(u_rxreg_N24),
    .d2(u_rxreg_N25),
    .o1(u_rxreg_counter[2]),
    .o2(u_rxreg_counter[3]),
    .si1(net1273),
    .si2(net1274),
    .ssb(net1863));
 b15fqy203ar1n02x5 u_rxreg_counter_reg_4__u_rxreg_counter_reg_5_ (.rb(net369),
    .clk(clknet_1_0__leaf_u_rxreg_net857),
    .d1(u_rxreg_N26),
    .d2(u_rxreg_N27),
    .o1(u_rxreg_counter[4]),
    .o2(u_rxreg_counter[5]),
    .si1(net1275),
    .si2(net1276),
    .ssb(net1864));
 b15fqy203ar1n02x5 u_rxreg_counter_reg_6__u_rxreg_counter_reg_7_ (.rb(net363),
    .clk(clknet_1_1__leaf_u_rxreg_net857),
    .d1(u_rxreg_N28),
    .d2(u_rxreg_N29),
    .o1(u_rxreg_counter[6]),
    .o2(u_rxreg_counter[7]),
    .si1(net1277),
    .si2(net1278),
    .ssb(net1865));
 b15fqy00car1n02x5 u_rxreg_counter_trgt_reg_0_ (.clk(clknet_1_1__leaf_u_rxreg_net873),
    .d(u_rxreg_counter_trgt_next[0]),
    .o(u_rxreg_counter_trgt[0]),
    .psb(n3777),
    .si(net1279),
    .ssb(net1866));
 b15fqy203ar1n02x5 u_rxreg_counter_trgt_reg_1__u_rxreg_counter_trgt_reg_2_ (.rb(net363),
    .clk(clknet_1_0__leaf_u_rxreg_net873),
    .d1(u_rxreg_counter_trgt_next[1]),
    .d2(u_rxreg_counter_trgt_next[2]),
    .o1(u_rxreg_counter_trgt[1]),
    .o2(u_rxreg_counter_trgt[2]),
    .si1(net1280),
    .si2(net1281),
    .ssb(net1867));
 b15fqy203ar1n02x5 u_rxreg_counter_trgt_reg_3__u_rxreg_counter_trgt_reg_4_ (.rb(net363),
    .clk(clknet_1_1__leaf_u_rxreg_net873),
    .d1(u_rxreg_counter_trgt_next[3]),
    .d2(u_rxreg_counter_trgt_next[4]),
    .o1(u_rxreg_counter_trgt[3]),
    .o2(u_rxreg_counter_trgt[4]),
    .si1(net1282),
    .si2(net1283),
    .ssb(net1868));
 b15fqy203ar1n02x5 u_rxreg_counter_trgt_reg_5__u_rxreg_counter_trgt_reg_6_ (.rb(net363),
    .clk(clknet_1_0__leaf_u_rxreg_net873),
    .d1(u_rxreg_counter_trgt_next[5]),
    .d2(u_rxreg_counter_trgt_next[6]),
    .o1(u_rxreg_counter_trgt[5]),
    .o2(u_rxreg_counter_trgt[6]),
    .si1(net1284),
    .si2(net1285),
    .ssb(net1869));
 b15fqy003ar1n02x5 u_rxreg_counter_trgt_reg_7_ (.rb(net363),
    .clk(clknet_1_0__leaf_u_rxreg_net873),
    .d(u_rxreg_counter_trgt_next[7]),
    .o(u_rxreg_counter_trgt[7]),
    .si(net1286),
    .ssb(net1870));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_0__u_rxreg_data_int_reg_1_ (.rb(n3774),
    .clk(clknet_1_0__leaf_u_rxreg_net863),
    .d1(net3),
    .d2(u_rxreg_N30),
    .o1(u_rxreg_data_int[0]),
    .o2(u_rxreg_data_int[1]),
    .si1(net1287),
    .si2(net1288),
    .ssb(net1871));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_10__u_rxreg_data_int_reg_11_ (.rb(n3773),
    .clk(clknet_1_0__leaf_u_rxreg_net863),
    .d1(u_rxreg_N39),
    .d2(u_rxreg_N40),
    .o1(u_rxreg_data_int[10]),
    .o2(u_rxreg_data_int[11]),
    .si1(net1289),
    .si2(net1290),
    .ssb(net1872));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_12__u_rxreg_data_int_reg_13_ (.rb(n3773),
    .clk(clknet_1_1__leaf_u_rxreg_net863),
    .d1(u_rxreg_N41),
    .d2(u_rxreg_N42),
    .o1(u_rxreg_data_int[12]),
    .o2(u_rxreg_data_int[13]),
    .si1(net1291),
    .si2(net1292),
    .ssb(net1873));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_14__u_rxreg_data_int_reg_15_ (.rb(n3773),
    .clk(clknet_1_0__leaf_u_rxreg_net863),
    .d1(u_rxreg_N43),
    .d2(u_rxreg_N44),
    .o1(u_rxreg_data_int[14]),
    .o2(u_rxreg_data_int[15]),
    .si1(net1293),
    .si2(net1294),
    .ssb(net1874));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_16__u_rxreg_data_int_reg_17_ (.rb(n3773),
    .clk(clknet_1_0__leaf_u_rxreg_net868),
    .d1(u_rxreg_N45),
    .d2(u_rxreg_N46),
    .o1(u_rxreg_data_int[16]),
    .o2(u_rxreg_data_int[17]),
    .si1(net1295),
    .si2(net1296),
    .ssb(net1875));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_18__u_rxreg_data_int_reg_19_ (.rb(n3773),
    .clk(clknet_1_0__leaf_u_rxreg_net868),
    .d1(u_rxreg_N47),
    .d2(u_rxreg_N48),
    .o1(u_rxreg_data_int[18]),
    .o2(u_rxreg_data_int[19]),
    .si1(net1297),
    .si2(net1298),
    .ssb(net1876));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_20__u_rxreg_data_int_reg_21_ (.rb(n3773),
    .clk(clknet_1_1__leaf_u_rxreg_net868),
    .d1(u_rxreg_N49),
    .d2(u_rxreg_N50),
    .o1(u_rxreg_data_int[20]),
    .o2(u_rxreg_data_int[21]),
    .si1(net1299),
    .si2(net1300),
    .ssb(net1877));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_22__u_rxreg_data_int_reg_23_ (.rb(n3773),
    .clk(clknet_1_1__leaf_u_rxreg_net868),
    .d1(u_rxreg_N51),
    .d2(u_rxreg_N52),
    .o1(u_rxreg_data_int[22]),
    .o2(u_rxreg_data_int[23]),
    .si1(net1301),
    .si2(net1302),
    .ssb(net1878));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_24__u_rxreg_data_int_reg_25_ (.rb(n3773),
    .clk(clknet_1_1__leaf_u_rxreg_net868),
    .d1(u_rxreg_N53),
    .d2(u_rxreg_N54),
    .o1(u_rxreg_data_int[24]),
    .o2(u_rxreg_data_int[25]),
    .si1(net1303),
    .si2(net1304),
    .ssb(net1879));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_26__u_rxreg_data_int_reg_27_ (.rb(n3773),
    .clk(clknet_1_0__leaf_u_rxreg_net868),
    .d1(u_rxreg_N55),
    .d2(u_rxreg_N56),
    .o1(u_rxreg_data_int[26]),
    .o2(u_rxreg_data_int[27]),
    .si1(net1305),
    .si2(net1306),
    .ssb(net1880));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_28__u_rxreg_data_int_reg_29_ (.rb(n3773),
    .clk(clknet_1_0__leaf_u_rxreg_net868),
    .d1(u_rxreg_N57),
    .d2(u_rxreg_N58),
    .o1(u_rxreg_data_int[28]),
    .o2(u_rxreg_data_int[29]),
    .si1(net1307),
    .si2(net1308),
    .ssb(net1881));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_2__u_rxreg_data_int_reg_3_ (.rb(n3774),
    .clk(clknet_1_0__leaf_u_rxreg_net863),
    .d1(u_rxreg_N31),
    .d2(u_rxreg_N32),
    .o1(u_rxreg_data_int[2]),
    .o2(u_rxreg_data_int[3]),
    .si1(net1309),
    .si2(net1310),
    .ssb(net1882));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_30__u_rxreg_data_int_reg_31_ (.rb(n3773),
    .clk(clknet_1_1__leaf_u_rxreg_net868),
    .d1(u_rxreg_N59),
    .d2(u_rxreg_N60),
    .o1(u_rxreg_data_int[30]),
    .o2(u_rxreg_data_int[31]),
    .si1(net1311),
    .si2(net1312),
    .ssb(net1883));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_4__u_rxreg_data_int_reg_5_ (.rb(n3778),
    .clk(clknet_1_1__leaf_u_rxreg_net863),
    .d1(u_rxreg_N33),
    .d2(u_rxreg_N34),
    .o1(u_rxreg_data_int[4]),
    .o2(u_rxreg_data_int[5]),
    .si1(net1313),
    .si2(net1314),
    .ssb(net1884));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_6__u_rxreg_data_int_reg_7_ (.rb(n3774),
    .clk(clknet_1_1__leaf_u_rxreg_net863),
    .d1(u_rxreg_N35),
    .d2(u_rxreg_N36),
    .o1(u_rxreg_data_int[6]),
    .o2(u_rxreg_data_int[7]),
    .si1(net1315),
    .si2(net1316),
    .ssb(net1885));
 b15fqy203ar1n02x5 u_rxreg_data_int_reg_8__u_rxreg_data_int_reg_9_ (.rb(n3773),
    .clk(clknet_1_1__leaf_u_rxreg_net863),
    .d1(u_rxreg_N37),
    .d2(u_rxreg_N38),
    .o1(u_rxreg_data_int[8]),
    .o2(u_rxreg_data_int[9]),
    .si1(net1317),
    .si2(net1318),
    .ssb(net1886));
 b15fqy043ar1n02x5 u_rxreg_running_reg (.clk(clknet_3_2__leaf_spi_sclk),
    .d(n2656),
    .den(u_rxreg_N9),
    .o(n1869),
    .rb(n3774),
    .si(net1319),
    .ssb(net1887));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_0__u_spi_device_tlul_plug_addr_reg_1_ (.rb(net455),
    .clk(clknet_1_0__leaf_u_spi_device_tlul_plug_net611),
    .d1(net2344),
    .d2(net2334),
    .si1(net1320),
    .si2(net1321),
    .ssb(net1888));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_10__u_spi_device_tlul_plug_addr_reg_11_ (.rb(net461),
    .clk(clknet_1_1__leaf_u_spi_device_tlul_plug_net611),
    .d1(addr_sync[10]),
    .d2(addr_sync[11]),
    .o1(net108),
    .o2(net109),
    .si1(net1322),
    .si2(net1323),
    .ssb(net1889));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_12__u_spi_device_tlul_plug_addr_reg_13_ (.rb(net461),
    .clk(clknet_1_0__leaf_u_spi_device_tlul_plug_net611),
    .d1(net2340),
    .d2(net2328),
    .o1(net110),
    .o2(net111),
    .si1(net1324),
    .si2(net1325),
    .ssb(net1890));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_14__u_spi_device_tlul_plug_addr_reg_15_ (.rb(net461),
    .clk(clknet_1_0__leaf_u_spi_device_tlul_plug_net611),
    .d1(net2368),
    .d2(net2361),
    .o1(net112),
    .o2(net113),
    .si1(net1326),
    .si2(net1327),
    .ssb(net1891));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_16__u_spi_device_tlul_plug_addr_reg_17_ (.rb(net461),
    .clk(clknet_1_0__leaf_u_spi_device_tlul_plug_net617),
    .d1(net2335),
    .d2(net2324),
    .o1(net114),
    .o2(net115),
    .si1(net1328),
    .si2(net1329),
    .ssb(net1892));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_18__u_spi_device_tlul_plug_addr_reg_19_ (.rb(net455),
    .clk(clknet_1_0__leaf_u_spi_device_tlul_plug_net617),
    .d1(addr_sync[18]),
    .d2(addr_sync[19]),
    .o1(net116),
    .o2(net117),
    .si1(net1330),
    .si2(net1331),
    .ssb(net1893));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_20__u_spi_device_tlul_plug_addr_reg_21_ (.rb(net461),
    .clk(clknet_1_0__leaf_u_spi_device_tlul_plug_net617),
    .d1(net2359),
    .d2(net2343),
    .o1(net118),
    .o2(net119),
    .si1(net1332),
    .si2(net1333),
    .ssb(net1894));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_22__u_spi_device_tlul_plug_addr_reg_23_ (.rb(net461),
    .clk(clknet_1_0__leaf_u_spi_device_tlul_plug_net617),
    .d1(net2321),
    .d2(net2318),
    .o1(net120),
    .o2(net121),
    .si1(net1334),
    .si2(net1335),
    .ssb(net1895));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_24__u_spi_device_tlul_plug_addr_reg_25_ (.rb(net461),
    .clk(clknet_1_1__leaf_u_spi_device_tlul_plug_net617),
    .d1(net2357),
    .d2(net2341),
    .o1(net122),
    .o2(net123),
    .si1(net1336),
    .si2(net1337),
    .ssb(net1896));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_26__u_spi_device_tlul_plug_addr_reg_27_ (.rb(net461),
    .clk(clknet_1_1__leaf_u_spi_device_tlul_plug_net617),
    .d1(net2369),
    .d2(net2363),
    .o1(net124),
    .o2(net125),
    .si1(net1338),
    .si2(net1339),
    .ssb(net1897));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_28__u_spi_device_tlul_plug_addr_reg_29_ (.rb(net461),
    .clk(clknet_1_1__leaf_u_spi_device_tlul_plug_net617),
    .d1(net2336),
    .d2(net2325),
    .o1(net126),
    .o2(net127),
    .si1(net1340),
    .si2(net1341),
    .ssb(net1898));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_2__u_spi_device_tlul_plug_addr_reg_3_ (.rb(net461),
    .clk(clknet_1_1__leaf_u_spi_device_tlul_plug_net611),
    .d1(addr_sync[2]),
    .d2(addr_sync[3]),
    .o1(net100),
    .o2(net101),
    .si1(net1342),
    .si2(net1343),
    .ssb(net1899));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_30__u_spi_device_tlul_plug_addr_reg_31_ (.rb(net463),
    .clk(clknet_1_1__leaf_u_spi_device_tlul_plug_net617),
    .d1(net2367),
    .d2(net2358),
    .o1(net129),
    .o2(net130),
    .si1(net1344),
    .si2(net1345),
    .ssb(net1900));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_4__u_spi_device_tlul_plug_addr_reg_5_ (.rb(net463),
    .clk(clknet_1_1__leaf_u_spi_device_tlul_plug_net611),
    .d1(addr_sync[4]),
    .d2(addr_sync[5]),
    .o1(net102),
    .o2(net103),
    .si1(net1346),
    .si2(net1347),
    .ssb(net1901));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_6__u_spi_device_tlul_plug_addr_reg_7_ (.rb(net463),
    .clk(clknet_1_1__leaf_u_spi_device_tlul_plug_net611),
    .d1(addr_sync[6]),
    .d2(addr_sync[7]),
    .o1(net104),
    .o2(net105),
    .si1(net1348),
    .si2(net1349),
    .ssb(net1902));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_addr_reg_8__u_spi_device_tlul_plug_addr_reg_9_ (.rb(net455),
    .clk(clknet_1_0__leaf_u_spi_device_tlul_plug_net611),
    .d1(net2331),
    .d2(net2323),
    .o1(net106),
    .o2(net107),
    .si1(net1350),
    .si2(net1351),
    .ssb(net1903));
 b15cilb05ah1n02x3 u_spi_device_tlul_plug_clk_gate_addr_reg_0_latch (.clk(clknet_2_3_0_clk_i),
    .clkout(u_spi_device_tlul_plug_net617),
    .en(u_spi_device_tlul_plug_N61),
    .te(net1352));
 b15cilb05ah1n02x3 u_spi_device_tlul_plug_clk_gate_addr_reg_latch (.clk(clknet_2_3_0_clk_i),
    .clkout(u_spi_device_tlul_plug_net611),
    .en(u_spi_device_tlul_plug_N61),
    .te(net1353));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_state_reg_1__u_spi_device_tlul_plug_u_tlul_adapter_host_g_multiple_reqs_source_q_reg_0_ (.rb(net438),
    .clk(clknet_2_1_0_clk_i),
    .d1(net2348),
    .d2(n604),
    .o1(u_spi_device_tlul_plug_state[1]),
    .o2(net131),
    .si1(net1354),
    .si2(net1355),
    .ssb(net1904));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_u_tlul_adapter_host_intg_err_q_reg_u_spi_device_tlul_plug_wdata_reg_0_ (.rb(net448),
    .clk(clknet_2_1_0_clk_i),
    .d1(n1456),
    .d2(u_spi_device_tlul_plug_wdata_next[0]),
    .o1(n1455),
    .o2(net68),
    .si1(net1356),
    .si2(net1357),
    .ssb(net1905));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_11__u_spi_device_tlul_plug_wdata_reg_12_ (.rb(net441),
    .clk(clknet_2_1_0_clk_i),
    .d1(u_spi_device_tlul_plug_wdata_next[11]),
    .d2(u_spi_device_tlul_plug_wdata_next[12]),
    .o1(net79),
    .o2(net80),
    .si1(net1358),
    .si2(net1359),
    .ssb(net1906));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_13__u_spi_device_tlul_plug_wdata_reg_14_ (.rb(net449),
    .clk(clknet_2_2_0_clk_i),
    .d1(u_spi_device_tlul_plug_wdata_next[13]),
    .d2(u_spi_device_tlul_plug_wdata_next[14]),
    .o1(net81),
    .o2(net82),
    .si1(net1360),
    .si2(net1361),
    .ssb(net1907));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_15__u_spi_device_tlul_plug_wdata_reg_16_ (.rb(net451),
    .clk(clknet_2_3_0_clk_i),
    .d1(u_spi_device_tlul_plug_wdata_next[15]),
    .d2(u_spi_device_tlul_plug_wdata_next[16]),
    .o1(net83),
    .o2(net84),
    .si1(net1362),
    .si2(net1363),
    .ssb(net1908));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_17__u_spi_device_tlul_plug_wdata_reg_18_ (.rb(net451),
    .clk(clknet_2_3_0_clk_i),
    .d1(u_spi_device_tlul_plug_wdata_next[17]),
    .d2(u_spi_device_tlul_plug_wdata_next[18]),
    .o1(net85),
    .o2(net86),
    .si1(net1364),
    .si2(net1365),
    .ssb(net1909));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_19__u_spi_device_tlul_plug_wdata_reg_20_ (.rb(net449),
    .clk(clknet_2_3_0_clk_i),
    .d1(u_spi_device_tlul_plug_wdata_next[19]),
    .d2(u_spi_device_tlul_plug_wdata_next[20]),
    .o1(net87),
    .o2(net88),
    .si1(net1366),
    .si2(net1367),
    .ssb(net1910));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_1__u_spi_device_tlul_plug_wdata_reg_2_ (.rb(net452),
    .clk(clknet_2_3_0_clk_i),
    .d1(u_spi_device_tlul_plug_wdata_next[1]),
    .d2(u_spi_device_tlul_plug_wdata_next[2]),
    .o1(net69),
    .o2(net70),
    .si1(net1368),
    .si2(net1369),
    .ssb(net1911));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_21__u_spi_device_tlul_plug_wdata_reg_22_ (.rb(net452),
    .clk(clknet_2_3_0_clk_i),
    .d1(u_spi_device_tlul_plug_wdata_next[21]),
    .d2(u_spi_device_tlul_plug_wdata_next[22]),
    .o1(net89),
    .o2(net90),
    .si1(net1370),
    .si2(net1371),
    .ssb(net1912));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_23__u_spi_device_tlul_plug_wdata_reg_24_ (.rb(net456),
    .clk(clknet_2_2_0_clk_i),
    .d1(net141),
    .d2(u_spi_device_tlul_plug_wdata_next[24]),
    .o1(net91),
    .o2(net92),
    .si1(net1372),
    .si2(net1373),
    .ssb(net1913));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_25__u_spi_device_tlul_plug_wdata_reg_26_ (.rb(net456),
    .clk(clknet_2_2_0_clk_i),
    .d1(u_spi_device_tlul_plug_wdata_next[25]),
    .d2(u_spi_device_tlul_plug_wdata_next[26]),
    .o1(net93),
    .o2(net94),
    .si1(net1374),
    .si2(net1375),
    .ssb(net1914));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_27__u_spi_device_tlul_plug_wdata_reg_28_ (.rb(net452),
    .clk(clknet_2_3_0_clk_i),
    .d1(u_spi_device_tlul_plug_wdata_next[27]),
    .d2(u_spi_device_tlul_plug_wdata_next[28]),
    .o1(net95),
    .o2(net96),
    .si1(net1376),
    .si2(net1377),
    .ssb(net1915));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_29__u_spi_device_tlul_plug_wdata_reg_30_ (.rb(net452),
    .clk(clknet_2_3_0_clk_i),
    .d1(u_spi_device_tlul_plug_wdata_next[29]),
    .d2(u_spi_device_tlul_plug_wdata_next[30]),
    .o1(net97),
    .o2(net98),
    .si1(net1378),
    .si2(net1379),
    .ssb(net1916));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_31__u_spi_device_tlul_plug_we_reg (.rb(net452),
    .clk(clknet_2_3_0_clk_i),
    .d1(u_spi_device_tlul_plug_wdata_next[31]),
    .d2(net168),
    .o1(net99),
    .o2(u_spi_device_tlul_plug_we),
    .si1(net1380),
    .si2(net1381),
    .ssb(net1917));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_3__u_spi_device_tlul_plug_wdata_reg_4_ (.rb(net441),
    .clk(clknet_2_1_0_clk_i),
    .d1(u_spi_device_tlul_plug_wdata_next[3]),
    .d2(u_spi_device_tlul_plug_wdata_next[4]),
    .o1(net71),
    .o2(net72),
    .si1(net1382),
    .si2(net1383),
    .ssb(net1918));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_5__u_spi_device_tlul_plug_wdata_reg_6_ (.rb(net438),
    .clk(clknet_2_1_0_clk_i),
    .d1(net142),
    .d2(u_spi_device_tlul_plug_wdata_next[6]),
    .o1(net73),
    .o2(net74),
    .si1(net1384),
    .si2(net1385),
    .ssb(net1919));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_7__u_spi_device_tlul_plug_wdata_reg_8_ (.rb(net449),
    .clk(clknet_2_2_0_clk_i),
    .d1(u_spi_device_tlul_plug_wdata_next[7]),
    .d2(u_spi_device_tlul_plug_wdata_next[8]),
    .o1(net75),
    .o2(net76),
    .si1(net1386),
    .si2(net1387),
    .ssb(net1920));
 b15fqy203ar1n02x5 u_spi_device_tlul_plug_wdata_reg_9__u_spi_device_tlul_plug_wdata_reg_10_ (.rb(net452),
    .clk(clknet_2_3_0_clk_i),
    .d1(u_spi_device_tlul_plug_wdata_next[9]),
    .d2(u_spi_device_tlul_plug_wdata_next[10]),
    .o1(net77),
    .o2(net78),
    .si1(net1388),
    .si2(net1389),
    .ssb(net1921));
 b15fqy00car1n02x5 u_syncro_cs_reg_reg_0_ (.clk(clknet_2_1_0_clk_i),
    .d(net427),
    .o(u_syncro_cs_reg_0_),
    .psb(net448),
    .si(net1390),
    .ssb(net1922));
 b15fqy00car1n06x5 u_syncro_cs_reg_reg_1_ (.clk(clknet_2_1_0_clk_i),
    .d(net2233),
    .psb(net448),
    .si(net1391),
    .ssb(net1923));
 b15fqy203ar1n02x5 u_syncro_rdwr_reg_reg_0__u_syncro_rdwr_reg_reg_1_ (.rb(net440),
    .clk(clknet_2_0_0_clk_i),
    .d1(net140),
    .d2(net2287),
    .o1(u_syncro_rdwr_reg_0_),
    .o2(rd_wr_sync),
    .si1(net1392),
    .si2(net1393),
    .ssb(net1924));
 b15fqy203ar1n02x5 u_syncro_valid_reg_reg_0__u_syncro_valid_reg_reg_1_ (.rb(net441),
    .clk(clknet_2_1_0_clk_i),
    .d1(ctrl_addr_valid),
    .d2(net2283),
    .o1(u_syncro_valid_reg[0]),
    .o2(u_syncro_valid_reg[1]),
    .si1(net1394),
    .si2(net1395),
    .ssb(net1925));
 b15fqy003ar1n02x5 u_syncro_valid_reg_reg_2_ (.rb(net441),
    .clk(clknet_2_1_0_clk_i),
    .d(net2319),
    .o(u_syncro_valid_reg[2]),
    .si(net1396),
    .ssb(net1926));
 b15cilb05ah1n02x3 u_txreg_clk_gate_counter_reg_latch (.clk(clknet_1_0__leaf_u_txreg_sclk_test),
    .clkout(u_txreg_net824),
    .en(u_txreg_N11),
    .te(net1397));
 b15cilb05ah1n02x3 u_txreg_clk_gate_counter_trgt_reg_latch (.clk(clknet_1_1__leaf_u_txreg_sclk_test),
    .clkout(u_txreg_net840),
    .en(net2337),
    .te(net1398));
 b15cilb05ah1n02x3 u_txreg_clk_gate_data_int_reg_0_latch (.clk(clknet_1_1__leaf_u_txreg_sclk_test),
    .clkout(u_txreg_net835),
    .en(u_txreg_N11),
    .te(net1399));
 b15cilb05ah1n02x3 u_txreg_clk_gate_data_int_reg_latch (.clk(clknet_1_0__leaf_u_txreg_sclk_test),
    .clkout(u_txreg_net830),
    .en(u_txreg_N11),
    .te(net1400));
 b15fqy203ar1n02x5 u_txreg_counter_reg_0__u_txreg_counter_reg_1_ (.rb(n3769),
    .clk(clknet_1_1__leaf_u_txreg_net824),
    .d1(u_txreg_N24),
    .d2(u_txreg_N25),
    .o1(u_txreg_counter[0]),
    .o2(u_txreg_counter[1]),
    .si1(net1401),
    .si2(net1402),
    .ssb(net1927));
 b15fqy203ar1n02x5 u_txreg_counter_reg_2__u_txreg_counter_reg_3_ (.rb(n3769),
    .clk(clknet_1_0__leaf_u_txreg_net824),
    .d1(u_txreg_N26),
    .d2(u_txreg_N27),
    .o1(u_txreg_counter[2]),
    .o2(u_txreg_counter[3]),
    .si1(net1403),
    .si2(net1404),
    .ssb(net1928));
 b15fqy203ar1n02x5 u_txreg_counter_reg_4__u_txreg_counter_reg_5_ (.rb(n3769),
    .clk(clknet_1_1__leaf_u_txreg_net824),
    .d1(u_txreg_N28),
    .d2(u_txreg_N29),
    .o1(u_txreg_counter[4]),
    .o2(u_txreg_counter[5]),
    .si1(net1405),
    .si2(net1406),
    .ssb(net1929));
 b15fqy203ar1n02x5 u_txreg_counter_reg_6__u_txreg_counter_reg_7_ (.rb(n3769),
    .clk(clknet_1_0__leaf_u_txreg_net824),
    .d1(u_txreg_N30),
    .d2(u_txreg_N31),
    .o1(u_txreg_counter[6]),
    .o2(u_txreg_counter[7]),
    .si1(net1407),
    .si2(net1408),
    .ssb(net1930));
 b15fqy00car1n02x5 u_txreg_counter_trgt_reg_0_ (.clk(clknet_1_0__leaf_u_txreg_net840),
    .d(net2494),
    .o(u_txreg_counter_trgt[0]),
    .psb(n3769),
    .si(net1409),
    .ssb(net1931));
 b15fqy00car1n02x5 u_txreg_counter_trgt_reg_1_ (.clk(clknet_1_0__leaf_u_txreg_net840),
    .d(net2480),
    .o(u_txreg_counter_trgt[1]),
    .psb(n3769),
    .si(net1410),
    .ssb(net1932));
 b15fqy00car1n02x5 u_txreg_counter_trgt_reg_2_ (.clk(clknet_1_0__leaf_u_txreg_net840),
    .d(net2492),
    .o(u_txreg_counter_trgt[2]),
    .psb(n3769),
    .si(net1411),
    .ssb(net1933));
 b15fqy203ar1n02x5 u_txreg_counter_trgt_reg_3__u_txreg_counter_trgt_reg_4_ (.rb(n3769),
    .clk(clknet_1_1__leaf_u_txreg_net840),
    .d1(net2216),
    .d2(net2490),
    .o1(u_txreg_counter_trgt[3]),
    .o2(u_txreg_counter_trgt[4]),
    .si1(net1412),
    .si2(net1413),
    .ssb(net1934));
 b15fqy203ar1n02x5 u_txreg_counter_trgt_reg_5__u_txreg_counter_trgt_reg_6_ (.rb(n3769),
    .clk(clknet_1_1__leaf_u_txreg_net840),
    .d1(net2486),
    .d2(net2482),
    .o1(u_txreg_counter_trgt[5]),
    .o2(u_txreg_counter_trgt[6]),
    .si1(net1414),
    .si2(net1415),
    .ssb(net1935));
 b15fqy003ar1n02x5 u_txreg_counter_trgt_reg_7_ (.rb(n3769),
    .clk(clknet_1_1__leaf_u_txreg_net840),
    .d(net2446),
    .o(u_txreg_counter_trgt[7]),
    .si(net1416),
    .ssb(net1936));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_0__u_txreg_data_int_reg_1_ (.rb(n3778),
    .clk(clknet_1_0__leaf_u_txreg_net830),
    .d1(net2197),
    .d2(net2313),
    .o1(u_txreg_data_int[0]),
    .o2(u_txreg_data_int[1]),
    .si1(net1417),
    .si2(net1418),
    .ssb(net1937));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_10__u_txreg_data_int_reg_11_ (.rb(n3772),
    .clk(clknet_1_1__leaf_u_txreg_net830),
    .d1(u_txreg_N44),
    .d2(net2175),
    .o1(u_txreg_data_int[10]),
    .o2(u_txreg_data_int[11]),
    .si1(net1419),
    .si2(net1420),
    .ssb(net1938));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_12__u_txreg_data_int_reg_13_ (.rb(n3773),
    .clk(clknet_1_1__leaf_u_txreg_net830),
    .d1(net2178),
    .d2(net2185),
    .o1(u_txreg_data_int[12]),
    .o2(u_txreg_data_int[13]),
    .si1(net1421),
    .si2(net1422),
    .ssb(net1939));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_14__u_txreg_data_int_reg_15_ (.rb(n3773),
    .clk(clknet_1_1__leaf_u_txreg_net830),
    .d1(net2203),
    .d2(net2191),
    .o1(u_txreg_data_int[14]),
    .o2(u_txreg_data_int[15]),
    .si1(net1423),
    .si2(net1424),
    .ssb(net1940));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_16__u_txreg_data_int_reg_17_ (.rb(n3771),
    .clk(clknet_1_0__leaf_u_txreg_net835),
    .d1(net2154),
    .d2(net2200),
    .o1(u_txreg_data_int[16]),
    .o2(u_txreg_data_int[17]),
    .si1(net1425),
    .si2(net1426),
    .ssb(net1941));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_18__u_txreg_data_int_reg_19_ (.rb(n3771),
    .clk(clknet_1_1__leaf_u_txreg_net835),
    .d1(net2157),
    .d2(net2143),
    .o1(u_txreg_data_int[18]),
    .o2(u_txreg_data_int[19]),
    .si1(net1427),
    .si2(net1428),
    .ssb(net1942));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_20__u_txreg_data_int_reg_21_ (.rb(n3771),
    .clk(clknet_1_1__leaf_u_txreg_net835),
    .d1(net2172),
    .d2(net2188),
    .o1(u_txreg_data_int[20]),
    .o2(u_txreg_data_int[21]),
    .si1(net1429),
    .si2(net1430),
    .ssb(net1943));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_22__u_txreg_data_int_reg_23_ (.rb(n3771),
    .clk(clknet_1_0__leaf_u_txreg_net835),
    .d1(u_txreg_N56),
    .d2(net2211),
    .o1(u_txreg_data_int[22]),
    .o2(u_txreg_data_int[23]),
    .si1(net1431),
    .si2(net1432),
    .ssb(net1944));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_24__u_txreg_data_int_reg_25_ (.rb(n3771),
    .clk(clknet_1_1__leaf_u_txreg_net835),
    .d1(net2146),
    .d2(net2165),
    .o1(u_txreg_data_int[24]),
    .o2(u_txreg_data_int[25]),
    .si1(net1433),
    .si2(net1434),
    .ssb(net1945));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_26__u_txreg_data_int_reg_27_ (.rb(n3771),
    .clk(clknet_1_0__leaf_u_txreg_net835),
    .d1(net2181),
    .d2(net2168),
    .o1(u_txreg_data_int[26]),
    .o2(u_txreg_data_int[27]),
    .si1(net1435),
    .si2(net1436),
    .ssb(net1946));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_28__u_txreg_data_int_reg_29_ (.rb(n3771),
    .clk(clknet_1_0__leaf_u_txreg_net835),
    .d1(net2236),
    .d2(net2301),
    .o1(u_txreg_data_int[28]),
    .o2(u_txreg_data_int[29]),
    .si1(net1437),
    .si2(net1438),
    .ssb(net1947));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_2__u_txreg_data_int_reg_3_ (.rb(n3778),
    .clk(clknet_1_0__leaf_u_txreg_net830),
    .d1(net2316),
    .d2(net2215),
    .o1(u_txreg_data_int[2]),
    .o2(u_txreg_data_int[3]),
    .si1(net1439),
    .si2(net1440),
    .ssb(net1948));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_30__u_txreg_data_int_reg_31_ (.rb(n3773),
    .clk(clknet_1_1__leaf_u_txreg_net835),
    .d1(u_txreg_N64),
    .d2(u_txreg_N65),
    .o1(u_txreg_data_int[30]),
    .o2(u_txreg_data_int[31]),
    .si1(net1441),
    .si2(net1442),
    .ssb(net1949));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_4__u_txreg_data_int_reg_5_ (.rb(n3772),
    .clk(clknet_1_0__leaf_u_txreg_net830),
    .d1(u_txreg_N38),
    .d2(net2224),
    .o1(u_txreg_data_int[4]),
    .o2(u_txreg_data_int[5]),
    .si1(net1443),
    .si2(net1444),
    .ssb(net1950));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_6__u_txreg_data_int_reg_7_ (.rb(n3772),
    .clk(clknet_1_0__leaf_u_txreg_net830),
    .d1(net2221),
    .d2(net2227),
    .o1(u_txreg_data_int[6]),
    .o2(u_txreg_data_int[7]),
    .si1(net1445),
    .si2(net1446),
    .ssb(net1951));
 b15fqy203ar1n02x5 u_txreg_data_int_reg_8__u_txreg_data_int_reg_9_ (.rb(n3772),
    .clk(clknet_1_1__leaf_u_txreg_net830),
    .d1(net2240),
    .d2(net2194),
    .o1(u_txreg_data_int[8]),
    .o2(u_txreg_data_int[9]),
    .si1(net1447),
    .si2(net1448),
    .ssb(net1952));
 b15fqy043ar1n02x5 u_txreg_running_reg (.clk(clknet_1_1__leaf_u_txreg_sclk_test),
    .d(tx_counter_upd),
    .den(u_txreg_N10),
    .o(u_txreg_running),
    .rb(net365),
    .si(net1449),
    .ssb(net1953));
 b15tihi00an1n03x5 U3029_1450 (.o(net1450));
 b15inv000ar1n03x5 U3002_1 (.a(clknet_3_0__leaf_spi_sclk),
    .o1(net1954));
 b15ztpn00an1n08x5 PHY_96 ();
 b15ztpn00an1n08x5 PHY_97 ();
 b15ztpn00an1n08x5 PHY_98 ();
 b15ztpn00an1n08x5 PHY_99 ();
 b15ztpn00an1n08x5 PHY_100 ();
 b15ztpn00an1n08x5 PHY_101 ();
 b15ztpn00an1n08x5 PHY_102 ();
 b15ztpn00an1n08x5 PHY_103 ();
 b15ztpn00an1n08x5 PHY_104 ();
 b15ztpn00an1n08x5 PHY_105 ();
 b15ztpn00an1n08x5 PHY_106 ();
 b15ztpn00an1n08x5 PHY_107 ();
 b15ztpn00an1n08x5 PHY_108 ();
 b15ztpn00an1n08x5 PHY_109 ();
 b15ztpn00an1n08x5 PHY_110 ();
 b15ztpn00an1n08x5 PHY_111 ();
 b15ztpn00an1n08x5 PHY_112 ();
 b15ztpn00an1n08x5 PHY_113 ();
 b15ztpn00an1n08x5 PHY_114 ();
 b15ztpn00an1n08x5 PHY_115 ();
 b15ztpn00an1n08x5 PHY_116 ();
 b15ztpn00an1n08x5 PHY_117 ();
 b15ztpn00an1n08x5 PHY_118 ();
 b15ztpn00an1n08x5 PHY_119 ();
 b15ztpn00an1n08x5 PHY_120 ();
 b15ztpn00an1n08x5 PHY_121 ();
 b15ztpn00an1n08x5 PHY_122 ();
 b15ztpn00an1n08x5 PHY_123 ();
 b15ztpn00an1n08x5 PHY_124 ();
 b15ztpn00an1n08x5 PHY_125 ();
 b15ztpn00an1n08x5 PHY_126 ();
 b15ztpn00an1n08x5 PHY_127 ();
 b15ztpn00an1n08x5 PHY_128 ();
 b15ztpn00an1n08x5 PHY_129 ();
 b15ztpn00an1n08x5 PHY_130 ();
 b15ztpn00an1n08x5 PHY_131 ();
 b15ztpn00an1n08x5 PHY_132 ();
 b15ztpn00an1n08x5 PHY_133 ();
 b15ztpn00an1n08x5 PHY_134 ();
 b15ztpn00an1n08x5 PHY_135 ();
 b15ztpn00an1n08x5 PHY_136 ();
 b15ztpn00an1n08x5 PHY_137 ();
 b15ztpn00an1n08x5 PHY_138 ();
 b15ztpn00an1n08x5 PHY_139 ();
 b15ztpn00an1n08x5 PHY_140 ();
 b15ztpn00an1n08x5 PHY_141 ();
 b15ztpn00an1n08x5 PHY_142 ();
 b15ztpn00an1n08x5 PHY_143 ();
 b15ztpn00an1n08x5 PHY_144 ();
 b15ztpn00an1n08x5 PHY_145 ();
 b15ztpn00an1n08x5 PHY_146 ();
 b15ztpn00an1n08x5 PHY_147 ();
 b15ztpn00an1n08x5 PHY_148 ();
 b15ztpn00an1n08x5 PHY_149 ();
 b15ztpn00an1n08x5 PHY_150 ();
 b15ztpn00an1n08x5 PHY_151 ();
 b15ztpn00an1n08x5 PHY_152 ();
 b15ztpn00an1n08x5 PHY_153 ();
 b15ztpn00an1n08x5 PHY_154 ();
 b15ztpn00an1n08x5 PHY_155 ();
 b15ztpn00an1n08x5 PHY_156 ();
 b15ztpn00an1n08x5 PHY_157 ();
 b15ztpn00an1n08x5 PHY_158 ();
 b15ztpn00an1n08x5 PHY_159 ();
 b15ztpn00an1n08x5 PHY_160 ();
 b15ztpn00an1n08x5 PHY_161 ();
 b15ztpn00an1n08x5 PHY_162 ();
 b15ztpn00an1n08x5 PHY_163 ();
 b15ztpn00an1n08x5 PHY_164 ();
 b15ztpn00an1n08x5 PHY_165 ();
 b15ztpn00an1n08x5 PHY_166 ();
 b15ztpn00an1n08x5 PHY_167 ();
 b15ztpn00an1n08x5 PHY_168 ();
 b15ztpn00an1n08x5 PHY_169 ();
 b15ztpn00an1n08x5 PHY_170 ();
 b15ztpn00an1n08x5 PHY_171 ();
 b15ztpn00an1n08x5 PHY_172 ();
 b15ztpn00an1n08x5 PHY_173 ();
 b15ztpn00an1n08x5 PHY_174 ();
 b15ztpn00an1n08x5 PHY_175 ();
 b15ztpn00an1n08x5 PHY_176 ();
 b15ztpn00an1n08x5 PHY_177 ();
 b15ztpn00an1n08x5 PHY_178 ();
 b15ztpn00an1n08x5 PHY_179 ();
 b15ztpn00an1n08x5 PHY_180 ();
 b15ztpn00an1n08x5 PHY_181 ();
 b15ztpn00an1n08x5 PHY_182 ();
 b15ztpn00an1n08x5 PHY_183 ();
 b15ztpn00an1n08x5 PHY_184 ();
 b15ztpn00an1n08x5 PHY_185 ();
 b15ztpn00an1n08x5 PHY_186 ();
 b15ztpn00an1n08x5 PHY_187 ();
 b15ztpn00an1n08x5 PHY_188 ();
 b15ztpn00an1n08x5 PHY_189 ();
 b15ztpn00an1n08x5 PHY_190 ();
 b15ztpn00an1n08x5 PHY_191 ();
 b15ztpn00an1n08x5 PHY_192 ();
 b15ztpn00an1n08x5 PHY_193 ();
 b15ztpn00an1n08x5 PHY_194 ();
 b15ztpn00an1n08x5 PHY_195 ();
 b15ztpn00an1n08x5 PHY_196 ();
 b15ztpn00an1n08x5 PHY_197 ();
 b15ztpn00an1n08x5 PHY_198 ();
 b15ztpn00an1n08x5 PHY_199 ();
 b15ztpn00an1n08x5 PHY_200 ();
 b15ztpn00an1n08x5 PHY_201 ();
 b15ztpn00an1n08x5 PHY_202 ();
 b15ztpn00an1n08x5 PHY_203 ();
 b15ztpn00an1n08x5 PHY_204 ();
 b15ztpn00an1n08x5 PHY_205 ();
 b15ztpn00an1n08x5 PHY_206 ();
 b15ztpn00an1n08x5 PHY_207 ();
 b15ztpn00an1n08x5 PHY_208 ();
 b15ztpn00an1n08x5 PHY_209 ();
 b15ztpn00an1n08x5 PHY_210 ();
 b15ztpn00an1n08x5 PHY_211 ();
 b15ztpn00an1n08x5 PHY_212 ();
 b15ztpn00an1n08x5 PHY_213 ();
 b15ztpn00an1n08x5 PHY_214 ();
 b15ztpn00an1n08x5 PHY_215 ();
 b15ztpn00an1n08x5 PHY_216 ();
 b15ztpn00an1n08x5 PHY_217 ();
 b15ztpn00an1n08x5 PHY_218 ();
 b15ztpn00an1n08x5 PHY_219 ();
 b15ztpn00an1n08x5 PHY_220 ();
 b15ztpn00an1n08x5 PHY_221 ();
 b15ztpn00an1n08x5 PHY_222 ();
 b15ztpn00an1n08x5 PHY_223 ();
 b15ztpn00an1n08x5 PHY_224 ();
 b15ztpn00an1n08x5 PHY_225 ();
 b15ztpn00an1n08x5 PHY_226 ();
 b15ztpn00an1n08x5 PHY_227 ();
 b15ztpn00an1n08x5 PHY_228 ();
 b15ztpn00an1n08x5 PHY_229 ();
 b15ztpn00an1n08x5 PHY_230 ();
 b15ztpn00an1n08x5 PHY_231 ();
 b15ztpn00an1n08x5 PHY_232 ();
 b15ztpn00an1n08x5 PHY_233 ();
 b15ztpn00an1n08x5 PHY_234 ();
 b15ztpn00an1n08x5 PHY_235 ();
 b15ztpn00an1n08x5 PHY_236 ();
 b15ztpn00an1n08x5 PHY_237 ();
 b15ztpn00an1n08x5 PHY_238 ();
 b15ztpn00an1n08x5 PHY_239 ();
 b15ztpn00an1n08x5 PHY_240 ();
 b15ztpn00an1n08x5 PHY_241 ();
 b15ztpn00an1n08x5 PHY_242 ();
 b15ztpn00an1n08x5 PHY_243 ();
 b15ztpn00an1n08x5 PHY_244 ();
 b15ztpn00an1n08x5 PHY_245 ();
 b15ztpn00an1n08x5 PHY_246 ();
 b15ztpn00an1n08x5 PHY_247 ();
 b15ztpn00an1n08x5 PHY_248 ();
 b15ztpn00an1n08x5 PHY_249 ();
 b15ztpn00an1n08x5 PHY_250 ();
 b15ztpn00an1n08x5 PHY_251 ();
 b15ztpn00an1n08x5 PHY_252 ();
 b15ztpn00an1n08x5 PHY_253 ();
 b15ztpn00an1n08x5 PHY_254 ();
 b15ztpn00an1n08x5 PHY_255 ();
 b15ztpn00an1n08x5 PHY_256 ();
 b15ztpn00an1n08x5 PHY_257 ();
 b15ztpn00an1n08x5 PHY_258 ();
 b15ztpn00an1n08x5 PHY_259 ();
 b15ztpn00an1n08x5 PHY_260 ();
 b15ztpn00an1n08x5 PHY_261 ();
 b15ztpn00an1n08x5 PHY_262 ();
 b15ztpn00an1n08x5 PHY_263 ();
 b15ztpn00an1n08x5 PHY_264 ();
 b15ztpn00an1n08x5 PHY_265 ();
 b15ztpn00an1n08x5 PHY_266 ();
 b15ztpn00an1n08x5 PHY_267 ();
 b15ztpn00an1n08x5 PHY_268 ();
 b15ztpn00an1n08x5 PHY_269 ();
 b15ztpn00an1n08x5 PHY_270 ();
 b15ztpn00an1n08x5 PHY_271 ();
 b15ztpn00an1n08x5 PHY_272 ();
 b15ztpn00an1n08x5 PHY_273 ();
 b15ztpn00an1n08x5 PHY_274 ();
 b15ztpn00an1n08x5 PHY_275 ();
 b15ztpn00an1n08x5 PHY_276 ();
 b15ztpn00an1n08x5 PHY_277 ();
 b15ztpn00an1n08x5 PHY_278 ();
 b15ztpn00an1n08x5 PHY_279 ();
 b15ztpn00an1n08x5 PHY_280 ();
 b15ztpn00an1n08x5 PHY_281 ();
 b15ztpn00an1n08x5 PHY_282 ();
 b15ztpn00an1n08x5 PHY_283 ();
 b15ztpn00an1n08x5 PHY_284 ();
 b15ztpn00an1n08x5 PHY_285 ();
 b15ztpn00an1n08x5 PHY_286 ();
 b15ztpn00an1n08x5 PHY_287 ();
 b15ztpn00an1n08x5 PHY_288 ();
 b15ztpn00an1n08x5 PHY_289 ();
 b15ztpn00an1n08x5 PHY_290 ();
 b15ztpn00an1n08x5 PHY_291 ();
 b15ztpn00an1n08x5 PHY_292 ();
 b15ztpn00an1n08x5 PHY_293 ();
 b15ztpn00an1n08x5 PHY_294 ();
 b15ztpn00an1n08x5 PHY_295 ();
 b15ztpn00an1n08x5 PHY_296 ();
 b15ztpn00an1n08x5 PHY_297 ();
 b15ztpn00an1n08x5 PHY_298 ();
 b15ztpn00an1n08x5 PHY_299 ();
 b15ztpn00an1n08x5 PHY_300 ();
 b15ztpn00an1n08x5 PHY_301 ();
 b15ztpn00an1n08x5 PHY_302 ();
 b15ztpn00an1n08x5 PHY_303 ();
 b15ztpn00an1n08x5 PHY_304 ();
 b15ztpn00an1n08x5 PHY_305 ();
 b15ztpn00an1n08x5 PHY_306 ();
 b15ztpn00an1n08x5 PHY_307 ();
 b15ztpn00an1n08x5 PHY_308 ();
 b15ztpn00an1n08x5 PHY_309 ();
 b15ztpn00an1n08x5 PHY_310 ();
 b15ztpn00an1n08x5 PHY_311 ();
 b15ztpn00an1n08x5 PHY_312 ();
 b15ztpn00an1n08x5 PHY_313 ();
 b15ztpn00an1n08x5 PHY_314 ();
 b15ztpn00an1n08x5 PHY_315 ();
 b15ztpn00an1n08x5 PHY_316 ();
 b15ztpn00an1n08x5 PHY_317 ();
 b15ztpn00an1n08x5 PHY_318 ();
 b15ztpn00an1n08x5 PHY_319 ();
 b15ztpn00an1n08x5 PHY_320 ();
 b15ztpn00an1n08x5 PHY_321 ();
 b15ztpn00an1n08x5 PHY_322 ();
 b15ztpn00an1n08x5 PHY_323 ();
 b15ztpn00an1n08x5 PHY_324 ();
 b15ztpn00an1n08x5 PHY_325 ();
 b15ztpn00an1n08x5 PHY_326 ();
 b15ztpn00an1n08x5 PHY_327 ();
 b15ztpn00an1n08x5 PHY_328 ();
 b15ztpn00an1n08x5 PHY_329 ();
 b15ztpn00an1n08x5 PHY_330 ();
 b15ztpn00an1n08x5 PHY_331 ();
 b15ztpn00an1n08x5 PHY_332 ();
 b15ztpn00an1n08x5 PHY_333 ();
 b15ztpn00an1n08x5 PHY_334 ();
 b15ztpn00an1n08x5 PHY_335 ();
 b15ztpn00an1n08x5 PHY_336 ();
 b15ztpn00an1n08x5 PHY_337 ();
 b15ztpn00an1n08x5 PHY_338 ();
 b15ztpn00an1n08x5 PHY_339 ();
 b15ztpn00an1n08x5 PHY_340 ();
 b15ztpn00an1n08x5 PHY_341 ();
 b15ztpn00an1n08x5 PHY_342 ();
 b15ztpn00an1n08x5 PHY_343 ();
 b15ztpn00an1n08x5 PHY_344 ();
 b15ztpn00an1n08x5 PHY_345 ();
 b15ztpn00an1n08x5 PHY_346 ();
 b15ztpn00an1n08x5 PHY_347 ();
 b15ztpn00an1n08x5 PHY_348 ();
 b15ztpn00an1n08x5 PHY_349 ();
 b15ztpn00an1n08x5 PHY_350 ();
 b15ztpn00an1n08x5 PHY_351 ();
 b15ztpn00an1n08x5 PHY_352 ();
 b15ztpn00an1n08x5 PHY_353 ();
 b15ztpn00an1n08x5 PHY_354 ();
 b15ztpn00an1n08x5 PHY_355 ();
 b15ztpn00an1n08x5 PHY_356 ();
 b15ztpn00an1n08x5 PHY_357 ();
 b15ztpn00an1n08x5 PHY_358 ();
 b15ztpn00an1n08x5 PHY_359 ();
 b15ztpn00an1n08x5 PHY_360 ();
 b15ztpn00an1n08x5 PHY_361 ();
 b15ztpn00an1n08x5 PHY_362 ();
 b15ztpn00an1n08x5 PHY_363 ();
 b15ztpn00an1n08x5 PHY_364 ();
 b15ztpn00an1n08x5 PHY_365 ();
 b15ztpn00an1n08x5 PHY_366 ();
 b15ztpn00an1n08x5 PHY_367 ();
 b15ztpn00an1n08x5 PHY_368 ();
 b15ztpn00an1n08x5 PHY_369 ();
 b15ztpn00an1n08x5 PHY_370 ();
 b15ztpn00an1n08x5 PHY_371 ();
 b15ztpn00an1n08x5 PHY_372 ();
 b15ztpn00an1n08x5 PHY_373 ();
 b15ztpn00an1n08x5 PHY_374 ();
 b15ztpn00an1n08x5 PHY_375 ();
 b15ztpn00an1n08x5 PHY_376 ();
 b15ztpn00an1n08x5 PHY_377 ();
 b15ztpn00an1n08x5 PHY_378 ();
 b15ztpn00an1n08x5 PHY_379 ();
 b15ztpn00an1n08x5 PHY_380 ();
 b15ztpn00an1n08x5 PHY_381 ();
 b15ztpn00an1n08x5 PHY_382 ();
 b15ztpn00an1n08x5 PHY_383 ();
 b15ztpn00an1n08x5 PHY_384 ();
 b15ztpn00an1n08x5 PHY_385 ();
 b15ztpn00an1n08x5 PHY_386 ();
 b15ztpn00an1n08x5 PHY_387 ();
 b15ztpn00an1n08x5 PHY_388 ();
 b15ztpn00an1n08x5 PHY_389 ();
 b15ztpn00an1n08x5 TAP_390 ();
 b15ztpn00an1n08x5 TAP_391 ();
 b15ztpn00an1n08x5 TAP_392 ();
 b15ztpn00an1n08x5 TAP_393 ();
 b15ztpn00an1n08x5 TAP_394 ();
 b15ztpn00an1n08x5 TAP_395 ();
 b15ztpn00an1n08x5 TAP_396 ();
 b15ztpn00an1n08x5 TAP_397 ();
 b15ztpn00an1n08x5 TAP_398 ();
 b15ztpn00an1n08x5 TAP_399 ();
 b15ztpn00an1n08x5 TAP_400 ();
 b15ztpn00an1n08x5 TAP_401 ();
 b15ztpn00an1n08x5 TAP_402 ();
 b15ztpn00an1n08x5 TAP_403 ();
 b15ztpn00an1n08x5 TAP_404 ();
 b15ztpn00an1n08x5 TAP_405 ();
 b15ztpn00an1n08x5 TAP_406 ();
 b15ztpn00an1n08x5 TAP_407 ();
 b15ztpn00an1n08x5 TAP_408 ();
 b15ztpn00an1n08x5 TAP_409 ();
 b15ztpn00an1n08x5 TAP_410 ();
 b15ztpn00an1n08x5 TAP_411 ();
 b15ztpn00an1n08x5 TAP_412 ();
 b15ztpn00an1n08x5 TAP_413 ();
 b15ztpn00an1n08x5 TAP_414 ();
 b15ztpn00an1n08x5 TAP_415 ();
 b15ztpn00an1n08x5 TAP_416 ();
 b15ztpn00an1n08x5 TAP_417 ();
 b15ztpn00an1n08x5 TAP_418 ();
 b15ztpn00an1n08x5 TAP_419 ();
 b15ztpn00an1n08x5 TAP_420 ();
 b15ztpn00an1n08x5 TAP_421 ();
 b15ztpn00an1n08x5 TAP_422 ();
 b15ztpn00an1n08x5 TAP_423 ();
 b15ztpn00an1n08x5 TAP_424 ();
 b15ztpn00an1n08x5 TAP_425 ();
 b15ztpn00an1n08x5 TAP_426 ();
 b15ztpn00an1n08x5 TAP_427 ();
 b15ztpn00an1n08x5 TAP_428 ();
 b15ztpn00an1n08x5 TAP_429 ();
 b15ztpn00an1n08x5 TAP_430 ();
 b15ztpn00an1n08x5 TAP_431 ();
 b15ztpn00an1n08x5 TAP_432 ();
 b15ztpn00an1n08x5 TAP_433 ();
 b15ztpn00an1n08x5 TAP_434 ();
 b15ztpn00an1n08x5 TAP_435 ();
 b15ztpn00an1n08x5 TAP_436 ();
 b15ztpn00an1n08x5 TAP_437 ();
 b15ztpn00an1n08x5 TAP_438 ();
 b15ztpn00an1n08x5 TAP_439 ();
 b15ztpn00an1n08x5 TAP_440 ();
 b15ztpn00an1n08x5 TAP_441 ();
 b15ztpn00an1n08x5 TAP_442 ();
 b15ztpn00an1n08x5 TAP_443 ();
 b15ztpn00an1n08x5 TAP_444 ();
 b15ztpn00an1n08x5 TAP_445 ();
 b15ztpn00an1n08x5 TAP_446 ();
 b15ztpn00an1n08x5 TAP_447 ();
 b15ztpn00an1n08x5 TAP_448 ();
 b15ztpn00an1n08x5 TAP_449 ();
 b15ztpn00an1n08x5 TAP_450 ();
 b15ztpn00an1n08x5 TAP_451 ();
 b15ztpn00an1n08x5 TAP_452 ();
 b15ztpn00an1n08x5 TAP_453 ();
 b15ztpn00an1n08x5 TAP_454 ();
 b15ztpn00an1n08x5 TAP_455 ();
 b15ztpn00an1n08x5 TAP_456 ();
 b15ztpn00an1n08x5 TAP_457 ();
 b15ztpn00an1n08x5 TAP_458 ();
 b15ztpn00an1n08x5 TAP_459 ();
 b15ztpn00an1n08x5 TAP_460 ();
 b15ztpn00an1n08x5 TAP_461 ();
 b15ztpn00an1n08x5 TAP_462 ();
 b15ztpn00an1n08x5 TAP_463 ();
 b15ztpn00an1n08x5 TAP_464 ();
 b15ztpn00an1n08x5 TAP_465 ();
 b15ztpn00an1n08x5 TAP_466 ();
 b15ztpn00an1n08x5 TAP_467 ();
 b15ztpn00an1n08x5 TAP_468 ();
 b15ztpn00an1n08x5 TAP_469 ();
 b15ztpn00an1n08x5 TAP_470 ();
 b15ztpn00an1n08x5 TAP_471 ();
 b15ztpn00an1n08x5 TAP_472 ();
 b15ztpn00an1n08x5 TAP_473 ();
 b15ztpn00an1n08x5 TAP_474 ();
 b15ztpn00an1n08x5 TAP_475 ();
 b15ztpn00an1n08x5 TAP_476 ();
 b15ztpn00an1n08x5 TAP_477 ();
 b15ztpn00an1n08x5 TAP_478 ();
 b15ztpn00an1n08x5 TAP_479 ();
 b15ztpn00an1n08x5 TAP_480 ();
 b15ztpn00an1n08x5 TAP_481 ();
 b15ztpn00an1n08x5 TAP_482 ();
 b15ztpn00an1n08x5 TAP_483 ();
 b15ztpn00an1n08x5 TAP_484 ();
 b15ztpn00an1n08x5 TAP_485 ();
 b15ztpn00an1n08x5 TAP_486 ();
 b15ztpn00an1n08x5 TAP_487 ();
 b15ztpn00an1n08x5 TAP_488 ();
 b15ztpn00an1n08x5 TAP_489 ();
 b15ztpn00an1n08x5 TAP_490 ();
 b15ztpn00an1n08x5 TAP_491 ();
 b15ztpn00an1n08x5 TAP_492 ();
 b15ztpn00an1n08x5 TAP_493 ();
 b15ztpn00an1n08x5 TAP_494 ();
 b15ztpn00an1n08x5 TAP_495 ();
 b15ztpn00an1n08x5 TAP_496 ();
 b15ztpn00an1n08x5 TAP_497 ();
 b15ztpn00an1n08x5 TAP_498 ();
 b15ztpn00an1n08x5 TAP_499 ();
 b15ztpn00an1n08x5 TAP_500 ();
 b15ztpn00an1n08x5 TAP_501 ();
 b15ztpn00an1n08x5 TAP_502 ();
 b15ztpn00an1n08x5 TAP_503 ();
 b15ztpn00an1n08x5 TAP_504 ();
 b15ztpn00an1n08x5 TAP_505 ();
 b15ztpn00an1n08x5 TAP_506 ();
 b15ztpn00an1n08x5 TAP_507 ();
 b15ztpn00an1n08x5 TAP_508 ();
 b15ztpn00an1n08x5 TAP_509 ();
 b15ztpn00an1n08x5 TAP_510 ();
 b15ztpn00an1n08x5 TAP_511 ();
 b15ztpn00an1n08x5 TAP_512 ();
 b15ztpn00an1n08x5 TAP_513 ();
 b15ztpn00an1n08x5 TAP_514 ();
 b15ztpn00an1n08x5 TAP_515 ();
 b15ztpn00an1n08x5 TAP_516 ();
 b15ztpn00an1n08x5 TAP_517 ();
 b15ztpn00an1n08x5 TAP_518 ();
 b15ztpn00an1n08x5 TAP_519 ();
 b15ztpn00an1n08x5 TAP_520 ();
 b15ztpn00an1n08x5 TAP_521 ();
 b15ztpn00an1n08x5 TAP_522 ();
 b15ztpn00an1n08x5 TAP_523 ();
 b15ztpn00an1n08x5 TAP_524 ();
 b15ztpn00an1n08x5 TAP_525 ();
 b15ztpn00an1n08x5 TAP_526 ();
 b15ztpn00an1n08x5 TAP_527 ();
 b15ztpn00an1n08x5 TAP_528 ();
 b15ztpn00an1n08x5 TAP_529 ();
 b15ztpn00an1n08x5 TAP_530 ();
 b15ztpn00an1n08x5 TAP_531 ();
 b15ztpn00an1n08x5 TAP_532 ();
 b15ztpn00an1n08x5 TAP_533 ();
 b15ztpn00an1n08x5 TAP_534 ();
 b15ztpn00an1n08x5 TAP_535 ();
 b15ztpn00an1n08x5 TAP_536 ();
 b15ztpn00an1n08x5 TAP_537 ();
 b15ztpn00an1n08x5 TAP_538 ();
 b15ztpn00an1n08x5 TAP_539 ();
 b15ztpn00an1n08x5 TAP_540 ();
 b15ztpn00an1n08x5 TAP_541 ();
 b15ztpn00an1n08x5 TAP_542 ();
 b15ztpn00an1n08x5 TAP_543 ();
 b15ztpn00an1n08x5 TAP_544 ();
 b15ztpn00an1n08x5 TAP_545 ();
 b15ztpn00an1n08x5 TAP_546 ();
 b15ztpn00an1n08x5 TAP_547 ();
 b15ztpn00an1n08x5 TAP_548 ();
 b15ztpn00an1n08x5 TAP_549 ();
 b15ztpn00an1n08x5 TAP_550 ();
 b15ztpn00an1n08x5 TAP_551 ();
 b15ztpn00an1n08x5 TAP_552 ();
 b15ztpn00an1n08x5 TAP_553 ();
 b15ztpn00an1n08x5 TAP_554 ();
 b15ztpn00an1n08x5 TAP_555 ();
 b15ztpn00an1n08x5 TAP_556 ();
 b15ztpn00an1n08x5 TAP_557 ();
 b15ztpn00an1n08x5 TAP_558 ();
 b15ztpn00an1n08x5 TAP_559 ();
 b15ztpn00an1n08x5 TAP_560 ();
 b15ztpn00an1n08x5 TAP_561 ();
 b15ztpn00an1n08x5 TAP_562 ();
 b15ztpn00an1n08x5 TAP_563 ();
 b15ztpn00an1n08x5 TAP_564 ();
 b15ztpn00an1n08x5 TAP_565 ();
 b15ztpn00an1n08x5 TAP_566 ();
 b15ztpn00an1n08x5 TAP_567 ();
 b15ztpn00an1n08x5 TAP_568 ();
 b15ztpn00an1n08x5 TAP_569 ();
 b15ztpn00an1n08x5 TAP_570 ();
 b15ztpn00an1n08x5 TAP_571 ();
 b15ztpn00an1n08x5 TAP_572 ();
 b15ztpn00an1n08x5 TAP_573 ();
 b15ztpn00an1n08x5 TAP_574 ();
 b15ztpn00an1n08x5 TAP_575 ();
 b15ztpn00an1n08x5 TAP_576 ();
 b15ztpn00an1n08x5 TAP_577 ();
 b15ztpn00an1n08x5 TAP_578 ();
 b15ztpn00an1n08x5 TAP_579 ();
 b15ztpn00an1n08x5 TAP_580 ();
 b15ztpn00an1n08x5 TAP_581 ();
 b15ztpn00an1n08x5 TAP_582 ();
 b15ztpn00an1n08x5 TAP_583 ();
 b15ztpn00an1n08x5 TAP_584 ();
 b15ztpn00an1n08x5 TAP_585 ();
 b15ztpn00an1n08x5 TAP_586 ();
 b15ztpn00an1n08x5 TAP_587 ();
 b15ztpn00an1n08x5 TAP_588 ();
 b15ztpn00an1n08x5 TAP_589 ();
 b15ztpn00an1n08x5 TAP_590 ();
 b15ztpn00an1n08x5 TAP_591 ();
 b15ztpn00an1n08x5 TAP_592 ();
 b15ztpn00an1n08x5 TAP_593 ();
 b15ztpn00an1n08x5 TAP_594 ();
 b15ztpn00an1n08x5 TAP_595 ();
 b15ztpn00an1n08x5 TAP_596 ();
 b15ztpn00an1n08x5 TAP_597 ();
 b15ztpn00an1n08x5 TAP_598 ();
 b15ztpn00an1n08x5 TAP_599 ();
 b15ztpn00an1n08x5 TAP_600 ();
 b15ztpn00an1n08x5 TAP_601 ();
 b15ztpn00an1n08x5 TAP_602 ();
 b15ztpn00an1n08x5 TAP_603 ();
 b15ztpn00an1n08x5 TAP_604 ();
 b15ztpn00an1n08x5 TAP_605 ();
 b15ztpn00an1n08x5 TAP_606 ();
 b15ztpn00an1n08x5 TAP_607 ();
 b15ztpn00an1n08x5 TAP_608 ();
 b15ztpn00an1n08x5 TAP_609 ();
 b15ztpn00an1n08x5 TAP_610 ();
 b15ztpn00an1n08x5 TAP_611 ();
 b15ztpn00an1n08x5 TAP_612 ();
 b15ztpn00an1n08x5 TAP_613 ();
 b15ztpn00an1n08x5 TAP_614 ();
 b15ztpn00an1n08x5 TAP_615 ();
 b15ztpn00an1n08x5 TAP_616 ();
 b15ztpn00an1n08x5 TAP_617 ();
 b15ztpn00an1n08x5 TAP_618 ();
 b15ztpn00an1n08x5 TAP_619 ();
 b15ztpn00an1n08x5 TAP_620 ();
 b15ztpn00an1n08x5 TAP_621 ();
 b15ztpn00an1n08x5 TAP_622 ();
 b15ztpn00an1n08x5 TAP_623 ();
 b15ztpn00an1n08x5 TAP_624 ();
 b15ztpn00an1n08x5 TAP_625 ();
 b15ztpn00an1n08x5 TAP_626 ();
 b15ztpn00an1n08x5 TAP_627 ();
 b15ztpn00an1n08x5 TAP_628 ();
 b15ztpn00an1n08x5 TAP_629 ();
 b15ztpn00an1n08x5 TAP_630 ();
 b15ztpn00an1n08x5 TAP_631 ();
 b15ztpn00an1n08x5 TAP_632 ();
 b15ztpn00an1n08x5 TAP_633 ();
 b15ztpn00an1n08x5 TAP_634 ();
 b15ztpn00an1n08x5 TAP_635 ();
 b15ztpn00an1n08x5 TAP_636 ();
 b15ztpn00an1n08x5 TAP_637 ();
 b15ztpn00an1n08x5 TAP_638 ();
 b15ztpn00an1n08x5 TAP_639 ();
 b15ztpn00an1n08x5 TAP_640 ();
 b15ztpn00an1n08x5 TAP_641 ();
 b15ztpn00an1n08x5 TAP_642 ();
 b15ztpn00an1n08x5 TAP_643 ();
 b15ztpn00an1n08x5 TAP_644 ();
 b15ztpn00an1n08x5 TAP_645 ();
 b15ztpn00an1n08x5 TAP_646 ();
 b15ztpn00an1n08x5 TAP_647 ();
 b15ztpn00an1n08x5 TAP_648 ();
 b15ztpn00an1n08x5 TAP_649 ();
 b15ztpn00an1n08x5 TAP_650 ();
 b15ztpn00an1n08x5 TAP_651 ();
 b15ztpn00an1n08x5 TAP_652 ();
 b15ztpn00an1n08x5 TAP_653 ();
 b15ztpn00an1n08x5 TAP_654 ();
 b15ztpn00an1n08x5 TAP_655 ();
 b15ztpn00an1n08x5 TAP_656 ();
 b15ztpn00an1n08x5 TAP_657 ();
 b15ztpn00an1n08x5 TAP_658 ();
 b15ztpn00an1n08x5 TAP_659 ();
 b15ztpn00an1n08x5 TAP_660 ();
 b15ztpn00an1n08x5 TAP_661 ();
 b15ztpn00an1n08x5 TAP_662 ();
 b15ztpn00an1n08x5 TAP_663 ();
 b15ztpn00an1n08x5 TAP_664 ();
 b15ztpn00an1n08x5 TAP_665 ();
 b15ztpn00an1n08x5 TAP_666 ();
 b15ztpn00an1n08x5 TAP_667 ();
 b15ztpn00an1n08x5 TAP_668 ();
 b15ztpn00an1n08x5 TAP_669 ();
 b15ztpn00an1n08x5 TAP_670 ();
 b15ztpn00an1n08x5 TAP_671 ();
 b15ztpn00an1n08x5 TAP_672 ();
 b15ztpn00an1n08x5 TAP_673 ();
 b15ztpn00an1n08x5 TAP_674 ();
 b15ztpn00an1n08x5 TAP_675 ();
 b15ztpn00an1n08x5 TAP_676 ();
 b15ztpn00an1n08x5 TAP_677 ();
 b15ztpn00an1n08x5 TAP_678 ();
 b15ztpn00an1n08x5 TAP_679 ();
 b15ztpn00an1n08x5 TAP_680 ();
 b15ztpn00an1n08x5 TAP_681 ();
 b15ztpn00an1n08x5 TAP_682 ();
 b15ztpn00an1n08x5 TAP_683 ();
 b15ztpn00an1n08x5 TAP_684 ();
 b15ztpn00an1n08x5 TAP_685 ();
 b15ztpn00an1n08x5 TAP_686 ();
 b15ztpn00an1n08x5 TAP_687 ();
 b15ztpn00an1n08x5 TAP_688 ();
 b15ztpn00an1n08x5 TAP_689 ();
 b15ztpn00an1n08x5 TAP_690 ();
 b15ztpn00an1n08x5 TAP_691 ();
 b15ztpn00an1n08x5 TAP_692 ();
 b15ztpn00an1n08x5 TAP_693 ();
 b15ztpn00an1n08x5 TAP_694 ();
 b15ztpn00an1n08x5 TAP_695 ();
 b15ztpn00an1n08x5 TAP_696 ();
 b15ztpn00an1n08x5 TAP_697 ();
 b15ztpn00an1n08x5 TAP_698 ();
 b15ztpn00an1n08x5 TAP_699 ();
 b15ztpn00an1n08x5 TAP_700 ();
 b15ztpn00an1n08x5 TAP_701 ();
 b15ztpn00an1n08x5 TAP_702 ();
 b15ztpn00an1n08x5 TAP_703 ();
 b15ztpn00an1n08x5 TAP_704 ();
 b15ztpn00an1n08x5 TAP_705 ();
 b15ztpn00an1n08x5 TAP_706 ();
 b15ztpn00an1n08x5 TAP_707 ();
 b15ztpn00an1n08x5 TAP_708 ();
 b15ztpn00an1n08x5 TAP_709 ();
 b15ztpn00an1n08x5 TAP_710 ();
 b15ztpn00an1n08x5 TAP_711 ();
 b15ztpn00an1n08x5 TAP_712 ();
 b15ztpn00an1n08x5 TAP_713 ();
 b15ztpn00an1n08x5 TAP_714 ();
 b15ztpn00an1n08x5 TAP_715 ();
 b15ztpn00an1n08x5 TAP_716 ();
 b15ztpn00an1n08x5 TAP_717 ();
 b15ztpn00an1n08x5 TAP_718 ();
 b15ztpn00an1n08x5 TAP_719 ();
 b15ztpn00an1n08x5 TAP_720 ();
 b15ztpn00an1n08x5 TAP_721 ();
 b15ztpn00an1n08x5 TAP_722 ();
 b15ztpn00an1n08x5 TAP_723 ();
 b15ztpn00an1n08x5 TAP_724 ();
 b15ztpn00an1n08x5 TAP_725 ();
 b15ztpn00an1n08x5 TAP_726 ();
 b15ztpn00an1n08x5 TAP_727 ();
 b15ztpn00an1n08x5 TAP_728 ();
 b15ztpn00an1n08x5 TAP_729 ();
 b15ztpn00an1n08x5 TAP_730 ();
 b15ztpn00an1n08x5 TAP_731 ();
 b15ztpn00an1n08x5 TAP_732 ();
 b15ztpn00an1n08x5 TAP_733 ();
 b15ztpn00an1n08x5 TAP_734 ();
 b15ztpn00an1n08x5 TAP_735 ();
 b15ztpn00an1n08x5 TAP_736 ();
 b15ztpn00an1n08x5 TAP_737 ();
 b15ztpn00an1n08x5 TAP_738 ();
 b15ztpn00an1n08x5 TAP_739 ();
 b15ztpn00an1n08x5 TAP_740 ();
 b15ztpn00an1n08x5 TAP_741 ();
 b15ztpn00an1n08x5 TAP_742 ();
 b15ztpn00an1n08x5 TAP_743 ();
 b15ztpn00an1n08x5 TAP_744 ();
 b15ztpn00an1n08x5 TAP_745 ();
 b15ztpn00an1n08x5 TAP_746 ();
 b15ztpn00an1n08x5 TAP_747 ();
 b15ztpn00an1n08x5 TAP_748 ();
 b15ztpn00an1n08x5 TAP_749 ();
 b15ztpn00an1n08x5 TAP_750 ();
 b15ztpn00an1n08x5 TAP_751 ();
 b15ztpn00an1n08x5 TAP_752 ();
 b15ztpn00an1n08x5 TAP_753 ();
 b15ztpn00an1n08x5 TAP_754 ();
 b15ztpn00an1n08x5 TAP_755 ();
 b15ztpn00an1n08x5 TAP_756 ();
 b15ztpn00an1n08x5 TAP_757 ();
 b15ztpn00an1n08x5 TAP_758 ();
 b15ztpn00an1n08x5 TAP_759 ();
 b15ztpn00an1n08x5 TAP_760 ();
 b15ztpn00an1n08x5 TAP_761 ();
 b15ztpn00an1n08x5 TAP_762 ();
 b15ztpn00an1n08x5 TAP_763 ();
 b15ztpn00an1n08x5 TAP_764 ();
 b15ztpn00an1n08x5 TAP_765 ();
 b15ztpn00an1n08x5 TAP_766 ();
 b15ztpn00an1n08x5 TAP_767 ();
 b15ztpn00an1n08x5 TAP_768 ();
 b15ztpn00an1n08x5 TAP_769 ();
 b15ztpn00an1n08x5 TAP_770 ();
 b15ztpn00an1n08x5 TAP_771 ();
 b15ztpn00an1n08x5 TAP_772 ();
 b15ztpn00an1n08x5 TAP_773 ();
 b15ztpn00an1n08x5 TAP_774 ();
 b15ztpn00an1n08x5 TAP_775 ();
 b15ztpn00an1n08x5 TAP_776 ();
 b15ztpn00an1n08x5 TAP_777 ();
 b15ztpn00an1n08x5 TAP_778 ();
 b15ztpn00an1n08x5 TAP_779 ();
 b15ztpn00an1n08x5 TAP_780 ();
 b15bfn001ah1n24x5 input1 (.a(rst_ni),
    .o(net1));
 b15bfn001as1n64x5 input2 (.a(spi_cs),
    .o(net2));
 b15bfn001as1n16x5 input3 (.a(spi_sdi0),
    .o(net3));
 b15bfn001ah1n12x5 input4 (.a(spi_sdi1),
    .o(net4));
 b15bfn001as1n12x5 input5 (.a(spi_sdi2),
    .o(net5));
 b15bfn001as1n16x5 input6 (.a(spi_sdi3),
    .o(net6));
 b15bfn001as1n08x5 input7 (.a(test_mode),
    .o(net7));
 b15bfn000as1n04x5 input8 (.a(tl_i[0]),
    .o(net8));
 b15bfn000as1n02x5 input9 (.a(tl_i[10]),
    .o(net9));
 b15bfn000ah1n03x5 input10 (.a(tl_i[11]),
    .o(net10));
 b15bfn001aq1n06x5 input11 (.a(tl_i[12]),
    .o(net11));
 b15bfn000as1n02x5 input12 (.a(tl_i[13]),
    .o(net12));
 b15bfn000as1n02x5 input13 (.a(tl_i[14]),
    .o(net13));
 b15bfn000as1n02x5 input14 (.a(tl_i[15]),
    .o(net14));
 b15bfn001as1n32x5 input15 (.a(tl_i[16]),
    .o(net15));
 b15bfn001as1n32x5 input16 (.a(tl_i[17]),
    .o(net16));
 b15bfn001as1n24x5 input17 (.a(tl_i[18]),
    .o(net17));
 b15bfn001as1n24x5 input18 (.a(tl_i[19]),
    .o(net18));
 b15bfn000as1n02x5 input19 (.a(tl_i[1]),
    .o(net19));
 b15bfn001as1n32x5 input20 (.a(tl_i[20]),
    .o(net20));
 b15bfn001as1n32x5 input21 (.a(tl_i[21]),
    .o(net21));
 b15bfn001as1n32x5 input22 (.a(tl_i[22]),
    .o(net22));
 b15bfn001as1n32x5 input23 (.a(tl_i[23]),
    .o(net23));
 b15bfn001as1n32x5 input24 (.a(tl_i[24]),
    .o(net24));
 b15bfn001as1n32x5 input25 (.a(tl_i[25]),
    .o(net25));
 b15bfn001as1n24x5 input26 (.a(tl_i[26]),
    .o(net26));
 b15bfn001as1n24x5 input27 (.a(tl_i[27]),
    .o(net27));
 b15bfn001as1n32x5 input28 (.a(tl_i[28]),
    .o(net28));
 b15bfn001as1n32x5 input29 (.a(tl_i[29]),
    .o(net29));
 b15bfn001as1n32x5 input30 (.a(tl_i[30]),
    .o(net30));
 b15bfn001as1n32x5 input31 (.a(tl_i[31]),
    .o(net31));
 b15bfn001as1n24x5 input32 (.a(tl_i[32]),
    .o(net32));
 b15bfn001as1n24x5 input33 (.a(tl_i[33]),
    .o(net33));
 b15bfn001as1n32x5 input34 (.a(tl_i[34]),
    .o(net34));
 b15bfn001as1n32x5 input35 (.a(tl_i[35]),
    .o(net35));
 b15bfn001as1n32x5 input36 (.a(tl_i[36]),
    .o(net36));
 b15bfn001as1n32x5 input37 (.a(tl_i[37]),
    .o(net37));
 b15bfn001as1n32x5 input38 (.a(tl_i[38]),
    .o(net38));
 b15bfn001as1n32x5 input39 (.a(tl_i[39]),
    .o(net39));
 b15bfn001as1n32x5 input40 (.a(tl_i[40]),
    .o(net40));
 b15bfn001as1n32x5 input41 (.a(tl_i[41]),
    .o(net41));
 b15bfn001as1n32x5 input42 (.a(tl_i[42]),
    .o(net42));
 b15bfn001as1n32x5 input43 (.a(tl_i[43]),
    .o(net43));
 b15bfn001as1n16x5 input44 (.a(tl_i[44]),
    .o(net44));
 b15bfn001as1n16x5 input45 (.a(tl_i[45]),
    .o(net45));
 b15bfn001as1n12x5 input46 (.a(tl_i[46]),
    .o(net46));
 b15bfn001as1n12x5 input47 (.a(tl_i[47]),
    .o(net47));
 b15bfn001aq1n06x5 input48 (.a(tl_i[57]),
    .o(net48));
 b15qgbbf1an1n05x5 input49 (.a(tl_i[58]),
    .o(net49));
 b15bfn000ah1n06x5 input50 (.a(tl_i[62]),
    .o(net50));
 b15bfn001aq1n06x5 input51 (.a(tl_i[63]),
    .o(net51));
 b15bfn001ah1n08x5 input52 (.a(tl_i[64]),
    .o(net52));
 b15bfn001ah1n16x5 input53 (.a(tl_i[65]),
    .o(net53));
 b15bfn000aq1n02x5 input54 (.a(tl_i[9]),
    .o(net54));
 b15bfn000ah1n03x5 output55 (.a(net2080),
    .o(net2081));
 b15bfn000ah1n03x5 output56 (.a(net2092),
    .o(net2093));
 b15bfn000ah1n03x5 output57 (.a(net2229),
    .o(net2230));
 b15bfn000ah1n03x5 output58 (.a(net58),
    .o(spi_sdo1));
 b15bfn000ah1n03x5 output59 (.a(net59),
    .o(spi_sdo2));
 b15bfn000ah1n03x5 output60 (.a(net60),
    .o(spi_sdo3));
 b15bfn000ah1n03x5 output61 (.a(net2014),
    .o(net2015));
 b15bfn000ah1n03x5 output62 (.a(net1976),
    .o(net1977));
 b15bfn000ah1n03x5 output63 (.a(net2064),
    .o(net2065));
 b15bfn000ah1n03x5 output64 (.a(net2161),
    .o(net2162));
 b15bfn000ah1n03x5 output65 (.a(net2095),
    .o(net2096));
 b15bfn000ah1n03x5 output66 (.a(net2074),
    .o(net2075));
 b15bfn000ah1n03x5 output67 (.a(net2130),
    .o(net2131));
 b15bfn000ah1n03x5 output68 (.a(net2434),
    .o(net2007));
 b15bfn000ah1n03x5 output69 (.a(net2448),
    .o(net2032));
 b15bfn000ah1n03x5 output70 (.a(net2450),
    .o(net2034));
 b15bfn000ah1n03x5 output71 (.a(net2431),
    .o(net2009));
 b15bfn000ah1n03x5 output72 (.a(net2428),
    .o(net2011));
 b15bfn000ah1n03x5 output73 (.a(net2374),
    .o(net1957));
 b15bfn000ah1n03x5 output74 (.a(net2383),
    .o(net1963));
 b15bfn000ah1n03x5 output75 (.a(net2419),
    .o(net2001));
 b15bfn000ah1n03x5 output76 (.a(net2416),
    .o(net1999));
 b15bfn000ah1n03x5 output77 (.a(net2407),
    .o(net1990));
 b15bfn000ah1n03x5 output78 (.a(net2398),
    .o(net1985));
 b15bfn000ah1n03x5 output79 (.a(net2404),
    .o(net1983));
 b15bfn000ah1n03x5 output80 (.a(net2401),
    .o(net1979));
 b15bfn000ah1n03x5 output81 (.a(net2380),
    .o(net1961));
 b15bfn000ah1n03x5 output82 (.a(net2377),
    .o(net1959));
 b15bfn000ah1n03x5 output83 (.a(net2422),
    .o(net2003));
 b15bfn000ah1n03x5 output84 (.a(net2425),
    .o(net2005));
 b15bfn000ah1n03x5 output85 (.a(net2442),
    .o(net2017));
 b15bfn000ah1n03x5 output86 (.a(net2440),
    .o(net2019));
 b15bfn000ah1n03x5 output87 (.a(net2410),
    .o(net1995));
 b15bfn000ah1n03x5 output88 (.a(net2413),
    .o(net1997));
 b15bfn000ah1n03x5 output89 (.a(net1987),
    .o(net1988));
 b15bfn000ah1n03x5 output90 (.a(net1992),
    .o(net1993));
 b15bfn000ah1n03x5 output91 (.a(net2386),
    .o(net1968));
 b15bfn000ah1n03x5 output92 (.a(net2389),
    .o(net1970));
 b15bfn000ah1n03x5 output93 (.a(net2395),
    .o(net1974));
 b15bfn000ah1n03x5 output94 (.a(net2392),
    .o(net1972));
 b15bfn000ah1n03x5 output95 (.a(net1965),
    .o(net1966));
 b15bfn000ah1n03x5 output96 (.a(net2463),
    .o(net2052));
 b15bfn000ah1n03x5 output97 (.a(net2452),
    .o(net2040));
 b15bfn000ah1n03x5 output98 (.a(net2437),
    .o(net2028));
 b15bfn000ah1n03x5 output99 (.a(net2444),
    .o(net2024));
 b15bfn000ah1n03x5 output100 (.a(net2474),
    .o(net2047));
 b15bfn000ah1n03x5 output101 (.a(net2104),
    .o(net2105));
 b15bfn000ah1n03x5 output102 (.a(net2123),
    .o(net2124));
 b15bfn000ah1n03x5 output103 (.a(net2151),
    .o(tl_o[65]));
 b15bfn000ah1n03x5 output104 (.a(net2128),
    .o(net2085));
 b15bfn000ah1n03x5 output105 (.a(net2499),
    .o(net2119));
 b15bfn000ah1n03x5 output106 (.a(net2484),
    .o(net2083));
 b15bfn000ah1n03x5 output107 (.a(net2044),
    .o(net2045));
 b15bfn000ah1n03x5 output108 (.a(net2101),
    .o(net2102));
 b15bfn000ah1n03x5 output109 (.a(net2476),
    .o(net2054));
 b15bfn000ah1n03x5 output110 (.a(net2147),
    .o(net2148));
 b15bfn000ah1n03x5 output111 (.a(net2488),
    .o(net2115));
 b15bfn000ah1n03x5 output112 (.a(net2137),
    .o(net2107));
 b15bfn000ah1n03x5 output113 (.a(net2116),
    .o(net2117));
 b15bfn000ah1n03x5 output114 (.a(net2049),
    .o(net2050));
 b15bfn000ah1n03x5 output115 (.a(net2505),
    .o(net2133));
 b15bfn000ah1n03x5 output116 (.a(net286),
    .o(tl_o[78]));
 b15bfn000ah1n03x5 output117 (.a(net2134),
    .o(net2135));
 b15bfn000ah1n03x5 output118 (.a(net2468),
    .o(net2026));
 b15bfn000ah1n03x5 output119 (.a(net2037),
    .o(net2038));
 b15bfn000ah1n03x5 output120 (.a(net2021),
    .o(net2022));
 b15bfn000ah1n03x5 output121 (.a(net2470),
    .o(net2042));
 b15bfn000ah1n03x5 output122 (.a(net2459),
    .o(net2056));
 b15bfn000ah1n03x5 output123 (.a(net2069),
    .o(net2070));
 b15bfn000ah1n03x5 output124 (.a(net2472),
    .o(net2126));
 b15bfn000ah1n03x5 output125 (.a(net2503),
    .o(net2121));
 b15bfn000ah1n03x5 output126 (.a(net2098),
    .o(net2099));
 b15bfn000ah1n03x5 output127 (.a(net2461),
    .o(net2058));
 b15bfn000ah1n03x5 output128 (.a(net2112),
    .o(net2113));
 b15bfn000ah1n03x5 output129 (.a(net2111),
    .o(net2109));
 b15bfn000ah1n03x5 output130 (.a(net2455),
    .o(net2030));
 b15bfn000ah1n03x5 output131 (.a(net2457),
    .o(net1981));
 b15bfn000ah1n03x5 output132 (.a(net2139),
    .o(net2140));
 b15bfn001as1n16x5 wire133 (.a(u_dcfifo_rx_u_din_buffer_N28),
    .o(net133));
 b15bfn001as1n24x5 wire134 (.a(u_dcfifo_rx_u_din_write_enable),
    .o(net134));
 b15bfn001as1n48x5 fanout135 (.a(net139),
    .o(net135));
 b15bfn001ah1n48x5 load_slew136 (.a(net135),
    .o(net136));
 b15bfn001ah1n32x5 fanout137 (.a(net139),
    .o(net137));
 b15bfn001ah1n48x5 fanout138 (.a(n3822),
    .o(net138));
 b15bfn001ah1n32x5 wire139 (.a(net138),
    .o(net139));
 b15bfn001ah1n32x5 wire140 (.a(ctrl_rd_wr),
    .o(net140));
 b15bfn001as1n16x5 wire141 (.a(u_spi_device_tlul_plug_wdata_next[23]),
    .o(net141));
 b15bfn001as1n16x5 wire142 (.a(u_spi_device_tlul_plug_wdata_next[5]),
    .o(net142));
 b15bfn001as1n16x5 wire143 (.a(n3536),
    .o(net143));
 b15bfn001ah1n24x5 wire144 (.a(n3464),
    .o(net144));
 b15bfn001as1n16x5 wire145 (.a(n3434),
    .o(net145));
 b15bfn001ah1n24x5 wire146 (.a(n3376),
    .o(net146));
 b15bfn001as1n16x5 wire147 (.a(net148),
    .o(net147));
 b15bfn001as1n16x5 max_length148 (.a(u_device_sm_sample_ADDR),
    .o(net148));
 b15bfn001as1n64x5 fanout149 (.a(net150),
    .o(net149));
 b15bfn001as1n80x5 fanout150 (.a(n3365),
    .o(net150));
 b15bfn001ah1n48x5 fanout151 (.a(n3356),
    .o(net151));
 b15bfn001ah1n64x5 fanout152 (.a(n3356),
    .o(net152));
 b15bfn001ah1n48x5 fanout153 (.a(n3353),
    .o(net153));
 b15bfn000ah1n48x5 fanout154 (.a(n3353),
    .o(net154));
 b15bfn001ah1n48x5 fanout155 (.a(n3347),
    .o(net155));
 b15bfn001ah1n48x5 fanout156 (.a(n3347),
    .o(net156));
 b15bfn001as1n16x5 wire157 (.a(u_dcfifo_rx_u_din_full_full_dn),
    .o(net157));
 b15bfn001ah1n64x5 fanout158 (.a(n3362),
    .o(net158));
 b15bfn001ah1n80x5 fanout159 (.a(n3362),
    .o(net159));
 b15bfn001as1n48x5 fanout160 (.a(n3359),
    .o(net160));
 b15bfn001ah1n80x5 fanout161 (.a(n3359),
    .o(net161));
 b15bfn001as1n48x5 fanout162 (.a(n3351),
    .o(net162));
 b15bfn001ah1n64x5 fanout163 (.a(n3351),
    .o(net163));
 b15bfn001ah1n48x5 fanout164 (.a(net165),
    .o(net164));
 b15bfn001as1n48x5 fanout165 (.a(n3349),
    .o(net165));
 b15bfn001as1n48x5 max_length166 (.a(net165),
    .o(net166));
 b15bfn001as1n24x5 fanout167 (.a(net168),
    .o(net167));
 b15bfn000as1n32x5 fanout168 (.a(n3309),
    .o(net168));
 b15bfn001as1n48x5 fanout169 (.a(net171),
    .o(net169));
 b15bfn001ah1n64x5 fanout170 (.a(net171),
    .o(net170));
 b15bfn001as1n32x5 wire171 (.a(n3020),
    .o(net171));
 b15bfn001as1n48x5 fanout172 (.a(n3018),
    .o(net172));
 b15bfn000ah1n48x5 fanout173 (.a(n3018),
    .o(net173));
 b15bfn001ah1n64x5 fanout174 (.a(n3015),
    .o(net174));
 b15bfn001ah1n48x5 fanout175 (.a(net176),
    .o(net175));
 b15bfn001ah1n24x5 wire176 (.a(n3015),
    .o(net176));
 b15bfn001ah1n64x5 fanout177 (.a(net179),
    .o(net177));
 b15bfn001ah1n48x5 fanout178 (.a(net179),
    .o(net178));
 b15bfn001as1n32x5 wire179 (.a(n3011),
    .o(net179));
 b15bfn001ah1n48x5 fanout180 (.a(n3009),
    .o(net180));
 b15bfn001as1n48x5 fanout181 (.a(n3009),
    .o(net181));
 b15bfn001ah1n48x5 fanout182 (.a(net184),
    .o(net182));
 b15bfn000ah1n48x5 fanout183 (.a(net184),
    .o(net183));
 b15bfn001ah1n32x5 wire184 (.a(n3006),
    .o(net184));
 b15bfn001ah1n64x5 fanout185 (.a(n3004),
    .o(net185));
 b15bfn001ah1n64x5 fanout186 (.a(net187),
    .o(net186));
 b15bfn001ah1n24x5 wire187 (.a(n3004),
    .o(net187));
 b15bfn001ah1n48x5 fanout188 (.a(n3002),
    .o(net188));
 b15bfn001ah1n48x5 fanout189 (.a(n3002),
    .o(net189));
 b15bfn001as1n24x5 wire190 (.a(n3820),
    .o(net190));
 b15bfn001ah1n24x5 wire191 (.a(n3820),
    .o(net191));
 b15bfn001ah1n32x5 wire192 (.a(ctrl_data_rx[15]),
    .o(net192));
 b15bfn001ah1n24x5 wire193 (.a(ctrl_data_rx[12]),
    .o(net193));
 b15bfn001as1n16x5 max_length194 (.a(ctrl_data_rx[12]),
    .o(net194));
 b15bfn001ah1n32x5 max_length195 (.a(net196),
    .o(net195));
 b15bfn001as1n24x5 wire196 (.a(ctrl_data_rx[21]),
    .o(net196));
 b15bfn001as1n24x5 wire197 (.a(net198),
    .o(net197));
 b15bfn001as1n24x5 wire198 (.a(ctrl_data_rx[24]),
    .o(net198));
 b15bfn001as1n16x5 max_length199 (.a(net200),
    .o(net199));
 b15bfn001ah1n24x5 max_length200 (.a(ctrl_data_rx[27]),
    .o(net200));
 b15bfn001as1n16x5 max_length201 (.a(net202),
    .o(net201));
 b15bfn001ah1n24x5 max_length202 (.a(ctrl_data_rx[26]),
    .o(net202));
 b15bfn001ah1n32x5 max_length203 (.a(net204),
    .o(net203));
 b15bfn001as1n24x5 wire204 (.a(ctrl_data_rx[18]),
    .o(net204));
 b15bfn001as1n24x5 max_length205 (.a(net206),
    .o(net205));
 b15bfn001as1n16x5 max_length206 (.a(ctrl_data_rx[28]),
    .o(net206));
 b15bfn001ah1n24x5 max_length207 (.a(net208),
    .o(net207));
 b15bfn001as1n24x5 max_length208 (.a(ctrl_data_rx[30]),
    .o(net208));
 b15bfn001as1n24x5 wire209 (.a(net210),
    .o(net209));
 b15bfn001as1n24x5 wire210 (.a(ctrl_data_rx[25]),
    .o(net210));
 b15bfn001ah1n24x5 max_length211 (.a(ctrl_data_rx[16]),
    .o(net211));
 b15bfn001ah1n24x5 max_length212 (.a(ctrl_data_rx[16]),
    .o(net212));
 b15bfn001ah1n24x5 wire213 (.a(ctrl_data_rx[13]),
    .o(net213));
 b15bfn001ah1n24x5 max_length214 (.a(ctrl_data_rx[13]),
    .o(net214));
 b15bfn001ah1n32x5 max_length215 (.a(net216),
    .o(net215));
 b15bfn001as1n24x5 wire216 (.a(ctrl_data_rx[19]),
    .o(net216));
 b15bfn001as1n24x5 wire217 (.a(ctrl_data_rx[10]),
    .o(net217));
 b15bfn001as1n24x5 wire218 (.a(net219),
    .o(net218));
 b15bfn001ah1n32x5 max_length219 (.a(ctrl_data_rx[22]),
    .o(net219));
 b15bfn001ah1n24x5 max_length220 (.a(net221),
    .o(net220));
 b15bfn001as1n24x5 max_length221 (.a(ctrl_data_rx[14]),
    .o(net221));
 b15bfn001as1n24x5 wire222 (.a(net223),
    .o(net222));
 b15bfn001as1n24x5 max_length223 (.a(ctrl_data_rx[23]),
    .o(net223));
 b15bfn001ah1n24x5 max_length224 (.a(net226),
    .o(net224));
 b15bfn001ah1n24x5 max_length225 (.a(ctrl_data_rx[17]),
    .o(net225));
 b15bfn001ah1n24x5 max_length226 (.a(ctrl_data_rx[17]),
    .o(net226));
 b15bfn001ah1n32x5 max_length227 (.a(net228),
    .o(net227));
 b15bfn001as1n24x5 wire228 (.a(ctrl_data_rx[20]),
    .o(net228));
 b15bfn001as1n24x5 wire229 (.a(ctrl_data_rx[11]),
    .o(net229));
 b15bfn001ah1n24x5 wire230 (.a(ctrl_data_rx[31]),
    .o(net230));
 b15bfn001as1n24x5 max_length231 (.a(net232),
    .o(net231));
 b15bfn001as1n24x5 max_length232 (.a(ctrl_data_rx[29]),
    .o(net232));
 b15bfn001ah1n32x5 wire233 (.a(ctrl_data_rx[4]),
    .o(net233));
 b15bfn000as1n32x5 wire234 (.a(ctrl_data_rx[4]),
    .o(net234));
 b15bfn000as1n32x5 wire235 (.a(net237),
    .o(net235));
 b15bfn001as1n16x5 max_length236 (.a(ctrl_data_rx[2]),
    .o(net236));
 b15bfn001ah1n32x5 max_length237 (.a(ctrl_data_rx[2]),
    .o(net237));
 b15bfn001ah1n32x5 wire238 (.a(ctrl_data_rx[1]),
    .o(net238));
 b15bfn001ah1n32x5 wire239 (.a(ctrl_data_rx[1]),
    .o(net239));
 b15bfn001as1n24x5 wire240 (.a(ctrl_data_rx[6]),
    .o(net240));
 b15bfn001as1n16x5 max_length241 (.a(net242),
    .o(net241));
 b15bfn001as1n24x5 wire242 (.a(ctrl_data_rx[6]),
    .o(net242));
 b15bfn001ah1n32x5 wire243 (.a(ctrl_data_rx[7]),
    .o(net243));
 b15bfn001as1n16x5 max_length244 (.a(net245),
    .o(net244));
 b15bfn001as1n24x5 wire245 (.a(ctrl_data_rx[7]),
    .o(net245));
 b15bfn001ah1n32x5 wire246 (.a(net247),
    .o(net246));
 b15bfn001as1n32x5 wire247 (.a(ctrl_data_rx[3]),
    .o(net247));
 b15bfn001as1n24x5 wire248 (.a(ctrl_data_rx[3]),
    .o(net248));
 b15bfn001ah1n12x5 load_slew249 (.a(net2242),
    .o(net249));
 b15bfn001as1n16x5 wire250 (.a(net2241),
    .o(net250));
 b15bfn001ah1n24x5 wire251 (.a(net252),
    .o(net251));
 b15bfn001ah1n12x5 wire252 (.a(net2296),
    .o(net252));
 b15bfn001ah1n24x5 wire253 (.a(net254),
    .o(net253));
 b15bfn001ah1n12x5 wire254 (.a(net2317),
    .o(net254));
 b15bfn001as1n12x5 wire255 (.a(net2228),
    .o(net255));
 b15bfn001as1n16x5 fanout256 (.a(n2919),
    .o(net256));
 b15bfn001as1n12x5 fanout257 (.a(n2919),
    .o(net257));
 b15bfn001ah1n24x5 wire258 (.a(n3818),
    .o(net258));
 b15bfn001as1n24x5 wire259 (.a(n3818),
    .o(net259));
 b15bfn001ah1n24x5 fanout260 (.a(net261),
    .o(net260));
 b15bfn001as1n24x5 fanout261 (.a(n2917),
    .o(net261));
 b15bfn001as1n24x5 wire262 (.a(n3815),
    .o(net262));
 b15bfn001ah1n64x5 wire263 (.a(n3813),
    .o(net263));
 b15bfn001ah1n32x5 wire264 (.a(n2783),
    .o(net264));
 b15bfn001ah1n12x5 wire265 (.a(net2043),
    .o(net265));
 b15bfn001ah1n12x5 wire266 (.a(net2043),
    .o(net266));
 b15bfn001as1n12x5 wire267 (.a(net2082),
    .o(net267));
 b15bfn001ah1n24x5 wire268 (.a(net2150),
    .o(net268));
 b15bfn001as1n08x5 wire269 (.a(net2149),
    .o(net269));
 b15bfn001ah1n12x5 load_slew270 (.a(net2122),
    .o(net270));
 b15bfn001as1n12x5 wire271 (.a(net2029),
    .o(net271));
 b15bfn001ah1n12x5 wire272 (.a(net2103),
    .o(net272));
 b15bfn001ah1n12x5 wire273 (.a(net2046),
    .o(net273));
 b15bfn001ah1n12x5 wire274 (.a(net2057),
    .o(net274));
 b15bfn001as1n16x5 wire275 (.a(net2057),
    .o(net275));
 b15bfn001ah1n12x5 load_slew276 (.a(net2068),
    .o(net276));
 b15bfn001as1n12x5 wire277 (.a(net2041),
    .o(net277));
 b15bfn001ah1n16x5 wire278 (.a(net279),
    .o(net278));
 b15bfn001ah1n12x5 wire279 (.a(net2021),
    .o(net279));
 b15bfn001as1n12x5 wire280 (.a(net2020),
    .o(net280));
 b15bfn001ah1n12x5 load_slew281 (.a(net2036),
    .o(net281));
 b15bfn001ah1n12x5 wire282 (.a(net2035),
    .o(net282));
 b15bfn001as1n08x5 wire283 (.a(net285),
    .o(net283));
 b15bfn000ah1n24x5 wire284 (.a(net285),
    .o(net284));
 b15bfn001as1n08x5 load_slew285 (.a(net2025),
    .o(net285));
 b15bfn001as1n12x5 max_cap286 (.a(net2060),
    .o(net286));
 b15bfn001ah1n12x5 load_slew287 (.a(net2067),
    .o(net287));
 b15bfn001ah1n12x5 load_slew288 (.a(net2049),
    .o(net288));
 b15bfn001ah1n12x5 load_slew289 (.a(net2048),
    .o(net289));
 b15bfn001as1n12x5 wire290 (.a(net2053),
    .o(net290));
 b15bfn001ah1n12x5 load_slew291 (.a(net2053),
    .o(net291));
 b15bfn001ah1n12x5 wire292 (.a(u_rxreg_data_int[8]),
    .o(net292));
 b15bfn001ah1n12x5 load_slew293 (.a(net294),
    .o(net293));
 b15bfn001ah1n12x5 wire294 (.a(net2349),
    .o(net294));
 b15bfn001as1n08x5 load_slew295 (.a(u_rxreg_data_int[14]),
    .o(net295));
 b15bfn001ah1n64x5 fanout296 (.a(net298),
    .o(net296));
 b15bfn001as1n24x5 fanout297 (.a(net298),
    .o(net297));
 b15bfn001as1n64x5 fanout298 (.a(net299),
    .o(net298));
 b15bfn001ah1n12x5 wire299 (.a(en_quad),
    .o(net299));
 b15bfn001ah1n12x5 load_slew300 (.a(net2506),
    .o(net300));
 b15bfn001ah1n12x5 wire301 (.a(net302),
    .o(net301));
 b15bfn001ah1n12x5 load_slew302 (.a(en_quad),
    .o(net302));
 b15bfn001as1n08x5 load_slew303 (.a(net304),
    .o(net303));
 b15bfn001ah1n12x5 load_slew304 (.a(u_dcfifo_tx_u_dout_read_token[7]),
    .o(net304));
 b15bfn001as1n12x5 max_cap305 (.a(u_dcfifo_tx_u_dout_read_token[3]),
    .o(net305));
 b15bfn001ah1n12x5 wire306 (.a(u_dcfifo_tx_u_dout_read_token[1]),
    .o(net306));
 b15bfn001as1n12x5 load_slew307 (.a(u_dcfifo_tx_u_dout_read_token[0]),
    .o(net307));
 b15bfn001ah1n12x5 wire308 (.a(net309),
    .o(net308));
 b15bfn001ah1n12x5 load_slew309 (.a(u_dcfifo_tx_write_token[7]),
    .o(net309));
 b15bfn001ah1n12x5 load_slew310 (.a(net311),
    .o(net310));
 b15bfn001ah1n12x5 load_slew311 (.a(net312),
    .o(net311));
 b15bfn001ah1n12x5 wire312 (.a(u_dcfifo_tx_write_token[6]),
    .o(net312));
 b15bfn001ah1n12x5 wire313 (.a(net314),
    .o(net313));
 b15bfn001ah1n12x5 wire314 (.a(u_dcfifo_tx_write_token[5]),
    .o(net314));
 b15bfn001as1n12x5 wire315 (.a(u_dcfifo_tx_write_token[4]),
    .o(net315));
 b15bfn001ah1n08x5 load_slew316 (.a(u_dcfifo_tx_write_token[4]),
    .o(net316));
 b15bfn001as1n08x5 load_slew317 (.a(net318),
    .o(net317));
 b15bfn001as1n12x5 wire318 (.a(u_dcfifo_tx_write_token[3]),
    .o(net318));
 b15bfn001as1n06x5 load_slew319 (.a(net320),
    .o(net319));
 b15bfn001as1n12x5 wire320 (.a(net2306),
    .o(net320));
 b15bfn001as1n12x5 wire321 (.a(net322),
    .o(net321));
 b15bfn001ah1n12x5 wire322 (.a(u_dcfifo_tx_write_token[1]),
    .o(net322));
 b15bfn001as1n08x5 load_slew323 (.a(net324),
    .o(net323));
 b15bfn001ah1n12x5 load_slew324 (.a(u_dcfifo_tx_write_token[0]),
    .o(net324));
 b15bfn001ah1n12x5 wire325 (.a(u_dcfifo_rx_u_dout_read_token[5]),
    .o(net325));
 b15bfn001ah1n12x5 wire326 (.a(u_dcfifo_rx_u_dout_read_token[3]),
    .o(net326));
 b15bfn001as1n08x5 load_slew327 (.a(u_dcfifo_rx_write_token[7]),
    .o(net327));
 b15bfn001ah1n08x5 load_slew328 (.a(net329),
    .o(net328));
 b15bfn001ah1n12x5 wire329 (.a(u_dcfifo_rx_write_token[5]),
    .o(net329));
 b15bfn001as1n12x5 wire330 (.a(u_dcfifo_rx_write_token[4]),
    .o(net330));
 b15bfn001ah1n16x5 max_cap331 (.a(net332),
    .o(net331));
 b15bfn001as1n12x5 wire332 (.a(u_dcfifo_rx_write_token[3]),
    .o(net332));
 b15bfn001as1n12x5 load_slew333 (.a(net334),
    .o(net333));
 b15bfn001as1n12x5 wire334 (.a(u_dcfifo_rx_write_token[2]),
    .o(net334));
 b15bfn001as1n12x5 load_slew335 (.a(net336),
    .o(net335));
 b15bfn001ah1n12x5 wire336 (.a(u_dcfifo_rx_write_token[1]),
    .o(net336));
 b15bfn001ah1n16x5 wire337 (.a(u_dcfifo_rx_u_din_buffer_data[94]),
    .o(net337));
 b15bfn001ah1n16x5 wire338 (.a(u_dcfifo_rx_u_din_buffer_data[44]),
    .o(net338));
 b15bfn001ah1n12x5 load_slew339 (.a(net2013),
    .o(net339));
 b15bfn001as1n16x5 wire340 (.a(net2012),
    .o(net340));
 b15bfn001ah1n16x5 wire341 (.a(net2478),
    .o(net341));
 b15bfn001as1n16x5 wire342 (.a(net1991),
    .o(net342));
 b15bfn001as1n16x5 wire343 (.a(net1986),
    .o(net343));
 b15bfn001ah1n16x5 wire344 (.a(net2464),
    .o(net344));
 b15bfn001as1n80x5 fanout345 (.a(net346),
    .o(net345));
 b15bfn001as1n80x5 fanout346 (.a(net349),
    .o(net346));
 b15bfn001as1n08x5 load_slew347 (.a(net348),
    .o(net347));
 b15bfn001as1n08x5 load_slew348 (.a(net349),
    .o(net348));
 b15bfn001ah1n16x5 wire349 (.a(net351),
    .o(net349));
 b15bfn001ah1n12x5 load_slew350 (.a(net351),
    .o(net350));
 b15bfn001as1n12x5 wire351 (.a(n1869),
    .o(net351));
 b15bfn001ah1n32x5 fanout352 (.a(net353),
    .o(net352));
 b15bfn001ah1n32x5 fanout353 (.a(net354),
    .o(net353));
 b15bfn001ah1n16x5 wire354 (.a(net2298),
    .o(net354));
 b15bfn001ah1n12x5 load_slew355 (.a(u_device_sm_state[2]),
    .o(net355));
 b15bfn001ah1n12x5 load_slew356 (.a(net2078),
    .o(net356));
 b15bfn001as1n12x5 max_cap357 (.a(net2077),
    .o(net357));
 b15bfn001ah1n12x5 wire358 (.a(net2076),
    .o(net358));
 b15bfn001as1n08x5 load_slew359 (.a(net2088),
    .o(net359));
 b15bfn001as1n12x5 wire360 (.a(net2087),
    .o(net360));
 b15bfn001ah1n12x5 load_slew361 (.a(net362),
    .o(net361));
 b15bfn001as1n12x5 max_cap362 (.a(net2347),
    .o(net362));
 b15bfn001ah1n48x5 wire363 (.a(n3778),
    .o(net363));
 b15bfn001ah1n48x5 max_length364 (.a(n3777),
    .o(net364));
 b15bfn001ah1n32x5 max_length365 (.a(n3777),
    .o(net365));
 b15bfn001as1n32x5 wire366 (.a(n3776),
    .o(net366));
 b15bfn001ah1n32x5 wire367 (.a(n3776),
    .o(net367));
 b15bfn001as1n32x5 wire368 (.a(n3772),
    .o(net368));
 b15bfn001as1n32x5 max_length369 (.a(n3772),
    .o(net369));
 b15bfn001ah1n24x5 max_length370 (.a(net371),
    .o(net370));
 b15bfn000as1n32x5 wire371 (.a(net47),
    .o(net371));
 b15bfn001ah1n24x5 max_length372 (.a(net373),
    .o(net372));
 b15bfn000as1n32x5 wire373 (.a(net46),
    .o(net373));
 b15bfn001as1n24x5 max_length374 (.a(net375),
    .o(net374));
 b15bfn001ah1n32x5 wire375 (.a(net45),
    .o(net375));
 b15bfn001as1n24x5 max_length376 (.a(net377),
    .o(net376));
 b15bfn001ah1n32x5 wire377 (.a(net44),
    .o(net377));
 b15bfn001ah1n24x5 max_length378 (.a(net379),
    .o(net378));
 b15bfn001ah1n32x5 wire379 (.a(net43),
    .o(net379));
 b15bfn001ah1n24x5 max_length380 (.a(net381),
    .o(net380));
 b15bfn001ah1n32x5 wire381 (.a(net42),
    .o(net381));
 b15bfn001as1n24x5 max_length382 (.a(net383),
    .o(net382));
 b15bfn001ah1n32x5 wire383 (.a(net41),
    .o(net383));
 b15bfn001as1n24x5 max_length384 (.a(net385),
    .o(net384));
 b15bfn001ah1n32x5 wire385 (.a(net40),
    .o(net385));
 b15bfn001as1n16x5 max_length386 (.a(net387),
    .o(net386));
 b15bfn001ah1n32x5 wire387 (.a(net39),
    .o(net387));
 b15bfn001as1n16x5 max_length388 (.a(net389),
    .o(net388));
 b15bfn001ah1n32x5 wire389 (.a(net38),
    .o(net389));
 b15bfn001ah1n24x5 max_length390 (.a(net391),
    .o(net390));
 b15bfn001as1n32x5 wire391 (.a(net37),
    .o(net391));
 b15bfn001ah1n24x5 max_length392 (.a(net393),
    .o(net392));
 b15bfn001as1n32x5 wire393 (.a(net36),
    .o(net393));
 b15bfn001as1n24x5 max_length394 (.a(net395),
    .o(net394));
 b15bfn001as1n32x5 wire395 (.a(net35),
    .o(net395));
 b15bfn001as1n24x5 max_length396 (.a(net397),
    .o(net396));
 b15bfn001as1n32x5 wire397 (.a(net34),
    .o(net397));
 b15bfn001ah1n24x5 max_length398 (.a(net399),
    .o(net398));
 b15bfn001as1n32x5 wire399 (.a(net33),
    .o(net399));
 b15bfn001ah1n24x5 max_length400 (.a(net401),
    .o(net400));
 b15bfn001as1n32x5 wire401 (.a(net32),
    .o(net401));
 b15bfn001ah1n24x5 max_length402 (.a(net403),
    .o(net402));
 b15bfn001ah1n48x5 wire403 (.a(net31),
    .o(net403));
 b15bfn001ah1n24x5 max_length404 (.a(net405),
    .o(net404));
 b15bfn001ah1n48x5 wire405 (.a(net30),
    .o(net405));
 b15bfn001ah1n24x5 wire406 (.a(net407),
    .o(net406));
 b15bfn001ah1n48x5 wire407 (.a(net29),
    .o(net407));
 b15bfn001ah1n24x5 wire408 (.a(net409),
    .o(net408));
 b15bfn001ah1n48x5 wire409 (.a(net28),
    .o(net409));
 b15bfn001ah1n24x5 max_length410 (.a(net411),
    .o(net410));
 b15bfn000ah1n48x5 wire411 (.a(net27),
    .o(net411));
 b15bfn001ah1n24x5 max_length412 (.a(net413),
    .o(net412));
 b15bfn000ah1n48x5 wire413 (.a(net26),
    .o(net413));
 b15bfn001ah1n24x5 wire414 (.a(net415),
    .o(net414));
 b15bfn001as1n32x5 wire415 (.a(net25),
    .o(net415));
 b15bfn001ah1n24x5 wire416 (.a(net417),
    .o(net416));
 b15bfn001as1n32x5 wire417 (.a(net24),
    .o(net417));
 b15bfn001ah1n24x5 max_length418 (.a(net419),
    .o(net418));
 b15bfn001ah1n48x5 wire419 (.a(net23),
    .o(net419));
 b15bfn001ah1n24x5 max_length420 (.a(net421),
    .o(net420));
 b15bfn001ah1n48x5 wire421 (.a(net22),
    .o(net421));
 b15bfn001ah1n32x5 max_length422 (.a(net423),
    .o(net422));
 b15bfn001ah1n48x5 wire423 (.a(net21),
    .o(net423));
 b15bfn001ah1n32x5 max_length424 (.a(net425),
    .o(net424));
 b15bfn001ah1n48x5 wire425 (.a(net20),
    .o(net425));
 b15bfn001ah1n64x5 wire426 (.a(net2),
    .o(net426));
 b15bfn001ah1n48x5 load_slew427 (.a(net2),
    .o(net427));
 b15bfn001as1n16x5 max_length428 (.a(net429),
    .o(net428));
 b15bfn000ah1n48x5 wire429 (.a(net18),
    .o(net429));
 b15bfn001as1n16x5 max_length430 (.a(net431),
    .o(net430));
 b15bfn000ah1n48x5 wire431 (.a(net17),
    .o(net431));
 b15bfn001ah1n32x5 max_length432 (.a(net433),
    .o(net432));
 b15bfn001ah1n48x5 wire433 (.a(net16),
    .o(net433));
 b15bfn001ah1n32x5 max_length434 (.a(net435),
    .o(net434));
 b15bfn001ah1n48x5 wire435 (.a(net15),
    .o(net435));
 b15bfn001as1n48x5 fanout436 (.a(net448),
    .o(net436));
 b15bfn001as1n32x5 fanout437 (.a(net448),
    .o(net437));
 b15bfn001as1n48x5 fanout438 (.a(net448),
    .o(net438));
 b15bfn001as1n48x5 fanout439 (.a(net440),
    .o(net439));
 b15bfn001as1n48x5 fanout440 (.a(net441),
    .o(net440));
 b15bfn001as1n32x5 fanout441 (.a(net448),
    .o(net441));
 b15bfn001ah1n48x5 fanout442 (.a(net446),
    .o(net442));
 b15bfn001as1n48x5 fanout443 (.a(net444),
    .o(net443));
 b15bfn001as1n48x5 fanout444 (.a(net446),
    .o(net444));
 b15bfn001as1n48x5 fanout445 (.a(net446),
    .o(net445));
 b15bfn001as1n48x5 fanout446 (.a(net447),
    .o(net446));
 b15bfn001as1n32x5 fanout447 (.a(net1),
    .o(net447));
 b15bfn001as1n48x5 wire448 (.a(net447),
    .o(net448));
 b15bfn001as1n48x5 fanout449 (.a(net465),
    .o(net449));
 b15bfn001as1n32x5 fanout450 (.a(net465),
    .o(net450));
 b15bfn001as1n48x5 fanout451 (.a(net452),
    .o(net451));
 b15bfn001as1n48x5 fanout452 (.a(net465),
    .o(net452));
 b15bfn001ah1n48x5 fanout453 (.a(net456),
    .o(net453));
 b15bfn001as1n48x5 fanout454 (.a(net456),
    .o(net454));
 b15bfn001as1n24x5 fanout455 (.a(net456),
    .o(net455));
 b15bfn001ah1n48x5 fanout456 (.a(net465),
    .o(net456));
 b15bfn001as1n48x5 fanout457 (.a(net458),
    .o(net457));
 b15bfn001ah1n48x5 fanout458 (.a(net464),
    .o(net458));
 b15bfn001as1n48x5 fanout459 (.a(net464),
    .o(net459));
 b15bfn001ah1n48x5 fanout460 (.a(net464),
    .o(net460));
 b15bfn001as1n48x5 fanout461 (.a(net463),
    .o(net461));
 b15bfn001as1n48x5 fanout462 (.a(net463),
    .o(net462));
 b15bfn001as1n32x5 fanout463 (.a(net464),
    .o(net463));
 b15bfn001as1n48x5 fanout464 (.a(net1),
    .o(net464));
 b15bfn001ah1n48x5 wire465 (.a(net464),
    .o(net465));
 b15tilo00an1n03x5 U2924_466 (.o(net466));
 b15tilo00an1n03x5 U3035_467 (.o(net467));
 b15tilo00an1n03x5 U3045_468 (.o(net468));
 b15tilo00an1n03x5 U3114_469 (.o(net469));
 b15tilo00an1n03x5 U3242_470 (.o(net470));
 b15tilo00an1n03x5 U3298_471 (.o(net471));
 b15tilo00an1n03x5 U3320_472 (.o(net472));
 b15tilo00an1n03x5 U3322_473 (.o(net473));
 b15tilo00an1n03x5 U3334_474 (.o(net474));
 b15tilo00an1n03x5 U3340_475 (.o(net475));
 b15tilo00an1n03x5 U3439_476 (.o(net476));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_0__0_latch_477 (.o(net477));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_0__latch_478 (.o(net478));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_1__0_latch_479 (.o(net479));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_1__latch_480 (.o(net480));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_2__0_latch_481 (.o(net481));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_2__latch_482 (.o(net482));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_3__0_latch_483 (.o(net483));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_3__latch_484 (.o(net484));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_4__0_latch_485 (.o(net485));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_4__latch_486 (.o(net486));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_5__0_latch_487 (.o(net487));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_5__latch_488 (.o(net488));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_6__0_latch_489 (.o(net489));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_6__latch_490 (.o(net490));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_7__0_latch_491 (.o(net491));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_clk_gate_data_reg_7__latch_492 (.o(net492));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__0__u_dcfifo_rx_u_din_buffer_data_reg_0__1__493 (.o(net493));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__0__u_dcfifo_rx_u_din_buffer_data_reg_0__1__494 (.o(net494));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__10__u_dcfifo_rx_u_din_buffer_data_reg_0__11__495 (.o(net495));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__10__u_dcfifo_rx_u_din_buffer_data_reg_0__11__496 (.o(net496));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__12__u_dcfifo_rx_u_din_buffer_data_reg_0__13__497 (.o(net497));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__12__u_dcfifo_rx_u_din_buffer_data_reg_0__13__498 (.o(net498));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__14__u_dcfifo_rx_u_din_buffer_data_reg_0__15__499 (.o(net499));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__14__u_dcfifo_rx_u_din_buffer_data_reg_0__15__500 (.o(net500));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__16__u_dcfifo_rx_u_din_buffer_data_reg_0__17__501 (.o(net501));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__16__u_dcfifo_rx_u_din_buffer_data_reg_0__17__502 (.o(net502));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__18__u_dcfifo_rx_u_din_buffer_data_reg_0__19__503 (.o(net503));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__18__u_dcfifo_rx_u_din_buffer_data_reg_0__19__504 (.o(net504));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__20__u_dcfifo_rx_u_din_buffer_data_reg_0__21__505 (.o(net505));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__20__u_dcfifo_rx_u_din_buffer_data_reg_0__21__506 (.o(net506));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__22__u_dcfifo_rx_u_din_buffer_data_reg_0__23__507 (.o(net507));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__22__u_dcfifo_rx_u_din_buffer_data_reg_0__23__508 (.o(net508));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__24__u_dcfifo_rx_u_din_buffer_data_reg_0__25__509 (.o(net509));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__24__u_dcfifo_rx_u_din_buffer_data_reg_0__25__510 (.o(net510));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__26__u_dcfifo_rx_u_din_buffer_data_reg_0__27__511 (.o(net511));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__26__u_dcfifo_rx_u_din_buffer_data_reg_0__27__512 (.o(net512));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__28__u_dcfifo_rx_u_din_buffer_data_reg_0__29__513 (.o(net513));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__28__u_dcfifo_rx_u_din_buffer_data_reg_0__29__514 (.o(net514));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__2__u_dcfifo_rx_u_din_buffer_data_reg_0__3__515 (.o(net515));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__2__u_dcfifo_rx_u_din_buffer_data_reg_0__3__516 (.o(net516));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__30__u_dcfifo_rx_u_din_buffer_data_reg_0__31__517 (.o(net517));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__30__u_dcfifo_rx_u_din_buffer_data_reg_0__31__518 (.o(net518));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__4__u_dcfifo_rx_u_din_buffer_data_reg_0__5__519 (.o(net519));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__4__u_dcfifo_rx_u_din_buffer_data_reg_0__5__520 (.o(net520));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__6__u_dcfifo_rx_u_din_buffer_data_reg_0__7__521 (.o(net521));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__6__u_dcfifo_rx_u_din_buffer_data_reg_0__7__522 (.o(net522));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__8__u_dcfifo_rx_u_din_buffer_data_reg_0__9__523 (.o(net523));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__8__u_dcfifo_rx_u_din_buffer_data_reg_0__9__524 (.o(net524));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__0__u_dcfifo_rx_u_din_buffer_data_reg_1__1__525 (.o(net525));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__0__u_dcfifo_rx_u_din_buffer_data_reg_1__1__526 (.o(net526));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__10__u_dcfifo_rx_u_din_buffer_data_reg_1__11__527 (.o(net527));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__10__u_dcfifo_rx_u_din_buffer_data_reg_1__11__528 (.o(net528));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__12__u_dcfifo_rx_u_din_buffer_data_reg_1__13__529 (.o(net529));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__12__u_dcfifo_rx_u_din_buffer_data_reg_1__13__530 (.o(net530));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__14__u_dcfifo_rx_u_din_buffer_data_reg_1__15__531 (.o(net531));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__14__u_dcfifo_rx_u_din_buffer_data_reg_1__15__532 (.o(net532));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__16__u_dcfifo_rx_u_din_buffer_data_reg_1__17__533 (.o(net533));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__16__u_dcfifo_rx_u_din_buffer_data_reg_1__17__534 (.o(net534));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__18__u_dcfifo_rx_u_din_buffer_data_reg_1__19__535 (.o(net535));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__18__u_dcfifo_rx_u_din_buffer_data_reg_1__19__536 (.o(net536));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__20__u_dcfifo_rx_u_din_buffer_data_reg_1__21__537 (.o(net537));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__20__u_dcfifo_rx_u_din_buffer_data_reg_1__21__538 (.o(net538));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__22__u_dcfifo_rx_u_din_buffer_data_reg_1__23__539 (.o(net539));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__22__u_dcfifo_rx_u_din_buffer_data_reg_1__23__540 (.o(net540));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__24__u_dcfifo_rx_u_din_buffer_data_reg_1__25__541 (.o(net541));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__24__u_dcfifo_rx_u_din_buffer_data_reg_1__25__542 (.o(net542));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__26__u_dcfifo_rx_u_din_buffer_data_reg_1__27__543 (.o(net543));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__26__u_dcfifo_rx_u_din_buffer_data_reg_1__27__544 (.o(net544));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__28__u_dcfifo_rx_u_din_buffer_data_reg_1__29__545 (.o(net545));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__28__u_dcfifo_rx_u_din_buffer_data_reg_1__29__546 (.o(net546));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__2__u_dcfifo_rx_u_din_buffer_data_reg_1__3__547 (.o(net547));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__2__u_dcfifo_rx_u_din_buffer_data_reg_1__3__548 (.o(net548));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__30__u_dcfifo_rx_u_din_buffer_data_reg_1__31__549 (.o(net549));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__30__u_dcfifo_rx_u_din_buffer_data_reg_1__31__550 (.o(net550));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__4__u_dcfifo_rx_u_din_buffer_data_reg_1__5__551 (.o(net551));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__4__u_dcfifo_rx_u_din_buffer_data_reg_1__5__552 (.o(net552));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__6__u_dcfifo_rx_u_din_buffer_data_reg_1__7__553 (.o(net553));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__6__u_dcfifo_rx_u_din_buffer_data_reg_1__7__554 (.o(net554));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__8__u_dcfifo_rx_u_din_buffer_data_reg_1__9__555 (.o(net555));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__8__u_dcfifo_rx_u_din_buffer_data_reg_1__9__556 (.o(net556));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__0__u_dcfifo_rx_u_din_buffer_data_reg_2__1__557 (.o(net557));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__0__u_dcfifo_rx_u_din_buffer_data_reg_2__1__558 (.o(net558));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__10__u_dcfifo_rx_u_din_buffer_data_reg_2__11__559 (.o(net559));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__10__u_dcfifo_rx_u_din_buffer_data_reg_2__11__560 (.o(net560));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__12__u_dcfifo_rx_u_din_buffer_data_reg_2__13__561 (.o(net561));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__12__u_dcfifo_rx_u_din_buffer_data_reg_2__13__562 (.o(net562));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__14__u_dcfifo_rx_u_din_buffer_data_reg_2__15__563 (.o(net563));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__14__u_dcfifo_rx_u_din_buffer_data_reg_2__15__564 (.o(net564));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__16__u_dcfifo_rx_u_din_buffer_data_reg_2__17__565 (.o(net565));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__16__u_dcfifo_rx_u_din_buffer_data_reg_2__17__566 (.o(net566));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__18__u_dcfifo_rx_u_din_buffer_data_reg_2__19__567 (.o(net567));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__18__u_dcfifo_rx_u_din_buffer_data_reg_2__19__568 (.o(net568));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__20__u_dcfifo_rx_u_din_buffer_data_reg_2__21__569 (.o(net569));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__20__u_dcfifo_rx_u_din_buffer_data_reg_2__21__570 (.o(net570));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__22__u_dcfifo_rx_u_din_buffer_data_reg_2__23__571 (.o(net571));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__22__u_dcfifo_rx_u_din_buffer_data_reg_2__23__572 (.o(net572));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__24__u_dcfifo_rx_u_din_buffer_data_reg_2__25__573 (.o(net573));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__24__u_dcfifo_rx_u_din_buffer_data_reg_2__25__574 (.o(net574));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__26__u_dcfifo_rx_u_din_buffer_data_reg_2__27__575 (.o(net575));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__26__u_dcfifo_rx_u_din_buffer_data_reg_2__27__576 (.o(net576));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__28__u_dcfifo_rx_u_din_buffer_data_reg_2__29__577 (.o(net577));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__28__u_dcfifo_rx_u_din_buffer_data_reg_2__29__578 (.o(net578));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__2__u_dcfifo_rx_u_din_buffer_data_reg_2__3__579 (.o(net579));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__2__u_dcfifo_rx_u_din_buffer_data_reg_2__3__580 (.o(net580));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__30__u_dcfifo_rx_u_din_buffer_data_reg_2__31__581 (.o(net581));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__30__u_dcfifo_rx_u_din_buffer_data_reg_2__31__582 (.o(net582));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__4__u_dcfifo_rx_u_din_buffer_data_reg_2__5__583 (.o(net583));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__4__u_dcfifo_rx_u_din_buffer_data_reg_2__5__584 (.o(net584));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__6__u_dcfifo_rx_u_din_buffer_data_reg_2__7__585 (.o(net585));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__6__u_dcfifo_rx_u_din_buffer_data_reg_2__7__586 (.o(net586));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__8__u_dcfifo_rx_u_din_buffer_data_reg_2__9__587 (.o(net587));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__8__u_dcfifo_rx_u_din_buffer_data_reg_2__9__588 (.o(net588));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__0__u_dcfifo_rx_u_din_buffer_data_reg_3__1__589 (.o(net589));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__0__u_dcfifo_rx_u_din_buffer_data_reg_3__1__590 (.o(net590));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__10__u_dcfifo_rx_u_din_buffer_data_reg_3__11__591 (.o(net591));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__10__u_dcfifo_rx_u_din_buffer_data_reg_3__11__592 (.o(net592));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__12__u_dcfifo_rx_u_din_buffer_data_reg_3__13__593 (.o(net593));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__12__u_dcfifo_rx_u_din_buffer_data_reg_3__13__594 (.o(net594));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__14__u_dcfifo_rx_u_din_buffer_data_reg_3__15__595 (.o(net595));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__14__u_dcfifo_rx_u_din_buffer_data_reg_3__15__596 (.o(net596));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__16__u_dcfifo_rx_u_din_buffer_data_reg_3__17__597 (.o(net597));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__16__u_dcfifo_rx_u_din_buffer_data_reg_3__17__598 (.o(net598));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__18__u_dcfifo_rx_u_din_buffer_data_reg_3__19__599 (.o(net599));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__18__u_dcfifo_rx_u_din_buffer_data_reg_3__19__600 (.o(net600));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__20__u_dcfifo_rx_u_din_buffer_data_reg_3__21__601 (.o(net601));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__20__u_dcfifo_rx_u_din_buffer_data_reg_3__21__602 (.o(net602));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__22__u_dcfifo_rx_u_din_buffer_data_reg_3__23__603 (.o(net603));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__22__u_dcfifo_rx_u_din_buffer_data_reg_3__23__604 (.o(net604));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__24__u_dcfifo_rx_u_din_buffer_data_reg_3__25__605 (.o(net605));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__24__u_dcfifo_rx_u_din_buffer_data_reg_3__25__606 (.o(net606));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__26__u_dcfifo_rx_u_din_buffer_data_reg_3__27__607 (.o(net607));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__26__u_dcfifo_rx_u_din_buffer_data_reg_3__27__608 (.o(net608));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__28__u_dcfifo_rx_u_din_buffer_data_reg_3__29__609 (.o(net609));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__28__u_dcfifo_rx_u_din_buffer_data_reg_3__29__610 (.o(net610));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__2__u_dcfifo_rx_u_din_buffer_data_reg_3__3__611 (.o(net611));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__2__u_dcfifo_rx_u_din_buffer_data_reg_3__3__612 (.o(net612));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__30__u_dcfifo_rx_u_din_buffer_data_reg_3__31__613 (.o(net613));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__30__u_dcfifo_rx_u_din_buffer_data_reg_3__31__614 (.o(net614));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__4__u_dcfifo_rx_u_din_buffer_data_reg_3__5__615 (.o(net615));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__4__u_dcfifo_rx_u_din_buffer_data_reg_3__5__616 (.o(net616));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__6__u_dcfifo_rx_u_din_buffer_data_reg_3__7__617 (.o(net617));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__6__u_dcfifo_rx_u_din_buffer_data_reg_3__7__618 (.o(net618));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__8__u_dcfifo_rx_u_din_buffer_data_reg_3__9__619 (.o(net619));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__8__u_dcfifo_rx_u_din_buffer_data_reg_3__9__620 (.o(net620));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__0__u_dcfifo_rx_u_din_buffer_data_reg_4__1__621 (.o(net621));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__0__u_dcfifo_rx_u_din_buffer_data_reg_4__1__622 (.o(net622));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__10__u_dcfifo_rx_u_din_buffer_data_reg_4__11__623 (.o(net623));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__10__u_dcfifo_rx_u_din_buffer_data_reg_4__11__624 (.o(net624));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__12__u_dcfifo_rx_u_din_buffer_data_reg_4__13__625 (.o(net625));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__12__u_dcfifo_rx_u_din_buffer_data_reg_4__13__626 (.o(net626));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__14__u_dcfifo_rx_u_din_buffer_data_reg_4__15__627 (.o(net627));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__14__u_dcfifo_rx_u_din_buffer_data_reg_4__15__628 (.o(net628));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__16__u_dcfifo_rx_u_din_buffer_data_reg_4__17__629 (.o(net629));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__16__u_dcfifo_rx_u_din_buffer_data_reg_4__17__630 (.o(net630));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__18__u_dcfifo_rx_u_din_buffer_data_reg_4__19__631 (.o(net631));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__18__u_dcfifo_rx_u_din_buffer_data_reg_4__19__632 (.o(net632));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__20__u_dcfifo_rx_u_din_buffer_data_reg_4__21__633 (.o(net633));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__20__u_dcfifo_rx_u_din_buffer_data_reg_4__21__634 (.o(net634));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__22__u_dcfifo_rx_u_din_buffer_data_reg_4__23__635 (.o(net635));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__22__u_dcfifo_rx_u_din_buffer_data_reg_4__23__636 (.o(net636));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__24__u_dcfifo_rx_u_din_buffer_data_reg_4__25__637 (.o(net637));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__24__u_dcfifo_rx_u_din_buffer_data_reg_4__25__638 (.o(net638));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__26__u_dcfifo_rx_u_din_buffer_data_reg_4__27__639 (.o(net639));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__26__u_dcfifo_rx_u_din_buffer_data_reg_4__27__640 (.o(net640));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__28__u_dcfifo_rx_u_din_buffer_data_reg_4__29__641 (.o(net641));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__28__u_dcfifo_rx_u_din_buffer_data_reg_4__29__642 (.o(net642));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__2__u_dcfifo_rx_u_din_buffer_data_reg_4__3__643 (.o(net643));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__2__u_dcfifo_rx_u_din_buffer_data_reg_4__3__644 (.o(net644));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__30__u_dcfifo_rx_u_din_buffer_data_reg_4__31__645 (.o(net645));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__30__u_dcfifo_rx_u_din_buffer_data_reg_4__31__646 (.o(net646));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__4__u_dcfifo_rx_u_din_buffer_data_reg_4__5__647 (.o(net647));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__4__u_dcfifo_rx_u_din_buffer_data_reg_4__5__648 (.o(net648));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__6__u_dcfifo_rx_u_din_buffer_data_reg_4__7__649 (.o(net649));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__6__u_dcfifo_rx_u_din_buffer_data_reg_4__7__650 (.o(net650));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__8__u_dcfifo_rx_u_din_buffer_data_reg_4__9__651 (.o(net651));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__8__u_dcfifo_rx_u_din_buffer_data_reg_4__9__652 (.o(net652));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__0__u_dcfifo_rx_u_din_buffer_data_reg_5__1__653 (.o(net653));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__0__u_dcfifo_rx_u_din_buffer_data_reg_5__1__654 (.o(net654));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__10__u_dcfifo_rx_u_din_buffer_data_reg_5__11__655 (.o(net655));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__10__u_dcfifo_rx_u_din_buffer_data_reg_5__11__656 (.o(net656));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__12__u_dcfifo_rx_u_din_buffer_data_reg_5__13__657 (.o(net657));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__12__u_dcfifo_rx_u_din_buffer_data_reg_5__13__658 (.o(net658));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__14__u_dcfifo_rx_u_din_buffer_data_reg_5__15__659 (.o(net659));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__14__u_dcfifo_rx_u_din_buffer_data_reg_5__15__660 (.o(net660));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__16__u_dcfifo_rx_u_din_buffer_data_reg_5__17__661 (.o(net661));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__16__u_dcfifo_rx_u_din_buffer_data_reg_5__17__662 (.o(net662));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__18__u_dcfifo_rx_u_din_buffer_data_reg_5__19__663 (.o(net663));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__18__u_dcfifo_rx_u_din_buffer_data_reg_5__19__664 (.o(net664));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__20__u_dcfifo_rx_u_din_buffer_data_reg_5__21__665 (.o(net665));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__20__u_dcfifo_rx_u_din_buffer_data_reg_5__21__666 (.o(net666));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__22__u_dcfifo_rx_u_din_buffer_data_reg_5__23__667 (.o(net667));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__22__u_dcfifo_rx_u_din_buffer_data_reg_5__23__668 (.o(net668));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__24__u_dcfifo_rx_u_din_buffer_data_reg_5__25__669 (.o(net669));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__24__u_dcfifo_rx_u_din_buffer_data_reg_5__25__670 (.o(net670));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__26__u_dcfifo_rx_u_din_buffer_data_reg_5__27__671 (.o(net671));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__26__u_dcfifo_rx_u_din_buffer_data_reg_5__27__672 (.o(net672));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__28__u_dcfifo_rx_u_din_buffer_data_reg_5__29__673 (.o(net673));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__28__u_dcfifo_rx_u_din_buffer_data_reg_5__29__674 (.o(net674));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__2__u_dcfifo_rx_u_din_buffer_data_reg_5__3__675 (.o(net675));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__2__u_dcfifo_rx_u_din_buffer_data_reg_5__3__676 (.o(net676));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__30__u_dcfifo_rx_u_din_buffer_data_reg_5__31__677 (.o(net677));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__30__u_dcfifo_rx_u_din_buffer_data_reg_5__31__678 (.o(net678));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__4__u_dcfifo_rx_u_din_buffer_data_reg_5__5__679 (.o(net679));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__4__u_dcfifo_rx_u_din_buffer_data_reg_5__5__680 (.o(net680));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__6__u_dcfifo_rx_u_din_buffer_data_reg_5__7__681 (.o(net681));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__6__u_dcfifo_rx_u_din_buffer_data_reg_5__7__682 (.o(net682));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__8__u_dcfifo_rx_u_din_buffer_data_reg_5__9__683 (.o(net683));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__8__u_dcfifo_rx_u_din_buffer_data_reg_5__9__684 (.o(net684));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__0__u_dcfifo_rx_u_din_buffer_data_reg_6__1__685 (.o(net685));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__0__u_dcfifo_rx_u_din_buffer_data_reg_6__1__686 (.o(net686));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__10__u_dcfifo_rx_u_din_buffer_data_reg_6__11__687 (.o(net687));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__10__u_dcfifo_rx_u_din_buffer_data_reg_6__11__688 (.o(net688));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__12__u_dcfifo_rx_u_din_buffer_data_reg_6__13__689 (.o(net689));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__12__u_dcfifo_rx_u_din_buffer_data_reg_6__13__690 (.o(net690));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__14__u_dcfifo_rx_u_din_buffer_data_reg_6__15__691 (.o(net691));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__14__u_dcfifo_rx_u_din_buffer_data_reg_6__15__692 (.o(net692));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__16__u_dcfifo_rx_u_din_buffer_data_reg_6__17__693 (.o(net693));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__16__u_dcfifo_rx_u_din_buffer_data_reg_6__17__694 (.o(net694));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__18__u_dcfifo_rx_u_din_buffer_data_reg_6__19__695 (.o(net695));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__18__u_dcfifo_rx_u_din_buffer_data_reg_6__19__696 (.o(net696));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__20__u_dcfifo_rx_u_din_buffer_data_reg_6__21__697 (.o(net697));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__20__u_dcfifo_rx_u_din_buffer_data_reg_6__21__698 (.o(net698));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__22__u_dcfifo_rx_u_din_buffer_data_reg_6__23__699 (.o(net699));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__22__u_dcfifo_rx_u_din_buffer_data_reg_6__23__700 (.o(net700));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__24__u_dcfifo_rx_u_din_buffer_data_reg_6__25__701 (.o(net701));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__24__u_dcfifo_rx_u_din_buffer_data_reg_6__25__702 (.o(net702));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__26__u_dcfifo_rx_u_din_buffer_data_reg_6__27__703 (.o(net703));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__26__u_dcfifo_rx_u_din_buffer_data_reg_6__27__704 (.o(net704));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__28__u_dcfifo_rx_u_din_buffer_data_reg_6__29__705 (.o(net705));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__28__u_dcfifo_rx_u_din_buffer_data_reg_6__29__706 (.o(net706));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__2__u_dcfifo_rx_u_din_buffer_data_reg_6__3__707 (.o(net707));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__2__u_dcfifo_rx_u_din_buffer_data_reg_6__3__708 (.o(net708));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__30__u_dcfifo_rx_u_din_buffer_data_reg_6__31__709 (.o(net709));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__30__u_dcfifo_rx_u_din_buffer_data_reg_6__31__710 (.o(net710));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__4__u_dcfifo_rx_u_din_buffer_data_reg_6__5__711 (.o(net711));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__4__u_dcfifo_rx_u_din_buffer_data_reg_6__5__712 (.o(net712));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__6__u_dcfifo_rx_u_din_buffer_data_reg_6__7__713 (.o(net713));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__6__u_dcfifo_rx_u_din_buffer_data_reg_6__7__714 (.o(net714));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__8__u_dcfifo_rx_u_din_buffer_data_reg_6__9__715 (.o(net715));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__8__u_dcfifo_rx_u_din_buffer_data_reg_6__9__716 (.o(net716));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__0__u_dcfifo_rx_u_din_buffer_data_reg_7__1__717 (.o(net717));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__0__u_dcfifo_rx_u_din_buffer_data_reg_7__1__718 (.o(net718));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__10__u_dcfifo_rx_u_din_buffer_data_reg_7__11__719 (.o(net719));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__10__u_dcfifo_rx_u_din_buffer_data_reg_7__11__720 (.o(net720));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__12__u_dcfifo_rx_u_din_buffer_data_reg_7__13__721 (.o(net721));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__12__u_dcfifo_rx_u_din_buffer_data_reg_7__13__722 (.o(net722));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__14__u_dcfifo_rx_u_din_buffer_data_reg_7__15__723 (.o(net723));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__14__u_dcfifo_rx_u_din_buffer_data_reg_7__15__724 (.o(net724));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__16__u_dcfifo_rx_u_din_buffer_data_reg_7__17__725 (.o(net725));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__16__u_dcfifo_rx_u_din_buffer_data_reg_7__17__726 (.o(net726));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__18__u_dcfifo_rx_u_din_buffer_data_reg_7__19__727 (.o(net727));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__18__u_dcfifo_rx_u_din_buffer_data_reg_7__19__728 (.o(net728));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__20__u_dcfifo_rx_u_din_buffer_data_reg_7__21__729 (.o(net729));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__20__u_dcfifo_rx_u_din_buffer_data_reg_7__21__730 (.o(net730));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__22__u_dcfifo_rx_u_din_buffer_data_reg_7__23__731 (.o(net731));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__22__u_dcfifo_rx_u_din_buffer_data_reg_7__23__732 (.o(net732));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__24__u_dcfifo_rx_u_din_buffer_data_reg_7__25__733 (.o(net733));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__24__u_dcfifo_rx_u_din_buffer_data_reg_7__25__734 (.o(net734));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__26__u_dcfifo_rx_u_din_buffer_data_reg_7__27__735 (.o(net735));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__26__u_dcfifo_rx_u_din_buffer_data_reg_7__27__736 (.o(net736));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__28__u_dcfifo_rx_u_din_buffer_data_reg_7__29__737 (.o(net737));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__28__u_dcfifo_rx_u_din_buffer_data_reg_7__29__738 (.o(net738));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__2__u_dcfifo_rx_u_din_buffer_data_reg_7__3__739 (.o(net739));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__2__u_dcfifo_rx_u_din_buffer_data_reg_7__3__740 (.o(net740));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__30__u_dcfifo_rx_u_din_buffer_data_reg_7__31__741 (.o(net741));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__30__u_dcfifo_rx_u_din_buffer_data_reg_7__31__742 (.o(net742));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__4__u_dcfifo_rx_u_din_buffer_data_reg_7__5__743 (.o(net743));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__4__u_dcfifo_rx_u_din_buffer_data_reg_7__5__744 (.o(net744));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__6__u_dcfifo_rx_u_din_buffer_data_reg_7__7__745 (.o(net745));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__6__u_dcfifo_rx_u_din_buffer_data_reg_7__7__746 (.o(net746));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__8__u_dcfifo_rx_u_din_buffer_data_reg_7__9__747 (.o(net747));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__8__u_dcfifo_rx_u_din_buffer_data_reg_7__9__748 (.o(net748));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_full_full_synch_d_middle_reg_0__u_dcfifo_rx_u_din_full_full_synch_d_out_reg_0__749 (.o(net749));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_full_full_synch_d_middle_reg_0__u_dcfifo_rx_u_din_full_full_synch_d_out_reg_0__750 (.o(net750));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_full_latched_full_s_reg_u_dcfifo_tx_u_dout_empty_synch_d_out_reg_1__751 (.o(net751));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_full_latched_full_s_reg_u_dcfifo_tx_u_dout_empty_synch_d_out_reg_1__752 (.o(net752));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_write_tr_clk_gate_state_reg_latch_753 (.o(net753));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_write_tr_state_reg_0__u_dcfifo_rx_u_din_write_tr_state_reg_1__754 (.o(net754));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_write_tr_state_reg_0__u_dcfifo_rx_u_din_write_tr_state_reg_1__755 (.o(net755));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_write_tr_state_reg_2__756 (.o(net756));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_write_tr_state_reg_3__757 (.o(net757));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_write_tr_state_reg_4__u_dcfifo_rx_u_din_write_tr_state_reg_5__758 (.o(net758));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_write_tr_state_reg_4__u_dcfifo_rx_u_din_write_tr_state_reg_5__759 (.o(net759));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_write_tr_state_reg_6__u_dcfifo_rx_u_din_write_tr_state_reg_7__760 (.o(net760));
 b15tilo00an1n03x5 u_dcfifo_rx_u_din_write_tr_state_reg_6__u_dcfifo_rx_u_din_write_tr_state_reg_7__761 (.o(net761));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_0__u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_1__762 (.o(net762));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_0__u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_1__763 (.o(net763));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_2__764 (.o(net764));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_3__765 (.o(net765));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_4__u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_5__766 (.o(net766));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_4__u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_5__767 (.o(net767));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_6__u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_7__768 (.o(net768));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_6__u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_7__769 (.o(net769));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_0__u_dcfifo_rx_u_dout_empty_synch_d_out_reg_1__770 (.o(net770));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_0__u_dcfifo_rx_u_dout_empty_synch_d_out_reg_1__771 (.o(net771));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_2__772 (.o(net772));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_3__773 (.o(net773));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_4__u_dcfifo_rx_u_dout_empty_synch_d_out_reg_5__774 (.o(net774));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_4__u_dcfifo_rx_u_dout_empty_synch_d_out_reg_5__775 (.o(net775));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_6__u_dcfifo_rx_u_dout_empty_synch_d_out_reg_7__776 (.o(net776));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_6__u_dcfifo_rx_u_dout_empty_synch_d_out_reg_7__777 (.o(net777));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_read_tr_clk_gate_state_reg_latch_778 (.o(net778));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_read_tr_state_reg_0__779 (.o(net779));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_read_tr_state_reg_1__780 (.o(net780));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_read_tr_state_reg_2__u_dcfifo_rx_u_dout_read_tr_state_reg_3__781 (.o(net781));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_read_tr_state_reg_2__u_dcfifo_rx_u_dout_read_tr_state_reg_3__782 (.o(net782));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_read_tr_state_reg_4__u_dcfifo_rx_u_dout_read_tr_state_reg_5__783 (.o(net783));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_read_tr_state_reg_4__u_dcfifo_rx_u_dout_read_tr_state_reg_5__784 (.o(net784));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_read_tr_state_reg_6__u_dcfifo_rx_u_dout_read_tr_state_reg_7__785 (.o(net785));
 b15tilo00an1n03x5 u_dcfifo_rx_u_dout_read_tr_state_reg_6__u_dcfifo_rx_u_dout_read_tr_state_reg_7__786 (.o(net786));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_0__0_latch_787 (.o(net787));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_0__latch_788 (.o(net788));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_1__0_latch_789 (.o(net789));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_1__latch_790 (.o(net790));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_2__0_latch_791 (.o(net791));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_2__latch_792 (.o(net792));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_3__0_latch_793 (.o(net793));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_3__latch_794 (.o(net794));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_4__0_latch_795 (.o(net795));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_4__latch_796 (.o(net796));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_5__0_latch_797 (.o(net797));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_5__latch_798 (.o(net798));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_6__0_latch_799 (.o(net799));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_6__latch_800 (.o(net800));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_7__0_latch_801 (.o(net801));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_clk_gate_data_reg_7__latch_802 (.o(net802));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__0__u_dcfifo_tx_u_din_buffer_data_reg_0__1__803 (.o(net803));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__0__u_dcfifo_tx_u_din_buffer_data_reg_0__1__804 (.o(net804));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__10__u_dcfifo_tx_u_din_buffer_data_reg_0__11__805 (.o(net805));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__10__u_dcfifo_tx_u_din_buffer_data_reg_0__11__806 (.o(net806));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__12__u_dcfifo_tx_u_din_buffer_data_reg_0__13__807 (.o(net807));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__12__u_dcfifo_tx_u_din_buffer_data_reg_0__13__808 (.o(net808));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__14__u_dcfifo_tx_u_din_buffer_data_reg_0__15__809 (.o(net809));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__14__u_dcfifo_tx_u_din_buffer_data_reg_0__15__810 (.o(net810));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__16__u_dcfifo_tx_u_din_buffer_data_reg_0__17__811 (.o(net811));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__16__u_dcfifo_tx_u_din_buffer_data_reg_0__17__812 (.o(net812));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__18__u_dcfifo_tx_u_din_buffer_data_reg_0__19__813 (.o(net813));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__18__u_dcfifo_tx_u_din_buffer_data_reg_0__19__814 (.o(net814));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__20__u_dcfifo_tx_u_din_buffer_data_reg_0__21__815 (.o(net815));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__20__u_dcfifo_tx_u_din_buffer_data_reg_0__21__816 (.o(net816));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__22__u_dcfifo_tx_u_din_buffer_data_reg_0__23__817 (.o(net817));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__22__u_dcfifo_tx_u_din_buffer_data_reg_0__23__818 (.o(net818));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__24__u_dcfifo_tx_u_din_buffer_data_reg_0__25__819 (.o(net819));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__24__u_dcfifo_tx_u_din_buffer_data_reg_0__25__820 (.o(net820));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__26__u_dcfifo_tx_u_din_buffer_data_reg_0__27__821 (.o(net821));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__26__u_dcfifo_tx_u_din_buffer_data_reg_0__27__822 (.o(net822));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__28__u_dcfifo_tx_u_din_buffer_data_reg_0__29__823 (.o(net823));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__28__u_dcfifo_tx_u_din_buffer_data_reg_0__29__824 (.o(net824));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__2__u_dcfifo_tx_u_din_buffer_data_reg_0__3__825 (.o(net825));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__2__u_dcfifo_tx_u_din_buffer_data_reg_0__3__826 (.o(net826));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__30__u_dcfifo_tx_u_din_buffer_data_reg_0__31__827 (.o(net827));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__30__u_dcfifo_tx_u_din_buffer_data_reg_0__31__828 (.o(net828));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__4__u_dcfifo_tx_u_din_buffer_data_reg_0__5__829 (.o(net829));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__4__u_dcfifo_tx_u_din_buffer_data_reg_0__5__830 (.o(net830));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__6__u_dcfifo_tx_u_din_buffer_data_reg_0__7__831 (.o(net831));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__6__u_dcfifo_tx_u_din_buffer_data_reg_0__7__832 (.o(net832));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__8__u_dcfifo_tx_u_din_buffer_data_reg_0__9__833 (.o(net833));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__8__u_dcfifo_tx_u_din_buffer_data_reg_0__9__834 (.o(net834));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__0__u_dcfifo_tx_u_din_buffer_data_reg_1__1__835 (.o(net835));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__0__u_dcfifo_tx_u_din_buffer_data_reg_1__1__836 (.o(net836));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__10__u_dcfifo_tx_u_din_buffer_data_reg_1__11__837 (.o(net837));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__10__u_dcfifo_tx_u_din_buffer_data_reg_1__11__838 (.o(net838));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__12__u_dcfifo_tx_u_din_buffer_data_reg_1__13__839 (.o(net839));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__12__u_dcfifo_tx_u_din_buffer_data_reg_1__13__840 (.o(net840));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__14__u_dcfifo_tx_u_din_buffer_data_reg_1__15__841 (.o(net841));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__14__u_dcfifo_tx_u_din_buffer_data_reg_1__15__842 (.o(net842));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__16__u_dcfifo_tx_u_din_buffer_data_reg_1__17__843 (.o(net843));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__16__u_dcfifo_tx_u_din_buffer_data_reg_1__17__844 (.o(net844));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__18__u_dcfifo_tx_u_din_buffer_data_reg_1__19__845 (.o(net845));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__18__u_dcfifo_tx_u_din_buffer_data_reg_1__19__846 (.o(net846));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__20__u_dcfifo_tx_u_din_buffer_data_reg_1__21__847 (.o(net847));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__20__u_dcfifo_tx_u_din_buffer_data_reg_1__21__848 (.o(net848));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__22__u_dcfifo_tx_u_din_buffer_data_reg_1__23__849 (.o(net849));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__22__u_dcfifo_tx_u_din_buffer_data_reg_1__23__850 (.o(net850));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__24__u_dcfifo_tx_u_din_buffer_data_reg_1__25__851 (.o(net851));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__24__u_dcfifo_tx_u_din_buffer_data_reg_1__25__852 (.o(net852));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__26__u_dcfifo_tx_u_din_buffer_data_reg_1__27__853 (.o(net853));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__26__u_dcfifo_tx_u_din_buffer_data_reg_1__27__854 (.o(net854));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__28__u_dcfifo_tx_u_din_buffer_data_reg_1__29__855 (.o(net855));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__28__u_dcfifo_tx_u_din_buffer_data_reg_1__29__856 (.o(net856));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__2__u_dcfifo_tx_u_din_buffer_data_reg_1__3__857 (.o(net857));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__2__u_dcfifo_tx_u_din_buffer_data_reg_1__3__858 (.o(net858));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__30__u_dcfifo_tx_u_din_buffer_data_reg_1__31__859 (.o(net859));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__30__u_dcfifo_tx_u_din_buffer_data_reg_1__31__860 (.o(net860));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__4__u_dcfifo_tx_u_din_buffer_data_reg_1__5__861 (.o(net861));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__4__u_dcfifo_tx_u_din_buffer_data_reg_1__5__862 (.o(net862));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__6__u_dcfifo_tx_u_din_buffer_data_reg_1__7__863 (.o(net863));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__6__u_dcfifo_tx_u_din_buffer_data_reg_1__7__864 (.o(net864));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__8__u_dcfifo_tx_u_din_buffer_data_reg_1__9__865 (.o(net865));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__8__u_dcfifo_tx_u_din_buffer_data_reg_1__9__866 (.o(net866));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__0__u_dcfifo_tx_u_din_buffer_data_reg_2__1__867 (.o(net867));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__0__u_dcfifo_tx_u_din_buffer_data_reg_2__1__868 (.o(net868));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__10__u_dcfifo_tx_u_din_buffer_data_reg_2__11__869 (.o(net869));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__10__u_dcfifo_tx_u_din_buffer_data_reg_2__11__870 (.o(net870));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__12__u_dcfifo_tx_u_din_buffer_data_reg_2__13__871 (.o(net871));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__12__u_dcfifo_tx_u_din_buffer_data_reg_2__13__872 (.o(net872));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__14__u_dcfifo_tx_u_din_buffer_data_reg_2__15__873 (.o(net873));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__14__u_dcfifo_tx_u_din_buffer_data_reg_2__15__874 (.o(net874));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__16__u_dcfifo_tx_u_din_buffer_data_reg_2__17__875 (.o(net875));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__16__u_dcfifo_tx_u_din_buffer_data_reg_2__17__876 (.o(net876));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__18__u_dcfifo_tx_u_din_buffer_data_reg_2__19__877 (.o(net877));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__18__u_dcfifo_tx_u_din_buffer_data_reg_2__19__878 (.o(net878));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__20__u_dcfifo_tx_u_din_buffer_data_reg_2__21__879 (.o(net879));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__20__u_dcfifo_tx_u_din_buffer_data_reg_2__21__880 (.o(net880));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__22__u_dcfifo_tx_u_din_buffer_data_reg_2__23__881 (.o(net881));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__22__u_dcfifo_tx_u_din_buffer_data_reg_2__23__882 (.o(net882));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__24__u_dcfifo_tx_u_din_buffer_data_reg_2__25__883 (.o(net883));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__24__u_dcfifo_tx_u_din_buffer_data_reg_2__25__884 (.o(net884));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__26__u_dcfifo_tx_u_din_buffer_data_reg_2__27__885 (.o(net885));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__26__u_dcfifo_tx_u_din_buffer_data_reg_2__27__886 (.o(net886));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__28__u_dcfifo_tx_u_din_buffer_data_reg_2__29__887 (.o(net887));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__28__u_dcfifo_tx_u_din_buffer_data_reg_2__29__888 (.o(net888));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__2__u_dcfifo_tx_u_din_buffer_data_reg_2__3__889 (.o(net889));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__2__u_dcfifo_tx_u_din_buffer_data_reg_2__3__890 (.o(net890));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__30__u_dcfifo_tx_u_din_buffer_data_reg_2__31__891 (.o(net891));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__30__u_dcfifo_tx_u_din_buffer_data_reg_2__31__892 (.o(net892));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__4__u_dcfifo_tx_u_din_buffer_data_reg_2__5__893 (.o(net893));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__4__u_dcfifo_tx_u_din_buffer_data_reg_2__5__894 (.o(net894));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__6__u_dcfifo_tx_u_din_buffer_data_reg_2__7__895 (.o(net895));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__6__u_dcfifo_tx_u_din_buffer_data_reg_2__7__896 (.o(net896));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__8__u_dcfifo_tx_u_din_buffer_data_reg_2__9__897 (.o(net897));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__8__u_dcfifo_tx_u_din_buffer_data_reg_2__9__898 (.o(net898));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__0__u_dcfifo_tx_u_din_buffer_data_reg_3__1__899 (.o(net899));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__0__u_dcfifo_tx_u_din_buffer_data_reg_3__1__900 (.o(net900));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__10__u_dcfifo_tx_u_din_buffer_data_reg_3__11__901 (.o(net901));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__10__u_dcfifo_tx_u_din_buffer_data_reg_3__11__902 (.o(net902));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__12__u_dcfifo_tx_u_din_buffer_data_reg_3__13__903 (.o(net903));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__12__u_dcfifo_tx_u_din_buffer_data_reg_3__13__904 (.o(net904));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__14__u_dcfifo_tx_u_din_buffer_data_reg_3__15__905 (.o(net905));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__14__u_dcfifo_tx_u_din_buffer_data_reg_3__15__906 (.o(net906));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__16__u_dcfifo_tx_u_din_buffer_data_reg_3__17__907 (.o(net907));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__16__u_dcfifo_tx_u_din_buffer_data_reg_3__17__908 (.o(net908));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__18__u_dcfifo_tx_u_din_buffer_data_reg_3__19__909 (.o(net909));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__18__u_dcfifo_tx_u_din_buffer_data_reg_3__19__910 (.o(net910));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__20__u_dcfifo_tx_u_din_buffer_data_reg_3__21__911 (.o(net911));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__20__u_dcfifo_tx_u_din_buffer_data_reg_3__21__912 (.o(net912));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__22__u_dcfifo_tx_u_din_buffer_data_reg_3__23__913 (.o(net913));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__22__u_dcfifo_tx_u_din_buffer_data_reg_3__23__914 (.o(net914));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__24__u_dcfifo_tx_u_din_buffer_data_reg_3__25__915 (.o(net915));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__24__u_dcfifo_tx_u_din_buffer_data_reg_3__25__916 (.o(net916));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__26__u_dcfifo_tx_u_din_buffer_data_reg_3__27__917 (.o(net917));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__26__u_dcfifo_tx_u_din_buffer_data_reg_3__27__918 (.o(net918));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__28__u_dcfifo_tx_u_din_buffer_data_reg_3__29__919 (.o(net919));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__28__u_dcfifo_tx_u_din_buffer_data_reg_3__29__920 (.o(net920));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__2__u_dcfifo_tx_u_din_buffer_data_reg_3__3__921 (.o(net921));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__2__u_dcfifo_tx_u_din_buffer_data_reg_3__3__922 (.o(net922));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__30__u_dcfifo_tx_u_din_buffer_data_reg_3__31__923 (.o(net923));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__30__u_dcfifo_tx_u_din_buffer_data_reg_3__31__924 (.o(net924));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__4__u_dcfifo_tx_u_din_buffer_data_reg_3__5__925 (.o(net925));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__4__u_dcfifo_tx_u_din_buffer_data_reg_3__5__926 (.o(net926));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__6__u_dcfifo_tx_u_din_buffer_data_reg_3__7__927 (.o(net927));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__6__u_dcfifo_tx_u_din_buffer_data_reg_3__7__928 (.o(net928));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__8__u_dcfifo_tx_u_din_buffer_data_reg_3__9__929 (.o(net929));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__8__u_dcfifo_tx_u_din_buffer_data_reg_3__9__930 (.o(net930));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__0__u_dcfifo_tx_u_din_buffer_data_reg_4__1__931 (.o(net931));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__0__u_dcfifo_tx_u_din_buffer_data_reg_4__1__932 (.o(net932));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__10__u_dcfifo_tx_u_din_buffer_data_reg_4__11__933 (.o(net933));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__10__u_dcfifo_tx_u_din_buffer_data_reg_4__11__934 (.o(net934));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__12__u_dcfifo_tx_u_din_buffer_data_reg_4__13__935 (.o(net935));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__12__u_dcfifo_tx_u_din_buffer_data_reg_4__13__936 (.o(net936));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__14__u_dcfifo_tx_u_din_buffer_data_reg_4__15__937 (.o(net937));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__14__u_dcfifo_tx_u_din_buffer_data_reg_4__15__938 (.o(net938));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__16__u_dcfifo_tx_u_din_buffer_data_reg_4__17__939 (.o(net939));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__16__u_dcfifo_tx_u_din_buffer_data_reg_4__17__940 (.o(net940));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__18__u_dcfifo_tx_u_din_buffer_data_reg_4__19__941 (.o(net941));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__18__u_dcfifo_tx_u_din_buffer_data_reg_4__19__942 (.o(net942));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__20__u_dcfifo_tx_u_din_buffer_data_reg_4__21__943 (.o(net943));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__20__u_dcfifo_tx_u_din_buffer_data_reg_4__21__944 (.o(net944));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__22__u_dcfifo_tx_u_din_buffer_data_reg_4__23__945 (.o(net945));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__22__u_dcfifo_tx_u_din_buffer_data_reg_4__23__946 (.o(net946));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__24__u_dcfifo_tx_u_din_buffer_data_reg_4__25__947 (.o(net947));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__24__u_dcfifo_tx_u_din_buffer_data_reg_4__25__948 (.o(net948));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__26__u_dcfifo_tx_u_din_buffer_data_reg_4__27__949 (.o(net949));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__26__u_dcfifo_tx_u_din_buffer_data_reg_4__27__950 (.o(net950));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__28__u_dcfifo_tx_u_din_buffer_data_reg_4__29__951 (.o(net951));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__28__u_dcfifo_tx_u_din_buffer_data_reg_4__29__952 (.o(net952));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__2__u_dcfifo_tx_u_din_buffer_data_reg_4__3__953 (.o(net953));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__2__u_dcfifo_tx_u_din_buffer_data_reg_4__3__954 (.o(net954));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__30__u_dcfifo_tx_u_din_buffer_data_reg_4__31__955 (.o(net955));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__30__u_dcfifo_tx_u_din_buffer_data_reg_4__31__956 (.o(net956));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__4__u_dcfifo_tx_u_din_buffer_data_reg_4__5__957 (.o(net957));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__4__u_dcfifo_tx_u_din_buffer_data_reg_4__5__958 (.o(net958));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__6__u_dcfifo_tx_u_din_buffer_data_reg_4__7__959 (.o(net959));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__6__u_dcfifo_tx_u_din_buffer_data_reg_4__7__960 (.o(net960));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__8__u_dcfifo_tx_u_din_buffer_data_reg_4__9__961 (.o(net961));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__8__u_dcfifo_tx_u_din_buffer_data_reg_4__9__962 (.o(net962));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__0__u_dcfifo_tx_u_din_buffer_data_reg_5__1__963 (.o(net963));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__0__u_dcfifo_tx_u_din_buffer_data_reg_5__1__964 (.o(net964));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__10__u_dcfifo_tx_u_din_buffer_data_reg_5__11__965 (.o(net965));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__10__u_dcfifo_tx_u_din_buffer_data_reg_5__11__966 (.o(net966));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__12__u_dcfifo_tx_u_din_buffer_data_reg_5__13__967 (.o(net967));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__12__u_dcfifo_tx_u_din_buffer_data_reg_5__13__968 (.o(net968));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__14__u_dcfifo_tx_u_din_buffer_data_reg_5__15__969 (.o(net969));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__14__u_dcfifo_tx_u_din_buffer_data_reg_5__15__970 (.o(net970));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__16__u_dcfifo_tx_u_din_buffer_data_reg_5__17__971 (.o(net971));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__16__u_dcfifo_tx_u_din_buffer_data_reg_5__17__972 (.o(net972));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__18__u_dcfifo_tx_u_din_buffer_data_reg_5__19__973 (.o(net973));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__18__u_dcfifo_tx_u_din_buffer_data_reg_5__19__974 (.o(net974));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__20__u_dcfifo_tx_u_din_buffer_data_reg_5__21__975 (.o(net975));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__20__u_dcfifo_tx_u_din_buffer_data_reg_5__21__976 (.o(net976));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__22__u_dcfifo_tx_u_din_buffer_data_reg_5__23__977 (.o(net977));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__22__u_dcfifo_tx_u_din_buffer_data_reg_5__23__978 (.o(net978));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__24__u_dcfifo_tx_u_din_buffer_data_reg_5__25__979 (.o(net979));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__24__u_dcfifo_tx_u_din_buffer_data_reg_5__25__980 (.o(net980));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__26__u_dcfifo_tx_u_din_buffer_data_reg_5__27__981 (.o(net981));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__26__u_dcfifo_tx_u_din_buffer_data_reg_5__27__982 (.o(net982));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__28__u_dcfifo_tx_u_din_buffer_data_reg_5__29__983 (.o(net983));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__28__u_dcfifo_tx_u_din_buffer_data_reg_5__29__984 (.o(net984));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__2__u_dcfifo_tx_u_din_buffer_data_reg_5__3__985 (.o(net985));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__2__u_dcfifo_tx_u_din_buffer_data_reg_5__3__986 (.o(net986));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__30__u_dcfifo_tx_u_din_buffer_data_reg_5__31__987 (.o(net987));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__30__u_dcfifo_tx_u_din_buffer_data_reg_5__31__988 (.o(net988));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__4__u_dcfifo_tx_u_din_buffer_data_reg_5__5__989 (.o(net989));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__4__u_dcfifo_tx_u_din_buffer_data_reg_5__5__990 (.o(net990));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__6__u_dcfifo_tx_u_din_buffer_data_reg_5__7__991 (.o(net991));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__6__u_dcfifo_tx_u_din_buffer_data_reg_5__7__992 (.o(net992));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__8__u_dcfifo_tx_u_din_buffer_data_reg_5__9__993 (.o(net993));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__8__u_dcfifo_tx_u_din_buffer_data_reg_5__9__994 (.o(net994));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__0__u_dcfifo_tx_u_din_buffer_data_reg_6__1__995 (.o(net995));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__0__u_dcfifo_tx_u_din_buffer_data_reg_6__1__996 (.o(net996));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__10__u_dcfifo_tx_u_din_buffer_data_reg_6__11__997 (.o(net997));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__10__u_dcfifo_tx_u_din_buffer_data_reg_6__11__998 (.o(net998));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__12__u_dcfifo_tx_u_din_buffer_data_reg_6__13__999 (.o(net999));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__12__u_dcfifo_tx_u_din_buffer_data_reg_6__13__1000 (.o(net1000));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__14__u_dcfifo_tx_u_din_buffer_data_reg_6__15__1001 (.o(net1001));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__14__u_dcfifo_tx_u_din_buffer_data_reg_6__15__1002 (.o(net1002));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__16__u_dcfifo_tx_u_din_buffer_data_reg_6__17__1003 (.o(net1003));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__16__u_dcfifo_tx_u_din_buffer_data_reg_6__17__1004 (.o(net1004));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__18__u_dcfifo_tx_u_din_buffer_data_reg_6__19__1005 (.o(net1005));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__18__u_dcfifo_tx_u_din_buffer_data_reg_6__19__1006 (.o(net1006));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__20__u_dcfifo_tx_u_din_buffer_data_reg_6__21__1007 (.o(net1007));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__20__u_dcfifo_tx_u_din_buffer_data_reg_6__21__1008 (.o(net1008));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__22__u_dcfifo_tx_u_din_buffer_data_reg_6__23__1009 (.o(net1009));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__22__u_dcfifo_tx_u_din_buffer_data_reg_6__23__1010 (.o(net1010));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__24__u_dcfifo_tx_u_din_buffer_data_reg_6__25__1011 (.o(net1011));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__24__u_dcfifo_tx_u_din_buffer_data_reg_6__25__1012 (.o(net1012));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__26__u_dcfifo_tx_u_din_buffer_data_reg_6__27__1013 (.o(net1013));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__26__u_dcfifo_tx_u_din_buffer_data_reg_6__27__1014 (.o(net1014));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__28__u_dcfifo_tx_u_din_buffer_data_reg_6__29__1015 (.o(net1015));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__28__u_dcfifo_tx_u_din_buffer_data_reg_6__29__1016 (.o(net1016));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__2__u_dcfifo_tx_u_din_buffer_data_reg_6__3__1017 (.o(net1017));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__2__u_dcfifo_tx_u_din_buffer_data_reg_6__3__1018 (.o(net1018));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__30__u_dcfifo_tx_u_din_buffer_data_reg_6__31__1019 (.o(net1019));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__30__u_dcfifo_tx_u_din_buffer_data_reg_6__31__1020 (.o(net1020));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__4__u_dcfifo_tx_u_din_buffer_data_reg_6__5__1021 (.o(net1021));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__4__u_dcfifo_tx_u_din_buffer_data_reg_6__5__1022 (.o(net1022));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__6__u_dcfifo_tx_u_din_buffer_data_reg_6__7__1023 (.o(net1023));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__6__u_dcfifo_tx_u_din_buffer_data_reg_6__7__1024 (.o(net1024));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__8__u_dcfifo_tx_u_din_buffer_data_reg_6__9__1025 (.o(net1025));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__8__u_dcfifo_tx_u_din_buffer_data_reg_6__9__1026 (.o(net1026));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__0__u_dcfifo_tx_u_din_buffer_data_reg_7__1__1027 (.o(net1027));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__0__u_dcfifo_tx_u_din_buffer_data_reg_7__1__1028 (.o(net1028));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__10__u_dcfifo_tx_u_din_buffer_data_reg_7__11__1029 (.o(net1029));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__10__u_dcfifo_tx_u_din_buffer_data_reg_7__11__1030 (.o(net1030));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__12__u_dcfifo_tx_u_din_buffer_data_reg_7__13__1031 (.o(net1031));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__12__u_dcfifo_tx_u_din_buffer_data_reg_7__13__1032 (.o(net1032));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__14__u_dcfifo_tx_u_din_buffer_data_reg_7__15__1033 (.o(net1033));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__14__u_dcfifo_tx_u_din_buffer_data_reg_7__15__1034 (.o(net1034));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__16__u_dcfifo_tx_u_din_buffer_data_reg_7__17__1035 (.o(net1035));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__16__u_dcfifo_tx_u_din_buffer_data_reg_7__17__1036 (.o(net1036));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__18__u_dcfifo_tx_u_din_buffer_data_reg_7__19__1037 (.o(net1037));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__18__u_dcfifo_tx_u_din_buffer_data_reg_7__19__1038 (.o(net1038));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__20__u_dcfifo_tx_u_din_buffer_data_reg_7__21__1039 (.o(net1039));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__20__u_dcfifo_tx_u_din_buffer_data_reg_7__21__1040 (.o(net1040));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__22__u_dcfifo_tx_u_din_buffer_data_reg_7__23__1041 (.o(net1041));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__22__u_dcfifo_tx_u_din_buffer_data_reg_7__23__1042 (.o(net1042));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__24__u_dcfifo_tx_u_din_buffer_data_reg_7__25__1043 (.o(net1043));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__24__u_dcfifo_tx_u_din_buffer_data_reg_7__25__1044 (.o(net1044));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__26__u_dcfifo_tx_u_din_buffer_data_reg_7__27__1045 (.o(net1045));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__26__u_dcfifo_tx_u_din_buffer_data_reg_7__27__1046 (.o(net1046));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__28__u_dcfifo_tx_u_din_buffer_data_reg_7__29__1047 (.o(net1047));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__28__u_dcfifo_tx_u_din_buffer_data_reg_7__29__1048 (.o(net1048));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__2__u_dcfifo_tx_u_din_buffer_data_reg_7__3__1049 (.o(net1049));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__2__u_dcfifo_tx_u_din_buffer_data_reg_7__3__1050 (.o(net1050));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__30__u_dcfifo_tx_u_din_buffer_data_reg_7__31__1051 (.o(net1051));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__30__u_dcfifo_tx_u_din_buffer_data_reg_7__31__1052 (.o(net1052));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__4__u_dcfifo_tx_u_din_buffer_data_reg_7__5__1053 (.o(net1053));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__4__u_dcfifo_tx_u_din_buffer_data_reg_7__5__1054 (.o(net1054));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__6__u_dcfifo_tx_u_din_buffer_data_reg_7__7__1055 (.o(net1055));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__6__u_dcfifo_tx_u_din_buffer_data_reg_7__7__1056 (.o(net1056));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__8__u_dcfifo_tx_u_din_buffer_data_reg_7__9__1057 (.o(net1057));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__8__u_dcfifo_tx_u_din_buffer_data_reg_7__9__1058 (.o(net1058));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_full_full_synch_d_middle_reg_0__u_dcfifo_tx_u_din_full_full_synch_d_out_reg_0__1059 (.o(net1059));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_full_full_synch_d_middle_reg_0__u_dcfifo_tx_u_din_full_full_synch_d_out_reg_0__1060 (.o(net1060));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_full_latched_full_s_reg_u_spi_device_tlul_plug_state_reg_0__1061 (.o(net1061));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_full_latched_full_s_reg_u_spi_device_tlul_plug_state_reg_0__1062 (.o(net1062));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_write_tr_clk_gate_state_reg_latch_1063 (.o(net1063));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_write_tr_state_reg_0__u_dcfifo_tx_u_din_write_tr_state_reg_1__1064 (.o(net1064));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_write_tr_state_reg_0__u_dcfifo_tx_u_din_write_tr_state_reg_1__1065 (.o(net1065));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_write_tr_state_reg_2__1066 (.o(net1066));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_write_tr_state_reg_3__1067 (.o(net1067));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_write_tr_state_reg_4__u_dcfifo_tx_u_din_write_tr_state_reg_5__1068 (.o(net1068));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_write_tr_state_reg_4__u_dcfifo_tx_u_din_write_tr_state_reg_5__1069 (.o(net1069));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_write_tr_state_reg_6__u_dcfifo_tx_u_din_write_tr_state_reg_7__1070 (.o(net1070));
 b15tilo00an1n03x5 u_dcfifo_tx_u_din_write_tr_state_reg_6__u_dcfifo_tx_u_din_write_tr_state_reg_7__1071 (.o(net1071));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_0__u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_1__1072 (.o(net1072));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_0__u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_1__1073 (.o(net1073));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_2__1074 (.o(net1074));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_3__1075 (.o(net1075));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_4__u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_5__1076 (.o(net1076));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_4__u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_5__1077 (.o(net1077));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_6__u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_7__1078 (.o(net1078));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_6__u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_7__1079 (.o(net1079));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_0__u_dcfifo_tx_u_dout_empty_synch_d_out_reg_5__1080 (.o(net1080));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_0__u_dcfifo_tx_u_dout_empty_synch_d_out_reg_5__1081 (.o(net1081));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_2__1082 (.o(net1082));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_3__1083 (.o(net1083));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_4__1084 (.o(net1084));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_6__u_dcfifo_tx_u_dout_empty_synch_d_out_reg_7__1085 (.o(net1085));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_6__u_dcfifo_tx_u_dout_empty_synch_d_out_reg_7__1086 (.o(net1086));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_read_tr_clk_gate_state_reg_latch_1087 (.o(net1087));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_read_tr_state_reg_0__1088 (.o(net1088));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_read_tr_state_reg_1__1089 (.o(net1089));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_read_tr_state_reg_2__u_dcfifo_tx_u_dout_read_tr_state_reg_3__1090 (.o(net1090));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_read_tr_state_reg_2__u_dcfifo_tx_u_dout_read_tr_state_reg_3__1091 (.o(net1091));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_read_tr_state_reg_4__u_dcfifo_tx_u_dout_read_tr_state_reg_5__1092 (.o(net1092));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_read_tr_state_reg_4__u_dcfifo_tx_u_dout_read_tr_state_reg_5__1093 (.o(net1093));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_read_tr_state_reg_6__u_dcfifo_tx_u_dout_read_tr_state_reg_7__1094 (.o(net1094));
 b15tilo00an1n03x5 u_dcfifo_tx_u_dout_read_tr_state_reg_6__u_dcfifo_tx_u_dout_read_tr_state_reg_7__1095 (.o(net1095));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_0__u_device_sm_addr_reg_reg_1__1096 (.o(net1096));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_0__u_device_sm_addr_reg_reg_1__1097 (.o(net1097));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_10__u_device_sm_addr_reg_reg_11__1098 (.o(net1098));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_10__u_device_sm_addr_reg_reg_11__1099 (.o(net1099));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_12__u_device_sm_addr_reg_reg_13__1100 (.o(net1100));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_12__u_device_sm_addr_reg_reg_13__1101 (.o(net1101));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_14__u_device_sm_addr_reg_reg_15__1102 (.o(net1102));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_14__u_device_sm_addr_reg_reg_15__1103 (.o(net1103));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_16__u_device_sm_addr_reg_reg_17__1104 (.o(net1104));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_16__u_device_sm_addr_reg_reg_17__1105 (.o(net1105));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_18__u_device_sm_addr_reg_reg_19__1106 (.o(net1106));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_18__u_device_sm_addr_reg_reg_19__1107 (.o(net1107));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_20__u_device_sm_addr_reg_reg_21__1108 (.o(net1108));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_20__u_device_sm_addr_reg_reg_21__1109 (.o(net1109));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_22__u_device_sm_addr_reg_reg_23__1110 (.o(net1110));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_22__u_device_sm_addr_reg_reg_23__1111 (.o(net1111));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_24__u_device_sm_addr_reg_reg_25__1112 (.o(net1112));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_24__u_device_sm_addr_reg_reg_25__1113 (.o(net1113));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_26__u_device_sm_addr_reg_reg_27__1114 (.o(net1114));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_26__u_device_sm_addr_reg_reg_27__1115 (.o(net1115));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_28__u_device_sm_addr_reg_reg_29__1116 (.o(net1116));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_28__u_device_sm_addr_reg_reg_29__1117 (.o(net1117));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_2__u_device_sm_addr_reg_reg_3__1118 (.o(net1118));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_2__u_device_sm_addr_reg_reg_3__1119 (.o(net1119));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_30__u_device_sm_addr_reg_reg_31__1120 (.o(net1120));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_30__u_device_sm_addr_reg_reg_31__1121 (.o(net1121));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_4__u_device_sm_addr_reg_reg_5__1122 (.o(net1122));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_4__u_device_sm_addr_reg_reg_5__1123 (.o(net1123));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_6__u_device_sm_addr_reg_reg_7__1124 (.o(net1124));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_6__u_device_sm_addr_reg_reg_7__1125 (.o(net1125));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_8__u_device_sm_addr_reg_reg_9__1126 (.o(net1126));
 b15tilo00an1n03x5 u_device_sm_addr_reg_reg_8__u_device_sm_addr_reg_reg_9__1127 (.o(net1127));
 b15tilo00an1n03x5 u_device_sm_clk_gate_addr_reg_reg_0_latch_1128 (.o(net1128));
 b15tilo00an1n03x5 u_device_sm_clk_gate_addr_reg_reg_latch_1129 (.o(net1129));
 b15tilo00an1n03x5 u_device_sm_clk_gate_cmd_reg_reg_latch_1130 (.o(net1130));
 b15tilo00an1n03x5 u_device_sm_cmd_reg_reg_0__u_device_sm_cmd_reg_reg_1__1131 (.o(net1131));
 b15tilo00an1n03x5 u_device_sm_cmd_reg_reg_0__u_device_sm_cmd_reg_reg_1__1132 (.o(net1132));
 b15tilo00an1n03x5 u_device_sm_cmd_reg_reg_2__u_device_sm_cmd_reg_reg_3__1133 (.o(net1133));
 b15tilo00an1n03x5 u_device_sm_cmd_reg_reg_2__u_device_sm_cmd_reg_reg_3__1134 (.o(net1134));
 b15tilo00an1n03x5 u_device_sm_cmd_reg_reg_4__u_device_sm_cmd_reg_reg_5__1135 (.o(net1135));
 b15tilo00an1n03x5 u_device_sm_cmd_reg_reg_4__u_device_sm_cmd_reg_reg_5__1136 (.o(net1136));
 b15tilo00an1n03x5 u_device_sm_cmd_reg_reg_6__u_device_sm_cmd_reg_reg_7__1137 (.o(net1137));
 b15tilo00an1n03x5 u_device_sm_cmd_reg_reg_6__u_device_sm_cmd_reg_reg_7__1138 (.o(net1138));
 b15tilo00an1n03x5 u_device_sm_ctrl_addr_valid_reg_u_device_sm_data_reg_reg_0__1139 (.o(net1139));
 b15tilo00an1n03x5 u_device_sm_ctrl_addr_valid_reg_u_device_sm_data_reg_reg_0__1140 (.o(net1140));
 b15tilo00an1n03x5 u_device_sm_ctrl_data_tx_ready_reg_u_device_sm_state_reg_1__1141 (.o(net1141));
 b15tilo00an1n03x5 u_device_sm_ctrl_data_tx_ready_reg_u_device_sm_state_reg_1__1142 (.o(net1142));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_10__u_device_sm_data_reg_reg_11__1143 (.o(net1143));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_10__u_device_sm_data_reg_reg_11__1144 (.o(net1144));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_12__u_device_sm_data_reg_reg_13__1145 (.o(net1145));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_12__u_device_sm_data_reg_reg_13__1146 (.o(net1146));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_14__u_device_sm_data_reg_reg_15__1147 (.o(net1147));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_14__u_device_sm_data_reg_reg_15__1148 (.o(net1148));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_16__u_device_sm_data_reg_reg_17__1149 (.o(net1149));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_16__u_device_sm_data_reg_reg_17__1150 (.o(net1150));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_18__u_device_sm_data_reg_reg_19__1151 (.o(net1151));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_18__u_device_sm_data_reg_reg_19__1152 (.o(net1152));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_1__u_device_sm_data_reg_reg_2__1153 (.o(net1153));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_1__u_device_sm_data_reg_reg_2__1154 (.o(net1154));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_20__u_device_sm_data_reg_reg_21__1155 (.o(net1155));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_20__u_device_sm_data_reg_reg_21__1156 (.o(net1156));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_22__u_device_sm_data_reg_reg_23__1157 (.o(net1157));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_22__u_device_sm_data_reg_reg_23__1158 (.o(net1158));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_24__u_device_sm_data_reg_reg_25__1159 (.o(net1159));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_24__u_device_sm_data_reg_reg_25__1160 (.o(net1160));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_26__u_device_sm_data_reg_reg_27__1161 (.o(net1161));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_26__u_device_sm_data_reg_reg_27__1162 (.o(net1162));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_28__u_device_sm_data_reg_reg_29__1163 (.o(net1163));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_28__u_device_sm_data_reg_reg_29__1164 (.o(net1164));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_30__u_device_sm_data_reg_reg_31__1165 (.o(net1165));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_30__u_device_sm_data_reg_reg_31__1166 (.o(net1166));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_3__u_device_sm_data_reg_reg_4__1167 (.o(net1167));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_3__u_device_sm_data_reg_reg_4__1168 (.o(net1168));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_5__u_device_sm_state_reg_0__1169 (.o(net1169));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_5__u_device_sm_state_reg_0__1170 (.o(net1170));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_6__u_device_sm_data_reg_reg_7__1171 (.o(net1171));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_6__u_device_sm_data_reg_reg_7__1172 (.o(net1172));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_8__u_device_sm_data_reg_reg_9__1173 (.o(net1173));
 b15tilo00an1n03x5 u_device_sm_data_reg_reg_8__u_device_sm_data_reg_reg_9__1174 (.o(net1174));
 b15tilo00an1n03x5 u_device_sm_mode_reg_reg_0__u_device_sm_mode_reg_reg_1__1175 (.o(net1175));
 b15tilo00an1n03x5 u_device_sm_mode_reg_reg_0__u_device_sm_mode_reg_reg_1__1176 (.o(net1176));
 b15tilo00an1n03x5 u_device_sm_mode_reg_reg_2__u_device_sm_mode_reg_reg_3__1177 (.o(net1177));
 b15tilo00an1n03x5 u_device_sm_mode_reg_reg_2__u_device_sm_mode_reg_reg_3__1178 (.o(net1178));
 b15tilo00an1n03x5 u_device_sm_mode_reg_reg_4__u_device_sm_mode_reg_reg_5__1179 (.o(net1179));
 b15tilo00an1n03x5 u_device_sm_mode_reg_reg_4__u_device_sm_mode_reg_reg_5__1180 (.o(net1180));
 b15tilo00an1n03x5 u_device_sm_mode_reg_reg_6__u_device_sm_mode_reg_reg_7__1181 (.o(net1181));
 b15tilo00an1n03x5 u_device_sm_mode_reg_reg_6__u_device_sm_mode_reg_reg_7__1182 (.o(net1182));
 b15tilo00an1n03x5 u_device_sm_pad_mode_next_reg_1__1183 (.o(net1183));
 b15tilo00an1n03x5 u_device_sm_state_reg_2__u_device_sm_tx_counter_reg_0__1184 (.o(net1184));
 b15tilo00an1n03x5 u_device_sm_state_reg_2__u_device_sm_tx_counter_reg_0__1185 (.o(net1185));
 b15tilo00an1n03x5 u_device_sm_tx_counter_reg_1__u_device_sm_tx_data_reg_0__1186 (.o(net1186));
 b15tilo00an1n03x5 u_device_sm_tx_counter_reg_1__u_device_sm_tx_data_reg_0__1187 (.o(net1187));
 b15tilo00an1n03x5 u_device_sm_tx_counter_reg_2__u_device_sm_tx_counter_reg_3__1188 (.o(net1188));
 b15tilo00an1n03x5 u_device_sm_tx_counter_reg_2__u_device_sm_tx_counter_reg_3__1189 (.o(net1189));
 b15tilo00an1n03x5 u_device_sm_tx_counter_reg_4__u_device_sm_tx_counter_upd_reg_1190 (.o(net1190));
 b15tilo00an1n03x5 u_device_sm_tx_counter_reg_4__u_device_sm_tx_counter_upd_reg_1191 (.o(net1191));
 b15tilo00an1n03x5 u_device_sm_tx_counter_reg_5__u_device_sm_tx_counter_reg_6__1192 (.o(net1192));
 b15tilo00an1n03x5 u_device_sm_tx_counter_reg_5__u_device_sm_tx_counter_reg_6__1193 (.o(net1193));
 b15tilo00an1n03x5 u_device_sm_tx_counter_reg_5__u_device_sm_tx_counter_reg_6__1194 (.o(net1194));
 b15tilo00an1n03x5 u_device_sm_tx_counter_reg_5__u_device_sm_tx_counter_reg_6__1195 (.o(net1195));
 b15tilo00an1n03x5 u_device_sm_tx_counter_reg_7__1196 (.o(net1196));
 b15tilo00an1n03x5 u_device_sm_tx_counter_reg_7__1197 (.o(net1197));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_11__u_device_sm_tx_data_reg_12__1198 (.o(net1198));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_11__u_device_sm_tx_data_reg_12__1199 (.o(net1199));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_13__u_device_sm_tx_data_reg_14__1200 (.o(net1200));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_13__u_device_sm_tx_data_reg_14__1201 (.o(net1201));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_15__1202 (.o(net1202));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_16__u_device_sm_tx_data_reg_17__1203 (.o(net1203));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_16__u_device_sm_tx_data_reg_17__1204 (.o(net1204));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_18__u_device_sm_tx_data_reg_19__1205 (.o(net1205));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_18__u_device_sm_tx_data_reg_19__1206 (.o(net1206));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_1__u_device_sm_tx_data_reg_2__1207 (.o(net1207));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_1__u_device_sm_tx_data_reg_2__1208 (.o(net1208));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_20__u_device_sm_tx_data_reg_21__1209 (.o(net1209));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_20__u_device_sm_tx_data_reg_21__1210 (.o(net1210));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_22__u_device_sm_tx_data_reg_23__1211 (.o(net1211));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_22__u_device_sm_tx_data_reg_23__1212 (.o(net1212));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_24__u_device_sm_tx_data_reg_25__1213 (.o(net1213));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_24__u_device_sm_tx_data_reg_25__1214 (.o(net1214));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_26__u_device_sm_tx_data_reg_27__1215 (.o(net1215));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_26__u_device_sm_tx_data_reg_27__1216 (.o(net1216));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_28__u_device_sm_tx_data_reg_29__1217 (.o(net1217));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_28__u_device_sm_tx_data_reg_29__1218 (.o(net1218));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_30__u_device_sm_tx_data_reg_31__1219 (.o(net1219));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_30__u_device_sm_tx_data_reg_31__1220 (.o(net1220));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_3__u_device_sm_tx_data_reg_4__1221 (.o(net1221));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_3__u_device_sm_tx_data_reg_4__1222 (.o(net1222));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_5__u_device_sm_tx_data_reg_6__1223 (.o(net1223));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_5__u_device_sm_tx_data_reg_6__1224 (.o(net1224));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_7__u_device_sm_tx_data_reg_8__1225 (.o(net1225));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_7__u_device_sm_tx_data_reg_8__1226 (.o(net1226));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_9__u_device_sm_tx_data_reg_10__1227 (.o(net1227));
 b15tilo00an1n03x5 u_device_sm_tx_data_reg_9__u_device_sm_tx_data_reg_10__1228 (.o(net1228));
 b15tilo00an1n03x5 u_device_sm_tx_data_valid_reg_u_device_sm_tx_done_reg_reg_1229 (.o(net1229));
 b15tilo00an1n03x5 u_device_sm_tx_data_valid_reg_u_device_sm_tx_done_reg_reg_1230 (.o(net1230));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_clk_gate_reg0_reg_latch_1231 (.o(net1231));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_clk_gate_reg1_reg_latch_1232 (.o(net1232));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_clk_gate_reg2_reg_latch_1233 (.o(net1233));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_clk_gate_reg3_reg_latch_1234 (.o(net1234));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg0_reg_0__u_device_sm_u_spiregs_reg0_reg_1__1235 (.o(net1235));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg0_reg_0__u_device_sm_u_spiregs_reg0_reg_1__1236 (.o(net1236));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg0_reg_2__u_device_sm_u_spiregs_reg0_reg_3__1237 (.o(net1237));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg0_reg_2__u_device_sm_u_spiregs_reg0_reg_3__1238 (.o(net1238));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg0_reg_4__u_device_sm_u_spiregs_reg0_reg_5__1239 (.o(net1239));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg0_reg_4__u_device_sm_u_spiregs_reg0_reg_5__1240 (.o(net1240));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg0_reg_6__u_device_sm_u_spiregs_reg0_reg_7__1241 (.o(net1241));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg0_reg_6__u_device_sm_u_spiregs_reg0_reg_7__1242 (.o(net1242));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg1_reg_0__u_device_sm_u_spiregs_reg1_reg_1__1243 (.o(net1243));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg1_reg_0__u_device_sm_u_spiregs_reg1_reg_1__1244 (.o(net1244));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg1_reg_2__u_device_sm_u_spiregs_reg1_reg_3__1245 (.o(net1245));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg1_reg_2__u_device_sm_u_spiregs_reg1_reg_3__1246 (.o(net1246));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg1_reg_4__u_device_sm_u_spiregs_reg1_reg_6__1247 (.o(net1247));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg1_reg_4__u_device_sm_u_spiregs_reg1_reg_6__1248 (.o(net1248));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg1_reg_5__1249 (.o(net1249));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg1_reg_7__1250 (.o(net1250));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg2_reg_0__u_device_sm_u_spiregs_reg2_reg_1__1251 (.o(net1251));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg2_reg_0__u_device_sm_u_spiregs_reg2_reg_1__1252 (.o(net1252));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg2_reg_2__u_device_sm_u_spiregs_reg2_reg_3__1253 (.o(net1253));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg2_reg_2__u_device_sm_u_spiregs_reg2_reg_3__1254 (.o(net1254));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg2_reg_4__u_device_sm_u_spiregs_reg2_reg_5__1255 (.o(net1255));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg2_reg_4__u_device_sm_u_spiregs_reg2_reg_5__1256 (.o(net1256));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg2_reg_6__u_device_sm_u_spiregs_reg2_reg_7__1257 (.o(net1257));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg2_reg_6__u_device_sm_u_spiregs_reg2_reg_7__1258 (.o(net1258));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg3_reg_0__u_device_sm_u_spiregs_reg3_reg_1__1259 (.o(net1259));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg3_reg_0__u_device_sm_u_spiregs_reg3_reg_1__1260 (.o(net1260));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg3_reg_2__u_device_sm_u_spiregs_reg3_reg_3__1261 (.o(net1261));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg3_reg_2__u_device_sm_u_spiregs_reg3_reg_3__1262 (.o(net1262));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg3_reg_4__u_device_sm_u_spiregs_reg3_reg_5__1263 (.o(net1263));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg3_reg_4__u_device_sm_u_spiregs_reg3_reg_5__1264 (.o(net1264));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg3_reg_6__u_device_sm_u_spiregs_reg3_reg_7__1265 (.o(net1265));
 b15tilo00an1n03x5 u_device_sm_u_spiregs_reg3_reg_6__u_device_sm_u_spiregs_reg3_reg_7__1266 (.o(net1266));
 b15tilo00an1n03x5 u_rxreg_clk_gate_counter_reg_latch_1267 (.o(net1267));
 b15tilo00an1n03x5 u_rxreg_clk_gate_counter_trgt_reg_latch_1268 (.o(net1268));
 b15tilo00an1n03x5 u_rxreg_clk_gate_data_int_reg_0_latch_1269 (.o(net1269));
 b15tilo00an1n03x5 u_rxreg_clk_gate_data_int_reg_latch_1270 (.o(net1270));
 b15tilo00an1n03x5 u_rxreg_counter_reg_0__u_rxreg_counter_reg_1__1271 (.o(net1271));
 b15tilo00an1n03x5 u_rxreg_counter_reg_0__u_rxreg_counter_reg_1__1272 (.o(net1272));
 b15tilo00an1n03x5 u_rxreg_counter_reg_2__u_rxreg_counter_reg_3__1273 (.o(net1273));
 b15tilo00an1n03x5 u_rxreg_counter_reg_2__u_rxreg_counter_reg_3__1274 (.o(net1274));
 b15tilo00an1n03x5 u_rxreg_counter_reg_4__u_rxreg_counter_reg_5__1275 (.o(net1275));
 b15tilo00an1n03x5 u_rxreg_counter_reg_4__u_rxreg_counter_reg_5__1276 (.o(net1276));
 b15tilo00an1n03x5 u_rxreg_counter_reg_6__u_rxreg_counter_reg_7__1277 (.o(net1277));
 b15tilo00an1n03x5 u_rxreg_counter_reg_6__u_rxreg_counter_reg_7__1278 (.o(net1278));
 b15tilo00an1n03x5 u_rxreg_counter_trgt_reg_0__1279 (.o(net1279));
 b15tilo00an1n03x5 u_rxreg_counter_trgt_reg_1__u_rxreg_counter_trgt_reg_2__1280 (.o(net1280));
 b15tilo00an1n03x5 u_rxreg_counter_trgt_reg_1__u_rxreg_counter_trgt_reg_2__1281 (.o(net1281));
 b15tilo00an1n03x5 u_rxreg_counter_trgt_reg_3__u_rxreg_counter_trgt_reg_4__1282 (.o(net1282));
 b15tilo00an1n03x5 u_rxreg_counter_trgt_reg_3__u_rxreg_counter_trgt_reg_4__1283 (.o(net1283));
 b15tilo00an1n03x5 u_rxreg_counter_trgt_reg_5__u_rxreg_counter_trgt_reg_6__1284 (.o(net1284));
 b15tilo00an1n03x5 u_rxreg_counter_trgt_reg_5__u_rxreg_counter_trgt_reg_6__1285 (.o(net1285));
 b15tilo00an1n03x5 u_rxreg_counter_trgt_reg_7__1286 (.o(net1286));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_0__u_rxreg_data_int_reg_1__1287 (.o(net1287));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_0__u_rxreg_data_int_reg_1__1288 (.o(net1288));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_10__u_rxreg_data_int_reg_11__1289 (.o(net1289));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_10__u_rxreg_data_int_reg_11__1290 (.o(net1290));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_12__u_rxreg_data_int_reg_13__1291 (.o(net1291));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_12__u_rxreg_data_int_reg_13__1292 (.o(net1292));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_14__u_rxreg_data_int_reg_15__1293 (.o(net1293));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_14__u_rxreg_data_int_reg_15__1294 (.o(net1294));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_16__u_rxreg_data_int_reg_17__1295 (.o(net1295));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_16__u_rxreg_data_int_reg_17__1296 (.o(net1296));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_18__u_rxreg_data_int_reg_19__1297 (.o(net1297));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_18__u_rxreg_data_int_reg_19__1298 (.o(net1298));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_20__u_rxreg_data_int_reg_21__1299 (.o(net1299));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_20__u_rxreg_data_int_reg_21__1300 (.o(net1300));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_22__u_rxreg_data_int_reg_23__1301 (.o(net1301));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_22__u_rxreg_data_int_reg_23__1302 (.o(net1302));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_24__u_rxreg_data_int_reg_25__1303 (.o(net1303));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_24__u_rxreg_data_int_reg_25__1304 (.o(net1304));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_26__u_rxreg_data_int_reg_27__1305 (.o(net1305));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_26__u_rxreg_data_int_reg_27__1306 (.o(net1306));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_28__u_rxreg_data_int_reg_29__1307 (.o(net1307));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_28__u_rxreg_data_int_reg_29__1308 (.o(net1308));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_2__u_rxreg_data_int_reg_3__1309 (.o(net1309));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_2__u_rxreg_data_int_reg_3__1310 (.o(net1310));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_30__u_rxreg_data_int_reg_31__1311 (.o(net1311));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_30__u_rxreg_data_int_reg_31__1312 (.o(net1312));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_4__u_rxreg_data_int_reg_5__1313 (.o(net1313));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_4__u_rxreg_data_int_reg_5__1314 (.o(net1314));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_6__u_rxreg_data_int_reg_7__1315 (.o(net1315));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_6__u_rxreg_data_int_reg_7__1316 (.o(net1316));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_8__u_rxreg_data_int_reg_9__1317 (.o(net1317));
 b15tilo00an1n03x5 u_rxreg_data_int_reg_8__u_rxreg_data_int_reg_9__1318 (.o(net1318));
 b15tilo00an1n03x5 u_rxreg_running_reg_1319 (.o(net1319));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_0__u_spi_device_tlul_plug_addr_reg_1__1320 (.o(net1320));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_0__u_spi_device_tlul_plug_addr_reg_1__1321 (.o(net1321));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_10__u_spi_device_tlul_plug_addr_reg_11__1322 (.o(net1322));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_10__u_spi_device_tlul_plug_addr_reg_11__1323 (.o(net1323));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_12__u_spi_device_tlul_plug_addr_reg_13__1324 (.o(net1324));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_12__u_spi_device_tlul_plug_addr_reg_13__1325 (.o(net1325));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_14__u_spi_device_tlul_plug_addr_reg_15__1326 (.o(net1326));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_14__u_spi_device_tlul_plug_addr_reg_15__1327 (.o(net1327));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_16__u_spi_device_tlul_plug_addr_reg_17__1328 (.o(net1328));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_16__u_spi_device_tlul_plug_addr_reg_17__1329 (.o(net1329));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_18__u_spi_device_tlul_plug_addr_reg_19__1330 (.o(net1330));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_18__u_spi_device_tlul_plug_addr_reg_19__1331 (.o(net1331));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_20__u_spi_device_tlul_plug_addr_reg_21__1332 (.o(net1332));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_20__u_spi_device_tlul_plug_addr_reg_21__1333 (.o(net1333));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_22__u_spi_device_tlul_plug_addr_reg_23__1334 (.o(net1334));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_22__u_spi_device_tlul_plug_addr_reg_23__1335 (.o(net1335));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_24__u_spi_device_tlul_plug_addr_reg_25__1336 (.o(net1336));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_24__u_spi_device_tlul_plug_addr_reg_25__1337 (.o(net1337));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_26__u_spi_device_tlul_plug_addr_reg_27__1338 (.o(net1338));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_26__u_spi_device_tlul_plug_addr_reg_27__1339 (.o(net1339));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_28__u_spi_device_tlul_plug_addr_reg_29__1340 (.o(net1340));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_28__u_spi_device_tlul_plug_addr_reg_29__1341 (.o(net1341));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_2__u_spi_device_tlul_plug_addr_reg_3__1342 (.o(net1342));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_2__u_spi_device_tlul_plug_addr_reg_3__1343 (.o(net1343));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_30__u_spi_device_tlul_plug_addr_reg_31__1344 (.o(net1344));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_30__u_spi_device_tlul_plug_addr_reg_31__1345 (.o(net1345));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_4__u_spi_device_tlul_plug_addr_reg_5__1346 (.o(net1346));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_4__u_spi_device_tlul_plug_addr_reg_5__1347 (.o(net1347));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_6__u_spi_device_tlul_plug_addr_reg_7__1348 (.o(net1348));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_6__u_spi_device_tlul_plug_addr_reg_7__1349 (.o(net1349));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_8__u_spi_device_tlul_plug_addr_reg_9__1350 (.o(net1350));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_addr_reg_8__u_spi_device_tlul_plug_addr_reg_9__1351 (.o(net1351));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_clk_gate_addr_reg_0_latch_1352 (.o(net1352));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_clk_gate_addr_reg_latch_1353 (.o(net1353));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_state_reg_1__u_spi_device_tlul_plug_u_tlul_adapter_host_g_multiple_reqs_source_q_reg_0__1354 (.o(net1354));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_state_reg_1__u_spi_device_tlul_plug_u_tlul_adapter_host_g_multiple_reqs_source_q_reg_0__1355 (.o(net1355));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_u_tlul_adapter_host_intg_err_q_reg_u_spi_device_tlul_plug_wdata_reg_0__1356 (.o(net1356));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_u_tlul_adapter_host_intg_err_q_reg_u_spi_device_tlul_plug_wdata_reg_0__1357 (.o(net1357));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_11__u_spi_device_tlul_plug_wdata_reg_12__1358 (.o(net1358));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_11__u_spi_device_tlul_plug_wdata_reg_12__1359 (.o(net1359));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_13__u_spi_device_tlul_plug_wdata_reg_14__1360 (.o(net1360));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_13__u_spi_device_tlul_plug_wdata_reg_14__1361 (.o(net1361));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_15__u_spi_device_tlul_plug_wdata_reg_16__1362 (.o(net1362));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_15__u_spi_device_tlul_plug_wdata_reg_16__1363 (.o(net1363));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_17__u_spi_device_tlul_plug_wdata_reg_18__1364 (.o(net1364));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_17__u_spi_device_tlul_plug_wdata_reg_18__1365 (.o(net1365));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_19__u_spi_device_tlul_plug_wdata_reg_20__1366 (.o(net1366));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_19__u_spi_device_tlul_plug_wdata_reg_20__1367 (.o(net1367));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_1__u_spi_device_tlul_plug_wdata_reg_2__1368 (.o(net1368));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_1__u_spi_device_tlul_plug_wdata_reg_2__1369 (.o(net1369));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_21__u_spi_device_tlul_plug_wdata_reg_22__1370 (.o(net1370));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_21__u_spi_device_tlul_plug_wdata_reg_22__1371 (.o(net1371));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_23__u_spi_device_tlul_plug_wdata_reg_24__1372 (.o(net1372));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_23__u_spi_device_tlul_plug_wdata_reg_24__1373 (.o(net1373));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_25__u_spi_device_tlul_plug_wdata_reg_26__1374 (.o(net1374));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_25__u_spi_device_tlul_plug_wdata_reg_26__1375 (.o(net1375));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_27__u_spi_device_tlul_plug_wdata_reg_28__1376 (.o(net1376));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_27__u_spi_device_tlul_plug_wdata_reg_28__1377 (.o(net1377));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_29__u_spi_device_tlul_plug_wdata_reg_30__1378 (.o(net1378));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_29__u_spi_device_tlul_plug_wdata_reg_30__1379 (.o(net1379));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_31__u_spi_device_tlul_plug_we_reg_1380 (.o(net1380));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_31__u_spi_device_tlul_plug_we_reg_1381 (.o(net1381));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_3__u_spi_device_tlul_plug_wdata_reg_4__1382 (.o(net1382));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_3__u_spi_device_tlul_plug_wdata_reg_4__1383 (.o(net1383));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_5__u_spi_device_tlul_plug_wdata_reg_6__1384 (.o(net1384));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_5__u_spi_device_tlul_plug_wdata_reg_6__1385 (.o(net1385));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_7__u_spi_device_tlul_plug_wdata_reg_8__1386 (.o(net1386));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_7__u_spi_device_tlul_plug_wdata_reg_8__1387 (.o(net1387));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_9__u_spi_device_tlul_plug_wdata_reg_10__1388 (.o(net1388));
 b15tilo00an1n03x5 u_spi_device_tlul_plug_wdata_reg_9__u_spi_device_tlul_plug_wdata_reg_10__1389 (.o(net1389));
 b15tilo00an1n03x5 u_syncro_cs_reg_reg_0__1390 (.o(net1390));
 b15tilo00an1n03x5 u_syncro_cs_reg_reg_1__1391 (.o(net1391));
 b15tilo00an1n03x5 u_syncro_rdwr_reg_reg_0__u_syncro_rdwr_reg_reg_1__1392 (.o(net1392));
 b15tilo00an1n03x5 u_syncro_rdwr_reg_reg_0__u_syncro_rdwr_reg_reg_1__1393 (.o(net1393));
 b15tilo00an1n03x5 u_syncro_valid_reg_reg_0__u_syncro_valid_reg_reg_1__1394 (.o(net1394));
 b15tilo00an1n03x5 u_syncro_valid_reg_reg_0__u_syncro_valid_reg_reg_1__1395 (.o(net1395));
 b15tilo00an1n03x5 u_syncro_valid_reg_reg_2__1396 (.o(net1396));
 b15tilo00an1n03x5 u_txreg_clk_gate_counter_reg_latch_1397 (.o(net1397));
 b15tilo00an1n03x5 u_txreg_clk_gate_counter_trgt_reg_latch_1398 (.o(net1398));
 b15tilo00an1n03x5 u_txreg_clk_gate_data_int_reg_0_latch_1399 (.o(net1399));
 b15tilo00an1n03x5 u_txreg_clk_gate_data_int_reg_latch_1400 (.o(net1400));
 b15tilo00an1n03x5 u_txreg_counter_reg_0__u_txreg_counter_reg_1__1401 (.o(net1401));
 b15tilo00an1n03x5 u_txreg_counter_reg_0__u_txreg_counter_reg_1__1402 (.o(net1402));
 b15tilo00an1n03x5 u_txreg_counter_reg_2__u_txreg_counter_reg_3__1403 (.o(net1403));
 b15tilo00an1n03x5 u_txreg_counter_reg_2__u_txreg_counter_reg_3__1404 (.o(net1404));
 b15tilo00an1n03x5 u_txreg_counter_reg_4__u_txreg_counter_reg_5__1405 (.o(net1405));
 b15tilo00an1n03x5 u_txreg_counter_reg_4__u_txreg_counter_reg_5__1406 (.o(net1406));
 b15tilo00an1n03x5 u_txreg_counter_reg_6__u_txreg_counter_reg_7__1407 (.o(net1407));
 b15tilo00an1n03x5 u_txreg_counter_reg_6__u_txreg_counter_reg_7__1408 (.o(net1408));
 b15tilo00an1n03x5 u_txreg_counter_trgt_reg_0__1409 (.o(net1409));
 b15tilo00an1n03x5 u_txreg_counter_trgt_reg_1__1410 (.o(net1410));
 b15tilo00an1n03x5 u_txreg_counter_trgt_reg_2__1411 (.o(net1411));
 b15tilo00an1n03x5 u_txreg_counter_trgt_reg_3__u_txreg_counter_trgt_reg_4__1412 (.o(net1412));
 b15tilo00an1n03x5 u_txreg_counter_trgt_reg_3__u_txreg_counter_trgt_reg_4__1413 (.o(net1413));
 b15tilo00an1n03x5 u_txreg_counter_trgt_reg_5__u_txreg_counter_trgt_reg_6__1414 (.o(net1414));
 b15tilo00an1n03x5 u_txreg_counter_trgt_reg_5__u_txreg_counter_trgt_reg_6__1415 (.o(net1415));
 b15tilo00an1n03x5 u_txreg_counter_trgt_reg_7__1416 (.o(net1416));
 b15tilo00an1n03x5 u_txreg_data_int_reg_0__u_txreg_data_int_reg_1__1417 (.o(net1417));
 b15tilo00an1n03x5 u_txreg_data_int_reg_0__u_txreg_data_int_reg_1__1418 (.o(net1418));
 b15tilo00an1n03x5 u_txreg_data_int_reg_10__u_txreg_data_int_reg_11__1419 (.o(net1419));
 b15tilo00an1n03x5 u_txreg_data_int_reg_10__u_txreg_data_int_reg_11__1420 (.o(net1420));
 b15tilo00an1n03x5 u_txreg_data_int_reg_12__u_txreg_data_int_reg_13__1421 (.o(net1421));
 b15tilo00an1n03x5 u_txreg_data_int_reg_12__u_txreg_data_int_reg_13__1422 (.o(net1422));
 b15tilo00an1n03x5 u_txreg_data_int_reg_14__u_txreg_data_int_reg_15__1423 (.o(net1423));
 b15tilo00an1n03x5 u_txreg_data_int_reg_14__u_txreg_data_int_reg_15__1424 (.o(net1424));
 b15tilo00an1n03x5 u_txreg_data_int_reg_16__u_txreg_data_int_reg_17__1425 (.o(net1425));
 b15tilo00an1n03x5 u_txreg_data_int_reg_16__u_txreg_data_int_reg_17__1426 (.o(net1426));
 b15tilo00an1n03x5 u_txreg_data_int_reg_18__u_txreg_data_int_reg_19__1427 (.o(net1427));
 b15tilo00an1n03x5 u_txreg_data_int_reg_18__u_txreg_data_int_reg_19__1428 (.o(net1428));
 b15tilo00an1n03x5 u_txreg_data_int_reg_20__u_txreg_data_int_reg_21__1429 (.o(net1429));
 b15tilo00an1n03x5 u_txreg_data_int_reg_20__u_txreg_data_int_reg_21__1430 (.o(net1430));
 b15tilo00an1n03x5 u_txreg_data_int_reg_22__u_txreg_data_int_reg_23__1431 (.o(net1431));
 b15tilo00an1n03x5 u_txreg_data_int_reg_22__u_txreg_data_int_reg_23__1432 (.o(net1432));
 b15tilo00an1n03x5 u_txreg_data_int_reg_24__u_txreg_data_int_reg_25__1433 (.o(net1433));
 b15tilo00an1n03x5 u_txreg_data_int_reg_24__u_txreg_data_int_reg_25__1434 (.o(net1434));
 b15tilo00an1n03x5 u_txreg_data_int_reg_26__u_txreg_data_int_reg_27__1435 (.o(net1435));
 b15tilo00an1n03x5 u_txreg_data_int_reg_26__u_txreg_data_int_reg_27__1436 (.o(net1436));
 b15tilo00an1n03x5 u_txreg_data_int_reg_28__u_txreg_data_int_reg_29__1437 (.o(net1437));
 b15tilo00an1n03x5 u_txreg_data_int_reg_28__u_txreg_data_int_reg_29__1438 (.o(net1438));
 b15tilo00an1n03x5 u_txreg_data_int_reg_2__u_txreg_data_int_reg_3__1439 (.o(net1439));
 b15tilo00an1n03x5 u_txreg_data_int_reg_2__u_txreg_data_int_reg_3__1440 (.o(net1440));
 b15tilo00an1n03x5 u_txreg_data_int_reg_30__u_txreg_data_int_reg_31__1441 (.o(net1441));
 b15tilo00an1n03x5 u_txreg_data_int_reg_30__u_txreg_data_int_reg_31__1442 (.o(net1442));
 b15tilo00an1n03x5 u_txreg_data_int_reg_4__u_txreg_data_int_reg_5__1443 (.o(net1443));
 b15tilo00an1n03x5 u_txreg_data_int_reg_4__u_txreg_data_int_reg_5__1444 (.o(net1444));
 b15tilo00an1n03x5 u_txreg_data_int_reg_6__u_txreg_data_int_reg_7__1445 (.o(net1445));
 b15tilo00an1n03x5 u_txreg_data_int_reg_6__u_txreg_data_int_reg_7__1446 (.o(net1446));
 b15tilo00an1n03x5 u_txreg_data_int_reg_8__u_txreg_data_int_reg_9__1447 (.o(net1447));
 b15tilo00an1n03x5 u_txreg_data_int_reg_8__u_txreg_data_int_reg_9__1448 (.o(net1448));
 b15tilo00an1n03x5 u_txreg_running_reg_1449 (.o(net1449));
 b15tihi00an1n03x5 U3043_1451 (.o(net1451));
 b15tihi00an1n03x5 U3047_1452 (.o(net1452));
 b15tihi00an1n03x5 U3164_1453 (.o(net1453));
 b15tihi00an1n03x5 U3292_1454 (.o(net1454));
 b15tihi00an1n03x5 U3294_1455 (.o(net1455));
 b15tihi00an1n03x5 U3300_1456 (.o(net1456));
 b15tihi00an1n03x5 U3302_1457 (.o(net1457));
 b15tihi00an1n03x5 U3304_1458 (.o(net1458));
 b15tihi00an1n03x5 U3306_1459 (.o(net1459));
 b15tihi00an1n03x5 U3314_1460 (.o(net1460));
 b15tihi00an1n03x5 U3419_1461 (.o(net1461));
 b15tihi00an1n03x5 U3421_1462 (.o(net1462));
 b15tihi00an1n03x5 U3423_1463 (.o(net1463));
 b15tihi00an1n03x5 U3425_1464 (.o(net1464));
 b15tihi00an1n03x5 U3427_1465 (.o(net1465));
 b15tihi00an1n03x5 U3429_1466 (.o(net1466));
 b15tihi00an1n03x5 U3431_1467 (.o(net1467));
 b15tihi00an1n03x5 U3433_1468 (.o(net1468));
 b15tihi00an1n03x5 U3435_1469 (.o(net1469));
 b15tihi00an1n03x5 U3437_1470 (.o(net1470));
 b15tihi00an1n03x5 U3441_1471 (.o(net1471));
 b15tihi00an1n03x5 U3443_1472 (.o(net1472));
 b15tihi00an1n03x5 U3445_1473 (.o(net1473));
 b15tihi00an1n03x5 U3447_1474 (.o(net1474));
 b15tihi00an1n03x5 U3449_1475 (.o(net1475));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__0__u_dcfifo_rx_u_din_buffer_data_reg_0__1__1476 (.o(net1476));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__10__u_dcfifo_rx_u_din_buffer_data_reg_0__11__1477 (.o(net1477));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__12__u_dcfifo_rx_u_din_buffer_data_reg_0__13__1478 (.o(net1478));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__14__u_dcfifo_rx_u_din_buffer_data_reg_0__15__1479 (.o(net1479));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__16__u_dcfifo_rx_u_din_buffer_data_reg_0__17__1480 (.o(net1480));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__18__u_dcfifo_rx_u_din_buffer_data_reg_0__19__1481 (.o(net1481));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__20__u_dcfifo_rx_u_din_buffer_data_reg_0__21__1482 (.o(net1482));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__22__u_dcfifo_rx_u_din_buffer_data_reg_0__23__1483 (.o(net1483));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__24__u_dcfifo_rx_u_din_buffer_data_reg_0__25__1484 (.o(net1484));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__26__u_dcfifo_rx_u_din_buffer_data_reg_0__27__1485 (.o(net1485));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__28__u_dcfifo_rx_u_din_buffer_data_reg_0__29__1486 (.o(net1486));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__2__u_dcfifo_rx_u_din_buffer_data_reg_0__3__1487 (.o(net1487));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__30__u_dcfifo_rx_u_din_buffer_data_reg_0__31__1488 (.o(net1488));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__4__u_dcfifo_rx_u_din_buffer_data_reg_0__5__1489 (.o(net1489));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__6__u_dcfifo_rx_u_din_buffer_data_reg_0__7__1490 (.o(net1490));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_0__8__u_dcfifo_rx_u_din_buffer_data_reg_0__9__1491 (.o(net1491));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__0__u_dcfifo_rx_u_din_buffer_data_reg_1__1__1492 (.o(net1492));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__10__u_dcfifo_rx_u_din_buffer_data_reg_1__11__1493 (.o(net1493));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__12__u_dcfifo_rx_u_din_buffer_data_reg_1__13__1494 (.o(net1494));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__14__u_dcfifo_rx_u_din_buffer_data_reg_1__15__1495 (.o(net1495));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__16__u_dcfifo_rx_u_din_buffer_data_reg_1__17__1496 (.o(net1496));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__18__u_dcfifo_rx_u_din_buffer_data_reg_1__19__1497 (.o(net1497));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__20__u_dcfifo_rx_u_din_buffer_data_reg_1__21__1498 (.o(net1498));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__22__u_dcfifo_rx_u_din_buffer_data_reg_1__23__1499 (.o(net1499));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__24__u_dcfifo_rx_u_din_buffer_data_reg_1__25__1500 (.o(net1500));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__26__u_dcfifo_rx_u_din_buffer_data_reg_1__27__1501 (.o(net1501));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__28__u_dcfifo_rx_u_din_buffer_data_reg_1__29__1502 (.o(net1502));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__2__u_dcfifo_rx_u_din_buffer_data_reg_1__3__1503 (.o(net1503));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__30__u_dcfifo_rx_u_din_buffer_data_reg_1__31__1504 (.o(net1504));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__4__u_dcfifo_rx_u_din_buffer_data_reg_1__5__1505 (.o(net1505));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__6__u_dcfifo_rx_u_din_buffer_data_reg_1__7__1506 (.o(net1506));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_1__8__u_dcfifo_rx_u_din_buffer_data_reg_1__9__1507 (.o(net1507));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__0__u_dcfifo_rx_u_din_buffer_data_reg_2__1__1508 (.o(net1508));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__10__u_dcfifo_rx_u_din_buffer_data_reg_2__11__1509 (.o(net1509));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__12__u_dcfifo_rx_u_din_buffer_data_reg_2__13__1510 (.o(net1510));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__14__u_dcfifo_rx_u_din_buffer_data_reg_2__15__1511 (.o(net1511));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__16__u_dcfifo_rx_u_din_buffer_data_reg_2__17__1512 (.o(net1512));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__18__u_dcfifo_rx_u_din_buffer_data_reg_2__19__1513 (.o(net1513));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__20__u_dcfifo_rx_u_din_buffer_data_reg_2__21__1514 (.o(net1514));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__22__u_dcfifo_rx_u_din_buffer_data_reg_2__23__1515 (.o(net1515));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__24__u_dcfifo_rx_u_din_buffer_data_reg_2__25__1516 (.o(net1516));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__26__u_dcfifo_rx_u_din_buffer_data_reg_2__27__1517 (.o(net1517));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__28__u_dcfifo_rx_u_din_buffer_data_reg_2__29__1518 (.o(net1518));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__2__u_dcfifo_rx_u_din_buffer_data_reg_2__3__1519 (.o(net1519));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__30__u_dcfifo_rx_u_din_buffer_data_reg_2__31__1520 (.o(net1520));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__4__u_dcfifo_rx_u_din_buffer_data_reg_2__5__1521 (.o(net1521));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__6__u_dcfifo_rx_u_din_buffer_data_reg_2__7__1522 (.o(net1522));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_2__8__u_dcfifo_rx_u_din_buffer_data_reg_2__9__1523 (.o(net1523));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__0__u_dcfifo_rx_u_din_buffer_data_reg_3__1__1524 (.o(net1524));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__10__u_dcfifo_rx_u_din_buffer_data_reg_3__11__1525 (.o(net1525));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__12__u_dcfifo_rx_u_din_buffer_data_reg_3__13__1526 (.o(net1526));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__14__u_dcfifo_rx_u_din_buffer_data_reg_3__15__1527 (.o(net1527));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__16__u_dcfifo_rx_u_din_buffer_data_reg_3__17__1528 (.o(net1528));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__18__u_dcfifo_rx_u_din_buffer_data_reg_3__19__1529 (.o(net1529));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__20__u_dcfifo_rx_u_din_buffer_data_reg_3__21__1530 (.o(net1530));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__22__u_dcfifo_rx_u_din_buffer_data_reg_3__23__1531 (.o(net1531));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__24__u_dcfifo_rx_u_din_buffer_data_reg_3__25__1532 (.o(net1532));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__26__u_dcfifo_rx_u_din_buffer_data_reg_3__27__1533 (.o(net1533));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__28__u_dcfifo_rx_u_din_buffer_data_reg_3__29__1534 (.o(net1534));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__2__u_dcfifo_rx_u_din_buffer_data_reg_3__3__1535 (.o(net1535));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__30__u_dcfifo_rx_u_din_buffer_data_reg_3__31__1536 (.o(net1536));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__4__u_dcfifo_rx_u_din_buffer_data_reg_3__5__1537 (.o(net1537));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__6__u_dcfifo_rx_u_din_buffer_data_reg_3__7__1538 (.o(net1538));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_3__8__u_dcfifo_rx_u_din_buffer_data_reg_3__9__1539 (.o(net1539));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__0__u_dcfifo_rx_u_din_buffer_data_reg_4__1__1540 (.o(net1540));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__10__u_dcfifo_rx_u_din_buffer_data_reg_4__11__1541 (.o(net1541));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__12__u_dcfifo_rx_u_din_buffer_data_reg_4__13__1542 (.o(net1542));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__14__u_dcfifo_rx_u_din_buffer_data_reg_4__15__1543 (.o(net1543));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__16__u_dcfifo_rx_u_din_buffer_data_reg_4__17__1544 (.o(net1544));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__18__u_dcfifo_rx_u_din_buffer_data_reg_4__19__1545 (.o(net1545));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__20__u_dcfifo_rx_u_din_buffer_data_reg_4__21__1546 (.o(net1546));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__22__u_dcfifo_rx_u_din_buffer_data_reg_4__23__1547 (.o(net1547));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__24__u_dcfifo_rx_u_din_buffer_data_reg_4__25__1548 (.o(net1548));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__26__u_dcfifo_rx_u_din_buffer_data_reg_4__27__1549 (.o(net1549));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__28__u_dcfifo_rx_u_din_buffer_data_reg_4__29__1550 (.o(net1550));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__2__u_dcfifo_rx_u_din_buffer_data_reg_4__3__1551 (.o(net1551));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__30__u_dcfifo_rx_u_din_buffer_data_reg_4__31__1552 (.o(net1552));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__4__u_dcfifo_rx_u_din_buffer_data_reg_4__5__1553 (.o(net1553));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__6__u_dcfifo_rx_u_din_buffer_data_reg_4__7__1554 (.o(net1554));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_4__8__u_dcfifo_rx_u_din_buffer_data_reg_4__9__1555 (.o(net1555));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__0__u_dcfifo_rx_u_din_buffer_data_reg_5__1__1556 (.o(net1556));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__10__u_dcfifo_rx_u_din_buffer_data_reg_5__11__1557 (.o(net1557));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__12__u_dcfifo_rx_u_din_buffer_data_reg_5__13__1558 (.o(net1558));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__14__u_dcfifo_rx_u_din_buffer_data_reg_5__15__1559 (.o(net1559));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__16__u_dcfifo_rx_u_din_buffer_data_reg_5__17__1560 (.o(net1560));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__18__u_dcfifo_rx_u_din_buffer_data_reg_5__19__1561 (.o(net1561));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__20__u_dcfifo_rx_u_din_buffer_data_reg_5__21__1562 (.o(net1562));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__22__u_dcfifo_rx_u_din_buffer_data_reg_5__23__1563 (.o(net1563));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__24__u_dcfifo_rx_u_din_buffer_data_reg_5__25__1564 (.o(net1564));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__26__u_dcfifo_rx_u_din_buffer_data_reg_5__27__1565 (.o(net1565));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__28__u_dcfifo_rx_u_din_buffer_data_reg_5__29__1566 (.o(net1566));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__2__u_dcfifo_rx_u_din_buffer_data_reg_5__3__1567 (.o(net1567));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__30__u_dcfifo_rx_u_din_buffer_data_reg_5__31__1568 (.o(net1568));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__4__u_dcfifo_rx_u_din_buffer_data_reg_5__5__1569 (.o(net1569));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__6__u_dcfifo_rx_u_din_buffer_data_reg_5__7__1570 (.o(net1570));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_5__8__u_dcfifo_rx_u_din_buffer_data_reg_5__9__1571 (.o(net1571));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__0__u_dcfifo_rx_u_din_buffer_data_reg_6__1__1572 (.o(net1572));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__10__u_dcfifo_rx_u_din_buffer_data_reg_6__11__1573 (.o(net1573));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__12__u_dcfifo_rx_u_din_buffer_data_reg_6__13__1574 (.o(net1574));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__14__u_dcfifo_rx_u_din_buffer_data_reg_6__15__1575 (.o(net1575));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__16__u_dcfifo_rx_u_din_buffer_data_reg_6__17__1576 (.o(net1576));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__18__u_dcfifo_rx_u_din_buffer_data_reg_6__19__1577 (.o(net1577));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__20__u_dcfifo_rx_u_din_buffer_data_reg_6__21__1578 (.o(net1578));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__22__u_dcfifo_rx_u_din_buffer_data_reg_6__23__1579 (.o(net1579));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__24__u_dcfifo_rx_u_din_buffer_data_reg_6__25__1580 (.o(net1580));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__26__u_dcfifo_rx_u_din_buffer_data_reg_6__27__1581 (.o(net1581));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__28__u_dcfifo_rx_u_din_buffer_data_reg_6__29__1582 (.o(net1582));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__2__u_dcfifo_rx_u_din_buffer_data_reg_6__3__1583 (.o(net1583));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__30__u_dcfifo_rx_u_din_buffer_data_reg_6__31__1584 (.o(net1584));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__4__u_dcfifo_rx_u_din_buffer_data_reg_6__5__1585 (.o(net1585));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__6__u_dcfifo_rx_u_din_buffer_data_reg_6__7__1586 (.o(net1586));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_6__8__u_dcfifo_rx_u_din_buffer_data_reg_6__9__1587 (.o(net1587));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__0__u_dcfifo_rx_u_din_buffer_data_reg_7__1__1588 (.o(net1588));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__10__u_dcfifo_rx_u_din_buffer_data_reg_7__11__1589 (.o(net1589));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__12__u_dcfifo_rx_u_din_buffer_data_reg_7__13__1590 (.o(net1590));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__14__u_dcfifo_rx_u_din_buffer_data_reg_7__15__1591 (.o(net1591));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__16__u_dcfifo_rx_u_din_buffer_data_reg_7__17__1592 (.o(net1592));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__18__u_dcfifo_rx_u_din_buffer_data_reg_7__19__1593 (.o(net1593));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__20__u_dcfifo_rx_u_din_buffer_data_reg_7__21__1594 (.o(net1594));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__22__u_dcfifo_rx_u_din_buffer_data_reg_7__23__1595 (.o(net1595));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__24__u_dcfifo_rx_u_din_buffer_data_reg_7__25__1596 (.o(net1596));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__26__u_dcfifo_rx_u_din_buffer_data_reg_7__27__1597 (.o(net1597));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__28__u_dcfifo_rx_u_din_buffer_data_reg_7__29__1598 (.o(net1598));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__2__u_dcfifo_rx_u_din_buffer_data_reg_7__3__1599 (.o(net1599));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__30__u_dcfifo_rx_u_din_buffer_data_reg_7__31__1600 (.o(net1600));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__4__u_dcfifo_rx_u_din_buffer_data_reg_7__5__1601 (.o(net1601));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__6__u_dcfifo_rx_u_din_buffer_data_reg_7__7__1602 (.o(net1602));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_buffer_data_reg_7__8__u_dcfifo_rx_u_din_buffer_data_reg_7__9__1603 (.o(net1603));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_full_full_synch_d_middle_reg_0__u_dcfifo_rx_u_din_full_full_synch_d_out_reg_0__1604 (.o(net1604));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_full_latched_full_s_reg_u_dcfifo_tx_u_dout_empty_synch_d_out_reg_1__1605 (.o(net1605));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_write_tr_state_reg_0__u_dcfifo_rx_u_din_write_tr_state_reg_1__1606 (.o(net1606));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_write_tr_state_reg_2__1607 (.o(net1607));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_write_tr_state_reg_3__1608 (.o(net1608));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_write_tr_state_reg_4__u_dcfifo_rx_u_din_write_tr_state_reg_5__1609 (.o(net1609));
 b15tihi00an1n03x5 u_dcfifo_rx_u_din_write_tr_state_reg_6__u_dcfifo_rx_u_din_write_tr_state_reg_7__1610 (.o(net1610));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_0__u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_1__1611 (.o(net1611));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_2__1612 (.o(net1612));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_3__1613 (.o(net1613));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_4__u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_5__1614 (.o(net1614));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_6__u_dcfifo_rx_u_dout_empty_synch_d_middle_reg_7__1615 (.o(net1615));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_0__u_dcfifo_rx_u_dout_empty_synch_d_out_reg_1__1616 (.o(net1616));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_2__1617 (.o(net1617));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_3__1618 (.o(net1618));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_4__u_dcfifo_rx_u_dout_empty_synch_d_out_reg_5__1619 (.o(net1619));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_empty_synch_d_out_reg_6__u_dcfifo_rx_u_dout_empty_synch_d_out_reg_7__1620 (.o(net1620));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_read_tr_state_reg_0__1621 (.o(net1621));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_read_tr_state_reg_1__1622 (.o(net1622));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_read_tr_state_reg_2__u_dcfifo_rx_u_dout_read_tr_state_reg_3__1623 (.o(net1623));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_read_tr_state_reg_4__u_dcfifo_rx_u_dout_read_tr_state_reg_5__1624 (.o(net1624));
 b15tihi00an1n03x5 u_dcfifo_rx_u_dout_read_tr_state_reg_6__u_dcfifo_rx_u_dout_read_tr_state_reg_7__1625 (.o(net1625));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__0__u_dcfifo_tx_u_din_buffer_data_reg_0__1__1626 (.o(net1626));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__10__u_dcfifo_tx_u_din_buffer_data_reg_0__11__1627 (.o(net1627));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__12__u_dcfifo_tx_u_din_buffer_data_reg_0__13__1628 (.o(net1628));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__14__u_dcfifo_tx_u_din_buffer_data_reg_0__15__1629 (.o(net1629));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__16__u_dcfifo_tx_u_din_buffer_data_reg_0__17__1630 (.o(net1630));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__18__u_dcfifo_tx_u_din_buffer_data_reg_0__19__1631 (.o(net1631));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__20__u_dcfifo_tx_u_din_buffer_data_reg_0__21__1632 (.o(net1632));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__22__u_dcfifo_tx_u_din_buffer_data_reg_0__23__1633 (.o(net1633));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__24__u_dcfifo_tx_u_din_buffer_data_reg_0__25__1634 (.o(net1634));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__26__u_dcfifo_tx_u_din_buffer_data_reg_0__27__1635 (.o(net1635));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__28__u_dcfifo_tx_u_din_buffer_data_reg_0__29__1636 (.o(net1636));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__2__u_dcfifo_tx_u_din_buffer_data_reg_0__3__1637 (.o(net1637));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__30__u_dcfifo_tx_u_din_buffer_data_reg_0__31__1638 (.o(net1638));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__4__u_dcfifo_tx_u_din_buffer_data_reg_0__5__1639 (.o(net1639));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__6__u_dcfifo_tx_u_din_buffer_data_reg_0__7__1640 (.o(net1640));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_0__8__u_dcfifo_tx_u_din_buffer_data_reg_0__9__1641 (.o(net1641));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__0__u_dcfifo_tx_u_din_buffer_data_reg_1__1__1642 (.o(net1642));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__10__u_dcfifo_tx_u_din_buffer_data_reg_1__11__1643 (.o(net1643));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__12__u_dcfifo_tx_u_din_buffer_data_reg_1__13__1644 (.o(net1644));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__14__u_dcfifo_tx_u_din_buffer_data_reg_1__15__1645 (.o(net1645));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__16__u_dcfifo_tx_u_din_buffer_data_reg_1__17__1646 (.o(net1646));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__18__u_dcfifo_tx_u_din_buffer_data_reg_1__19__1647 (.o(net1647));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__20__u_dcfifo_tx_u_din_buffer_data_reg_1__21__1648 (.o(net1648));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__22__u_dcfifo_tx_u_din_buffer_data_reg_1__23__1649 (.o(net1649));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__24__u_dcfifo_tx_u_din_buffer_data_reg_1__25__1650 (.o(net1650));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__26__u_dcfifo_tx_u_din_buffer_data_reg_1__27__1651 (.o(net1651));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__28__u_dcfifo_tx_u_din_buffer_data_reg_1__29__1652 (.o(net1652));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__2__u_dcfifo_tx_u_din_buffer_data_reg_1__3__1653 (.o(net1653));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__30__u_dcfifo_tx_u_din_buffer_data_reg_1__31__1654 (.o(net1654));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__4__u_dcfifo_tx_u_din_buffer_data_reg_1__5__1655 (.o(net1655));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__6__u_dcfifo_tx_u_din_buffer_data_reg_1__7__1656 (.o(net1656));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_1__8__u_dcfifo_tx_u_din_buffer_data_reg_1__9__1657 (.o(net1657));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__0__u_dcfifo_tx_u_din_buffer_data_reg_2__1__1658 (.o(net1658));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__10__u_dcfifo_tx_u_din_buffer_data_reg_2__11__1659 (.o(net1659));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__12__u_dcfifo_tx_u_din_buffer_data_reg_2__13__1660 (.o(net1660));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__14__u_dcfifo_tx_u_din_buffer_data_reg_2__15__1661 (.o(net1661));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__16__u_dcfifo_tx_u_din_buffer_data_reg_2__17__1662 (.o(net1662));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__18__u_dcfifo_tx_u_din_buffer_data_reg_2__19__1663 (.o(net1663));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__20__u_dcfifo_tx_u_din_buffer_data_reg_2__21__1664 (.o(net1664));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__22__u_dcfifo_tx_u_din_buffer_data_reg_2__23__1665 (.o(net1665));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__24__u_dcfifo_tx_u_din_buffer_data_reg_2__25__1666 (.o(net1666));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__26__u_dcfifo_tx_u_din_buffer_data_reg_2__27__1667 (.o(net1667));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__28__u_dcfifo_tx_u_din_buffer_data_reg_2__29__1668 (.o(net1668));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__2__u_dcfifo_tx_u_din_buffer_data_reg_2__3__1669 (.o(net1669));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__30__u_dcfifo_tx_u_din_buffer_data_reg_2__31__1670 (.o(net1670));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__4__u_dcfifo_tx_u_din_buffer_data_reg_2__5__1671 (.o(net1671));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__6__u_dcfifo_tx_u_din_buffer_data_reg_2__7__1672 (.o(net1672));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_2__8__u_dcfifo_tx_u_din_buffer_data_reg_2__9__1673 (.o(net1673));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__0__u_dcfifo_tx_u_din_buffer_data_reg_3__1__1674 (.o(net1674));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__10__u_dcfifo_tx_u_din_buffer_data_reg_3__11__1675 (.o(net1675));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__12__u_dcfifo_tx_u_din_buffer_data_reg_3__13__1676 (.o(net1676));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__14__u_dcfifo_tx_u_din_buffer_data_reg_3__15__1677 (.o(net1677));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__16__u_dcfifo_tx_u_din_buffer_data_reg_3__17__1678 (.o(net1678));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__18__u_dcfifo_tx_u_din_buffer_data_reg_3__19__1679 (.o(net1679));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__20__u_dcfifo_tx_u_din_buffer_data_reg_3__21__1680 (.o(net1680));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__22__u_dcfifo_tx_u_din_buffer_data_reg_3__23__1681 (.o(net1681));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__24__u_dcfifo_tx_u_din_buffer_data_reg_3__25__1682 (.o(net1682));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__26__u_dcfifo_tx_u_din_buffer_data_reg_3__27__1683 (.o(net1683));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__28__u_dcfifo_tx_u_din_buffer_data_reg_3__29__1684 (.o(net1684));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__2__u_dcfifo_tx_u_din_buffer_data_reg_3__3__1685 (.o(net1685));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__30__u_dcfifo_tx_u_din_buffer_data_reg_3__31__1686 (.o(net1686));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__4__u_dcfifo_tx_u_din_buffer_data_reg_3__5__1687 (.o(net1687));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__6__u_dcfifo_tx_u_din_buffer_data_reg_3__7__1688 (.o(net1688));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_3__8__u_dcfifo_tx_u_din_buffer_data_reg_3__9__1689 (.o(net1689));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__0__u_dcfifo_tx_u_din_buffer_data_reg_4__1__1690 (.o(net1690));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__10__u_dcfifo_tx_u_din_buffer_data_reg_4__11__1691 (.o(net1691));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__12__u_dcfifo_tx_u_din_buffer_data_reg_4__13__1692 (.o(net1692));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__14__u_dcfifo_tx_u_din_buffer_data_reg_4__15__1693 (.o(net1693));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__16__u_dcfifo_tx_u_din_buffer_data_reg_4__17__1694 (.o(net1694));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__18__u_dcfifo_tx_u_din_buffer_data_reg_4__19__1695 (.o(net1695));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__20__u_dcfifo_tx_u_din_buffer_data_reg_4__21__1696 (.o(net1696));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__22__u_dcfifo_tx_u_din_buffer_data_reg_4__23__1697 (.o(net1697));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__24__u_dcfifo_tx_u_din_buffer_data_reg_4__25__1698 (.o(net1698));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__26__u_dcfifo_tx_u_din_buffer_data_reg_4__27__1699 (.o(net1699));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__28__u_dcfifo_tx_u_din_buffer_data_reg_4__29__1700 (.o(net1700));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__2__u_dcfifo_tx_u_din_buffer_data_reg_4__3__1701 (.o(net1701));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__30__u_dcfifo_tx_u_din_buffer_data_reg_4__31__1702 (.o(net1702));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__4__u_dcfifo_tx_u_din_buffer_data_reg_4__5__1703 (.o(net1703));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__6__u_dcfifo_tx_u_din_buffer_data_reg_4__7__1704 (.o(net1704));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_4__8__u_dcfifo_tx_u_din_buffer_data_reg_4__9__1705 (.o(net1705));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__0__u_dcfifo_tx_u_din_buffer_data_reg_5__1__1706 (.o(net1706));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__10__u_dcfifo_tx_u_din_buffer_data_reg_5__11__1707 (.o(net1707));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__12__u_dcfifo_tx_u_din_buffer_data_reg_5__13__1708 (.o(net1708));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__14__u_dcfifo_tx_u_din_buffer_data_reg_5__15__1709 (.o(net1709));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__16__u_dcfifo_tx_u_din_buffer_data_reg_5__17__1710 (.o(net1710));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__18__u_dcfifo_tx_u_din_buffer_data_reg_5__19__1711 (.o(net1711));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__20__u_dcfifo_tx_u_din_buffer_data_reg_5__21__1712 (.o(net1712));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__22__u_dcfifo_tx_u_din_buffer_data_reg_5__23__1713 (.o(net1713));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__24__u_dcfifo_tx_u_din_buffer_data_reg_5__25__1714 (.o(net1714));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__26__u_dcfifo_tx_u_din_buffer_data_reg_5__27__1715 (.o(net1715));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__28__u_dcfifo_tx_u_din_buffer_data_reg_5__29__1716 (.o(net1716));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__2__u_dcfifo_tx_u_din_buffer_data_reg_5__3__1717 (.o(net1717));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__30__u_dcfifo_tx_u_din_buffer_data_reg_5__31__1718 (.o(net1718));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__4__u_dcfifo_tx_u_din_buffer_data_reg_5__5__1719 (.o(net1719));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__6__u_dcfifo_tx_u_din_buffer_data_reg_5__7__1720 (.o(net1720));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_5__8__u_dcfifo_tx_u_din_buffer_data_reg_5__9__1721 (.o(net1721));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__0__u_dcfifo_tx_u_din_buffer_data_reg_6__1__1722 (.o(net1722));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__10__u_dcfifo_tx_u_din_buffer_data_reg_6__11__1723 (.o(net1723));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__12__u_dcfifo_tx_u_din_buffer_data_reg_6__13__1724 (.o(net1724));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__14__u_dcfifo_tx_u_din_buffer_data_reg_6__15__1725 (.o(net1725));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__16__u_dcfifo_tx_u_din_buffer_data_reg_6__17__1726 (.o(net1726));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__18__u_dcfifo_tx_u_din_buffer_data_reg_6__19__1727 (.o(net1727));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__20__u_dcfifo_tx_u_din_buffer_data_reg_6__21__1728 (.o(net1728));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__22__u_dcfifo_tx_u_din_buffer_data_reg_6__23__1729 (.o(net1729));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__24__u_dcfifo_tx_u_din_buffer_data_reg_6__25__1730 (.o(net1730));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__26__u_dcfifo_tx_u_din_buffer_data_reg_6__27__1731 (.o(net1731));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__28__u_dcfifo_tx_u_din_buffer_data_reg_6__29__1732 (.o(net1732));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__2__u_dcfifo_tx_u_din_buffer_data_reg_6__3__1733 (.o(net1733));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__30__u_dcfifo_tx_u_din_buffer_data_reg_6__31__1734 (.o(net1734));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__4__u_dcfifo_tx_u_din_buffer_data_reg_6__5__1735 (.o(net1735));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__6__u_dcfifo_tx_u_din_buffer_data_reg_6__7__1736 (.o(net1736));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_6__8__u_dcfifo_tx_u_din_buffer_data_reg_6__9__1737 (.o(net1737));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__0__u_dcfifo_tx_u_din_buffer_data_reg_7__1__1738 (.o(net1738));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__10__u_dcfifo_tx_u_din_buffer_data_reg_7__11__1739 (.o(net1739));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__12__u_dcfifo_tx_u_din_buffer_data_reg_7__13__1740 (.o(net1740));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__14__u_dcfifo_tx_u_din_buffer_data_reg_7__15__1741 (.o(net1741));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__16__u_dcfifo_tx_u_din_buffer_data_reg_7__17__1742 (.o(net1742));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__18__u_dcfifo_tx_u_din_buffer_data_reg_7__19__1743 (.o(net1743));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__20__u_dcfifo_tx_u_din_buffer_data_reg_7__21__1744 (.o(net1744));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__22__u_dcfifo_tx_u_din_buffer_data_reg_7__23__1745 (.o(net1745));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__24__u_dcfifo_tx_u_din_buffer_data_reg_7__25__1746 (.o(net1746));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__26__u_dcfifo_tx_u_din_buffer_data_reg_7__27__1747 (.o(net1747));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__28__u_dcfifo_tx_u_din_buffer_data_reg_7__29__1748 (.o(net1748));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__2__u_dcfifo_tx_u_din_buffer_data_reg_7__3__1749 (.o(net1749));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__30__u_dcfifo_tx_u_din_buffer_data_reg_7__31__1750 (.o(net1750));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__4__u_dcfifo_tx_u_din_buffer_data_reg_7__5__1751 (.o(net1751));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__6__u_dcfifo_tx_u_din_buffer_data_reg_7__7__1752 (.o(net1752));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_buffer_data_reg_7__8__u_dcfifo_tx_u_din_buffer_data_reg_7__9__1753 (.o(net1753));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_full_full_synch_d_middle_reg_0__u_dcfifo_tx_u_din_full_full_synch_d_out_reg_0__1754 (.o(net1754));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_full_latched_full_s_reg_u_spi_device_tlul_plug_state_reg_0__1755 (.o(net1755));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_write_tr_state_reg_0__u_dcfifo_tx_u_din_write_tr_state_reg_1__1756 (.o(net1756));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_write_tr_state_reg_2__1757 (.o(net1757));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_write_tr_state_reg_3__1758 (.o(net1758));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_write_tr_state_reg_4__u_dcfifo_tx_u_din_write_tr_state_reg_5__1759 (.o(net1759));
 b15tihi00an1n03x5 u_dcfifo_tx_u_din_write_tr_state_reg_6__u_dcfifo_tx_u_din_write_tr_state_reg_7__1760 (.o(net1760));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_0__u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_1__1761 (.o(net1761));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_2__1762 (.o(net1762));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_3__1763 (.o(net1763));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_4__u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_5__1764 (.o(net1764));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_6__u_dcfifo_tx_u_dout_empty_synch_d_middle_reg_7__1765 (.o(net1765));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_0__u_dcfifo_tx_u_dout_empty_synch_d_out_reg_5__1766 (.o(net1766));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_2__1767 (.o(net1767));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_3__1768 (.o(net1768));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_4__1769 (.o(net1769));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_empty_synch_d_out_reg_6__u_dcfifo_tx_u_dout_empty_synch_d_out_reg_7__1770 (.o(net1770));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_read_tr_state_reg_0__1771 (.o(net1771));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_read_tr_state_reg_1__1772 (.o(net1772));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_read_tr_state_reg_2__u_dcfifo_tx_u_dout_read_tr_state_reg_3__1773 (.o(net1773));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_read_tr_state_reg_4__u_dcfifo_tx_u_dout_read_tr_state_reg_5__1774 (.o(net1774));
 b15tihi00an1n03x5 u_dcfifo_tx_u_dout_read_tr_state_reg_6__u_dcfifo_tx_u_dout_read_tr_state_reg_7__1775 (.o(net1775));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_0__u_device_sm_addr_reg_reg_1__1776 (.o(net1776));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_10__u_device_sm_addr_reg_reg_11__1777 (.o(net1777));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_12__u_device_sm_addr_reg_reg_13__1778 (.o(net1778));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_14__u_device_sm_addr_reg_reg_15__1779 (.o(net1779));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_16__u_device_sm_addr_reg_reg_17__1780 (.o(net1780));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_18__u_device_sm_addr_reg_reg_19__1781 (.o(net1781));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_20__u_device_sm_addr_reg_reg_21__1782 (.o(net1782));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_22__u_device_sm_addr_reg_reg_23__1783 (.o(net1783));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_24__u_device_sm_addr_reg_reg_25__1784 (.o(net1784));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_26__u_device_sm_addr_reg_reg_27__1785 (.o(net1785));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_28__u_device_sm_addr_reg_reg_29__1786 (.o(net1786));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_2__u_device_sm_addr_reg_reg_3__1787 (.o(net1787));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_30__u_device_sm_addr_reg_reg_31__1788 (.o(net1788));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_4__u_device_sm_addr_reg_reg_5__1789 (.o(net1789));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_6__u_device_sm_addr_reg_reg_7__1790 (.o(net1790));
 b15tihi00an1n03x5 u_device_sm_addr_reg_reg_8__u_device_sm_addr_reg_reg_9__1791 (.o(net1791));
 b15tihi00an1n03x5 u_device_sm_cmd_reg_reg_0__u_device_sm_cmd_reg_reg_1__1792 (.o(net1792));
 b15tihi00an1n03x5 u_device_sm_cmd_reg_reg_2__u_device_sm_cmd_reg_reg_3__1793 (.o(net1793));
 b15tihi00an1n03x5 u_device_sm_cmd_reg_reg_4__u_device_sm_cmd_reg_reg_5__1794 (.o(net1794));
 b15tihi00an1n03x5 u_device_sm_cmd_reg_reg_6__u_device_sm_cmd_reg_reg_7__1795 (.o(net1795));
 b15tihi00an1n03x5 u_device_sm_ctrl_addr_valid_reg_u_device_sm_data_reg_reg_0__1796 (.o(net1796));
 b15tihi00an1n03x5 u_device_sm_ctrl_data_tx_ready_reg_u_device_sm_state_reg_1__1797 (.o(net1797));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_10__u_device_sm_data_reg_reg_11__1798 (.o(net1798));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_12__u_device_sm_data_reg_reg_13__1799 (.o(net1799));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_14__u_device_sm_data_reg_reg_15__1800 (.o(net1800));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_16__u_device_sm_data_reg_reg_17__1801 (.o(net1801));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_18__u_device_sm_data_reg_reg_19__1802 (.o(net1802));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_1__u_device_sm_data_reg_reg_2__1803 (.o(net1803));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_20__u_device_sm_data_reg_reg_21__1804 (.o(net1804));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_22__u_device_sm_data_reg_reg_23__1805 (.o(net1805));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_24__u_device_sm_data_reg_reg_25__1806 (.o(net1806));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_26__u_device_sm_data_reg_reg_27__1807 (.o(net1807));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_28__u_device_sm_data_reg_reg_29__1808 (.o(net1808));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_30__u_device_sm_data_reg_reg_31__1809 (.o(net1809));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_3__u_device_sm_data_reg_reg_4__1810 (.o(net1810));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_5__u_device_sm_state_reg_0__1811 (.o(net1811));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_6__u_device_sm_data_reg_reg_7__1812 (.o(net1812));
 b15tihi00an1n03x5 u_device_sm_data_reg_reg_8__u_device_sm_data_reg_reg_9__1813 (.o(net1813));
 b15tihi00an1n03x5 u_device_sm_mode_reg_reg_0__u_device_sm_mode_reg_reg_1__1814 (.o(net1814));
 b15tihi00an1n03x5 u_device_sm_mode_reg_reg_2__u_device_sm_mode_reg_reg_3__1815 (.o(net1815));
 b15tihi00an1n03x5 u_device_sm_mode_reg_reg_4__u_device_sm_mode_reg_reg_5__1816 (.o(net1816));
 b15tihi00an1n03x5 u_device_sm_mode_reg_reg_6__u_device_sm_mode_reg_reg_7__1817 (.o(net1817));
 b15tihi00an1n03x5 u_device_sm_pad_mode_next_reg_0__1818 (.o(net1818));
 b15tihi00an1n03x5 u_device_sm_state_reg_2__u_device_sm_tx_counter_reg_0__1819 (.o(net1819));
 b15tihi00an1n03x5 u_device_sm_state_reg_2__u_device_sm_tx_counter_reg_0__1820 (.o(net1820));
 b15tihi00an1n03x5 u_device_sm_tx_counter_reg_1__u_device_sm_tx_data_reg_0__1821 (.o(net1821));
 b15tihi00an1n03x5 u_device_sm_tx_counter_reg_1__u_device_sm_tx_data_reg_0__1822 (.o(net1822));
 b15tihi00an1n03x5 u_device_sm_tx_counter_reg_2__u_device_sm_tx_counter_reg_3__1823 (.o(net1823));
 b15tihi00an1n03x5 u_device_sm_tx_counter_reg_2__u_device_sm_tx_counter_reg_3__1824 (.o(net1824));
 b15tihi00an1n03x5 u_device_sm_tx_counter_reg_4__u_device_sm_tx_counter_upd_reg_1825 (.o(net1825));
 b15tihi00an1n03x5 u_device_sm_tx_counter_reg_5__u_device_sm_tx_counter_reg_6__1826 (.o(net1826));
 b15tihi00an1n03x5 u_device_sm_tx_counter_reg_7__1827 (.o(net1827));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_11__u_device_sm_tx_data_reg_12__1828 (.o(net1828));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_13__u_device_sm_tx_data_reg_14__1829 (.o(net1829));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_15__1830 (.o(net1830));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_16__u_device_sm_tx_data_reg_17__1831 (.o(net1831));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_18__u_device_sm_tx_data_reg_19__1832 (.o(net1832));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_1__u_device_sm_tx_data_reg_2__1833 (.o(net1833));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_20__u_device_sm_tx_data_reg_21__1834 (.o(net1834));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_22__u_device_sm_tx_data_reg_23__1835 (.o(net1835));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_24__u_device_sm_tx_data_reg_25__1836 (.o(net1836));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_26__u_device_sm_tx_data_reg_27__1837 (.o(net1837));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_28__u_device_sm_tx_data_reg_29__1838 (.o(net1838));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_30__u_device_sm_tx_data_reg_31__1839 (.o(net1839));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_3__u_device_sm_tx_data_reg_4__1840 (.o(net1840));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_5__u_device_sm_tx_data_reg_6__1841 (.o(net1841));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_7__u_device_sm_tx_data_reg_8__1842 (.o(net1842));
 b15tihi00an1n03x5 u_device_sm_tx_data_reg_9__u_device_sm_tx_data_reg_10__1843 (.o(net1843));
 b15tihi00an1n03x5 u_device_sm_tx_data_valid_reg_u_device_sm_tx_done_reg_reg_1844 (.o(net1844));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg0_reg_0__u_device_sm_u_spiregs_reg0_reg_1__1845 (.o(net1845));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg0_reg_2__u_device_sm_u_spiregs_reg0_reg_3__1846 (.o(net1846));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg0_reg_4__u_device_sm_u_spiregs_reg0_reg_5__1847 (.o(net1847));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg0_reg_6__u_device_sm_u_spiregs_reg0_reg_7__1848 (.o(net1848));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg1_reg_0__u_device_sm_u_spiregs_reg1_reg_1__1849 (.o(net1849));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg1_reg_2__u_device_sm_u_spiregs_reg1_reg_3__1850 (.o(net1850));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg1_reg_4__u_device_sm_u_spiregs_reg1_reg_6__1851 (.o(net1851));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg1_reg_5__1852 (.o(net1852));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg1_reg_7__1853 (.o(net1853));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg2_reg_0__u_device_sm_u_spiregs_reg2_reg_1__1854 (.o(net1854));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg2_reg_2__u_device_sm_u_spiregs_reg2_reg_3__1855 (.o(net1855));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg2_reg_4__u_device_sm_u_spiregs_reg2_reg_5__1856 (.o(net1856));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg2_reg_6__u_device_sm_u_spiregs_reg2_reg_7__1857 (.o(net1857));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg3_reg_0__u_device_sm_u_spiregs_reg3_reg_1__1858 (.o(net1858));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg3_reg_2__u_device_sm_u_spiregs_reg3_reg_3__1859 (.o(net1859));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg3_reg_4__u_device_sm_u_spiregs_reg3_reg_5__1860 (.o(net1860));
 b15tihi00an1n03x5 u_device_sm_u_spiregs_reg3_reg_6__u_device_sm_u_spiregs_reg3_reg_7__1861 (.o(net1861));
 b15tihi00an1n03x5 u_rxreg_counter_reg_0__u_rxreg_counter_reg_1__1862 (.o(net1862));
 b15tihi00an1n03x5 u_rxreg_counter_reg_2__u_rxreg_counter_reg_3__1863 (.o(net1863));
 b15tihi00an1n03x5 u_rxreg_counter_reg_4__u_rxreg_counter_reg_5__1864 (.o(net1864));
 b15tihi00an1n03x5 u_rxreg_counter_reg_6__u_rxreg_counter_reg_7__1865 (.o(net1865));
 b15tihi00an1n03x5 u_rxreg_counter_trgt_reg_0__1866 (.o(net1866));
 b15tihi00an1n03x5 u_rxreg_counter_trgt_reg_1__u_rxreg_counter_trgt_reg_2__1867 (.o(net1867));
 b15tihi00an1n03x5 u_rxreg_counter_trgt_reg_3__u_rxreg_counter_trgt_reg_4__1868 (.o(net1868));
 b15tihi00an1n03x5 u_rxreg_counter_trgt_reg_5__u_rxreg_counter_trgt_reg_6__1869 (.o(net1869));
 b15tihi00an1n03x5 u_rxreg_counter_trgt_reg_7__1870 (.o(net1870));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_0__u_rxreg_data_int_reg_1__1871 (.o(net1871));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_10__u_rxreg_data_int_reg_11__1872 (.o(net1872));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_12__u_rxreg_data_int_reg_13__1873 (.o(net1873));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_14__u_rxreg_data_int_reg_15__1874 (.o(net1874));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_16__u_rxreg_data_int_reg_17__1875 (.o(net1875));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_18__u_rxreg_data_int_reg_19__1876 (.o(net1876));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_20__u_rxreg_data_int_reg_21__1877 (.o(net1877));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_22__u_rxreg_data_int_reg_23__1878 (.o(net1878));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_24__u_rxreg_data_int_reg_25__1879 (.o(net1879));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_26__u_rxreg_data_int_reg_27__1880 (.o(net1880));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_28__u_rxreg_data_int_reg_29__1881 (.o(net1881));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_2__u_rxreg_data_int_reg_3__1882 (.o(net1882));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_30__u_rxreg_data_int_reg_31__1883 (.o(net1883));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_4__u_rxreg_data_int_reg_5__1884 (.o(net1884));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_6__u_rxreg_data_int_reg_7__1885 (.o(net1885));
 b15tihi00an1n03x5 u_rxreg_data_int_reg_8__u_rxreg_data_int_reg_9__1886 (.o(net1886));
 b15tihi00an1n03x5 u_rxreg_running_reg_1887 (.o(net1887));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_0__u_spi_device_tlul_plug_addr_reg_1__1888 (.o(net1888));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_10__u_spi_device_tlul_plug_addr_reg_11__1889 (.o(net1889));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_12__u_spi_device_tlul_plug_addr_reg_13__1890 (.o(net1890));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_14__u_spi_device_tlul_plug_addr_reg_15__1891 (.o(net1891));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_16__u_spi_device_tlul_plug_addr_reg_17__1892 (.o(net1892));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_18__u_spi_device_tlul_plug_addr_reg_19__1893 (.o(net1893));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_20__u_spi_device_tlul_plug_addr_reg_21__1894 (.o(net1894));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_22__u_spi_device_tlul_plug_addr_reg_23__1895 (.o(net1895));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_24__u_spi_device_tlul_plug_addr_reg_25__1896 (.o(net1896));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_26__u_spi_device_tlul_plug_addr_reg_27__1897 (.o(net1897));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_28__u_spi_device_tlul_plug_addr_reg_29__1898 (.o(net1898));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_2__u_spi_device_tlul_plug_addr_reg_3__1899 (.o(net1899));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_30__u_spi_device_tlul_plug_addr_reg_31__1900 (.o(net1900));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_4__u_spi_device_tlul_plug_addr_reg_5__1901 (.o(net1901));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_6__u_spi_device_tlul_plug_addr_reg_7__1902 (.o(net1902));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_addr_reg_8__u_spi_device_tlul_plug_addr_reg_9__1903 (.o(net1903));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_state_reg_1__u_spi_device_tlul_plug_u_tlul_adapter_host_g_multiple_reqs_source_q_reg_0__1904 (.o(net1904));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_u_tlul_adapter_host_intg_err_q_reg_u_spi_device_tlul_plug_wdata_reg_0__1905 (.o(net1905));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_11__u_spi_device_tlul_plug_wdata_reg_12__1906 (.o(net1906));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_13__u_spi_device_tlul_plug_wdata_reg_14__1907 (.o(net1907));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_15__u_spi_device_tlul_plug_wdata_reg_16__1908 (.o(net1908));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_17__u_spi_device_tlul_plug_wdata_reg_18__1909 (.o(net1909));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_19__u_spi_device_tlul_plug_wdata_reg_20__1910 (.o(net1910));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_1__u_spi_device_tlul_plug_wdata_reg_2__1911 (.o(net1911));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_21__u_spi_device_tlul_plug_wdata_reg_22__1912 (.o(net1912));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_23__u_spi_device_tlul_plug_wdata_reg_24__1913 (.o(net1913));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_25__u_spi_device_tlul_plug_wdata_reg_26__1914 (.o(net1914));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_27__u_spi_device_tlul_plug_wdata_reg_28__1915 (.o(net1915));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_29__u_spi_device_tlul_plug_wdata_reg_30__1916 (.o(net1916));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_31__u_spi_device_tlul_plug_we_reg_1917 (.o(net1917));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_3__u_spi_device_tlul_plug_wdata_reg_4__1918 (.o(net1918));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_5__u_spi_device_tlul_plug_wdata_reg_6__1919 (.o(net1919));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_7__u_spi_device_tlul_plug_wdata_reg_8__1920 (.o(net1920));
 b15tihi00an1n03x5 u_spi_device_tlul_plug_wdata_reg_9__u_spi_device_tlul_plug_wdata_reg_10__1921 (.o(net1921));
 b15tihi00an1n03x5 u_syncro_cs_reg_reg_0__1922 (.o(net1922));
 b15tihi00an1n03x5 u_syncro_cs_reg_reg_1__1923 (.o(net1923));
 b15tihi00an1n03x5 u_syncro_rdwr_reg_reg_0__u_syncro_rdwr_reg_reg_1__1924 (.o(net1924));
 b15tihi00an1n03x5 u_syncro_valid_reg_reg_0__u_syncro_valid_reg_reg_1__1925 (.o(net1925));
 b15tihi00an1n03x5 u_syncro_valid_reg_reg_2__1926 (.o(net1926));
 b15tihi00an1n03x5 u_txreg_counter_reg_0__u_txreg_counter_reg_1__1927 (.o(net1927));
 b15tihi00an1n03x5 u_txreg_counter_reg_2__u_txreg_counter_reg_3__1928 (.o(net1928));
 b15tihi00an1n03x5 u_txreg_counter_reg_4__u_txreg_counter_reg_5__1929 (.o(net1929));
 b15tihi00an1n03x5 u_txreg_counter_reg_6__u_txreg_counter_reg_7__1930 (.o(net1930));
 b15tihi00an1n03x5 u_txreg_counter_trgt_reg_0__1931 (.o(net1931));
 b15tihi00an1n03x5 u_txreg_counter_trgt_reg_1__1932 (.o(net1932));
 b15tihi00an1n03x5 u_txreg_counter_trgt_reg_2__1933 (.o(net1933));
 b15tihi00an1n03x5 u_txreg_counter_trgt_reg_3__u_txreg_counter_trgt_reg_4__1934 (.o(net1934));
 b15tihi00an1n03x5 u_txreg_counter_trgt_reg_5__u_txreg_counter_trgt_reg_6__1935 (.o(net1935));
 b15tihi00an1n03x5 u_txreg_counter_trgt_reg_7__1936 (.o(net1936));
 b15tihi00an1n03x5 u_txreg_data_int_reg_0__u_txreg_data_int_reg_1__1937 (.o(net1937));
 b15tihi00an1n03x5 u_txreg_data_int_reg_10__u_txreg_data_int_reg_11__1938 (.o(net1938));
 b15tihi00an1n03x5 u_txreg_data_int_reg_12__u_txreg_data_int_reg_13__1939 (.o(net1939));
 b15tihi00an1n03x5 u_txreg_data_int_reg_14__u_txreg_data_int_reg_15__1940 (.o(net1940));
 b15tihi00an1n03x5 u_txreg_data_int_reg_16__u_txreg_data_int_reg_17__1941 (.o(net1941));
 b15tihi00an1n03x5 u_txreg_data_int_reg_18__u_txreg_data_int_reg_19__1942 (.o(net1942));
 b15tihi00an1n03x5 u_txreg_data_int_reg_20__u_txreg_data_int_reg_21__1943 (.o(net1943));
 b15tihi00an1n03x5 u_txreg_data_int_reg_22__u_txreg_data_int_reg_23__1944 (.o(net1944));
 b15tihi00an1n03x5 u_txreg_data_int_reg_24__u_txreg_data_int_reg_25__1945 (.o(net1945));
 b15tihi00an1n03x5 u_txreg_data_int_reg_26__u_txreg_data_int_reg_27__1946 (.o(net1946));
 b15tihi00an1n03x5 u_txreg_data_int_reg_28__u_txreg_data_int_reg_29__1947 (.o(net1947));
 b15tihi00an1n03x5 u_txreg_data_int_reg_2__u_txreg_data_int_reg_3__1948 (.o(net1948));
 b15tihi00an1n03x5 u_txreg_data_int_reg_30__u_txreg_data_int_reg_31__1949 (.o(net1949));
 b15tihi00an1n03x5 u_txreg_data_int_reg_4__u_txreg_data_int_reg_5__1950 (.o(net1950));
 b15tihi00an1n03x5 u_txreg_data_int_reg_6__u_txreg_data_int_reg_7__1951 (.o(net1951));
 b15tihi00an1n03x5 u_txreg_data_int_reg_8__u_txreg_data_int_reg_9__1952 (.o(net1952));
 b15tihi00an1n03x5 u_txreg_running_reg_1953 (.o(net1953));
 b15cbf000an1n16x5 clkbuf_2_0_0_clk_i (.clk(clknet_0_clk_i),
    .clkout(clknet_2_0_0_clk_i));
 b15cbf000an1n16x5 clkbuf_2_1_0_clk_i (.clk(clknet_0_clk_i),
    .clkout(clknet_2_1_0_clk_i));
 b15cbf000an1n16x5 clkbuf_2_2_0_clk_i (.clk(clknet_0_clk_i),
    .clkout(clknet_2_2_0_clk_i));
 b15cbf000an1n16x5 clkbuf_2_3_0_clk_i (.clk(clknet_0_clk_i),
    .clkout(clknet_2_3_0_clk_i));
 b15cbf000an1n16x5 clkbuf_0_u_spi_device_tlul_plug_net611 (.clk(u_spi_device_tlul_plug_net611),
    .clkout(clknet_0_u_spi_device_tlul_plug_net611));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_spi_device_tlul_plug_net611 (.clk(clknet_0_u_spi_device_tlul_plug_net611),
    .clkout(clknet_1_0__leaf_u_spi_device_tlul_plug_net611));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_spi_device_tlul_plug_net611 (.clk(clknet_0_u_spi_device_tlul_plug_net611),
    .clkout(clknet_1_1__leaf_u_spi_device_tlul_plug_net611));
 b15cbf000an1n16x5 clkbuf_0_u_spi_device_tlul_plug_net617 (.clk(u_spi_device_tlul_plug_net617),
    .clkout(clknet_0_u_spi_device_tlul_plug_net617));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_spi_device_tlul_plug_net617 (.clk(clknet_0_u_spi_device_tlul_plug_net617),
    .clkout(clknet_1_0__leaf_u_spi_device_tlul_plug_net617));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_spi_device_tlul_plug_net617 (.clk(clknet_0_u_spi_device_tlul_plug_net617),
    .clkout(clknet_1_1__leaf_u_spi_device_tlul_plug_net617));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_write_tr_net652 (.clk(u_dcfifo_tx_u_din_write_tr_net652),
    .clkout(clknet_0_u_dcfifo_tx_u_din_write_tr_net652));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_write_tr_net652 (.clk(clknet_0_u_dcfifo_tx_u_din_write_tr_net652),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_write_tr_net652));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_write_tr_net652 (.clk(clknet_0_u_dcfifo_tx_u_din_write_tr_net652),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_write_tr_net652));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net670 (.clk(u_dcfifo_tx_u_din_buffer_net670),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net670));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net670 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net670),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net670));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net670 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net670),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net670));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net676 (.clk(u_dcfifo_tx_u_din_buffer_net676),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net676));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net676 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net676),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net676));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net676 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net676),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net676));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net681 (.clk(u_dcfifo_tx_u_din_buffer_net681),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net681));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net681 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net681),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net681));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net681 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net681),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net681));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net686 (.clk(u_dcfifo_tx_u_din_buffer_net686),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net686));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net686 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net686),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net686));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net686 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net686),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net686));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net691 (.clk(u_dcfifo_tx_u_din_buffer_net691),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net691));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net691 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net691),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net691));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net691 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net691),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net691));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net696 (.clk(u_dcfifo_tx_u_din_buffer_net696),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net696));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net696 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net696),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net696));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net696 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net696),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net696));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net701 (.clk(u_dcfifo_tx_u_din_buffer_net701),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net701));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net701 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net701),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net701));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net701 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net701),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net701));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net706 (.clk(u_dcfifo_tx_u_din_buffer_net706),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net706));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net706 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net706),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net706));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net706 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net706),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net706));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net711 (.clk(u_dcfifo_tx_u_din_buffer_net711),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net711));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net711 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net711),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net711));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net711 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net711),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net711));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net716 (.clk(u_dcfifo_tx_u_din_buffer_net716),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net716));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net716 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net716),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net716));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net716 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net716),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net716));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net721 (.clk(u_dcfifo_tx_u_din_buffer_net721),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net721));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net721 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net721),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net721));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net721 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net721),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net721));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net726 (.clk(u_dcfifo_tx_u_din_buffer_net726),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net726));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net726 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net726),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net726));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net726 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net726),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net726));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net731 (.clk(u_dcfifo_tx_u_din_buffer_net731),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net731));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net731 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net731),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net731));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net731 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net731),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net731));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net736 (.clk(u_dcfifo_tx_u_din_buffer_net736),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net736));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net736 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net736),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net736));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net736 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net736),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net736));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net741 (.clk(u_dcfifo_tx_u_din_buffer_net741),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net741));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net741 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net741),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net741));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net741 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net741),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net741));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_din_buffer_net746 (.clk(u_dcfifo_tx_u_din_buffer_net746),
    .clkout(clknet_0_u_dcfifo_tx_u_din_buffer_net746));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_din_buffer_net746 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net746),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_din_buffer_net746));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_din_buffer_net746 (.clk(clknet_0_u_dcfifo_tx_u_din_buffer_net746),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_din_buffer_net746));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_dout_read_tr_net634 (.clk(u_dcfifo_rx_u_dout_read_tr_net634),
    .clkout(clknet_0_u_dcfifo_rx_u_dout_read_tr_net634));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_dout_read_tr_net634 (.clk(clknet_0_u_dcfifo_rx_u_dout_read_tr_net634),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_dout_read_tr_net634));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_dout_read_tr_net634 (.clk(clknet_0_u_dcfifo_rx_u_dout_read_tr_net634),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_dout_read_tr_net634));
 b15cbf000an1n16x5 clkbuf_0_spi_sclk (.clk(net1955),
    .clkout(clknet_0_spi_sclk));
 b15cbf000an1n16x5 clkbuf_2_0_0_spi_sclk (.clk(clknet_0_spi_sclk),
    .clkout(clknet_2_0_0_spi_sclk));
 b15cbf000an1n16x5 clkbuf_2_1_0_spi_sclk (.clk(clknet_0_spi_sclk),
    .clkout(clknet_2_1_0_spi_sclk));
 b15cbf000an1n16x5 clkbuf_2_2_0_spi_sclk (.clk(clknet_0_spi_sclk),
    .clkout(clknet_2_2_0_spi_sclk));
 b15cbf000an1n16x5 clkbuf_2_3_0_spi_sclk (.clk(clknet_0_spi_sclk),
    .clkout(clknet_2_3_0_spi_sclk));
 b15cbf000an1n16x5 clkbuf_3_0__f_spi_sclk (.clk(clknet_2_0_0_spi_sclk),
    .clkout(clknet_3_0__leaf_spi_sclk));
 b15cbf000an1n16x5 clkbuf_3_1__f_spi_sclk (.clk(clknet_2_0_0_spi_sclk),
    .clkout(clknet_3_1__leaf_spi_sclk));
 b15cbf000an1n16x5 clkbuf_3_2__f_spi_sclk (.clk(clknet_2_1_0_spi_sclk),
    .clkout(clknet_3_2__leaf_spi_sclk));
 b15cbf000an1n16x5 clkbuf_3_3__f_spi_sclk (.clk(clknet_2_1_0_spi_sclk),
    .clkout(clknet_3_3__leaf_spi_sclk));
 b15cbf000an1n16x5 clkbuf_3_4__f_spi_sclk (.clk(clknet_2_2_0_spi_sclk),
    .clkout(clknet_3_4__leaf_spi_sclk));
 b15cbf000an1n16x5 clkbuf_3_5__f_spi_sclk (.clk(clknet_2_2_0_spi_sclk),
    .clkout(clknet_3_5__leaf_spi_sclk));
 b15cbf000an1n16x5 clkbuf_3_6__f_spi_sclk (.clk(clknet_2_3_0_spi_sclk),
    .clkout(clknet_3_6__leaf_spi_sclk));
 b15cbf000an1n16x5 clkbuf_3_7__f_spi_sclk (.clk(clknet_2_3_0_spi_sclk),
    .clkout(clknet_3_7__leaf_spi_sclk));
 b15cbf000an1n16x5 clkbuf_0_u_txreg_sclk_test (.clk(u_txreg_sclk_test),
    .clkout(clknet_0_u_txreg_sclk_test));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_txreg_sclk_test (.clk(clknet_0_u_txreg_sclk_test),
    .clkout(clknet_1_0__leaf_u_txreg_sclk_test));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_txreg_sclk_test (.clk(clknet_0_u_txreg_sclk_test),
    .clkout(clknet_1_1__leaf_u_txreg_sclk_test));
 b15cbf000an1n16x5 clkbuf_0_u_txreg_net830 (.clk(u_txreg_net830),
    .clkout(clknet_0_u_txreg_net830));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_txreg_net830 (.clk(clknet_0_u_txreg_net830),
    .clkout(clknet_1_0__leaf_u_txreg_net830));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_txreg_net830 (.clk(clknet_0_u_txreg_net830),
    .clkout(clknet_1_1__leaf_u_txreg_net830));
 b15cbf000an1n16x5 clkbuf_0_u_txreg_net835 (.clk(u_txreg_net835),
    .clkout(clknet_0_u_txreg_net835));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_txreg_net835 (.clk(clknet_0_u_txreg_net835),
    .clkout(clknet_1_0__leaf_u_txreg_net835));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_txreg_net835 (.clk(clknet_0_u_txreg_net835),
    .clkout(clknet_1_1__leaf_u_txreg_net835));
 b15cbf000an1n16x5 clkbuf_0_u_txreg_net840 (.clk(u_txreg_net840),
    .clkout(clknet_0_u_txreg_net840));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_txreg_net840 (.clk(clknet_0_u_txreg_net840),
    .clkout(clknet_1_0__leaf_u_txreg_net840));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_txreg_net840 (.clk(clknet_0_u_txreg_net840),
    .clkout(clknet_1_1__leaf_u_txreg_net840));
 b15cbf000an1n16x5 clkbuf_0_u_txreg_net824 (.clk(u_txreg_net824),
    .clkout(clknet_0_u_txreg_net824));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_txreg_net824 (.clk(clknet_0_u_txreg_net824),
    .clkout(clknet_1_0__leaf_u_txreg_net824));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_txreg_net824 (.clk(clknet_0_u_txreg_net824),
    .clkout(clknet_1_1__leaf_u_txreg_net824));
 b15cbf000an1n16x5 clkbuf_0_u_rxreg_net863 (.clk(u_rxreg_net863),
    .clkout(clknet_0_u_rxreg_net863));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_rxreg_net863 (.clk(clknet_0_u_rxreg_net863),
    .clkout(clknet_1_0__leaf_u_rxreg_net863));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_rxreg_net863 (.clk(clknet_0_u_rxreg_net863),
    .clkout(clknet_1_1__leaf_u_rxreg_net863));
 b15cbf000an1n16x5 clkbuf_0_u_rxreg_net868 (.clk(u_rxreg_net868),
    .clkout(clknet_0_u_rxreg_net868));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_rxreg_net868 (.clk(clknet_0_u_rxreg_net868),
    .clkout(clknet_1_0__leaf_u_rxreg_net868));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_rxreg_net868 (.clk(clknet_0_u_rxreg_net868),
    .clkout(clknet_1_1__leaf_u_rxreg_net868));
 b15cbf000an1n16x5 clkbuf_0_u_rxreg_net873 (.clk(u_rxreg_net873),
    .clkout(clknet_0_u_rxreg_net873));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_rxreg_net873 (.clk(clknet_0_u_rxreg_net873),
    .clkout(clknet_1_0__leaf_u_rxreg_net873));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_rxreg_net873 (.clk(clknet_0_u_rxreg_net873),
    .clkout(clknet_1_1__leaf_u_rxreg_net873));
 b15cbf000an1n16x5 clkbuf_0_u_rxreg_net857 (.clk(u_rxreg_net857),
    .clkout(clknet_0_u_rxreg_net857));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_rxreg_net857 (.clk(clknet_0_u_rxreg_net857),
    .clkout(clknet_1_0__leaf_u_rxreg_net857));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_rxreg_net857 (.clk(clknet_0_u_rxreg_net857),
    .clkout(clknet_1_1__leaf_u_rxreg_net857));
 b15cbf000an1n16x5 clkbuf_0_u_device_sm_u_spiregs_net791 (.clk(u_device_sm_u_spiregs_net791),
    .clkout(clknet_0_u_device_sm_u_spiregs_net791));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_device_sm_u_spiregs_net791 (.clk(clknet_0_u_device_sm_u_spiregs_net791),
    .clkout(clknet_1_0__leaf_u_device_sm_u_spiregs_net791));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_device_sm_u_spiregs_net791 (.clk(clknet_0_u_device_sm_u_spiregs_net791),
    .clkout(clknet_1_1__leaf_u_device_sm_u_spiregs_net791));
 b15cbf000an1n16x5 clkbuf_0_u_device_sm_u_spiregs_net807 (.clk(u_device_sm_u_spiregs_net807),
    .clkout(clknet_0_u_device_sm_u_spiregs_net807));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_device_sm_u_spiregs_net807 (.clk(clknet_0_u_device_sm_u_spiregs_net807),
    .clkout(clknet_1_0__leaf_u_device_sm_u_spiregs_net807));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_device_sm_u_spiregs_net807 (.clk(clknet_0_u_device_sm_u_spiregs_net807),
    .clkout(clknet_1_1__leaf_u_device_sm_u_spiregs_net807));
 b15cbf000an1n16x5 clkbuf_0_u_device_sm_u_spiregs_net802 (.clk(u_device_sm_u_spiregs_net802),
    .clkout(clknet_0_u_device_sm_u_spiregs_net802));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_device_sm_u_spiregs_net802 (.clk(clknet_0_u_device_sm_u_spiregs_net802),
    .clkout(clknet_1_0__leaf_u_device_sm_u_spiregs_net802));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_device_sm_u_spiregs_net802 (.clk(clknet_0_u_device_sm_u_spiregs_net802),
    .clkout(clknet_1_1__leaf_u_device_sm_u_spiregs_net802));
 b15cbf000an1n16x5 clkbuf_0_u_device_sm_u_spiregs_net797 (.clk(u_device_sm_u_spiregs_net797),
    .clkout(clknet_0_u_device_sm_u_spiregs_net797));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_device_sm_u_spiregs_net797 (.clk(clknet_0_u_device_sm_u_spiregs_net797),
    .clkout(clknet_1_0__leaf_u_device_sm_u_spiregs_net797));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_device_sm_u_spiregs_net797 (.clk(clknet_0_u_device_sm_u_spiregs_net797),
    .clkout(clknet_1_1__leaf_u_device_sm_u_spiregs_net797));
 b15cbf000an1n16x5 clkbuf_0_u_device_sm_net774 (.clk(u_device_sm_net774),
    .clkout(clknet_0_u_device_sm_net774));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_device_sm_net774 (.clk(clknet_0_u_device_sm_net774),
    .clkout(clknet_1_0__leaf_u_device_sm_net774));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_device_sm_net774 (.clk(clknet_0_u_device_sm_net774),
    .clkout(clknet_1_1__leaf_u_device_sm_net774));
 b15cbf000an1n16x5 clkbuf_0_u_device_sm_net763 (.clk(u_device_sm_net763),
    .clkout(clknet_0_u_device_sm_net763));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_device_sm_net763 (.clk(clknet_0_u_device_sm_net763),
    .clkout(clknet_1_0__leaf_u_device_sm_net763));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_device_sm_net763 (.clk(clknet_0_u_device_sm_net763),
    .clkout(clknet_1_1__leaf_u_device_sm_net763));
 b15cbf000an1n16x5 clkbuf_0_u_device_sm_net769 (.clk(u_device_sm_net769),
    .clkout(clknet_0_u_device_sm_net769));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_device_sm_net769 (.clk(clknet_0_u_device_sm_net769),
    .clkout(clknet_1_0__leaf_u_device_sm_net769));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_device_sm_net769 (.clk(clknet_0_u_device_sm_net769),
    .clkout(clknet_1_1__leaf_u_device_sm_net769));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_tx_u_dout_read_tr_net634 (.clk(u_dcfifo_tx_u_dout_read_tr_net634),
    .clkout(clknet_0_u_dcfifo_tx_u_dout_read_tr_net634));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_tx_u_dout_read_tr_net634 (.clk(clknet_0_u_dcfifo_tx_u_dout_read_tr_net634),
    .clkout(clknet_1_0__leaf_u_dcfifo_tx_u_dout_read_tr_net634));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_tx_u_dout_read_tr_net634 (.clk(clknet_0_u_dcfifo_tx_u_dout_read_tr_net634),
    .clkout(clknet_1_1__leaf_u_dcfifo_tx_u_dout_read_tr_net634));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_write_tr_net652 (.clk(u_dcfifo_rx_u_din_write_tr_net652),
    .clkout(clknet_0_u_dcfifo_rx_u_din_write_tr_net652));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_write_tr_net652 (.clk(clknet_0_u_dcfifo_rx_u_din_write_tr_net652),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_write_tr_net652));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_write_tr_net652 (.clk(clknet_0_u_dcfifo_rx_u_din_write_tr_net652),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_write_tr_net652));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net670 (.clk(u_dcfifo_rx_u_din_buffer_net670),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net670));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net670 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net670),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net670));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net670 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net670),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net670));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net676 (.clk(u_dcfifo_rx_u_din_buffer_net676),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net676));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net676 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net676),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net676));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net676 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net676),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net676));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net681 (.clk(u_dcfifo_rx_u_din_buffer_net681),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net681));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net681 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net681),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net681));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net681 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net681),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net681));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net686 (.clk(u_dcfifo_rx_u_din_buffer_net686),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net686));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net686 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net686),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net686));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net686 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net686),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net686));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net691 (.clk(u_dcfifo_rx_u_din_buffer_net691),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net691));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net691 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net691),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net691));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net691 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net691),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net691));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net696 (.clk(u_dcfifo_rx_u_din_buffer_net696),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net696));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net696 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net696),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net696));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net696 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net696),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net696));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net701 (.clk(u_dcfifo_rx_u_din_buffer_net701),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net701));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net701 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net701),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net701));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net701 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net701),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net701));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net706 (.clk(u_dcfifo_rx_u_din_buffer_net706),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net706));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net706 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net706),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net706));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net706 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net706),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net706));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net711 (.clk(u_dcfifo_rx_u_din_buffer_net711),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net711));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net711 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net711),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net711));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net711 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net711),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net711));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net716 (.clk(u_dcfifo_rx_u_din_buffer_net716),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net716));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net716 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net716),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net716));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net716 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net716),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net716));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net721 (.clk(u_dcfifo_rx_u_din_buffer_net721),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net721));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net721 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net721),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net721));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net721 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net721),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net721));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net726 (.clk(u_dcfifo_rx_u_din_buffer_net726),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net726));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net726 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net726),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net726));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net726 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net726),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net726));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net731 (.clk(u_dcfifo_rx_u_din_buffer_net731),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net731));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net731 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net731),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net731));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net731 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net731),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net731));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net736 (.clk(u_dcfifo_rx_u_din_buffer_net736),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net736));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net736 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net736),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net736));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net736 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net736),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net736));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net741 (.clk(u_dcfifo_rx_u_din_buffer_net741),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net741));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net741 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net741),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net741));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net741 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net741),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net741));
 b15cbf000an1n16x5 clkbuf_0_u_dcfifo_rx_u_din_buffer_net746 (.clk(u_dcfifo_rx_u_din_buffer_net746),
    .clkout(clknet_0_u_dcfifo_rx_u_din_buffer_net746));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_dcfifo_rx_u_din_buffer_net746 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net746),
    .clkout(clknet_1_0__leaf_u_dcfifo_rx_u_din_buffer_net746));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_dcfifo_rx_u_din_buffer_net746 (.clk(clknet_0_u_dcfifo_rx_u_din_buffer_net746),
    .clkout(clknet_1_1__leaf_u_dcfifo_rx_u_din_buffer_net746));
 b15bfn001as1n16x5 wire2 (.a(spi_sclk),
    .o(net1955));
 b15cbf034ar1n64x5 hold3 (.clk(net2373),
    .clkout(net1956));
 b15cbf034ar1n64x5 hold4 (.clk(net2375),
    .clkout(tl_o[29]));
 b15cbf034ar1n64x5 hold5 (.clk(net2376),
    .clkout(net1958));
 b15cbf034ar1n64x5 hold6 (.clk(net2378),
    .clkout(tl_o[38]));
 b15cbf034ar1n64x5 hold7 (.clk(net2379),
    .clkout(net1960));
 b15cbf034ar1n64x5 hold8 (.clk(net2381),
    .clkout(tl_o[37]));
 b15cbf034ar1n64x5 hold9 (.clk(net2382),
    .clkout(net1962));
 b15cbf034ar1n64x5 hold10 (.clk(net2384),
    .clkout(tl_o[30]));
 b15cbf034ar1n64x5 hold11 (.clk(net2477),
    .clkout(net1964));
 b15cbf034ar1n64x5 hold12 (.clk(net341),
    .clkout(net1965));
 b15cbf034ar1n64x5 hold13 (.clk(net1966),
    .clkout(tl_o[51]));
 b15cbf034ar1n64x5 hold14 (.clk(net2385),
    .clkout(net1967));
 b15cbf034ar1n64x5 hold15 (.clk(net2387),
    .clkout(tl_o[47]));
 b15cbf034ar1n64x5 hold16 (.clk(net2388),
    .clkout(net1969));
 b15cbf034ar1n64x5 hold17 (.clk(net2390),
    .clkout(tl_o[48]));
 b15cbf034ar1n64x5 hold18 (.clk(net2391),
    .clkout(net1971));
 b15cbf034ar1n64x5 hold19 (.clk(net2393),
    .clkout(tl_o[50]));
 b15cbf034ar1n64x5 hold20 (.clk(net2394),
    .clkout(net1973));
 b15cbf034ar1n64x5 hold21 (.clk(net2396),
    .clkout(tl_o[49]));
 b15cbf034ar1n64x5 hold22 (.clk(net2347),
    .clkout(net1975));
 b15cbf034ar1n64x5 hold23 (.clk(net2466),
    .clkout(net1976));
 b15cbf034ar1n64x5 hold24 (.clk(net1977),
    .clkout(tl_o[108]));
 b15cbf034ar1n64x5 hold25 (.clk(net2400),
    .clkout(net1978));
 b15cbf034ar1n64x5 hold26 (.clk(net2402),
    .clkout(tl_o[36]));
 b15cbf034ar1n64x5 hold27 (.clk(net2456),
    .clkout(net1980));
 b15cbf034ar1n64x5 hold28 (.clk(net1981),
    .clkout(tl_o[92]));
 b15cbf034ar1n64x5 hold29 (.clk(net2403),
    .clkout(net1982));
 b15cbf034ar1n64x5 hold30 (.clk(net2405),
    .clkout(tl_o[35]));
 b15cbf034ar1n64x5 hold31 (.clk(net2397),
    .clkout(net1984));
 b15cbf034ar1n64x5 hold32 (.clk(net2399),
    .clkout(tl_o[34]));
 b15cbf034ar1n64x5 hold33 (.clk(net2495),
    .clkout(net1986));
 b15cbf034ar1n64x5 hold34 (.clk(net343),
    .clkout(net1987));
 b15cbf034ar1n64x5 hold35 (.clk(net1988),
    .clkout(tl_o[45]));
 b15cbf034ar1n64x5 hold36 (.clk(net2406),
    .clkout(net1989));
 b15cbf034ar1n64x5 hold37 (.clk(net2408),
    .clkout(tl_o[33]));
 b15cbf034ar1n64x5 hold38 (.clk(net2496),
    .clkout(net1991));
 b15cbf034ar1n64x5 hold39 (.clk(net342),
    .clkout(net1992));
 b15cbf034ar1n64x5 hold40 (.clk(net1993),
    .clkout(tl_o[46]));
 b15cbf034ar1n64x5 hold41 (.clk(net2409),
    .clkout(net1994));
 b15cbf034ar1n64x5 hold42 (.clk(net2411),
    .clkout(tl_o[43]));
 b15cbf034ar1n64x5 hold43 (.clk(net2412),
    .clkout(net1996));
 b15cbf034ar1n64x5 hold44 (.clk(net2414),
    .clkout(tl_o[44]));
 b15cbf034ar1n64x5 hold45 (.clk(net2415),
    .clkout(net1998));
 b15cbf034ar1n64x5 hold46 (.clk(net2417),
    .clkout(tl_o[32]));
 b15cbf034ar1n64x5 hold47 (.clk(net2418),
    .clkout(net2000));
 b15cbf034ar1n64x5 hold48 (.clk(net2420),
    .clkout(tl_o[31]));
 b15cbf034ar1n64x5 hold49 (.clk(net2421),
    .clkout(net2002));
 b15cbf034ar1n64x5 hold50 (.clk(net2423),
    .clkout(tl_o[39]));
 b15cbf034ar1n64x5 hold51 (.clk(net2424),
    .clkout(net2004));
 b15cbf034ar1n64x5 hold52 (.clk(net2426),
    .clkout(tl_o[40]));
 b15cbf034ar1n64x5 hold53 (.clk(net2433),
    .clkout(net2006));
 b15cbf034ar1n64x5 hold54 (.clk(net2435),
    .clkout(tl_o[24]));
 b15cbf034ar1n64x5 hold55 (.clk(net2430),
    .clkout(net2008));
 b15cbf034ar1n64x5 hold56 (.clk(net2432),
    .clkout(tl_o[27]));
 b15cbf034ar1n64x5 hold57 (.clk(net2427),
    .clkout(net2010));
 b15cbf034ar1n64x5 hold58 (.clk(net2429),
    .clkout(tl_o[28]));
 b15cbf034ar1n64x5 hold59 (.clk(u_spi_device_tlul_plug_we),
    .clkout(net2012));
 b15cbf034ar1n64x5 hold60 (.clk(net340),
    .clkout(net2013));
 b15cbf034ar1n64x5 hold61 (.clk(net61),
    .clkout(net2014));
 b15cbf034ar1n64x5 hold62 (.clk(net2015),
    .clkout(tl_o[107]));
 b15cbf034ar1n64x5 hold63 (.clk(net2441),
    .clkout(net2016));
 b15cbf034ar1n64x5 hold64 (.clk(net2017),
    .clkout(tl_o[41]));
 b15cbf034ar1n64x5 hold65 (.clk(net2439),
    .clkout(net2018));
 b15cbf034ar1n64x5 hold66 (.clk(net2019),
    .clkout(tl_o[42]));
 b15cbf034ar1n64x5 hold67 (.clk(net2508),
    .clkout(net2020));
 b15cbf034ar1n64x5 hold68 (.clk(net280),
    .clkout(net2021));
 b15cbf034ar1n64x5 hold69 (.clk(net2022),
    .clkout(tl_o[82]));
 b15cbf034ar1n64x5 hold70 (.clk(net2443),
    .clkout(net2023));
 b15cbf034ar1n64x5 hold71 (.clk(net2024),
    .clkout(tl_o[55]));
 b15cbf034ar1n64x5 hold72 (.clk(net2467),
    .clkout(net2025));
 b15cbf034ar1n64x5 hold73 (.clk(net2026),
    .clkout(tl_o[80]));
 b15cbf034ar1n64x5 hold74 (.clk(net2436),
    .clkout(net2027));
 b15cbf034ar1n64x5 hold75 (.clk(net2438),
    .clkout(tl_o[54]));
 b15cbf034ar1n64x5 hold76 (.clk(net2454),
    .clkout(net2029));
 b15cbf034ar1n64x5 hold77 (.clk(net2030),
    .clkout(tl_o[91]));
 b15cbf034ar1n64x5 hold78 (.clk(net2447),
    .clkout(net2031));
 b15cbf034ar1n64x5 hold79 (.clk(net2032),
    .clkout(tl_o[25]));
 b15cbf034ar1n64x5 hold80 (.clk(net2449),
    .clkout(net2033));
 b15cbf034ar1n64x5 hold81 (.clk(net2034),
    .clkout(tl_o[26]));
 b15cbf034ar1n64x5 hold82 (.clk(net119),
    .clkout(net2035));
 b15cbf034ar1n64x5 hold83 (.clk(net282),
    .clkout(net2036));
 b15cbf034ar1n64x5 hold84 (.clk(net281),
    .clkout(net2037));
 b15cbf034ar1n64x5 hold85 (.clk(net2038),
    .clkout(tl_o[81]));
 b15cbf034ar1n64x5 hold86 (.clk(net2451),
    .clkout(net2039));
 b15cbf034ar1n64x5 hold87 (.clk(net2453),
    .clkout(tl_o[53]));
 b15cbf034ar1n64x5 hold88 (.clk(net2469),
    .clkout(net2041));
 b15cbf034ar1n64x5 hold89 (.clk(net2042),
    .clkout(tl_o[83]));
 b15cbf034ar1n64x5 hold90 (.clk(net2511),
    .clkout(net2043));
 b15cbf034ar1n64x5 hold91 (.clk(net266),
    .clkout(net2044));
 b15cbf034ar1n64x5 hold92 (.clk(net2045),
    .clkout(tl_o[69]));
 b15cbf034ar1n64x5 hold93 (.clk(net2473),
    .clkout(net2046));
 b15cbf034ar1n64x5 hold94 (.clk(net2047),
    .clkout(tl_o[62]));
 b15cbf034ar1n64x5 hold95 (.clk(net2509),
    .clkout(net2048));
 b15cbf034ar1n64x5 hold96 (.clk(net289),
    .clkout(net2049));
 b15cbf034ar1n64x5 hold97 (.clk(net2050),
    .clkout(tl_o[76]));
 b15cbf034ar1n64x5 hold98 (.clk(net2462),
    .clkout(net2051));
 b15cbf034ar1n64x5 hold99 (.clk(net2052),
    .clkout(tl_o[52]));
 b15cbf034ar1n64x5 hold100 (.clk(net2475),
    .clkout(net2053));
 b15cbf034ar1n64x5 hold101 (.clk(net2054),
    .clkout(tl_o[71]));
 b15cbf034ar1n64x5 hold102 (.clk(net2458),
    .clkout(net2055));
 b15cbf034ar1n64x5 hold103 (.clk(net2056),
    .clkout(tl_o[84]));
 b15cbf034ar1n64x5 hold104 (.clk(net2460),
    .clkout(net2057));
 b15cbf034ar1n64x5 hold105 (.clk(net2058),
    .clkout(tl_o[89]));
 b15cbf034ar1n64x5 hold106 (.clk(net2066),
    .clkout(net2059));
 b15cbf034ar1n64x5 hold107 (.clk(net287),
    .clkout(net2060));
 b15cbf034ar1n64x5 hold108 (.clk(n3590),
    .clkout(net2061));
 b15cbf034ar1n64x5 hold109 (.clk(n3577),
    .clkout(net2062));
 b15cbf034ar1n64x5 hold110 (.clk(n3579),
    .clkout(net2063));
 b15cbf034ar1n64x5 hold111 (.clk(net63),
    .clkout(net2064));
 b15cbf034ar1n64x5 hold112 (.clk(net2065),
    .clkout(tl_o[10]));
 b15cbf034ar1n64x5 hold113 (.clk(net116),
    .clkout(net2066));
 b15cbf034ar1n64x5 hold114 (.clk(net2059),
    .clkout(net2067));
 b15cbf034ar1n64x5 hold115 (.clk(net2158),
    .clkout(net2068));
 b15cbf034ar1n64x5 hold116 (.clk(net276),
    .clkout(net2069));
 b15cbf034ar1n64x5 hold117 (.clk(net2070),
    .clkout(tl_o[85]));
 b15cbf034ar1n64x5 hold118 (.clk(net2100),
    .clkout(net2071));
 b15cbf034ar1n64x5 hold119 (.clk(n3562),
    .clkout(net2072));
 b15cbf034ar1n64x5 hold120 (.clk(n3327),
    .clkout(net2073));
 b15cbf034ar1n64x5 hold121 (.clk(net66),
    .clkout(net2074));
 b15cbf034ar1n64x5 hold122 (.clk(net2075),
    .clkout(tl_o[13]));
 b15cbf034ar1n64x5 hold123 (.clk(u_device_sm_state[0]),
    .clkout(net2076));
 b15cbf034ar1n64x5 hold124 (.clk(net358),
    .clkout(net2077));
 b15cbf034ar1n64x5 hold125 (.clk(net357),
    .clkout(net2078));
 b15cbf034ar1n64x5 hold126 (.clk(n3619),
    .clkout(net2079));
 b15cbf034ar1n64x5 hold127 (.clk(net55),
    .clkout(net2080));
 b15cbf034ar1n64x5 hold128 (.clk(net2081),
    .clkout(spi_mode[0]));
 b15cbf034ar1n64x5 hold129 (.clk(net2483),
    .clkout(net2082));
 b15cbf034ar1n64x5 hold130 (.clk(net2083),
    .clkout(tl_o[68]));
 b15cbf034ar1n64x5 hold131 (.clk(net2127),
    .clkout(net2084));
 b15cbf034ar1n64x5 hold132 (.clk(net2085),
    .clkout(tl_o[66]));
 b15cbf034ar1n64x5 hold133 (.clk(net2445),
    .clkout(net2086));
 b15cbf034ar1n64x5 hold134 (.clk(u_device_sm_state[1]),
    .clkout(net2087));
 b15cbf034ar1n64x5 hold135 (.clk(net360),
    .clkout(net2088));
 b15cbf034ar1n64x5 hold136 (.clk(net359),
    .clkout(net2089));
 b15cbf034ar1n64x5 hold137 (.clk(n2842),
    .clkout(net2090));
 b15cbf034ar1n64x5 hold138 (.clk(n2860),
    .clkout(net2091));
 b15cbf034ar1n64x5 hold139 (.clk(net56),
    .clkout(net2092));
 b15cbf034ar1n64x5 hold140 (.clk(net2093),
    .clkout(spi_mode[1]));
 b15cbf034ar1n64x5 hold141 (.clk(net2097),
    .clkout(net2094));
 b15cbf034ar1n64x5 hold142 (.clk(net65),
    .clkout(net2095));
 b15cbf034ar1n64x5 hold143 (.clk(net2096),
    .clkout(tl_o[12]));
 b15cbf034ar1n64x5 hold144 (.clk(net126),
    .clkout(net2097));
 b15cbf034ar1n64x5 hold145 (.clk(net2094),
    .clkout(net2098));
 b15cbf034ar1n64x5 hold146 (.clk(net2099),
    .clkout(tl_o[88]));
 b15cbf034ar1n64x5 hold147 (.clk(net108),
    .clkout(net2100));
 b15cbf034ar1n64x5 hold148 (.clk(net2071),
    .clkout(net2101));
 b15cbf034ar1n64x5 hold149 (.clk(net2102),
    .clkout(tl_o[70]));
 b15cbf034ar1n64x5 hold150 (.clk(net2510),
    .clkout(net2103));
 b15cbf034ar1n64x5 hold151 (.clk(net272),
    .clkout(net2104));
 b15cbf034ar1n64x5 hold152 (.clk(net2105),
    .clkout(tl_o[63]));
 b15cbf034ar1n64x5 hold153 (.clk(net2136),
    .clkout(net2106));
 b15cbf034ar1n64x5 hold154 (.clk(net2107),
    .clkout(tl_o[74]));
 b15cbf034ar1n64x5 hold155 (.clk(net2110),
    .clkout(net2108));
 b15cbf034ar1n64x5 hold156 (.clk(net2109),
    .clkout(tl_o[90]));
 b15cbf034ar1n64x5 hold157 (.clk(net129),
    .clkout(net2110));
 b15cbf034ar1n64x5 hold158 (.clk(net2108),
    .clkout(net2111));
 b15cbf034ar1n64x5 hold159 (.clk(net128),
    .clkout(net2112));
 b15cbf034ar1n64x5 hold160 (.clk(net2113),
    .clkout(tl_o[8]));
 b15cbf034ar1n64x5 hold161 (.clk(net2487),
    .clkout(net2114));
 b15cbf034ar1n64x5 hold162 (.clk(net2115),
    .clkout(tl_o[73]));
 b15cbf034ar1n64x5 hold163 (.clk(net2497),
    .clkout(net2116));
 b15cbf034ar1n64x5 hold164 (.clk(net2117),
    .clkout(tl_o[75]));
 b15cbf034ar1n64x5 hold165 (.clk(net2498),
    .clkout(net2118));
 b15cbf034ar1n64x5 hold166 (.clk(net2119),
    .clkout(tl_o[67]));
 b15cbf034ar1n64x5 hold167 (.clk(net2502),
    .clkout(net2120));
 b15cbf034ar1n64x5 hold168 (.clk(net2121),
    .clkout(tl_o[87]));
 b15cbf034ar1n64x5 hold169 (.clk(net2516),
    .clkout(net2122));
 b15cbf034ar1n64x5 hold170 (.clk(net270),
    .clkout(net2123));
 b15cbf034ar1n64x5 hold171 (.clk(net2124),
    .clkout(tl_o[64]));
 b15cbf034ar1n64x5 hold172 (.clk(net2471),
    .clkout(net2125));
 b15cbf034ar1n64x5 hold173 (.clk(net2126),
    .clkout(tl_o[86]));
 b15cbf034ar1n64x5 hold174 (.clk(net104),
    .clkout(net2127));
 b15cbf034ar1n64x5 hold175 (.clk(net2084),
    .clkout(net2128));
 b15cbf034ar1n64x5 hold176 (.clk(n3343),
    .clkout(net2129));
 b15cbf034ar1n64x5 hold177 (.clk(net67),
    .clkout(net2130));
 b15cbf034ar1n64x5 hold178 (.clk(net2131),
    .clkout(tl_o[14]));
 b15cbf034ar1n64x5 hold179 (.clk(net2504),
    .clkout(net2132));
 b15cbf034ar1n64x5 hold180 (.clk(net2133),
    .clkout(tl_o[77]));
 b15cbf034ar1n64x5 hold181 (.clk(net2507),
    .clkout(net2134));
 b15cbf034ar1n64x5 hold182 (.clk(net2135),
    .clkout(tl_o[79]));
 b15cbf034ar1n64x5 hold183 (.clk(net112),
    .clkout(net2136));
 b15cbf034ar1n64x5 hold184 (.clk(net2106),
    .clkout(net2137));
 b15cbf034ar1n64x5 hold185 (.clk(n3605),
    .clkout(net2138));
 b15cbf034ar1n64x5 hold186 (.clk(net132),
    .clkout(net2139));
 b15cbf034ar1n64x5 hold187 (.clk(net2140),
    .clkout(tl_o[9]));
 b15cbf034ar1n64x5 hold188 (.clk(tx_data[19]),
    .clkout(net2141));
 b15cbf034ar1n64x5 hold189 (.clk(n2928),
    .clkout(net2142));
 b15cbf034ar1n64x5 hold190 (.clk(u_txreg_N53),
    .clkout(net2143));
 b15cbf034ar1n64x5 hold191 (.clk(tx_data[24]),
    .clkout(net2144));
 b15cbf034ar1n64x5 hold192 (.clk(n2945),
    .clkout(net2145));
 b15cbf034ar1n64x5 hold193 (.clk(u_txreg_N58),
    .clkout(net2146));
 b15cbf034ar1n64x5 hold194 (.clk(net2501),
    .clkout(net2147));
 b15cbf034ar1n64x5 hold195 (.clk(net2148),
    .clkout(tl_o[72]));
 b15cbf034ar1n64x5 hold196 (.clk(net103),
    .clkout(net2149));
 b15cbf034ar1n64x5 hold197 (.clk(net269),
    .clkout(net2150));
 b15cbf034ar1n64x5 hold198 (.clk(net268),
    .clkout(net2151));
 b15cbf034ar1n64x5 hold199 (.clk(tx_data[16]),
    .clkout(net2152));
 b15cbf034ar1n64x5 hold200 (.clk(n2940),
    .clkout(net2153));
 b15cbf034ar1n64x5 hold201 (.clk(u_txreg_N50),
    .clkout(net2154));
 b15cbf034ar1n64x5 hold202 (.clk(tx_data[18]),
    .clkout(net2155));
 b15cbf034ar1n64x5 hold203 (.clk(n2938),
    .clkout(net2156));
 b15cbf034ar1n64x5 hold204 (.clk(u_txreg_N52),
    .clkout(net2157));
 b15cbf034ar1n64x5 hold205 (.clk(net123),
    .clkout(net2158));
 b15cbf034ar1n64x5 hold206 (.clk(net2068),
    .clkout(net2159));
 b15cbf034ar1n64x5 hold207 (.clk(n3608),
    .clkout(net2160));
 b15cbf034ar1n64x5 hold208 (.clk(net64),
    .clkout(net2161));
 b15cbf034ar1n64x5 hold209 (.clk(net2162),
    .clkout(tl_o[11]));
 b15cbf034ar1n64x5 hold210 (.clk(tx_data[25]),
    .clkout(net2163));
 b15cbf034ar1n64x5 hold211 (.clk(n2920),
    .clkout(net2164));
 b15cbf034ar1n64x5 hold212 (.clk(u_txreg_N59),
    .clkout(net2165));
 b15cbf034ar1n64x5 hold213 (.clk(tx_data[27]),
    .clkout(net2166));
 b15cbf034ar1n64x5 hold214 (.clk(n2922),
    .clkout(net2167));
 b15cbf034ar1n64x5 hold215 (.clk(u_txreg_N61),
    .clkout(net2168));
 b15cbf034ar1n64x5 hold216 (.clk(net2481),
    .clkout(net2169));
 b15cbf034ar1n64x5 hold217 (.clk(tx_data[20]),
    .clkout(net2170));
 b15cbf034ar1n64x5 hold218 (.clk(n2927),
    .clkout(net2171));
 b15cbf034ar1n64x5 hold219 (.clk(u_txreg_N54),
    .clkout(net2172));
 b15cbf034ar1n64x5 hold220 (.clk(tx_data[11]),
    .clkout(net2173));
 b15cbf034ar1n64x5 hold221 (.clk(n2939),
    .clkout(net2174));
 b15cbf034ar1n64x5 hold222 (.clk(u_txreg_N45),
    .clkout(net2175));
 b15cbf034ar1n64x5 hold223 (.clk(tx_data[12]),
    .clkout(net2176));
 b15cbf034ar1n64x5 hold224 (.clk(n2929),
    .clkout(net2177));
 b15cbf034ar1n64x5 hold225 (.clk(u_txreg_N46),
    .clkout(net2178));
 b15cbf034ar1n64x5 hold226 (.clk(tx_data[26]),
    .clkout(net2179));
 b15cbf034ar1n64x5 hold227 (.clk(n2925),
    .clkout(net2180));
 b15cbf034ar1n64x5 hold228 (.clk(u_txreg_N60),
    .clkout(net2181));
 b15cbf034ar1n64x5 hold229 (.clk(net2479),
    .clkout(net2182));
 b15cbf034ar1n64x5 hold230 (.clk(tx_data[13]),
    .clkout(net2183));
 b15cbf034ar1n64x5 hold231 (.clk(n2935),
    .clkout(net2184));
 b15cbf034ar1n64x5 hold232 (.clk(u_txreg_N47),
    .clkout(net2185));
 b15cbf034ar1n64x5 hold233 (.clk(tx_data[21]),
    .clkout(net2186));
 b15cbf034ar1n64x5 hold234 (.clk(n2941),
    .clkout(net2187));
 b15cbf034ar1n64x5 hold235 (.clk(u_txreg_N55),
    .clkout(net2188));
 b15cbf034ar1n64x5 hold236 (.clk(tx_data[15]),
    .clkout(net2189));
 b15cbf034ar1n64x5 hold237 (.clk(n2931),
    .clkout(net2190));
 b15cbf034ar1n64x5 hold238 (.clk(u_txreg_N49),
    .clkout(net2191));
 b15cbf034ar1n64x5 hold239 (.clk(tx_data[9]),
    .clkout(net2192));
 b15cbf034ar1n64x5 hold240 (.clk(n2936),
    .clkout(net2193));
 b15cbf034ar1n64x5 hold241 (.clk(u_txreg_N43),
    .clkout(net2194));
 b15cbf034ar1n64x5 hold242 (.clk(net2485),
    .clkout(net2195));
 b15cbf034ar1n64x5 hold243 (.clk(tx_data[0]),
    .clkout(net2196));
 b15cbf034ar1n64x5 hold244 (.clk(u_txreg_N34),
    .clkout(net2197));
 b15cbf034ar1n64x5 hold245 (.clk(tx_data[17]),
    .clkout(net2198));
 b15cbf034ar1n64x5 hold246 (.clk(n2937),
    .clkout(net2199));
 b15cbf034ar1n64x5 hold247 (.clk(u_txreg_N51),
    .clkout(net2200));
 b15cbf034ar1n64x5 hold248 (.clk(tx_data[14]),
    .clkout(net2201));
 b15cbf034ar1n64x5 hold249 (.clk(n2933),
    .clkout(net2202));
 b15cbf034ar1n64x5 hold250 (.clk(u_txreg_N48),
    .clkout(net2203));
 b15cbf034ar1n64x5 hold251 (.clk(tx_data[10]),
    .clkout(net2204));
 b15cbf034ar1n64x5 hold252 (.clk(n2932),
    .clkout(net2205));
 b15cbf034ar1n64x5 hold253 (.clk(tx_data[22]),
    .clkout(net2206));
 b15cbf034ar1n64x5 hold254 (.clk(n2943),
    .clkout(net2207));
 b15cbf034ar1n64x5 hold255 (.clk(net2489),
    .clkout(net2208));
 b15cbf034ar1n64x5 hold256 (.clk(tx_data[23]),
    .clkout(net2209));
 b15cbf034ar1n64x5 hold257 (.clk(n2934),
    .clkout(net2210));
 b15cbf034ar1n64x5 hold258 (.clk(u_txreg_N57),
    .clkout(net2211));
 b15cbf034ar1n64x5 hold259 (.clk(net2493),
    .clkout(net2212));
 b15cbf034ar1n64x5 hold260 (.clk(net2491),
    .clkout(net2213));
 b15cbf034ar1n64x5 hold261 (.clk(tx_data[3]),
    .clkout(net2214));
 b15cbf034ar1n64x5 hold262 (.clk(u_txreg_N37),
    .clkout(net2215));
 b15cbf034ar1n64x5 hold263 (.clk(net2500),
    .clkout(net2216));
 b15cbf034ar1n64x5 hold264 (.clk(tx_data[4]),
    .clkout(net2217));
 b15cbf034ar1n64x5 hold265 (.clk(n3688),
    .clkout(net2218));
 b15cbf034ar1n64x5 hold266 (.clk(tx_data[6]),
    .clkout(net2219));
 b15cbf034ar1n64x5 hold267 (.clk(n2946),
    .clkout(net2220));
 b15cbf034ar1n64x5 hold268 (.clk(u_txreg_N40),
    .clkout(net2221));
 b15cbf034ar1n64x5 hold269 (.clk(tx_data[5]),
    .clkout(net2222));
 b15cbf034ar1n64x5 hold270 (.clk(n3685),
    .clkout(net2223));
 b15cbf034ar1n64x5 hold271 (.clk(u_txreg_N39),
    .clkout(net2224));
 b15cbf034ar1n64x5 hold272 (.clk(tx_data[7]),
    .clkout(net2225));
 b15cbf034ar1n64x5 hold273 (.clk(n2948),
    .clkout(net2226));
 b15cbf034ar1n64x5 hold274 (.clk(u_txreg_N41),
    .clkout(net2227));
 b15cbf034ar1n64x5 hold275 (.clk(u_txreg_data_int[28]),
    .clkout(net2228));
 b15cbf034ar1n64x5 hold276 (.clk(net57),
    .clkout(net2229));
 b15cbf034ar1n64x5 hold277 (.clk(net2230),
    .clkout(spi_sdo0));
 b15cbf034ar1n64x5 hold278 (.clk(tx_data[30]),
    .clkout(net2231));
 b15cbf034ar1n64x5 hold279 (.clk(n2923),
    .clkout(net2232));
 b15cbf034ar1n64x5 hold280 (.clk(net2515),
    .clkout(net2233));
 b15cbf034ar1n64x5 hold281 (.clk(tx_data[28]),
    .clkout(net2234));
 b15cbf034ar1n64x5 hold282 (.clk(n2951),
    .clkout(net2235));
 b15cbf034ar1n64x5 hold283 (.clk(u_txreg_N62),
    .clkout(net2236));
 b15cbf034ar1n64x5 hold284 (.clk(u_dcfifo_tx_u_dout_empty_synch_d_middle[3]),
    .clkout(net2237));
 b15cbf034ar1n64x5 hold285 (.clk(tx_data[8]),
    .clkout(net2238));
 b15cbf034ar1n64x5 hold286 (.clk(n2942),
    .clkout(net2239));
 b15cbf034ar1n64x5 hold287 (.clk(u_txreg_N42),
    .clkout(net2240));
 b15cbf034ar1n64x5 hold288 (.clk(u_txreg_data_int[31]),
    .clkout(net2241));
 b15cbf034ar1n64x5 hold289 (.clk(net250),
    .clkout(net2242));
 b15cbf034ar1n64x5 hold290 (.clk(n1739),
    .clkout(net2243));
 b15cbf034ar1n64x5 hold291 (.clk(n1757),
    .clkout(net2244));
 b15cbf034ar1n64x5 hold292 (.clk(u_dcfifo_rx_u_dout_empty_synch_d_middle[7]),
    .clkout(net2245));
 b15cbf034ar1n64x5 hold293 (.clk(n1733),
    .clkout(net2246));
 b15cbf034ar1n64x5 hold294 (.clk(n1769),
    .clkout(net2247));
 b15cbf034ar1n64x5 hold295 (.clk(n1751),
    .clkout(net2248));
 b15cbf034ar1n64x5 hold296 (.clk(n1878),
    .clkout(net2249));
 b15cbf034ar1n64x5 hold297 (.clk(n1727),
    .clkout(net2250));
 b15cbf034ar1n64x5 hold298 (.clk(n1730),
    .clkout(net2251));
 b15cbf034ar1n64x5 hold299 (.clk(n1793),
    .clkout(net2252));
 b15cbf034ar1n64x5 hold300 (.clk(n1712),
    .clkout(net2253));
 b15cbf034ar1n64x5 hold301 (.clk(n1745),
    .clkout(net2254));
 b15cbf034ar1n64x5 hold302 (.clk(n1775),
    .clkout(net2255));
 b15cbf034ar1n64x5 hold303 (.clk(n1715),
    .clkout(net2256));
 b15cbf034ar1n64x5 hold304 (.clk(n1787),
    .clkout(net2257));
 b15cbf034ar1n64x5 hold305 (.clk(n1706),
    .clkout(net2258));
 b15cbf034ar1n64x5 hold306 (.clk(n1781),
    .clkout(net2259));
 b15cbf034ar1n64x5 hold307 (.clk(n1763),
    .clkout(net2260));
 b15cbf034ar1n64x5 hold308 (.clk(n1799),
    .clkout(net2261));
 b15cbf034ar1n64x5 hold309 (.clk(n1691),
    .clkout(net2262));
 b15cbf034ar1n64x5 hold310 (.clk(n1700),
    .clkout(net2263));
 b15cbf034ar1n64x5 hold311 (.clk(n1742),
    .clkout(net2264));
 b15cbf034ar1n64x5 hold312 (.clk(n1760),
    .clkout(net2265));
 b15cbf034ar1n64x5 hold313 (.clk(n1736),
    .clkout(net2266));
 b15cbf034ar1n64x5 hold314 (.clk(n1772),
    .clkout(net2267));
 b15cbf034ar1n64x5 hold315 (.clk(n1754),
    .clkout(net2268));
 b15cbf034ar1n64x5 hold316 (.clk(n1703),
    .clkout(net2269));
 b15cbf034ar1n64x5 hold317 (.clk(n1721),
    .clkout(net2270));
 b15cbf034ar1n64x5 hold318 (.clk(n1724),
    .clkout(net2271));
 b15cbf034ar1n64x5 hold319 (.clk(n1796),
    .clkout(net2272));
 b15cbf034ar1n64x5 hold320 (.clk(n1748),
    .clkout(net2273));
 b15cbf034ar1n64x5 hold321 (.clk(n1778),
    .clkout(net2274));
 b15cbf034ar1n64x5 hold322 (.clk(n1709),
    .clkout(net2275));
 b15cbf034ar1n64x5 hold323 (.clk(n1694),
    .clkout(net2276));
 b15cbf034ar1n64x5 hold324 (.clk(n1784),
    .clkout(net2277));
 b15cbf034ar1n64x5 hold325 (.clk(n1802),
    .clkout(net2278));
 b15cbf034ar1n64x5 hold326 (.clk(n1697),
    .clkout(net2279));
 b15cbf034ar1n64x5 hold327 (.clk(n1790),
    .clkout(net2280));
 b15cbf034ar1n64x5 hold328 (.clk(n1766),
    .clkout(net2281));
 b15cbf034ar1n64x5 hold329 (.clk(n1718),
    .clkout(net2282));
 b15cbf034ar1n64x5 hold330 (.clk(u_syncro_valid_reg[0]),
    .clkout(net2283));
 b15cbf034ar1n64x5 hold331 (.clk(u_dcfifo_tx_u_din_full_full_synch_d_middle_0_),
    .clkout(net2284));
 b15cbf034ar1n64x5 hold332 (.clk(u_dcfifo_rx_u_din_full_full_synch_d_middle_0_),
    .clkout(net2285));
 b15cbf034ar1n64x5 hold333 (.clk(n1881),
    .clkout(net2286));
 b15cbf034ar1n64x5 hold334 (.clk(u_syncro_rdwr_reg_0_),
    .clkout(net2287));
 b15cbf034ar1n64x5 hold335 (.clk(tx_data[31]),
    .clkout(net2288));
 b15cbf034ar1n64x5 hold336 (.clk(n2930),
    .clkout(net2289));
 b15cbf034ar1n64x5 hold337 (.clk(u_dcfifo_rx_write_token[1]),
    .clkout(net2290));
 b15cbf034ar1n64x5 hold338 (.clk(u_dcfifo_rx_u_dout_empty_synch_d_middle[6]),
    .clkout(net2291));
 b15cbf034ar1n64x5 hold339 (.clk(u_dcfifo_tx_u_dout_empty_synch_d_middle[7]),
    .clkout(net2292));
 b15cbf034ar1n64x5 hold340 (.clk(u_dcfifo_tx_u_dout_empty_synch_d_middle[1]),
    .clkout(net2293));
 b15cbf034ar1n64x5 hold341 (.clk(u_dcfifo_tx_u_dout_empty_synch_d_middle[0]),
    .clkout(net2294));
 b15cbf034ar1n64x5 hold342 (.clk(u_dcfifo_rx_u_dout_empty_synch_d_middle[2]),
    .clkout(net2295));
 b15cbf034ar1n64x5 hold343 (.clk(u_txreg_data_int[30]),
    .clkout(net2296));
 b15cbf034ar1n64x5 hold344 (.clk(u_dcfifo_rx_u_dout_empty_synch_d_middle[3]),
    .clkout(net2297));
 b15cbf034ar1n64x5 hold345 (.clk(tx_data_valid),
    .clkout(net2298));
 b15cbf034ar1n64x5 hold346 (.clk(net354),
    .clkout(net2299));
 b15cbf034ar1n64x5 hold347 (.clk(n2921),
    .clkout(net2300));
 b15cbf034ar1n64x5 hold348 (.clk(u_txreg_N63),
    .clkout(net2301));
 b15cbf034ar1n64x5 hold349 (.clk(u_dcfifo_tx_u_dout_read_token[7]),
    .clkout(net2302));
 b15cbf034ar1n64x5 hold350 (.clk(u_dcfifo_rx_u_dout_empty_synch_d_middle[4]),
    .clkout(net2303));
 b15cbf034ar1n64x5 hold351 (.clk(u_dcfifo_tx_write_token[1]),
    .clkout(net2304));
 b15cbf034ar1n64x5 hold352 (.clk(u_dcfifo_tx_u_dout_empty_synch_d_middle[6]),
    .clkout(net2305));
 b15cbf034ar1n64x5 hold353 (.clk(u_dcfifo_tx_write_token[2]),
    .clkout(net2306));
 b15cbf034ar1n64x5 hold354 (.clk(u_dcfifo_rx_write_token[2]),
    .clkout(net2307));
 b15cbf034ar1n64x5 hold355 (.clk(u_dcfifo_tx_write_token[0]),
    .clkout(net2308));
 b15cbf034ar1n64x5 hold356 (.clk(u_dcfifo_rx_u_dout_empty_synch_d_middle[0]),
    .clkout(net2309));
 b15cbf034ar1n64x5 hold357 (.clk(u_dcfifo_rx_u_dout_empty_synch_d_middle[5]),
    .clkout(net2310));
 b15cbf034ar1n64x5 hold358 (.clk(u_dcfifo_tx_write_token[6]),
    .clkout(net2311));
 b15cbf034ar1n64x5 hold359 (.clk(tx_data[1]),
    .clkout(net2312));
 b15cbf034ar1n64x5 hold360 (.clk(u_txreg_N35),
    .clkout(net2313));
 b15cbf034ar1n64x5 hold361 (.clk(u_dcfifo_rx_u_dout_empty_synch_d_middle[1]),
    .clkout(net2314));
 b15cbf034ar1n64x5 hold362 (.clk(tx_data[2]),
    .clkout(net2315));
 b15cbf034ar1n64x5 hold363 (.clk(u_txreg_N36),
    .clkout(net2316));
 b15cbf034ar1n64x5 hold364 (.clk(u_txreg_data_int[29]),
    .clkout(net2317));
 b15cbf034ar1n64x5 hold365 (.clk(addr_sync[23]),
    .clkout(net2318));
 b15cbf034ar1n64x5 hold366 (.clk(u_syncro_valid_reg[1]),
    .clkout(net2319));
 b15cbf034ar1n64x5 hold367 (.clk(n1455),
    .clkout(net2320));
 b15cbf034ar1n64x5 hold368 (.clk(addr_sync[22]),
    .clkout(net2321));
 b15cbf034ar1n64x5 hold369 (.clk(u_dcfifo_tx_u_dout_empty_synch_d_middle[4]),
    .clkout(net2322));
 b15cbf034ar1n64x5 hold370 (.clk(addr_sync[9]),
    .clkout(net2323));
 b15cbf034ar1n64x5 hold371 (.clk(addr_sync[17]),
    .clkout(net2324));
 b15cbf034ar1n64x5 hold372 (.clk(addr_sync[29]),
    .clkout(net2325));
 b15cbf034ar1n64x5 hold373 (.clk(u_dcfifo_tx_u_dout_empty_synch_d_middle[5]),
    .clkout(net2326));
 b15cbf034ar1n64x5 hold374 (.clk(u_dcfifo_rx_u_dout_read_token[7]),
    .clkout(net2327));
 b15cbf034ar1n64x5 hold375 (.clk(addr_sync[13]),
    .clkout(net2328));
 b15cbf034ar1n64x5 hold376 (.clk(u_dcfifo_tx_u_din_full_latched_full_s),
    .clkout(net2329));
 b15cbf034ar1n64x5 hold377 (.clk(u_dcfifo_rx_write_token[4]),
    .clkout(net2330));
 b15cbf034ar1n64x5 hold378 (.clk(addr_sync[8]),
    .clkout(net2331));
 b15cbf034ar1n64x5 hold379 (.clk(u_device_sm_s_dummy_cycles[5]),
    .clkout(net2332));
 b15cbf034ar1n64x5 hold380 (.clk(u_rxreg_data_int[12]),
    .clkout(net2333));
 b15cbf034ar1n64x5 hold381 (.clk(addr_sync[1]),
    .clkout(net2334));
 b15cbf034ar1n64x5 hold382 (.clk(addr_sync[16]),
    .clkout(net2335));
 b15cbf034ar1n64x5 hold383 (.clk(addr_sync[28]),
    .clkout(net2336));
 b15cbf034ar1n64x5 hold384 (.clk(tx_counter_upd),
    .clkout(net2337));
 b15cbf034ar1n64x5 hold385 (.clk(u_dcfifo_rx_u_dout_read_token[3]),
    .clkout(net2338));
 b15cbf034ar1n64x5 hold386 (.clk(u_rxreg_data_int[9]),
    .clkout(net2339));
 b15cbf034ar1n64x5 hold387 (.clk(addr_sync[12]),
    .clkout(net2340));
 b15cbf034ar1n64x5 hold388 (.clk(addr_sync[25]),
    .clkout(net2341));
 b15cbf034ar1n64x5 hold389 (.clk(u_rxreg_data_int[30]),
    .clkout(net2342));
 b15cbf034ar1n64x5 hold390 (.clk(addr_sync[21]),
    .clkout(net2343));
 b15cbf034ar1n64x5 hold391 (.clk(addr_sync[0]),
    .clkout(net2344));
 b15cbf034ar1n64x5 hold392 (.clk(u_dcfifo_rx_u_dout_read_token[6]),
    .clkout(net2345));
 b15cbf034ar1n64x5 hold393 (.clk(u_device_sm_s_dummy_cycles[2]),
    .clkout(net2346));
 b15cbf034ar1n64x5 hold394 (.clk(u_spi_device_tlul_plug_state[0]),
    .clkout(net2347));
 b15cbf034ar1n64x5 hold395 (.clk(u_spi_device_tlul_plug_state_next[1]),
    .clkout(net2348));
 b15cbf034ar1n64x5 hold396 (.clk(u_rxreg_data_int[5]),
    .clkout(net2349));
 b15cbf034ar1n64x5 hold397 (.clk(u_rxreg_data_int[6]),
    .clkout(net2350));
 b15cbf034ar1n64x5 hold398 (.clk(u_dcfifo_tx_u_dout_write_token_dn[0]),
    .clkout(net2351));
 b15cbf034ar1n64x5 hold399 (.clk(n2773),
    .clkout(net2352));
 b15cbf034ar1n64x5 hold400 (.clk(u_dcfifo_tx_u_dout_read_enable),
    .clkout(net2353));
 b15cbf034ar1n64x5 hold401 (.clk(u_rxreg_data_int[24]),
    .clkout(net2354));
 b15cbf034ar1n64x5 hold402 (.clk(u_dcfifo_rx_write_token[5]),
    .clkout(net2355));
 b15cbf034ar1n64x5 hold403 (.clk(u_dcfifo_tx_write_token[5]),
    .clkout(net2356));
 b15cbf034ar1n64x5 hold404 (.clk(addr_sync[24]),
    .clkout(net2357));
 b15cbf034ar1n64x5 hold405 (.clk(addr_sync[31]),
    .clkout(net2358));
 b15cbf034ar1n64x5 hold406 (.clk(addr_sync[20]),
    .clkout(net2359));
 b15cbf034ar1n64x5 hold407 (.clk(u_dcfifo_rx_write_token[7]),
    .clkout(net2360));
 b15cbf034ar1n64x5 hold408 (.clk(addr_sync[15]),
    .clkout(net2361));
 b15cbf034ar1n64x5 hold409 (.clk(u_dcfifo_rx_u_dout_read_token[5]),
    .clkout(net2362));
 b15cbf034ar1n64x5 hold410 (.clk(addr_sync[27]),
    .clkout(net2363));
 b15cbf034ar1n64x5 hold411 (.clk(u_rxreg_data_int[1]),
    .clkout(net2364));
 b15cbf034ar1n64x5 hold412 (.clk(u_dcfifo_tx_u_dout_read_token[1]),
    .clkout(net2365));
 b15cbf034ar1n64x5 hold413 (.clk(u_dcfifo_rx_u_dout_write_token_dn[1]),
    .clkout(net2366));
 b15cbf034ar1n64x5 hold414 (.clk(addr_sync[30]),
    .clkout(net2367));
 b15cbf034ar1n64x5 hold415 (.clk(addr_sync[14]),
    .clkout(net2368));
 b15cbf034ar1n64x5 hold416 (.clk(addr_sync[26]),
    .clkout(net2369));
 b15cbf034ar1n64x5 hold417 (.clk(u_rxreg_counter[7]),
    .clkout(net2370));
 b15cbf034ar1n64x5 hold418 (.clk(u_dcfifo_rx_write_token[3]),
    .clkout(net2371));
 b15cbf034ar1n64x5 hold419 (.clk(u_txreg_counter[2]),
    .clkout(net2372));
 b15cbf034ar1n64x5 hold420 (.clk(net73),
    .clkout(net2373));
 b15cbf034ar1n64x5 hold421 (.clk(net1956),
    .clkout(net2374));
 b15cbf034ar1n64x5 hold422 (.clk(net1957),
    .clkout(net2375));
 b15cbf034ar1n64x5 hold423 (.clk(net82),
    .clkout(net2376));
 b15cbf034ar1n64x5 hold424 (.clk(net1958),
    .clkout(net2377));
 b15cbf034ar1n64x5 hold425 (.clk(net1959),
    .clkout(net2378));
 b15cbf034ar1n64x5 hold426 (.clk(net81),
    .clkout(net2379));
 b15cbf034ar1n64x5 hold427 (.clk(net1960),
    .clkout(net2380));
 b15cbf034ar1n64x5 hold428 (.clk(net1961),
    .clkout(net2381));
 b15cbf034ar1n64x5 hold429 (.clk(net74),
    .clkout(net2382));
 b15cbf034ar1n64x5 hold430 (.clk(net1962),
    .clkout(net2383));
 b15cbf034ar1n64x5 hold431 (.clk(net1963),
    .clkout(net2384));
 b15cbf034ar1n64x5 hold432 (.clk(net91),
    .clkout(net2385));
 b15cbf034ar1n64x5 hold433 (.clk(net1967),
    .clkout(net2386));
 b15cbf034ar1n64x5 hold434 (.clk(net1968),
    .clkout(net2387));
 b15cbf034ar1n64x5 hold435 (.clk(net92),
    .clkout(net2388));
 b15cbf034ar1n64x5 hold436 (.clk(net1969),
    .clkout(net2389));
 b15cbf034ar1n64x5 hold437 (.clk(net1970),
    .clkout(net2390));
 b15cbf034ar1n64x5 hold438 (.clk(net94),
    .clkout(net2391));
 b15cbf034ar1n64x5 hold439 (.clk(net1971),
    .clkout(net2392));
 b15cbf034ar1n64x5 hold440 (.clk(net1972),
    .clkout(net2393));
 b15cbf034ar1n64x5 hold441 (.clk(net93),
    .clkout(net2394));
 b15cbf034ar1n64x5 hold442 (.clk(net1973),
    .clkout(net2395));
 b15cbf034ar1n64x5 hold443 (.clk(net1974),
    .clkout(net2396));
 b15cbf034ar1n64x5 hold444 (.clk(net78),
    .clkout(net2397));
 b15cbf034ar1n64x5 hold445 (.clk(net1984),
    .clkout(net2398));
 b15cbf034ar1n64x5 hold446 (.clk(net1985),
    .clkout(net2399));
 b15cbf034ar1n64x5 hold447 (.clk(net80),
    .clkout(net2400));
 b15cbf034ar1n64x5 hold448 (.clk(net1978),
    .clkout(net2401));
 b15cbf034ar1n64x5 hold449 (.clk(net1979),
    .clkout(net2402));
 b15cbf034ar1n64x5 hold450 (.clk(net79),
    .clkout(net2403));
 b15cbf034ar1n64x5 hold451 (.clk(net1982),
    .clkout(net2404));
 b15cbf034ar1n64x5 hold452 (.clk(net1983),
    .clkout(net2405));
 b15cbf034ar1n64x5 hold453 (.clk(net77),
    .clkout(net2406));
 b15cbf034ar1n64x5 hold454 (.clk(net1989),
    .clkout(net2407));
 b15cbf034ar1n64x5 hold455 (.clk(net1990),
    .clkout(net2408));
 b15cbf034ar1n64x5 hold456 (.clk(net87),
    .clkout(net2409));
 b15cbf034ar1n64x5 hold457 (.clk(net1994),
    .clkout(net2410));
 b15cbf034ar1n64x5 hold458 (.clk(net1995),
    .clkout(net2411));
 b15cbf034ar1n64x5 hold459 (.clk(net88),
    .clkout(net2412));
 b15cbf034ar1n64x5 hold460 (.clk(net1996),
    .clkout(net2413));
 b15cbf034ar1n64x5 hold461 (.clk(net1997),
    .clkout(net2414));
 b15cbf034ar1n64x5 hold462 (.clk(net76),
    .clkout(net2415));
 b15cbf034ar1n64x5 hold463 (.clk(net1998),
    .clkout(net2416));
 b15cbf034ar1n64x5 hold464 (.clk(net1999),
    .clkout(net2417));
 b15cbf034ar1n64x5 hold465 (.clk(net75),
    .clkout(net2418));
 b15cbf034ar1n64x5 hold466 (.clk(net2000),
    .clkout(net2419));
 b15cbf034ar1n64x5 hold467 (.clk(net2001),
    .clkout(net2420));
 b15cbf034ar1n64x5 hold468 (.clk(net83),
    .clkout(net2421));
 b15cbf034ar1n64x5 hold469 (.clk(net2002),
    .clkout(net2422));
 b15cbf034ar1n64x5 hold470 (.clk(net2003),
    .clkout(net2423));
 b15cbf034ar1n64x5 hold471 (.clk(net84),
    .clkout(net2424));
 b15cbf034ar1n64x5 hold472 (.clk(net2004),
    .clkout(net2425));
 b15cbf034ar1n64x5 hold473 (.clk(net2005),
    .clkout(net2426));
 b15cbf034ar1n64x5 hold474 (.clk(net72),
    .clkout(net2427));
 b15cbf034ar1n64x5 hold475 (.clk(net2010),
    .clkout(net2428));
 b15cbf034ar1n64x5 hold476 (.clk(net2011),
    .clkout(net2429));
 b15cbf034ar1n64x5 hold477 (.clk(net71),
    .clkout(net2430));
 b15cbf034ar1n64x5 hold478 (.clk(net2008),
    .clkout(net2431));
 b15cbf034ar1n64x5 hold479 (.clk(net2009),
    .clkout(net2432));
 b15cbf034ar1n64x5 hold480 (.clk(net68),
    .clkout(net2433));
 b15cbf034ar1n64x5 hold481 (.clk(net2006),
    .clkout(net2434));
 b15cbf034ar1n64x5 hold482 (.clk(net2007),
    .clkout(net2435));
 b15cbf034ar1n64x5 hold483 (.clk(net98),
    .clkout(net2436));
 b15cbf034ar1n64x5 hold484 (.clk(net2027),
    .clkout(net2437));
 b15cbf034ar1n64x5 hold485 (.clk(net2028),
    .clkout(net2438));
 b15cbf034ar1n64x5 hold486 (.clk(net86),
    .clkout(net2439));
 b15cbf034ar1n64x5 hold487 (.clk(net2018),
    .clkout(net2440));
 b15cbf034ar1n64x5 hold488 (.clk(net85),
    .clkout(net2441));
 b15cbf034ar1n64x5 hold489 (.clk(net2016),
    .clkout(net2442));
 b15cbf034ar1n64x5 hold490 (.clk(net99),
    .clkout(net2443));
 b15cbf034ar1n64x5 hold491 (.clk(net2023),
    .clkout(net2444));
 b15cbf034ar1n64x5 hold492 (.clk(tx_counter[7]),
    .clkout(net2445));
 b15cbf034ar1n64x5 hold493 (.clk(net2086),
    .clkout(net2446));
 b15cbf034ar1n64x5 hold494 (.clk(net69),
    .clkout(net2447));
 b15cbf034ar1n64x5 hold495 (.clk(net2031),
    .clkout(net2448));
 b15cbf034ar1n64x5 hold496 (.clk(net70),
    .clkout(net2449));
 b15cbf034ar1n64x5 hold497 (.clk(net2033),
    .clkout(net2450));
 b15cbf034ar1n64x5 hold498 (.clk(net97),
    .clkout(net2451));
 b15cbf034ar1n64x5 hold499 (.clk(net2039),
    .clkout(net2452));
 b15cbf034ar1n64x5 hold500 (.clk(net2040),
    .clkout(net2453));
 b15cbf034ar1n64x5 hold501 (.clk(net130),
    .clkout(net2454));
 b15cbf034ar1n64x5 hold502 (.clk(net2029),
    .clkout(net2455));
 b15cbf034ar1n64x5 hold503 (.clk(net131),
    .clkout(net2456));
 b15cbf034ar1n64x5 hold504 (.clk(net1980),
    .clkout(net2457));
 b15cbf034ar1n64x5 hold505 (.clk(net122),
    .clkout(net2458));
 b15cbf034ar1n64x5 hold506 (.clk(net2055),
    .clkout(net2459));
 b15cbf034ar1n64x5 hold507 (.clk(net127),
    .clkout(net2460));
 b15cbf034ar1n64x5 hold508 (.clk(net2057),
    .clkout(net2461));
 b15cbf034ar1n64x5 hold509 (.clk(net96),
    .clkout(net2462));
 b15cbf034ar1n64x5 hold510 (.clk(net2051),
    .clkout(net2463));
 b15cbf034ar1n64x5 hold511 (.clk(u_spi_device_tlul_plug_state[1]),
    .clkout(net2464));
 b15cbf034ar1n64x5 hold512 (.clk(net344),
    .clkout(net2465));
 b15cbf034ar1n64x5 hold513 (.clk(net62),
    .clkout(net2466));
 b15cbf034ar1n64x5 hold514 (.clk(net118),
    .clkout(net2467));
 b15cbf034ar1n64x5 hold515 (.clk(net2025),
    .clkout(net2468));
 b15cbf034ar1n64x5 hold516 (.clk(net121),
    .clkout(net2469));
 b15cbf034ar1n64x5 hold517 (.clk(net2041),
    .clkout(net2470));
 b15cbf034ar1n64x5 hold518 (.clk(net124),
    .clkout(net2471));
 b15cbf034ar1n64x5 hold519 (.clk(net2125),
    .clkout(net2472));
 b15cbf034ar1n64x5 hold520 (.clk(net100),
    .clkout(net2473));
 b15cbf034ar1n64x5 hold521 (.clk(net2046),
    .clkout(net2474));
 b15cbf034ar1n64x5 hold522 (.clk(net109),
    .clkout(net2475));
 b15cbf034ar1n64x5 hold523 (.clk(net2053),
    .clkout(net2476));
 b15cbf034ar1n64x5 hold524 (.clk(net95),
    .clkout(net2477));
 b15cbf034ar1n64x5 hold525 (.clk(net1964),
    .clkout(net2478));
 b15cbf034ar1n64x5 hold526 (.clk(tx_counter[1]),
    .clkout(net2479));
 b15cbf034ar1n64x5 hold527 (.clk(net2182),
    .clkout(net2480));
 b15cbf034ar1n64x5 hold528 (.clk(tx_counter[6]),
    .clkout(net2481));
 b15cbf034ar1n64x5 hold529 (.clk(net2169),
    .clkout(net2482));
 b15cbf034ar1n64x5 hold530 (.clk(net106),
    .clkout(net2483));
 b15cbf034ar1n64x5 hold531 (.clk(net2082),
    .clkout(net2484));
 b15cbf034ar1n64x5 hold532 (.clk(tx_counter[5]),
    .clkout(net2485));
 b15cbf034ar1n64x5 hold533 (.clk(net2195),
    .clkout(net2486));
 b15cbf034ar1n64x5 hold534 (.clk(net111),
    .clkout(net2487));
 b15cbf034ar1n64x5 hold535 (.clk(net2114),
    .clkout(net2488));
 b15cbf034ar1n64x5 hold536 (.clk(tx_counter[4]),
    .clkout(net2489));
 b15cbf034ar1n64x5 hold537 (.clk(net2208),
    .clkout(net2490));
 b15cbf034ar1n64x5 hold538 (.clk(tx_counter[2]),
    .clkout(net2491));
 b15cbf034ar1n64x5 hold539 (.clk(net2213),
    .clkout(net2492));
 b15cbf034ar1n64x5 hold540 (.clk(tx_counter[0]),
    .clkout(net2493));
 b15cbf034ar1n64x5 hold541 (.clk(net2212),
    .clkout(net2494));
 b15cbf034ar1n64x5 hold542 (.clk(net89),
    .clkout(net2495));
 b15cbf034ar1n64x5 hold543 (.clk(net90),
    .clkout(net2496));
 b15cbf034ar1n64x5 hold544 (.clk(net113),
    .clkout(net2497));
 b15cbf034ar1n64x5 hold545 (.clk(net105),
    .clkout(net2498));
 b15cbf034ar1n64x5 hold546 (.clk(net2118),
    .clkout(net2499));
 b15cbf034ar1n64x5 hold547 (.clk(tx_counter[3]),
    .clkout(net2500));
 b15cbf034ar1n64x5 hold548 (.clk(net110),
    .clkout(net2501));
 b15cbf034ar1n64x5 hold549 (.clk(net125),
    .clkout(net2502));
 b15cbf034ar1n64x5 hold550 (.clk(net2120),
    .clkout(net2503));
 b15cbf034ar1n64x5 hold551 (.clk(net115),
    .clkout(net2504));
 b15cbf034ar1n64x5 hold552 (.clk(net2132),
    .clkout(net2505));
 b15cbf034ar1n64x5 hold553 (.clk(en_quad),
    .clkout(net2506));
 b15cbf034ar1n64x5 hold554 (.clk(net117),
    .clkout(net2507));
 b15cbf034ar1n64x5 hold555 (.clk(net120),
    .clkout(net2508));
 b15cbf034ar1n64x5 hold556 (.clk(net114),
    .clkout(net2509));
 b15cbf034ar1n64x5 hold557 (.clk(net101),
    .clkout(net2510));
 b15cbf034ar1n64x5 hold558 (.clk(net107),
    .clkout(net2511));
 b15cbf034ar1n64x5 hold559 (.clk(net102),
    .clkout(net2512));
 b15cbf034ar1n64x5 hold560 (.clk(n3316),
    .clkout(net2513));
 b15cbf034ar1n64x5 hold561 (.clk(u_rxreg_data_int[30]),
    .clkout(net2514));
 b15cbf034ar1n64x5 hold562 (.clk(u_syncro_cs_reg_0_),
    .clkout(net2515));
 b15cbf034ar1n64x5 hold563 (.clk(net102),
    .clkout(net2516));
 b15zdnd11an1n64x5 FILLER_0_8 ();
 b15zdnd11an1n64x5 FILLER_0_72 ();
 b15zdnd11an1n64x5 FILLER_0_136 ();
 b15zdnd11an1n64x5 FILLER_0_200 ();
 b15zdnd11an1n64x5 FILLER_0_264 ();
 b15zdnd11an1n64x5 FILLER_0_328 ();
 b15zdnd11an1n64x5 FILLER_0_392 ();
 b15zdnd11an1n64x5 FILLER_0_456 ();
 b15zdnd11an1n16x5 FILLER_0_520 ();
 b15zdnd11an1n04x5 FILLER_0_540 ();
 b15zdnd11an1n64x5 FILLER_0_586 ();
 b15zdnd11an1n64x5 FILLER_0_650 ();
 b15zdnd11an1n04x5 FILLER_0_714 ();
 b15zdnd11an1n64x5 FILLER_0_726 ();
 b15zdnd11an1n16x5 FILLER_0_790 ();
 b15zdnd11an1n08x5 FILLER_0_806 ();
 b15zdnd11an1n04x5 FILLER_0_814 ();
 b15zdnd00an1n02x5 FILLER_0_818 ();
 b15zdnd11an1n04x5 FILLER_0_862 ();
 b15zdnd11an1n16x5 FILLER_0_908 ();
 b15zdnd11an1n08x5 FILLER_0_966 ();
 b15zdnd11an1n04x5 FILLER_0_978 ();
 b15zdnd11an1n04x5 FILLER_0_1024 ();
 b15zdnd00an1n02x5 FILLER_0_1028 ();
 b15zdnd00an1n01x5 FILLER_0_1030 ();
 b15zdnd11an1n04x5 FILLER_0_1073 ();
 b15zdnd00an1n01x5 FILLER_0_1077 ();
 b15zdnd11an1n64x5 FILLER_0_1120 ();
 b15zdnd11an1n16x5 FILLER_0_1184 ();
 b15zdnd11an1n04x5 FILLER_0_1204 ();
 b15zdnd11an1n16x5 FILLER_0_1250 ();
 b15zdnd11an1n04x5 FILLER_0_1266 ();
 b15zdnd00an1n01x5 FILLER_0_1270 ();
 b15zdnd11an1n16x5 FILLER_0_1313 ();
 b15zdnd11an1n04x5 FILLER_0_1333 ();
 b15zdnd11an1n08x5 FILLER_0_1379 ();
 b15zdnd11an1n04x5 FILLER_0_1429 ();
 b15zdnd00an1n02x5 FILLER_0_1433 ();
 b15zdnd00an1n01x5 FILLER_0_1435 ();
 b15zdnd00an1n02x5 FILLER_0_1444 ();
 b15zdnd11an1n08x5 FILLER_0_1488 ();
 b15zdnd00an1n02x5 FILLER_0_1496 ();
 b15zdnd11an1n04x5 FILLER_0_1540 ();
 b15zdnd00an1n02x5 FILLER_0_1544 ();
 b15zdnd00an1n01x5 FILLER_0_1546 ();
 b15zdnd11an1n08x5 FILLER_0_1589 ();
 b15zdnd11an1n04x5 FILLER_0_1639 ();
 b15zdnd11an1n04x5 FILLER_0_1685 ();
 b15zdnd11an1n64x5 FILLER_0_1731 ();
 b15zdnd11an1n32x5 FILLER_0_1795 ();
 b15zdnd11an1n16x5 FILLER_0_1827 ();
 b15zdnd11an1n08x5 FILLER_0_1843 ();
 b15zdnd11an1n04x5 FILLER_0_1851 ();
 b15zdnd00an1n02x5 FILLER_0_1855 ();
 b15zdnd11an1n04x5 FILLER_0_1861 ();
 b15zdnd00an1n02x5 FILLER_0_1865 ();
 b15zdnd11an1n04x5 FILLER_0_1909 ();
 b15zdnd00an1n01x5 FILLER_0_1913 ();
 b15zdnd11an1n04x5 FILLER_0_1956 ();
 b15zdnd11an1n64x5 FILLER_0_2002 ();
 b15zdnd11an1n64x5 FILLER_0_2066 ();
 b15zdnd11an1n16x5 FILLER_0_2130 ();
 b15zdnd11an1n08x5 FILLER_0_2146 ();
 b15zdnd11an1n64x5 FILLER_0_2162 ();
 b15zdnd11an1n32x5 FILLER_0_2226 ();
 b15zdnd11an1n16x5 FILLER_0_2258 ();
 b15zdnd00an1n02x5 FILLER_0_2274 ();
 b15zdnd11an1n64x5 FILLER_1_0 ();
 b15zdnd11an1n64x5 FILLER_1_64 ();
 b15zdnd11an1n64x5 FILLER_1_128 ();
 b15zdnd11an1n64x5 FILLER_1_192 ();
 b15zdnd11an1n64x5 FILLER_1_256 ();
 b15zdnd11an1n64x5 FILLER_1_320 ();
 b15zdnd11an1n64x5 FILLER_1_384 ();
 b15zdnd11an1n64x5 FILLER_1_448 ();
 b15zdnd11an1n32x5 FILLER_1_512 ();
 b15zdnd00an1n01x5 FILLER_1_544 ();
 b15zdnd11an1n64x5 FILLER_1_587 ();
 b15zdnd11an1n64x5 FILLER_1_651 ();
 b15zdnd11an1n64x5 FILLER_1_715 ();
 b15zdnd11an1n32x5 FILLER_1_779 ();
 b15zdnd11an1n16x5 FILLER_1_811 ();
 b15zdnd11an1n04x5 FILLER_1_827 ();
 b15zdnd00an1n01x5 FILLER_1_831 ();
 b15zdnd11an1n32x5 FILLER_1_836 ();
 b15zdnd00an1n02x5 FILLER_1_868 ();
 b15zdnd11an1n16x5 FILLER_1_874 ();
 b15zdnd11an1n08x5 FILLER_1_890 ();
 b15zdnd00an1n02x5 FILLER_1_898 ();
 b15zdnd11an1n08x5 FILLER_1_908 ();
 b15zdnd11an1n04x5 FILLER_1_916 ();
 b15zdnd00an1n01x5 FILLER_1_920 ();
 b15zdnd11an1n04x5 FILLER_1_928 ();
 b15zdnd11an1n04x5 FILLER_1_974 ();
 b15zdnd00an1n02x5 FILLER_1_978 ();
 b15zdnd11an1n04x5 FILLER_1_984 ();
 b15zdnd11an1n08x5 FILLER_1_1030 ();
 b15zdnd00an1n01x5 FILLER_1_1038 ();
 b15zdnd11an1n04x5 FILLER_1_1081 ();
 b15zdnd00an1n02x5 FILLER_1_1085 ();
 b15zdnd11an1n64x5 FILLER_1_1129 ();
 b15zdnd11an1n16x5 FILLER_1_1193 ();
 b15zdnd00an1n01x5 FILLER_1_1209 ();
 b15zdnd11an1n16x5 FILLER_1_1252 ();
 b15zdnd11an1n08x5 FILLER_1_1268 ();
 b15zdnd11an1n04x5 FILLER_1_1276 ();
 b15zdnd11an1n16x5 FILLER_1_1322 ();
 b15zdnd00an1n01x5 FILLER_1_1338 ();
 b15zdnd11an1n08x5 FILLER_1_1381 ();
 b15zdnd11an1n08x5 FILLER_1_1431 ();
 b15zdnd00an1n01x5 FILLER_1_1439 ();
 b15zdnd11an1n04x5 FILLER_1_1482 ();
 b15zdnd00an1n02x5 FILLER_1_1486 ();
 b15zdnd11an1n04x5 FILLER_1_1492 ();
 b15zdnd11an1n04x5 FILLER_1_1538 ();
 b15zdnd11an1n32x5 FILLER_1_1546 ();
 b15zdnd11an1n08x5 FILLER_1_1578 ();
 b15zdnd11an1n04x5 FILLER_1_1586 ();
 b15zdnd00an1n01x5 FILLER_1_1590 ();
 b15zdnd11an1n16x5 FILLER_1_1595 ();
 b15zdnd11an1n04x5 FILLER_1_1611 ();
 b15zdnd00an1n02x5 FILLER_1_1615 ();
 b15zdnd11an1n04x5 FILLER_1_1621 ();
 b15zdnd00an1n02x5 FILLER_1_1625 ();
 b15zdnd11an1n04x5 FILLER_1_1669 ();
 b15zdnd11an1n04x5 FILLER_1_1677 ();
 b15zdnd11an1n64x5 FILLER_1_1723 ();
 b15zdnd11an1n64x5 FILLER_1_1787 ();
 b15zdnd11an1n32x5 FILLER_1_1851 ();
 b15zdnd11an1n16x5 FILLER_1_1883 ();
 b15zdnd00an1n02x5 FILLER_1_1899 ();
 b15zdnd00an1n01x5 FILLER_1_1901 ();
 b15zdnd11an1n08x5 FILLER_1_1906 ();
 b15zdnd11an1n04x5 FILLER_1_1956 ();
 b15zdnd11an1n64x5 FILLER_1_2002 ();
 b15zdnd11an1n64x5 FILLER_1_2066 ();
 b15zdnd11an1n64x5 FILLER_1_2130 ();
 b15zdnd11an1n64x5 FILLER_1_2194 ();
 b15zdnd11an1n16x5 FILLER_1_2258 ();
 b15zdnd11an1n08x5 FILLER_1_2274 ();
 b15zdnd00an1n02x5 FILLER_1_2282 ();
 b15zdnd11an1n64x5 FILLER_2_8 ();
 b15zdnd11an1n64x5 FILLER_2_72 ();
 b15zdnd11an1n64x5 FILLER_2_136 ();
 b15zdnd11an1n64x5 FILLER_2_200 ();
 b15zdnd11an1n64x5 FILLER_2_264 ();
 b15zdnd11an1n64x5 FILLER_2_328 ();
 b15zdnd11an1n64x5 FILLER_2_392 ();
 b15zdnd11an1n64x5 FILLER_2_456 ();
 b15zdnd11an1n64x5 FILLER_2_520 ();
 b15zdnd11an1n64x5 FILLER_2_584 ();
 b15zdnd11an1n64x5 FILLER_2_648 ();
 b15zdnd11an1n04x5 FILLER_2_712 ();
 b15zdnd00an1n02x5 FILLER_2_716 ();
 b15zdnd11an1n64x5 FILLER_2_726 ();
 b15zdnd11an1n64x5 FILLER_2_790 ();
 b15zdnd11an1n64x5 FILLER_2_854 ();
 b15zdnd11an1n16x5 FILLER_2_918 ();
 b15zdnd00an1n02x5 FILLER_2_934 ();
 b15zdnd11an1n32x5 FILLER_2_940 ();
 b15zdnd11an1n04x5 FILLER_2_972 ();
 b15zdnd11an1n04x5 FILLER_2_1018 ();
 b15zdnd00an1n02x5 FILLER_2_1022 ();
 b15zdnd00an1n01x5 FILLER_2_1024 ();
 b15zdnd11an1n04x5 FILLER_2_1067 ();
 b15zdnd11an1n08x5 FILLER_2_1079 ();
 b15zdnd11an1n04x5 FILLER_2_1087 ();
 b15zdnd11an1n64x5 FILLER_2_1095 ();
 b15zdnd11an1n64x5 FILLER_2_1159 ();
 b15zdnd11an1n32x5 FILLER_2_1223 ();
 b15zdnd11an1n16x5 FILLER_2_1255 ();
 b15zdnd11an1n08x5 FILLER_2_1271 ();
 b15zdnd11an1n04x5 FILLER_2_1279 ();
 b15zdnd00an1n01x5 FILLER_2_1283 ();
 b15zdnd11an1n64x5 FILLER_2_1288 ();
 b15zdnd11an1n32x5 FILLER_2_1352 ();
 b15zdnd00an1n02x5 FILLER_2_1384 ();
 b15zdnd00an1n01x5 FILLER_2_1386 ();
 b15zdnd11an1n32x5 FILLER_2_1391 ();
 b15zdnd11an1n04x5 FILLER_2_1423 ();
 b15zdnd00an1n02x5 FILLER_2_1427 ();
 b15zdnd00an1n01x5 FILLER_2_1429 ();
 b15zdnd11an1n64x5 FILLER_2_1434 ();
 b15zdnd11an1n64x5 FILLER_2_1498 ();
 b15zdnd11an1n64x5 FILLER_2_1562 ();
 b15zdnd11an1n64x5 FILLER_2_1626 ();
 b15zdnd11an1n64x5 FILLER_2_1690 ();
 b15zdnd11an1n64x5 FILLER_2_1754 ();
 b15zdnd11an1n64x5 FILLER_2_1818 ();
 b15zdnd11an1n32x5 FILLER_2_1882 ();
 b15zdnd11an1n04x5 FILLER_2_1914 ();
 b15zdnd00an1n02x5 FILLER_2_1918 ();
 b15zdnd00an1n01x5 FILLER_2_1920 ();
 b15zdnd11an1n64x5 FILLER_2_1963 ();
 b15zdnd11an1n64x5 FILLER_2_2027 ();
 b15zdnd11an1n32x5 FILLER_2_2091 ();
 b15zdnd11an1n16x5 FILLER_2_2123 ();
 b15zdnd11an1n08x5 FILLER_2_2139 ();
 b15zdnd11an1n04x5 FILLER_2_2147 ();
 b15zdnd00an1n02x5 FILLER_2_2151 ();
 b15zdnd00an1n01x5 FILLER_2_2153 ();
 b15zdnd11an1n64x5 FILLER_2_2162 ();
 b15zdnd11an1n32x5 FILLER_2_2226 ();
 b15zdnd11an1n16x5 FILLER_2_2258 ();
 b15zdnd00an1n02x5 FILLER_2_2274 ();
 b15zdnd11an1n64x5 FILLER_3_0 ();
 b15zdnd11an1n64x5 FILLER_3_64 ();
 b15zdnd11an1n64x5 FILLER_3_128 ();
 b15zdnd11an1n64x5 FILLER_3_192 ();
 b15zdnd11an1n64x5 FILLER_3_256 ();
 b15zdnd11an1n64x5 FILLER_3_320 ();
 b15zdnd11an1n64x5 FILLER_3_384 ();
 b15zdnd11an1n64x5 FILLER_3_448 ();
 b15zdnd11an1n64x5 FILLER_3_512 ();
 b15zdnd11an1n64x5 FILLER_3_576 ();
 b15zdnd11an1n64x5 FILLER_3_640 ();
 b15zdnd11an1n64x5 FILLER_3_704 ();
 b15zdnd11an1n64x5 FILLER_3_768 ();
 b15zdnd11an1n64x5 FILLER_3_832 ();
 b15zdnd11an1n64x5 FILLER_3_896 ();
 b15zdnd11an1n08x5 FILLER_3_960 ();
 b15zdnd00an1n01x5 FILLER_3_968 ();
 b15zdnd11an1n08x5 FILLER_3_1011 ();
 b15zdnd00an1n02x5 FILLER_3_1019 ();
 b15zdnd11an1n64x5 FILLER_3_1063 ();
 b15zdnd11an1n64x5 FILLER_3_1127 ();
 b15zdnd11an1n64x5 FILLER_3_1191 ();
 b15zdnd11an1n64x5 FILLER_3_1255 ();
 b15zdnd11an1n64x5 FILLER_3_1319 ();
 b15zdnd11an1n64x5 FILLER_3_1383 ();
 b15zdnd11an1n64x5 FILLER_3_1447 ();
 b15zdnd11an1n64x5 FILLER_3_1511 ();
 b15zdnd11an1n64x5 FILLER_3_1575 ();
 b15zdnd11an1n64x5 FILLER_3_1639 ();
 b15zdnd11an1n64x5 FILLER_3_1703 ();
 b15zdnd11an1n64x5 FILLER_3_1767 ();
 b15zdnd11an1n64x5 FILLER_3_1831 ();
 b15zdnd11an1n16x5 FILLER_3_1895 ();
 b15zdnd11an1n08x5 FILLER_3_1911 ();
 b15zdnd00an1n02x5 FILLER_3_1919 ();
 b15zdnd00an1n01x5 FILLER_3_1921 ();
 b15zdnd11an1n16x5 FILLER_3_1926 ();
 b15zdnd11an1n08x5 FILLER_3_1942 ();
 b15zdnd11an1n64x5 FILLER_3_1954 ();
 b15zdnd11an1n08x5 FILLER_3_2018 ();
 b15zdnd11an1n64x5 FILLER_3_2068 ();
 b15zdnd11an1n64x5 FILLER_3_2132 ();
 b15zdnd11an1n64x5 FILLER_3_2196 ();
 b15zdnd11an1n16x5 FILLER_3_2260 ();
 b15zdnd11an1n08x5 FILLER_3_2276 ();
 b15zdnd11an1n64x5 FILLER_4_8 ();
 b15zdnd11an1n64x5 FILLER_4_72 ();
 b15zdnd11an1n64x5 FILLER_4_136 ();
 b15zdnd11an1n64x5 FILLER_4_200 ();
 b15zdnd11an1n64x5 FILLER_4_264 ();
 b15zdnd11an1n64x5 FILLER_4_328 ();
 b15zdnd11an1n64x5 FILLER_4_392 ();
 b15zdnd11an1n64x5 FILLER_4_456 ();
 b15zdnd11an1n64x5 FILLER_4_520 ();
 b15zdnd11an1n64x5 FILLER_4_584 ();
 b15zdnd11an1n64x5 FILLER_4_648 ();
 b15zdnd11an1n04x5 FILLER_4_712 ();
 b15zdnd00an1n02x5 FILLER_4_716 ();
 b15zdnd11an1n64x5 FILLER_4_726 ();
 b15zdnd11an1n64x5 FILLER_4_790 ();
 b15zdnd11an1n64x5 FILLER_4_854 ();
 b15zdnd11an1n64x5 FILLER_4_918 ();
 b15zdnd11an1n16x5 FILLER_4_982 ();
 b15zdnd11an1n08x5 FILLER_4_998 ();
 b15zdnd00an1n01x5 FILLER_4_1006 ();
 b15zdnd11an1n08x5 FILLER_4_1014 ();
 b15zdnd00an1n02x5 FILLER_4_1022 ();
 b15zdnd00an1n01x5 FILLER_4_1024 ();
 b15zdnd11an1n08x5 FILLER_4_1029 ();
 b15zdnd11an1n04x5 FILLER_4_1037 ();
 b15zdnd11an1n64x5 FILLER_4_1045 ();
 b15zdnd11an1n64x5 FILLER_4_1109 ();
 b15zdnd11an1n64x5 FILLER_4_1173 ();
 b15zdnd11an1n64x5 FILLER_4_1237 ();
 b15zdnd11an1n64x5 FILLER_4_1301 ();
 b15zdnd11an1n64x5 FILLER_4_1365 ();
 b15zdnd11an1n64x5 FILLER_4_1429 ();
 b15zdnd11an1n64x5 FILLER_4_1493 ();
 b15zdnd11an1n64x5 FILLER_4_1557 ();
 b15zdnd11an1n64x5 FILLER_4_1621 ();
 b15zdnd11an1n64x5 FILLER_4_1685 ();
 b15zdnd11an1n64x5 FILLER_4_1749 ();
 b15zdnd11an1n64x5 FILLER_4_1813 ();
 b15zdnd11an1n64x5 FILLER_4_1877 ();
 b15zdnd11an1n32x5 FILLER_4_1941 ();
 b15zdnd11an1n16x5 FILLER_4_1973 ();
 b15zdnd11an1n04x5 FILLER_4_1989 ();
 b15zdnd11an1n64x5 FILLER_4_2035 ();
 b15zdnd11an1n32x5 FILLER_4_2099 ();
 b15zdnd11an1n16x5 FILLER_4_2131 ();
 b15zdnd11an1n04x5 FILLER_4_2147 ();
 b15zdnd00an1n02x5 FILLER_4_2151 ();
 b15zdnd00an1n01x5 FILLER_4_2153 ();
 b15zdnd11an1n64x5 FILLER_4_2162 ();
 b15zdnd11an1n32x5 FILLER_4_2226 ();
 b15zdnd11an1n16x5 FILLER_4_2258 ();
 b15zdnd00an1n02x5 FILLER_4_2274 ();
 b15zdnd11an1n64x5 FILLER_5_0 ();
 b15zdnd11an1n64x5 FILLER_5_64 ();
 b15zdnd11an1n64x5 FILLER_5_128 ();
 b15zdnd11an1n64x5 FILLER_5_192 ();
 b15zdnd11an1n64x5 FILLER_5_256 ();
 b15zdnd11an1n64x5 FILLER_5_320 ();
 b15zdnd11an1n64x5 FILLER_5_384 ();
 b15zdnd11an1n64x5 FILLER_5_448 ();
 b15zdnd11an1n64x5 FILLER_5_512 ();
 b15zdnd11an1n64x5 FILLER_5_576 ();
 b15zdnd11an1n64x5 FILLER_5_640 ();
 b15zdnd11an1n64x5 FILLER_5_704 ();
 b15zdnd11an1n64x5 FILLER_5_768 ();
 b15zdnd11an1n64x5 FILLER_5_832 ();
 b15zdnd11an1n64x5 FILLER_5_896 ();
 b15zdnd11an1n64x5 FILLER_5_960 ();
 b15zdnd11an1n64x5 FILLER_5_1024 ();
 b15zdnd11an1n64x5 FILLER_5_1088 ();
 b15zdnd11an1n64x5 FILLER_5_1152 ();
 b15zdnd11an1n64x5 FILLER_5_1216 ();
 b15zdnd11an1n64x5 FILLER_5_1280 ();
 b15zdnd11an1n64x5 FILLER_5_1344 ();
 b15zdnd11an1n64x5 FILLER_5_1408 ();
 b15zdnd11an1n64x5 FILLER_5_1472 ();
 b15zdnd11an1n64x5 FILLER_5_1536 ();
 b15zdnd11an1n64x5 FILLER_5_1600 ();
 b15zdnd11an1n64x5 FILLER_5_1664 ();
 b15zdnd11an1n64x5 FILLER_5_1728 ();
 b15zdnd11an1n64x5 FILLER_5_1792 ();
 b15zdnd11an1n64x5 FILLER_5_1856 ();
 b15zdnd11an1n64x5 FILLER_5_1920 ();
 b15zdnd11an1n64x5 FILLER_5_1984 ();
 b15zdnd11an1n64x5 FILLER_5_2048 ();
 b15zdnd11an1n64x5 FILLER_5_2112 ();
 b15zdnd11an1n64x5 FILLER_5_2176 ();
 b15zdnd11an1n32x5 FILLER_5_2240 ();
 b15zdnd11an1n08x5 FILLER_5_2272 ();
 b15zdnd11an1n04x5 FILLER_5_2280 ();
 b15zdnd11an1n64x5 FILLER_6_8 ();
 b15zdnd11an1n64x5 FILLER_6_72 ();
 b15zdnd11an1n64x5 FILLER_6_136 ();
 b15zdnd11an1n64x5 FILLER_6_200 ();
 b15zdnd11an1n64x5 FILLER_6_264 ();
 b15zdnd11an1n64x5 FILLER_6_328 ();
 b15zdnd11an1n64x5 FILLER_6_392 ();
 b15zdnd11an1n64x5 FILLER_6_456 ();
 b15zdnd11an1n64x5 FILLER_6_520 ();
 b15zdnd11an1n64x5 FILLER_6_584 ();
 b15zdnd11an1n64x5 FILLER_6_648 ();
 b15zdnd11an1n04x5 FILLER_6_712 ();
 b15zdnd00an1n02x5 FILLER_6_716 ();
 b15zdnd11an1n64x5 FILLER_6_726 ();
 b15zdnd11an1n64x5 FILLER_6_790 ();
 b15zdnd11an1n64x5 FILLER_6_854 ();
 b15zdnd11an1n64x5 FILLER_6_918 ();
 b15zdnd11an1n64x5 FILLER_6_982 ();
 b15zdnd11an1n64x5 FILLER_6_1046 ();
 b15zdnd11an1n64x5 FILLER_6_1110 ();
 b15zdnd11an1n64x5 FILLER_6_1174 ();
 b15zdnd11an1n64x5 FILLER_6_1238 ();
 b15zdnd11an1n64x5 FILLER_6_1302 ();
 b15zdnd11an1n64x5 FILLER_6_1366 ();
 b15zdnd11an1n64x5 FILLER_6_1430 ();
 b15zdnd11an1n64x5 FILLER_6_1494 ();
 b15zdnd11an1n64x5 FILLER_6_1558 ();
 b15zdnd11an1n64x5 FILLER_6_1622 ();
 b15zdnd11an1n64x5 FILLER_6_1686 ();
 b15zdnd11an1n64x5 FILLER_6_1750 ();
 b15zdnd11an1n64x5 FILLER_6_1814 ();
 b15zdnd11an1n64x5 FILLER_6_1878 ();
 b15zdnd11an1n64x5 FILLER_6_1942 ();
 b15zdnd11an1n16x5 FILLER_6_2006 ();
 b15zdnd11an1n04x5 FILLER_6_2022 ();
 b15zdnd00an1n02x5 FILLER_6_2026 ();
 b15zdnd00an1n01x5 FILLER_6_2028 ();
 b15zdnd11an1n04x5 FILLER_6_2071 ();
 b15zdnd11an1n32x5 FILLER_6_2117 ();
 b15zdnd11an1n04x5 FILLER_6_2149 ();
 b15zdnd00an1n01x5 FILLER_6_2153 ();
 b15zdnd11an1n64x5 FILLER_6_2162 ();
 b15zdnd11an1n32x5 FILLER_6_2226 ();
 b15zdnd11an1n16x5 FILLER_6_2258 ();
 b15zdnd00an1n02x5 FILLER_6_2274 ();
 b15zdnd11an1n64x5 FILLER_7_0 ();
 b15zdnd11an1n64x5 FILLER_7_64 ();
 b15zdnd11an1n32x5 FILLER_7_128 ();
 b15zdnd11an1n08x5 FILLER_7_160 ();
 b15zdnd00an1n02x5 FILLER_7_168 ();
 b15zdnd00an1n01x5 FILLER_7_170 ();
 b15zdnd11an1n64x5 FILLER_7_174 ();
 b15zdnd11an1n08x5 FILLER_7_238 ();
 b15zdnd11an1n04x5 FILLER_7_246 ();
 b15zdnd00an1n02x5 FILLER_7_250 ();
 b15zdnd00an1n01x5 FILLER_7_252 ();
 b15zdnd11an1n08x5 FILLER_7_256 ();
 b15zdnd11an1n64x5 FILLER_7_267 ();
 b15zdnd11an1n64x5 FILLER_7_331 ();
 b15zdnd11an1n64x5 FILLER_7_395 ();
 b15zdnd11an1n64x5 FILLER_7_459 ();
 b15zdnd11an1n64x5 FILLER_7_523 ();
 b15zdnd11an1n64x5 FILLER_7_587 ();
 b15zdnd11an1n64x5 FILLER_7_651 ();
 b15zdnd11an1n64x5 FILLER_7_715 ();
 b15zdnd11an1n64x5 FILLER_7_779 ();
 b15zdnd11an1n64x5 FILLER_7_843 ();
 b15zdnd11an1n64x5 FILLER_7_907 ();
 b15zdnd11an1n64x5 FILLER_7_971 ();
 b15zdnd11an1n64x5 FILLER_7_1035 ();
 b15zdnd11an1n64x5 FILLER_7_1099 ();
 b15zdnd11an1n64x5 FILLER_7_1163 ();
 b15zdnd11an1n64x5 FILLER_7_1227 ();
 b15zdnd11an1n64x5 FILLER_7_1291 ();
 b15zdnd11an1n64x5 FILLER_7_1355 ();
 b15zdnd11an1n64x5 FILLER_7_1419 ();
 b15zdnd11an1n64x5 FILLER_7_1483 ();
 b15zdnd11an1n64x5 FILLER_7_1547 ();
 b15zdnd11an1n64x5 FILLER_7_1611 ();
 b15zdnd11an1n64x5 FILLER_7_1675 ();
 b15zdnd11an1n64x5 FILLER_7_1739 ();
 b15zdnd11an1n64x5 FILLER_7_1803 ();
 b15zdnd11an1n64x5 FILLER_7_1867 ();
 b15zdnd11an1n64x5 FILLER_7_1931 ();
 b15zdnd11an1n64x5 FILLER_7_1995 ();
 b15zdnd11an1n64x5 FILLER_7_2059 ();
 b15zdnd11an1n64x5 FILLER_7_2123 ();
 b15zdnd11an1n64x5 FILLER_7_2187 ();
 b15zdnd11an1n32x5 FILLER_7_2251 ();
 b15zdnd00an1n01x5 FILLER_7_2283 ();
 b15zdnd11an1n64x5 FILLER_8_8 ();
 b15zdnd11an1n64x5 FILLER_8_72 ();
 b15zdnd11an1n32x5 FILLER_8_136 ();
 b15zdnd00an1n01x5 FILLER_8_168 ();
 b15zdnd11an1n64x5 FILLER_8_172 ();
 b15zdnd11an1n16x5 FILLER_8_236 ();
 b15zdnd00an1n02x5 FILLER_8_252 ();
 b15zdnd00an1n01x5 FILLER_8_254 ();
 b15zdnd11an1n08x5 FILLER_8_258 ();
 b15zdnd11an1n64x5 FILLER_8_269 ();
 b15zdnd11an1n64x5 FILLER_8_333 ();
 b15zdnd11an1n64x5 FILLER_8_397 ();
 b15zdnd11an1n64x5 FILLER_8_461 ();
 b15zdnd11an1n64x5 FILLER_8_525 ();
 b15zdnd11an1n64x5 FILLER_8_589 ();
 b15zdnd11an1n64x5 FILLER_8_653 ();
 b15zdnd00an1n01x5 FILLER_8_717 ();
 b15zdnd11an1n64x5 FILLER_8_726 ();
 b15zdnd11an1n64x5 FILLER_8_790 ();
 b15zdnd11an1n64x5 FILLER_8_854 ();
 b15zdnd11an1n64x5 FILLER_8_918 ();
 b15zdnd11an1n64x5 FILLER_8_982 ();
 b15zdnd11an1n64x5 FILLER_8_1046 ();
 b15zdnd11an1n64x5 FILLER_8_1110 ();
 b15zdnd11an1n64x5 FILLER_8_1174 ();
 b15zdnd11an1n64x5 FILLER_8_1238 ();
 b15zdnd11an1n64x5 FILLER_8_1302 ();
 b15zdnd11an1n64x5 FILLER_8_1366 ();
 b15zdnd11an1n64x5 FILLER_8_1430 ();
 b15zdnd11an1n64x5 FILLER_8_1494 ();
 b15zdnd11an1n64x5 FILLER_8_1558 ();
 b15zdnd11an1n64x5 FILLER_8_1622 ();
 b15zdnd11an1n64x5 FILLER_8_1686 ();
 b15zdnd11an1n64x5 FILLER_8_1750 ();
 b15zdnd11an1n64x5 FILLER_8_1814 ();
 b15zdnd11an1n64x5 FILLER_8_1878 ();
 b15zdnd11an1n64x5 FILLER_8_1942 ();
 b15zdnd11an1n64x5 FILLER_8_2006 ();
 b15zdnd11an1n64x5 FILLER_8_2070 ();
 b15zdnd11an1n16x5 FILLER_8_2134 ();
 b15zdnd11an1n04x5 FILLER_8_2150 ();
 b15zdnd11an1n64x5 FILLER_8_2162 ();
 b15zdnd11an1n32x5 FILLER_8_2226 ();
 b15zdnd11an1n16x5 FILLER_8_2258 ();
 b15zdnd00an1n02x5 FILLER_8_2274 ();
 b15zdnd11an1n64x5 FILLER_9_0 ();
 b15zdnd11an1n64x5 FILLER_9_64 ();
 b15zdnd11an1n64x5 FILLER_9_128 ();
 b15zdnd11an1n64x5 FILLER_9_192 ();
 b15zdnd11an1n64x5 FILLER_9_256 ();
 b15zdnd11an1n64x5 FILLER_9_320 ();
 b15zdnd11an1n64x5 FILLER_9_384 ();
 b15zdnd11an1n64x5 FILLER_9_448 ();
 b15zdnd11an1n64x5 FILLER_9_512 ();
 b15zdnd11an1n64x5 FILLER_9_576 ();
 b15zdnd11an1n64x5 FILLER_9_640 ();
 b15zdnd11an1n64x5 FILLER_9_704 ();
 b15zdnd11an1n64x5 FILLER_9_768 ();
 b15zdnd11an1n64x5 FILLER_9_832 ();
 b15zdnd11an1n64x5 FILLER_9_896 ();
 b15zdnd11an1n64x5 FILLER_9_960 ();
 b15zdnd11an1n64x5 FILLER_9_1024 ();
 b15zdnd11an1n64x5 FILLER_9_1088 ();
 b15zdnd11an1n16x5 FILLER_9_1152 ();
 b15zdnd11an1n08x5 FILLER_9_1168 ();
 b15zdnd11an1n04x5 FILLER_9_1176 ();
 b15zdnd00an1n02x5 FILLER_9_1180 ();
 b15zdnd11an1n64x5 FILLER_9_1186 ();
 b15zdnd11an1n64x5 FILLER_9_1250 ();
 b15zdnd11an1n32x5 FILLER_9_1314 ();
 b15zdnd11an1n08x5 FILLER_9_1346 ();
 b15zdnd00an1n01x5 FILLER_9_1354 ();
 b15zdnd11an1n08x5 FILLER_9_1397 ();
 b15zdnd00an1n01x5 FILLER_9_1405 ();
 b15zdnd11an1n64x5 FILLER_9_1448 ();
 b15zdnd11an1n64x5 FILLER_9_1512 ();
 b15zdnd11an1n64x5 FILLER_9_1576 ();
 b15zdnd11an1n64x5 FILLER_9_1640 ();
 b15zdnd11an1n64x5 FILLER_9_1704 ();
 b15zdnd11an1n64x5 FILLER_9_1768 ();
 b15zdnd11an1n64x5 FILLER_9_1832 ();
 b15zdnd11an1n64x5 FILLER_9_1896 ();
 b15zdnd11an1n64x5 FILLER_9_1960 ();
 b15zdnd11an1n32x5 FILLER_9_2024 ();
 b15zdnd11an1n16x5 FILLER_9_2056 ();
 b15zdnd11an1n08x5 FILLER_9_2072 ();
 b15zdnd00an1n02x5 FILLER_9_2080 ();
 b15zdnd00an1n01x5 FILLER_9_2082 ();
 b15zdnd11an1n04x5 FILLER_9_2125 ();
 b15zdnd11an1n64x5 FILLER_9_2171 ();
 b15zdnd11an1n32x5 FILLER_9_2235 ();
 b15zdnd11an1n16x5 FILLER_9_2267 ();
 b15zdnd00an1n01x5 FILLER_9_2283 ();
 b15zdnd11an1n64x5 FILLER_10_8 ();
 b15zdnd11an1n64x5 FILLER_10_72 ();
 b15zdnd11an1n64x5 FILLER_10_136 ();
 b15zdnd11an1n64x5 FILLER_10_200 ();
 b15zdnd11an1n64x5 FILLER_10_264 ();
 b15zdnd11an1n64x5 FILLER_10_328 ();
 b15zdnd11an1n64x5 FILLER_10_392 ();
 b15zdnd11an1n64x5 FILLER_10_456 ();
 b15zdnd11an1n64x5 FILLER_10_520 ();
 b15zdnd11an1n64x5 FILLER_10_584 ();
 b15zdnd11an1n64x5 FILLER_10_648 ();
 b15zdnd11an1n04x5 FILLER_10_712 ();
 b15zdnd00an1n02x5 FILLER_10_716 ();
 b15zdnd11an1n64x5 FILLER_10_726 ();
 b15zdnd11an1n64x5 FILLER_10_790 ();
 b15zdnd11an1n64x5 FILLER_10_854 ();
 b15zdnd11an1n64x5 FILLER_10_918 ();
 b15zdnd11an1n64x5 FILLER_10_982 ();
 b15zdnd11an1n64x5 FILLER_10_1046 ();
 b15zdnd11an1n16x5 FILLER_10_1110 ();
 b15zdnd11an1n04x5 FILLER_10_1126 ();
 b15zdnd00an1n01x5 FILLER_10_1130 ();
 b15zdnd11an1n64x5 FILLER_10_1134 ();
 b15zdnd11an1n64x5 FILLER_10_1198 ();
 b15zdnd11an1n64x5 FILLER_10_1262 ();
 b15zdnd11an1n64x5 FILLER_10_1326 ();
 b15zdnd11an1n64x5 FILLER_10_1390 ();
 b15zdnd11an1n64x5 FILLER_10_1454 ();
 b15zdnd11an1n64x5 FILLER_10_1518 ();
 b15zdnd11an1n64x5 FILLER_10_1582 ();
 b15zdnd11an1n64x5 FILLER_10_1646 ();
 b15zdnd11an1n64x5 FILLER_10_1710 ();
 b15zdnd11an1n64x5 FILLER_10_1774 ();
 b15zdnd11an1n64x5 FILLER_10_1838 ();
 b15zdnd11an1n64x5 FILLER_10_1902 ();
 b15zdnd11an1n64x5 FILLER_10_1966 ();
 b15zdnd11an1n64x5 FILLER_10_2030 ();
 b15zdnd11an1n32x5 FILLER_10_2094 ();
 b15zdnd11an1n16x5 FILLER_10_2126 ();
 b15zdnd11an1n08x5 FILLER_10_2142 ();
 b15zdnd11an1n04x5 FILLER_10_2150 ();
 b15zdnd11an1n64x5 FILLER_10_2162 ();
 b15zdnd11an1n32x5 FILLER_10_2226 ();
 b15zdnd11an1n16x5 FILLER_10_2258 ();
 b15zdnd00an1n02x5 FILLER_10_2274 ();
 b15zdnd11an1n64x5 FILLER_11_0 ();
 b15zdnd11an1n64x5 FILLER_11_64 ();
 b15zdnd11an1n64x5 FILLER_11_128 ();
 b15zdnd11an1n64x5 FILLER_11_192 ();
 b15zdnd11an1n64x5 FILLER_11_256 ();
 b15zdnd11an1n64x5 FILLER_11_320 ();
 b15zdnd11an1n64x5 FILLER_11_384 ();
 b15zdnd11an1n64x5 FILLER_11_448 ();
 b15zdnd11an1n64x5 FILLER_11_512 ();
 b15zdnd11an1n64x5 FILLER_11_576 ();
 b15zdnd11an1n64x5 FILLER_11_640 ();
 b15zdnd11an1n64x5 FILLER_11_704 ();
 b15zdnd11an1n64x5 FILLER_11_768 ();
 b15zdnd11an1n64x5 FILLER_11_832 ();
 b15zdnd11an1n64x5 FILLER_11_896 ();
 b15zdnd11an1n64x5 FILLER_11_960 ();
 b15zdnd11an1n64x5 FILLER_11_1024 ();
 b15zdnd11an1n16x5 FILLER_11_1088 ();
 b15zdnd11an1n04x5 FILLER_11_1104 ();
 b15zdnd00an1n01x5 FILLER_11_1108 ();
 b15zdnd11an1n04x5 FILLER_11_1136 ();
 b15zdnd00an1n01x5 FILLER_11_1140 ();
 b15zdnd11an1n64x5 FILLER_11_1144 ();
 b15zdnd11an1n64x5 FILLER_11_1208 ();
 b15zdnd11an1n64x5 FILLER_11_1272 ();
 b15zdnd11an1n64x5 FILLER_11_1336 ();
 b15zdnd11an1n64x5 FILLER_11_1400 ();
 b15zdnd11an1n64x5 FILLER_11_1464 ();
 b15zdnd11an1n64x5 FILLER_11_1528 ();
 b15zdnd11an1n64x5 FILLER_11_1592 ();
 b15zdnd11an1n64x5 FILLER_11_1656 ();
 b15zdnd11an1n64x5 FILLER_11_1720 ();
 b15zdnd11an1n64x5 FILLER_11_1784 ();
 b15zdnd11an1n64x5 FILLER_11_1848 ();
 b15zdnd11an1n64x5 FILLER_11_1912 ();
 b15zdnd11an1n64x5 FILLER_11_1976 ();
 b15zdnd11an1n64x5 FILLER_11_2040 ();
 b15zdnd11an1n16x5 FILLER_11_2104 ();
 b15zdnd11an1n08x5 FILLER_11_2120 ();
 b15zdnd11an1n04x5 FILLER_11_2128 ();
 b15zdnd11an1n64x5 FILLER_11_2184 ();
 b15zdnd11an1n32x5 FILLER_11_2248 ();
 b15zdnd11an1n04x5 FILLER_11_2280 ();
 b15zdnd11an1n64x5 FILLER_12_8 ();
 b15zdnd11an1n64x5 FILLER_12_72 ();
 b15zdnd11an1n64x5 FILLER_12_136 ();
 b15zdnd11an1n64x5 FILLER_12_200 ();
 b15zdnd11an1n64x5 FILLER_12_264 ();
 b15zdnd11an1n64x5 FILLER_12_328 ();
 b15zdnd11an1n64x5 FILLER_12_392 ();
 b15zdnd11an1n64x5 FILLER_12_456 ();
 b15zdnd11an1n64x5 FILLER_12_520 ();
 b15zdnd11an1n64x5 FILLER_12_584 ();
 b15zdnd11an1n64x5 FILLER_12_648 ();
 b15zdnd11an1n04x5 FILLER_12_712 ();
 b15zdnd00an1n02x5 FILLER_12_716 ();
 b15zdnd11an1n64x5 FILLER_12_726 ();
 b15zdnd11an1n64x5 FILLER_12_790 ();
 b15zdnd11an1n64x5 FILLER_12_854 ();
 b15zdnd11an1n64x5 FILLER_12_918 ();
 b15zdnd11an1n64x5 FILLER_12_982 ();
 b15zdnd11an1n32x5 FILLER_12_1046 ();
 b15zdnd11an1n16x5 FILLER_12_1078 ();
 b15zdnd11an1n08x5 FILLER_12_1094 ();
 b15zdnd11an1n04x5 FILLER_12_1102 ();
 b15zdnd00an1n02x5 FILLER_12_1106 ();
 b15zdnd11an1n04x5 FILLER_12_1111 ();
 b15zdnd11an1n04x5 FILLER_12_1147 ();
 b15zdnd11an1n64x5 FILLER_12_1154 ();
 b15zdnd11an1n64x5 FILLER_12_1218 ();
 b15zdnd11an1n64x5 FILLER_12_1282 ();
 b15zdnd11an1n64x5 FILLER_12_1346 ();
 b15zdnd11an1n64x5 FILLER_12_1410 ();
 b15zdnd11an1n64x5 FILLER_12_1474 ();
 b15zdnd11an1n64x5 FILLER_12_1538 ();
 b15zdnd11an1n64x5 FILLER_12_1602 ();
 b15zdnd11an1n64x5 FILLER_12_1666 ();
 b15zdnd11an1n64x5 FILLER_12_1730 ();
 b15zdnd11an1n64x5 FILLER_12_1794 ();
 b15zdnd11an1n64x5 FILLER_12_1858 ();
 b15zdnd11an1n64x5 FILLER_12_1922 ();
 b15zdnd11an1n64x5 FILLER_12_1986 ();
 b15zdnd11an1n64x5 FILLER_12_2050 ();
 b15zdnd11an1n32x5 FILLER_12_2114 ();
 b15zdnd00an1n02x5 FILLER_12_2146 ();
 b15zdnd00an1n01x5 FILLER_12_2148 ();
 b15zdnd00an1n02x5 FILLER_12_2152 ();
 b15zdnd00an1n02x5 FILLER_12_2162 ();
 b15zdnd11an1n64x5 FILLER_12_2167 ();
 b15zdnd11an1n32x5 FILLER_12_2231 ();
 b15zdnd11an1n08x5 FILLER_12_2263 ();
 b15zdnd11an1n04x5 FILLER_12_2271 ();
 b15zdnd00an1n01x5 FILLER_12_2275 ();
 b15zdnd11an1n64x5 FILLER_13_0 ();
 b15zdnd11an1n64x5 FILLER_13_64 ();
 b15zdnd11an1n64x5 FILLER_13_128 ();
 b15zdnd11an1n64x5 FILLER_13_192 ();
 b15zdnd11an1n64x5 FILLER_13_256 ();
 b15zdnd11an1n32x5 FILLER_13_320 ();
 b15zdnd11an1n08x5 FILLER_13_352 ();
 b15zdnd11an1n64x5 FILLER_13_363 ();
 b15zdnd11an1n32x5 FILLER_13_427 ();
 b15zdnd11an1n08x5 FILLER_13_459 ();
 b15zdnd11an1n04x5 FILLER_13_467 ();
 b15zdnd00an1n02x5 FILLER_13_471 ();
 b15zdnd11an1n64x5 FILLER_13_476 ();
 b15zdnd11an1n64x5 FILLER_13_540 ();
 b15zdnd11an1n64x5 FILLER_13_604 ();
 b15zdnd11an1n64x5 FILLER_13_668 ();
 b15zdnd11an1n64x5 FILLER_13_732 ();
 b15zdnd11an1n64x5 FILLER_13_796 ();
 b15zdnd11an1n64x5 FILLER_13_860 ();
 b15zdnd11an1n64x5 FILLER_13_924 ();
 b15zdnd11an1n64x5 FILLER_13_988 ();
 b15zdnd11an1n32x5 FILLER_13_1052 ();
 b15zdnd11an1n16x5 FILLER_13_1084 ();
 b15zdnd11an1n04x5 FILLER_13_1100 ();
 b15zdnd00an1n01x5 FILLER_13_1104 ();
 b15zdnd11an1n64x5 FILLER_13_1157 ();
 b15zdnd11an1n64x5 FILLER_13_1221 ();
 b15zdnd11an1n64x5 FILLER_13_1285 ();
 b15zdnd11an1n64x5 FILLER_13_1349 ();
 b15zdnd11an1n64x5 FILLER_13_1413 ();
 b15zdnd11an1n64x5 FILLER_13_1477 ();
 b15zdnd11an1n64x5 FILLER_13_1541 ();
 b15zdnd11an1n64x5 FILLER_13_1605 ();
 b15zdnd11an1n64x5 FILLER_13_1669 ();
 b15zdnd11an1n64x5 FILLER_13_1733 ();
 b15zdnd11an1n64x5 FILLER_13_1797 ();
 b15zdnd11an1n64x5 FILLER_13_1861 ();
 b15zdnd11an1n64x5 FILLER_13_1925 ();
 b15zdnd11an1n64x5 FILLER_13_1989 ();
 b15zdnd11an1n64x5 FILLER_13_2053 ();
 b15zdnd11an1n08x5 FILLER_13_2117 ();
 b15zdnd00an1n02x5 FILLER_13_2125 ();
 b15zdnd11an1n64x5 FILLER_13_2179 ();
 b15zdnd11an1n32x5 FILLER_13_2243 ();
 b15zdnd11an1n08x5 FILLER_13_2275 ();
 b15zdnd00an1n01x5 FILLER_13_2283 ();
 b15zdnd11an1n64x5 FILLER_14_8 ();
 b15zdnd11an1n64x5 FILLER_14_72 ();
 b15zdnd11an1n64x5 FILLER_14_136 ();
 b15zdnd11an1n64x5 FILLER_14_200 ();
 b15zdnd11an1n64x5 FILLER_14_264 ();
 b15zdnd11an1n32x5 FILLER_14_328 ();
 b15zdnd11an1n32x5 FILLER_14_387 ();
 b15zdnd11an1n16x5 FILLER_14_419 ();
 b15zdnd11an1n08x5 FILLER_14_435 ();
 b15zdnd00an1n02x5 FILLER_14_443 ();
 b15zdnd00an1n01x5 FILLER_14_445 ();
 b15zdnd11an1n64x5 FILLER_14_498 ();
 b15zdnd11an1n64x5 FILLER_14_562 ();
 b15zdnd11an1n64x5 FILLER_14_626 ();
 b15zdnd11an1n16x5 FILLER_14_690 ();
 b15zdnd11an1n08x5 FILLER_14_706 ();
 b15zdnd11an1n04x5 FILLER_14_714 ();
 b15zdnd11an1n64x5 FILLER_14_726 ();
 b15zdnd11an1n64x5 FILLER_14_790 ();
 b15zdnd11an1n64x5 FILLER_14_854 ();
 b15zdnd11an1n64x5 FILLER_14_918 ();
 b15zdnd11an1n64x5 FILLER_14_982 ();
 b15zdnd11an1n64x5 FILLER_14_1046 ();
 b15zdnd00an1n02x5 FILLER_14_1110 ();
 b15zdnd00an1n01x5 FILLER_14_1112 ();
 b15zdnd11an1n04x5 FILLER_14_1145 ();
 b15zdnd11an1n64x5 FILLER_14_1152 ();
 b15zdnd11an1n64x5 FILLER_14_1216 ();
 b15zdnd11an1n64x5 FILLER_14_1280 ();
 b15zdnd00an1n02x5 FILLER_14_1344 ();
 b15zdnd11an1n64x5 FILLER_14_1349 ();
 b15zdnd11an1n64x5 FILLER_14_1413 ();
 b15zdnd11an1n64x5 FILLER_14_1477 ();
 b15zdnd11an1n64x5 FILLER_14_1541 ();
 b15zdnd11an1n64x5 FILLER_14_1605 ();
 b15zdnd11an1n64x5 FILLER_14_1669 ();
 b15zdnd11an1n64x5 FILLER_14_1733 ();
 b15zdnd11an1n64x5 FILLER_14_1797 ();
 b15zdnd11an1n64x5 FILLER_14_1861 ();
 b15zdnd11an1n64x5 FILLER_14_1925 ();
 b15zdnd11an1n64x5 FILLER_14_1989 ();
 b15zdnd11an1n64x5 FILLER_14_2053 ();
 b15zdnd11an1n16x5 FILLER_14_2117 ();
 b15zdnd11an1n08x5 FILLER_14_2133 ();
 b15zdnd00an1n01x5 FILLER_14_2141 ();
 b15zdnd11an1n04x5 FILLER_14_2145 ();
 b15zdnd00an1n02x5 FILLER_14_2152 ();
 b15zdnd00an1n02x5 FILLER_14_2162 ();
 b15zdnd11an1n32x5 FILLER_14_2167 ();
 b15zdnd11an1n08x5 FILLER_14_2199 ();
 b15zdnd00an1n02x5 FILLER_14_2207 ();
 b15zdnd00an1n01x5 FILLER_14_2209 ();
 b15zdnd11an1n32x5 FILLER_14_2218 ();
 b15zdnd11an1n16x5 FILLER_14_2250 ();
 b15zdnd11an1n08x5 FILLER_14_2266 ();
 b15zdnd00an1n02x5 FILLER_14_2274 ();
 b15zdnd11an1n64x5 FILLER_15_0 ();
 b15zdnd11an1n64x5 FILLER_15_64 ();
 b15zdnd11an1n64x5 FILLER_15_128 ();
 b15zdnd11an1n64x5 FILLER_15_192 ();
 b15zdnd11an1n64x5 FILLER_15_256 ();
 b15zdnd11an1n32x5 FILLER_15_320 ();
 b15zdnd11an1n16x5 FILLER_15_352 ();
 b15zdnd11an1n04x5 FILLER_15_368 ();
 b15zdnd00an1n01x5 FILLER_15_372 ();
 b15zdnd11an1n32x5 FILLER_15_425 ();
 b15zdnd11an1n16x5 FILLER_15_457 ();
 b15zdnd11an1n08x5 FILLER_15_476 ();
 b15zdnd00an1n02x5 FILLER_15_484 ();
 b15zdnd00an1n01x5 FILLER_15_486 ();
 b15zdnd11an1n04x5 FILLER_15_490 ();
 b15zdnd00an1n02x5 FILLER_15_494 ();
 b15zdnd00an1n01x5 FILLER_15_496 ();
 b15zdnd11an1n04x5 FILLER_15_500 ();
 b15zdnd00an1n02x5 FILLER_15_504 ();
 b15zdnd11an1n64x5 FILLER_15_509 ();
 b15zdnd11an1n64x5 FILLER_15_573 ();
 b15zdnd11an1n64x5 FILLER_15_637 ();
 b15zdnd11an1n64x5 FILLER_15_701 ();
 b15zdnd11an1n64x5 FILLER_15_765 ();
 b15zdnd11an1n64x5 FILLER_15_829 ();
 b15zdnd11an1n64x5 FILLER_15_893 ();
 b15zdnd11an1n64x5 FILLER_15_957 ();
 b15zdnd11an1n64x5 FILLER_15_1021 ();
 b15zdnd11an1n32x5 FILLER_15_1085 ();
 b15zdnd00an1n02x5 FILLER_15_1117 ();
 b15zdnd00an1n01x5 FILLER_15_1119 ();
 b15zdnd11an1n04x5 FILLER_15_1123 ();
 b15zdnd11an1n04x5 FILLER_15_1136 ();
 b15zdnd00an1n02x5 FILLER_15_1140 ();
 b15zdnd00an1n01x5 FILLER_15_1142 ();
 b15zdnd11an1n08x5 FILLER_15_1146 ();
 b15zdnd00an1n01x5 FILLER_15_1154 ();
 b15zdnd11an1n64x5 FILLER_15_1197 ();
 b15zdnd11an1n32x5 FILLER_15_1261 ();
 b15zdnd11an1n16x5 FILLER_15_1293 ();
 b15zdnd11an1n08x5 FILLER_15_1309 ();
 b15zdnd00an1n02x5 FILLER_15_1317 ();
 b15zdnd00an1n01x5 FILLER_15_1319 ();
 b15zdnd11an1n64x5 FILLER_15_1372 ();
 b15zdnd11an1n64x5 FILLER_15_1436 ();
 b15zdnd11an1n64x5 FILLER_15_1500 ();
 b15zdnd11an1n64x5 FILLER_15_1564 ();
 b15zdnd11an1n64x5 FILLER_15_1628 ();
 b15zdnd11an1n64x5 FILLER_15_1692 ();
 b15zdnd11an1n64x5 FILLER_15_1756 ();
 b15zdnd11an1n64x5 FILLER_15_1820 ();
 b15zdnd11an1n64x5 FILLER_15_1884 ();
 b15zdnd11an1n64x5 FILLER_15_1948 ();
 b15zdnd11an1n64x5 FILLER_15_2012 ();
 b15zdnd11an1n64x5 FILLER_15_2076 ();
 b15zdnd11an1n08x5 FILLER_15_2140 ();
 b15zdnd11an1n04x5 FILLER_15_2148 ();
 b15zdnd11an1n64x5 FILLER_15_2155 ();
 b15zdnd11an1n64x5 FILLER_15_2219 ();
 b15zdnd00an1n01x5 FILLER_15_2283 ();
 b15zdnd11an1n64x5 FILLER_16_8 ();
 b15zdnd11an1n64x5 FILLER_16_72 ();
 b15zdnd11an1n64x5 FILLER_16_136 ();
 b15zdnd11an1n64x5 FILLER_16_200 ();
 b15zdnd11an1n64x5 FILLER_16_264 ();
 b15zdnd11an1n64x5 FILLER_16_328 ();
 b15zdnd00an1n01x5 FILLER_16_392 ();
 b15zdnd11an1n04x5 FILLER_16_396 ();
 b15zdnd11an1n64x5 FILLER_16_403 ();
 b15zdnd11an1n08x5 FILLER_16_470 ();
 b15zdnd00an1n02x5 FILLER_16_478 ();
 b15zdnd00an1n01x5 FILLER_16_480 ();
 b15zdnd11an1n64x5 FILLER_16_533 ();
 b15zdnd11an1n64x5 FILLER_16_597 ();
 b15zdnd11an1n32x5 FILLER_16_661 ();
 b15zdnd11an1n16x5 FILLER_16_693 ();
 b15zdnd11an1n08x5 FILLER_16_709 ();
 b15zdnd00an1n01x5 FILLER_16_717 ();
 b15zdnd11an1n64x5 FILLER_16_726 ();
 b15zdnd11an1n64x5 FILLER_16_790 ();
 b15zdnd11an1n64x5 FILLER_16_854 ();
 b15zdnd11an1n64x5 FILLER_16_918 ();
 b15zdnd11an1n64x5 FILLER_16_982 ();
 b15zdnd11an1n32x5 FILLER_16_1046 ();
 b15zdnd11an1n16x5 FILLER_16_1078 ();
 b15zdnd11an1n08x5 FILLER_16_1094 ();
 b15zdnd00an1n02x5 FILLER_16_1102 ();
 b15zdnd11an1n64x5 FILLER_16_1146 ();
 b15zdnd11an1n64x5 FILLER_16_1210 ();
 b15zdnd11an1n64x5 FILLER_16_1274 ();
 b15zdnd11an1n04x5 FILLER_16_1338 ();
 b15zdnd00an1n02x5 FILLER_16_1342 ();
 b15zdnd00an1n01x5 FILLER_16_1344 ();
 b15zdnd11an1n04x5 FILLER_16_1348 ();
 b15zdnd11an1n08x5 FILLER_16_1355 ();
 b15zdnd00an1n01x5 FILLER_16_1363 ();
 b15zdnd11an1n64x5 FILLER_16_1406 ();
 b15zdnd11an1n64x5 FILLER_16_1470 ();
 b15zdnd11an1n64x5 FILLER_16_1534 ();
 b15zdnd11an1n32x5 FILLER_16_1598 ();
 b15zdnd11an1n64x5 FILLER_16_1654 ();
 b15zdnd11an1n64x5 FILLER_16_1718 ();
 b15zdnd11an1n64x5 FILLER_16_1782 ();
 b15zdnd11an1n64x5 FILLER_16_1846 ();
 b15zdnd11an1n64x5 FILLER_16_1910 ();
 b15zdnd11an1n64x5 FILLER_16_1974 ();
 b15zdnd11an1n64x5 FILLER_16_2038 ();
 b15zdnd11an1n32x5 FILLER_16_2102 ();
 b15zdnd11an1n16x5 FILLER_16_2134 ();
 b15zdnd11an1n04x5 FILLER_16_2150 ();
 b15zdnd11an1n64x5 FILLER_16_2162 ();
 b15zdnd11an1n32x5 FILLER_16_2226 ();
 b15zdnd11an1n16x5 FILLER_16_2258 ();
 b15zdnd00an1n02x5 FILLER_16_2274 ();
 b15zdnd11an1n64x5 FILLER_17_0 ();
 b15zdnd11an1n64x5 FILLER_17_64 ();
 b15zdnd11an1n64x5 FILLER_17_128 ();
 b15zdnd11an1n64x5 FILLER_17_192 ();
 b15zdnd11an1n64x5 FILLER_17_256 ();
 b15zdnd11an1n64x5 FILLER_17_320 ();
 b15zdnd11an1n08x5 FILLER_17_384 ();
 b15zdnd11an1n04x5 FILLER_17_392 ();
 b15zdnd00an1n02x5 FILLER_17_396 ();
 b15zdnd11an1n64x5 FILLER_17_401 ();
 b15zdnd11an1n64x5 FILLER_17_465 ();
 b15zdnd11an1n64x5 FILLER_17_529 ();
 b15zdnd11an1n64x5 FILLER_17_593 ();
 b15zdnd11an1n64x5 FILLER_17_657 ();
 b15zdnd11an1n64x5 FILLER_17_721 ();
 b15zdnd11an1n64x5 FILLER_17_785 ();
 b15zdnd11an1n64x5 FILLER_17_849 ();
 b15zdnd11an1n32x5 FILLER_17_913 ();
 b15zdnd11an1n08x5 FILLER_17_945 ();
 b15zdnd11an1n04x5 FILLER_17_956 ();
 b15zdnd11an1n64x5 FILLER_17_963 ();
 b15zdnd11an1n64x5 FILLER_17_1027 ();
 b15zdnd11an1n32x5 FILLER_17_1091 ();
 b15zdnd11an1n08x5 FILLER_17_1123 ();
 b15zdnd00an1n01x5 FILLER_17_1131 ();
 b15zdnd11an1n64x5 FILLER_17_1135 ();
 b15zdnd11an1n64x5 FILLER_17_1199 ();
 b15zdnd11an1n64x5 FILLER_17_1263 ();
 b15zdnd11an1n08x5 FILLER_17_1327 ();
 b15zdnd11an1n04x5 FILLER_17_1335 ();
 b15zdnd00an1n01x5 FILLER_17_1339 ();
 b15zdnd11an1n04x5 FILLER_17_1382 ();
 b15zdnd00an1n02x5 FILLER_17_1386 ();
 b15zdnd00an1n01x5 FILLER_17_1388 ();
 b15zdnd11an1n64x5 FILLER_17_1431 ();
 b15zdnd11an1n64x5 FILLER_17_1495 ();
 b15zdnd11an1n64x5 FILLER_17_1559 ();
 b15zdnd11an1n64x5 FILLER_17_1623 ();
 b15zdnd11an1n64x5 FILLER_17_1687 ();
 b15zdnd11an1n64x5 FILLER_17_1751 ();
 b15zdnd11an1n64x5 FILLER_17_1815 ();
 b15zdnd11an1n64x5 FILLER_17_1879 ();
 b15zdnd11an1n64x5 FILLER_17_1943 ();
 b15zdnd11an1n64x5 FILLER_17_2007 ();
 b15zdnd11an1n64x5 FILLER_17_2071 ();
 b15zdnd11an1n64x5 FILLER_17_2135 ();
 b15zdnd11an1n64x5 FILLER_17_2199 ();
 b15zdnd11an1n16x5 FILLER_17_2263 ();
 b15zdnd11an1n04x5 FILLER_17_2279 ();
 b15zdnd00an1n01x5 FILLER_17_2283 ();
 b15zdnd11an1n64x5 FILLER_18_8 ();
 b15zdnd11an1n64x5 FILLER_18_72 ();
 b15zdnd11an1n64x5 FILLER_18_136 ();
 b15zdnd11an1n64x5 FILLER_18_200 ();
 b15zdnd11an1n64x5 FILLER_18_264 ();
 b15zdnd11an1n64x5 FILLER_18_328 ();
 b15zdnd11an1n64x5 FILLER_18_392 ();
 b15zdnd11an1n64x5 FILLER_18_456 ();
 b15zdnd11an1n64x5 FILLER_18_520 ();
 b15zdnd11an1n64x5 FILLER_18_584 ();
 b15zdnd11an1n64x5 FILLER_18_648 ();
 b15zdnd11an1n04x5 FILLER_18_712 ();
 b15zdnd00an1n02x5 FILLER_18_716 ();
 b15zdnd11an1n64x5 FILLER_18_726 ();
 b15zdnd11an1n32x5 FILLER_18_790 ();
 b15zdnd11an1n16x5 FILLER_18_822 ();
 b15zdnd11an1n04x5 FILLER_18_838 ();
 b15zdnd00an1n02x5 FILLER_18_842 ();
 b15zdnd00an1n01x5 FILLER_18_844 ();
 b15zdnd11an1n04x5 FILLER_18_848 ();
 b15zdnd11an1n16x5 FILLER_18_904 ();
 b15zdnd11an1n08x5 FILLER_18_920 ();
 b15zdnd00an1n02x5 FILLER_18_928 ();
 b15zdnd11an1n64x5 FILLER_18_982 ();
 b15zdnd11an1n64x5 FILLER_18_1046 ();
 b15zdnd11an1n64x5 FILLER_18_1110 ();
 b15zdnd11an1n64x5 FILLER_18_1174 ();
 b15zdnd11an1n16x5 FILLER_18_1238 ();
 b15zdnd11an1n08x5 FILLER_18_1254 ();
 b15zdnd11an1n64x5 FILLER_18_1266 ();
 b15zdnd11an1n32x5 FILLER_18_1330 ();
 b15zdnd11an1n16x5 FILLER_18_1362 ();
 b15zdnd11an1n08x5 FILLER_18_1378 ();
 b15zdnd11an1n04x5 FILLER_18_1386 ();
 b15zdnd00an1n02x5 FILLER_18_1390 ();
 b15zdnd00an1n01x5 FILLER_18_1392 ();
 b15zdnd11an1n64x5 FILLER_18_1435 ();
 b15zdnd11an1n64x5 FILLER_18_1499 ();
 b15zdnd11an1n64x5 FILLER_18_1563 ();
 b15zdnd11an1n64x5 FILLER_18_1627 ();
 b15zdnd11an1n64x5 FILLER_18_1691 ();
 b15zdnd11an1n64x5 FILLER_18_1755 ();
 b15zdnd11an1n64x5 FILLER_18_1819 ();
 b15zdnd11an1n64x5 FILLER_18_1883 ();
 b15zdnd11an1n64x5 FILLER_18_1947 ();
 b15zdnd11an1n64x5 FILLER_18_2011 ();
 b15zdnd11an1n64x5 FILLER_18_2075 ();
 b15zdnd11an1n08x5 FILLER_18_2139 ();
 b15zdnd11an1n04x5 FILLER_18_2147 ();
 b15zdnd00an1n02x5 FILLER_18_2151 ();
 b15zdnd00an1n01x5 FILLER_18_2153 ();
 b15zdnd11an1n64x5 FILLER_18_2162 ();
 b15zdnd11an1n32x5 FILLER_18_2226 ();
 b15zdnd11an1n16x5 FILLER_18_2258 ();
 b15zdnd00an1n02x5 FILLER_18_2274 ();
 b15zdnd11an1n64x5 FILLER_19_0 ();
 b15zdnd11an1n64x5 FILLER_19_64 ();
 b15zdnd11an1n64x5 FILLER_19_128 ();
 b15zdnd11an1n64x5 FILLER_19_192 ();
 b15zdnd11an1n64x5 FILLER_19_256 ();
 b15zdnd11an1n64x5 FILLER_19_320 ();
 b15zdnd11an1n64x5 FILLER_19_384 ();
 b15zdnd11an1n64x5 FILLER_19_448 ();
 b15zdnd11an1n64x5 FILLER_19_512 ();
 b15zdnd11an1n64x5 FILLER_19_576 ();
 b15zdnd11an1n08x5 FILLER_19_640 ();
 b15zdnd11an1n04x5 FILLER_19_648 ();
 b15zdnd11an1n64x5 FILLER_19_683 ();
 b15zdnd11an1n64x5 FILLER_19_747 ();
 b15zdnd11an1n32x5 FILLER_19_811 ();
 b15zdnd00an1n01x5 FILLER_19_843 ();
 b15zdnd11an1n04x5 FILLER_19_847 ();
 b15zdnd11an1n16x5 FILLER_19_854 ();
 b15zdnd00an1n02x5 FILLER_19_870 ();
 b15zdnd11an1n04x5 FILLER_19_875 ();
 b15zdnd11an1n04x5 FILLER_19_882 ();
 b15zdnd11an1n64x5 FILLER_19_889 ();
 b15zdnd11an1n04x5 FILLER_19_953 ();
 b15zdnd11an1n64x5 FILLER_19_960 ();
 b15zdnd11an1n64x5 FILLER_19_1024 ();
 b15zdnd11an1n64x5 FILLER_19_1088 ();
 b15zdnd11an1n64x5 FILLER_19_1152 ();
 b15zdnd11an1n64x5 FILLER_19_1216 ();
 b15zdnd11an1n64x5 FILLER_19_1280 ();
 b15zdnd11an1n32x5 FILLER_19_1344 ();
 b15zdnd11an1n08x5 FILLER_19_1376 ();
 b15zdnd00an1n02x5 FILLER_19_1384 ();
 b15zdnd11an1n64x5 FILLER_19_1438 ();
 b15zdnd11an1n64x5 FILLER_19_1502 ();
 b15zdnd11an1n64x5 FILLER_19_1566 ();
 b15zdnd11an1n64x5 FILLER_19_1630 ();
 b15zdnd11an1n64x5 FILLER_19_1694 ();
 b15zdnd11an1n64x5 FILLER_19_1758 ();
 b15zdnd11an1n64x5 FILLER_19_1822 ();
 b15zdnd11an1n64x5 FILLER_19_1886 ();
 b15zdnd11an1n64x5 FILLER_19_1950 ();
 b15zdnd11an1n64x5 FILLER_19_2014 ();
 b15zdnd11an1n64x5 FILLER_19_2078 ();
 b15zdnd11an1n64x5 FILLER_19_2142 ();
 b15zdnd11an1n64x5 FILLER_19_2206 ();
 b15zdnd11an1n08x5 FILLER_19_2270 ();
 b15zdnd11an1n04x5 FILLER_19_2278 ();
 b15zdnd00an1n02x5 FILLER_19_2282 ();
 b15zdnd11an1n64x5 FILLER_20_8 ();
 b15zdnd11an1n64x5 FILLER_20_72 ();
 b15zdnd11an1n64x5 FILLER_20_136 ();
 b15zdnd11an1n64x5 FILLER_20_200 ();
 b15zdnd11an1n64x5 FILLER_20_264 ();
 b15zdnd11an1n64x5 FILLER_20_328 ();
 b15zdnd11an1n64x5 FILLER_20_392 ();
 b15zdnd11an1n64x5 FILLER_20_456 ();
 b15zdnd11an1n64x5 FILLER_20_520 ();
 b15zdnd11an1n64x5 FILLER_20_584 ();
 b15zdnd11an1n64x5 FILLER_20_648 ();
 b15zdnd11an1n04x5 FILLER_20_712 ();
 b15zdnd00an1n02x5 FILLER_20_716 ();
 b15zdnd11an1n64x5 FILLER_20_726 ();
 b15zdnd11an1n32x5 FILLER_20_790 ();
 b15zdnd00an1n02x5 FILLER_20_822 ();
 b15zdnd11an1n64x5 FILLER_20_876 ();
 b15zdnd11an1n64x5 FILLER_20_940 ();
 b15zdnd11an1n64x5 FILLER_20_1004 ();
 b15zdnd11an1n64x5 FILLER_20_1068 ();
 b15zdnd11an1n64x5 FILLER_20_1132 ();
 b15zdnd11an1n32x5 FILLER_20_1196 ();
 b15zdnd11an1n64x5 FILLER_20_1244 ();
 b15zdnd11an1n64x5 FILLER_20_1308 ();
 b15zdnd11an1n32x5 FILLER_20_1372 ();
 b15zdnd11an1n04x5 FILLER_20_1407 ();
 b15zdnd11an1n64x5 FILLER_20_1414 ();
 b15zdnd11an1n64x5 FILLER_20_1478 ();
 b15zdnd11an1n64x5 FILLER_20_1542 ();
 b15zdnd11an1n64x5 FILLER_20_1606 ();
 b15zdnd11an1n64x5 FILLER_20_1670 ();
 b15zdnd11an1n64x5 FILLER_20_1734 ();
 b15zdnd11an1n64x5 FILLER_20_1798 ();
 b15zdnd11an1n64x5 FILLER_20_1862 ();
 b15zdnd11an1n64x5 FILLER_20_1926 ();
 b15zdnd11an1n64x5 FILLER_20_1990 ();
 b15zdnd11an1n64x5 FILLER_20_2054 ();
 b15zdnd11an1n32x5 FILLER_20_2118 ();
 b15zdnd11an1n04x5 FILLER_20_2150 ();
 b15zdnd11an1n64x5 FILLER_20_2162 ();
 b15zdnd11an1n32x5 FILLER_20_2226 ();
 b15zdnd11an1n16x5 FILLER_20_2258 ();
 b15zdnd00an1n02x5 FILLER_20_2274 ();
 b15zdnd11an1n16x5 FILLER_21_0 ();
 b15zdnd11an1n04x5 FILLER_21_16 ();
 b15zdnd00an1n01x5 FILLER_21_20 ();
 b15zdnd11an1n64x5 FILLER_21_24 ();
 b15zdnd11an1n64x5 FILLER_21_88 ();
 b15zdnd11an1n64x5 FILLER_21_152 ();
 b15zdnd11an1n64x5 FILLER_21_216 ();
 b15zdnd11an1n64x5 FILLER_21_280 ();
 b15zdnd11an1n64x5 FILLER_21_344 ();
 b15zdnd11an1n16x5 FILLER_21_408 ();
 b15zdnd11an1n08x5 FILLER_21_424 ();
 b15zdnd11an1n64x5 FILLER_21_441 ();
 b15zdnd11an1n64x5 FILLER_21_505 ();
 b15zdnd11an1n32x5 FILLER_21_569 ();
 b15zdnd11an1n16x5 FILLER_21_601 ();
 b15zdnd11an1n04x5 FILLER_21_617 ();
 b15zdnd11an1n64x5 FILLER_21_645 ();
 b15zdnd11an1n64x5 FILLER_21_709 ();
 b15zdnd11an1n32x5 FILLER_21_773 ();
 b15zdnd11an1n16x5 FILLER_21_805 ();
 b15zdnd11an1n08x5 FILLER_21_821 ();
 b15zdnd11an1n04x5 FILLER_21_829 ();
 b15zdnd00an1n01x5 FILLER_21_833 ();
 b15zdnd11an1n64x5 FILLER_21_886 ();
 b15zdnd11an1n64x5 FILLER_21_950 ();
 b15zdnd11an1n64x5 FILLER_21_1014 ();
 b15zdnd11an1n32x5 FILLER_21_1078 ();
 b15zdnd11an1n16x5 FILLER_21_1110 ();
 b15zdnd11an1n08x5 FILLER_21_1126 ();
 b15zdnd00an1n01x5 FILLER_21_1134 ();
 b15zdnd11an1n64x5 FILLER_21_1177 ();
 b15zdnd11an1n08x5 FILLER_21_1241 ();
 b15zdnd11an1n64x5 FILLER_21_1272 ();
 b15zdnd11an1n64x5 FILLER_21_1336 ();
 b15zdnd11an1n08x5 FILLER_21_1400 ();
 b15zdnd00an1n01x5 FILLER_21_1408 ();
 b15zdnd11an1n64x5 FILLER_21_1412 ();
 b15zdnd11an1n64x5 FILLER_21_1476 ();
 b15zdnd11an1n64x5 FILLER_21_1540 ();
 b15zdnd11an1n64x5 FILLER_21_1604 ();
 b15zdnd11an1n64x5 FILLER_21_1668 ();
 b15zdnd11an1n64x5 FILLER_21_1732 ();
 b15zdnd11an1n64x5 FILLER_21_1796 ();
 b15zdnd11an1n64x5 FILLER_21_1860 ();
 b15zdnd11an1n64x5 FILLER_21_1924 ();
 b15zdnd11an1n64x5 FILLER_21_1988 ();
 b15zdnd11an1n64x5 FILLER_21_2052 ();
 b15zdnd11an1n64x5 FILLER_21_2116 ();
 b15zdnd11an1n64x5 FILLER_21_2180 ();
 b15zdnd11an1n32x5 FILLER_21_2244 ();
 b15zdnd11an1n08x5 FILLER_21_2276 ();
 b15zdnd11an1n08x5 FILLER_22_8 ();
 b15zdnd11an1n04x5 FILLER_22_16 ();
 b15zdnd00an1n02x5 FILLER_22_20 ();
 b15zdnd11an1n64x5 FILLER_22_25 ();
 b15zdnd11an1n64x5 FILLER_22_89 ();
 b15zdnd11an1n64x5 FILLER_22_153 ();
 b15zdnd11an1n64x5 FILLER_22_217 ();
 b15zdnd11an1n64x5 FILLER_22_281 ();
 b15zdnd11an1n64x5 FILLER_22_345 ();
 b15zdnd11an1n64x5 FILLER_22_409 ();
 b15zdnd11an1n64x5 FILLER_22_473 ();
 b15zdnd11an1n64x5 FILLER_22_537 ();
 b15zdnd11an1n64x5 FILLER_22_601 ();
 b15zdnd11an1n32x5 FILLER_22_665 ();
 b15zdnd11an1n16x5 FILLER_22_697 ();
 b15zdnd11an1n04x5 FILLER_22_713 ();
 b15zdnd00an1n01x5 FILLER_22_717 ();
 b15zdnd11an1n64x5 FILLER_22_726 ();
 b15zdnd11an1n64x5 FILLER_22_790 ();
 b15zdnd11an1n04x5 FILLER_22_857 ();
 b15zdnd11an1n64x5 FILLER_22_864 ();
 b15zdnd11an1n64x5 FILLER_22_928 ();
 b15zdnd11an1n64x5 FILLER_22_992 ();
 b15zdnd11an1n64x5 FILLER_22_1056 ();
 b15zdnd11an1n04x5 FILLER_22_1120 ();
 b15zdnd00an1n02x5 FILLER_22_1124 ();
 b15zdnd00an1n01x5 FILLER_22_1126 ();
 b15zdnd11an1n04x5 FILLER_22_1136 ();
 b15zdnd00an1n01x5 FILLER_22_1140 ();
 b15zdnd11an1n64x5 FILLER_22_1183 ();
 b15zdnd11an1n64x5 FILLER_22_1247 ();
 b15zdnd11an1n64x5 FILLER_22_1311 ();
 b15zdnd11an1n64x5 FILLER_22_1375 ();
 b15zdnd11an1n64x5 FILLER_22_1439 ();
 b15zdnd11an1n64x5 FILLER_22_1503 ();
 b15zdnd11an1n64x5 FILLER_22_1567 ();
 b15zdnd11an1n64x5 FILLER_22_1631 ();
 b15zdnd11an1n64x5 FILLER_22_1695 ();
 b15zdnd11an1n64x5 FILLER_22_1759 ();
 b15zdnd11an1n64x5 FILLER_22_1823 ();
 b15zdnd11an1n64x5 FILLER_22_1887 ();
 b15zdnd11an1n64x5 FILLER_22_1951 ();
 b15zdnd11an1n64x5 FILLER_22_2015 ();
 b15zdnd11an1n64x5 FILLER_22_2079 ();
 b15zdnd11an1n08x5 FILLER_22_2143 ();
 b15zdnd00an1n02x5 FILLER_22_2151 ();
 b15zdnd00an1n01x5 FILLER_22_2153 ();
 b15zdnd11an1n64x5 FILLER_22_2162 ();
 b15zdnd11an1n32x5 FILLER_22_2226 ();
 b15zdnd11an1n16x5 FILLER_22_2258 ();
 b15zdnd00an1n02x5 FILLER_22_2274 ();
 b15zdnd11an1n64x5 FILLER_23_0 ();
 b15zdnd11an1n64x5 FILLER_23_64 ();
 b15zdnd11an1n64x5 FILLER_23_128 ();
 b15zdnd11an1n64x5 FILLER_23_192 ();
 b15zdnd11an1n64x5 FILLER_23_256 ();
 b15zdnd11an1n64x5 FILLER_23_320 ();
 b15zdnd11an1n64x5 FILLER_23_384 ();
 b15zdnd11an1n64x5 FILLER_23_448 ();
 b15zdnd11an1n64x5 FILLER_23_512 ();
 b15zdnd11an1n64x5 FILLER_23_576 ();
 b15zdnd11an1n64x5 FILLER_23_640 ();
 b15zdnd11an1n64x5 FILLER_23_704 ();
 b15zdnd11an1n64x5 FILLER_23_768 ();
 b15zdnd11an1n16x5 FILLER_23_832 ();
 b15zdnd11an1n08x5 FILLER_23_848 ();
 b15zdnd00an1n02x5 FILLER_23_856 ();
 b15zdnd00an1n01x5 FILLER_23_858 ();
 b15zdnd11an1n64x5 FILLER_23_862 ();
 b15zdnd11an1n64x5 FILLER_23_926 ();
 b15zdnd11an1n64x5 FILLER_23_990 ();
 b15zdnd11an1n64x5 FILLER_23_1054 ();
 b15zdnd11an1n64x5 FILLER_23_1118 ();
 b15zdnd11an1n64x5 FILLER_23_1182 ();
 b15zdnd11an1n08x5 FILLER_23_1246 ();
 b15zdnd11an1n04x5 FILLER_23_1254 ();
 b15zdnd00an1n02x5 FILLER_23_1258 ();
 b15zdnd11an1n64x5 FILLER_23_1283 ();
 b15zdnd11an1n64x5 FILLER_23_1347 ();
 b15zdnd11an1n64x5 FILLER_23_1411 ();
 b15zdnd11an1n64x5 FILLER_23_1475 ();
 b15zdnd11an1n32x5 FILLER_23_1539 ();
 b15zdnd11an1n08x5 FILLER_23_1613 ();
 b15zdnd11an1n04x5 FILLER_23_1621 ();
 b15zdnd11an1n04x5 FILLER_23_1667 ();
 b15zdnd11an1n64x5 FILLER_23_1691 ();
 b15zdnd11an1n64x5 FILLER_23_1755 ();
 b15zdnd11an1n64x5 FILLER_23_1819 ();
 b15zdnd11an1n64x5 FILLER_23_1883 ();
 b15zdnd11an1n64x5 FILLER_23_1947 ();
 b15zdnd11an1n64x5 FILLER_23_2011 ();
 b15zdnd11an1n64x5 FILLER_23_2075 ();
 b15zdnd11an1n64x5 FILLER_23_2139 ();
 b15zdnd11an1n64x5 FILLER_23_2203 ();
 b15zdnd11an1n16x5 FILLER_23_2267 ();
 b15zdnd00an1n01x5 FILLER_23_2283 ();
 b15zdnd11an1n64x5 FILLER_24_8 ();
 b15zdnd11an1n64x5 FILLER_24_72 ();
 b15zdnd11an1n64x5 FILLER_24_136 ();
 b15zdnd11an1n64x5 FILLER_24_200 ();
 b15zdnd11an1n64x5 FILLER_24_264 ();
 b15zdnd11an1n64x5 FILLER_24_328 ();
 b15zdnd11an1n64x5 FILLER_24_392 ();
 b15zdnd11an1n64x5 FILLER_24_456 ();
 b15zdnd11an1n64x5 FILLER_24_520 ();
 b15zdnd11an1n64x5 FILLER_24_584 ();
 b15zdnd11an1n64x5 FILLER_24_648 ();
 b15zdnd11an1n04x5 FILLER_24_712 ();
 b15zdnd00an1n02x5 FILLER_24_716 ();
 b15zdnd11an1n64x5 FILLER_24_726 ();
 b15zdnd11an1n64x5 FILLER_24_790 ();
 b15zdnd11an1n64x5 FILLER_24_854 ();
 b15zdnd11an1n16x5 FILLER_24_918 ();
 b15zdnd11an1n08x5 FILLER_24_934 ();
 b15zdnd00an1n01x5 FILLER_24_942 ();
 b15zdnd11an1n64x5 FILLER_24_985 ();
 b15zdnd11an1n64x5 FILLER_24_1049 ();
 b15zdnd11an1n64x5 FILLER_24_1113 ();
 b15zdnd11an1n32x5 FILLER_24_1177 ();
 b15zdnd11an1n16x5 FILLER_24_1209 ();
 b15zdnd00an1n01x5 FILLER_24_1225 ();
 b15zdnd11an1n16x5 FILLER_24_1235 ();
 b15zdnd11an1n08x5 FILLER_24_1251 ();
 b15zdnd11an1n04x5 FILLER_24_1259 ();
 b15zdnd00an1n02x5 FILLER_24_1263 ();
 b15zdnd00an1n01x5 FILLER_24_1265 ();
 b15zdnd11an1n64x5 FILLER_24_1282 ();
 b15zdnd11an1n64x5 FILLER_24_1346 ();
 b15zdnd11an1n64x5 FILLER_24_1410 ();
 b15zdnd11an1n64x5 FILLER_24_1474 ();
 b15zdnd11an1n64x5 FILLER_24_1538 ();
 b15zdnd11an1n64x5 FILLER_24_1602 ();
 b15zdnd11an1n64x5 FILLER_24_1666 ();
 b15zdnd11an1n64x5 FILLER_24_1730 ();
 b15zdnd11an1n64x5 FILLER_24_1794 ();
 b15zdnd11an1n64x5 FILLER_24_1858 ();
 b15zdnd11an1n64x5 FILLER_24_1922 ();
 b15zdnd11an1n64x5 FILLER_24_1986 ();
 b15zdnd11an1n64x5 FILLER_24_2050 ();
 b15zdnd11an1n32x5 FILLER_24_2114 ();
 b15zdnd11an1n08x5 FILLER_24_2146 ();
 b15zdnd11an1n64x5 FILLER_24_2162 ();
 b15zdnd11an1n32x5 FILLER_24_2226 ();
 b15zdnd11an1n16x5 FILLER_24_2258 ();
 b15zdnd00an1n02x5 FILLER_24_2274 ();
 b15zdnd11an1n64x5 FILLER_25_0 ();
 b15zdnd11an1n64x5 FILLER_25_64 ();
 b15zdnd11an1n64x5 FILLER_25_128 ();
 b15zdnd11an1n64x5 FILLER_25_192 ();
 b15zdnd11an1n64x5 FILLER_25_256 ();
 b15zdnd11an1n64x5 FILLER_25_320 ();
 b15zdnd11an1n64x5 FILLER_25_384 ();
 b15zdnd11an1n64x5 FILLER_25_448 ();
 b15zdnd11an1n64x5 FILLER_25_512 ();
 b15zdnd11an1n64x5 FILLER_25_576 ();
 b15zdnd11an1n64x5 FILLER_25_640 ();
 b15zdnd11an1n16x5 FILLER_25_704 ();
 b15zdnd00an1n01x5 FILLER_25_720 ();
 b15zdnd11an1n64x5 FILLER_25_741 ();
 b15zdnd11an1n64x5 FILLER_25_805 ();
 b15zdnd11an1n64x5 FILLER_25_869 ();
 b15zdnd11an1n32x5 FILLER_25_933 ();
 b15zdnd11an1n16x5 FILLER_25_965 ();
 b15zdnd00an1n02x5 FILLER_25_981 ();
 b15zdnd11an1n32x5 FILLER_25_1025 ();
 b15zdnd11an1n08x5 FILLER_25_1057 ();
 b15zdnd00an1n01x5 FILLER_25_1065 ();
 b15zdnd11an1n16x5 FILLER_25_1108 ();
 b15zdnd11an1n04x5 FILLER_25_1124 ();
 b15zdnd11an1n64x5 FILLER_25_1170 ();
 b15zdnd11an1n64x5 FILLER_25_1234 ();
 b15zdnd11an1n64x5 FILLER_25_1298 ();
 b15zdnd11an1n64x5 FILLER_25_1362 ();
 b15zdnd11an1n64x5 FILLER_25_1426 ();
 b15zdnd11an1n64x5 FILLER_25_1490 ();
 b15zdnd11an1n64x5 FILLER_25_1554 ();
 b15zdnd11an1n64x5 FILLER_25_1618 ();
 b15zdnd11an1n64x5 FILLER_25_1682 ();
 b15zdnd11an1n64x5 FILLER_25_1746 ();
 b15zdnd11an1n64x5 FILLER_25_1810 ();
 b15zdnd11an1n64x5 FILLER_25_1874 ();
 b15zdnd11an1n64x5 FILLER_25_1938 ();
 b15zdnd11an1n64x5 FILLER_25_2002 ();
 b15zdnd11an1n64x5 FILLER_25_2066 ();
 b15zdnd11an1n64x5 FILLER_25_2130 ();
 b15zdnd11an1n64x5 FILLER_25_2194 ();
 b15zdnd11an1n16x5 FILLER_25_2258 ();
 b15zdnd11an1n08x5 FILLER_25_2274 ();
 b15zdnd00an1n02x5 FILLER_25_2282 ();
 b15zdnd11an1n64x5 FILLER_26_8 ();
 b15zdnd11an1n64x5 FILLER_26_72 ();
 b15zdnd11an1n64x5 FILLER_26_136 ();
 b15zdnd11an1n64x5 FILLER_26_200 ();
 b15zdnd11an1n64x5 FILLER_26_264 ();
 b15zdnd11an1n64x5 FILLER_26_328 ();
 b15zdnd11an1n08x5 FILLER_26_392 ();
 b15zdnd11an1n04x5 FILLER_26_400 ();
 b15zdnd00an1n01x5 FILLER_26_404 ();
 b15zdnd11an1n16x5 FILLER_26_414 ();
 b15zdnd11an1n08x5 FILLER_26_430 ();
 b15zdnd00an1n02x5 FILLER_26_438 ();
 b15zdnd00an1n01x5 FILLER_26_440 ();
 b15zdnd11an1n64x5 FILLER_26_450 ();
 b15zdnd11an1n64x5 FILLER_26_514 ();
 b15zdnd11an1n64x5 FILLER_26_578 ();
 b15zdnd11an1n64x5 FILLER_26_642 ();
 b15zdnd11an1n08x5 FILLER_26_706 ();
 b15zdnd11an1n04x5 FILLER_26_714 ();
 b15zdnd11an1n64x5 FILLER_26_726 ();
 b15zdnd11an1n64x5 FILLER_26_790 ();
 b15zdnd11an1n32x5 FILLER_26_854 ();
 b15zdnd11an1n16x5 FILLER_26_886 ();
 b15zdnd00an1n02x5 FILLER_26_902 ();
 b15zdnd00an1n01x5 FILLER_26_904 ();
 b15zdnd11an1n64x5 FILLER_26_914 ();
 b15zdnd11an1n64x5 FILLER_26_978 ();
 b15zdnd11an1n32x5 FILLER_26_1042 ();
 b15zdnd11an1n16x5 FILLER_26_1074 ();
 b15zdnd11an1n08x5 FILLER_26_1090 ();
 b15zdnd00an1n01x5 FILLER_26_1098 ();
 b15zdnd11an1n04x5 FILLER_26_1108 ();
 b15zdnd11an1n04x5 FILLER_26_1115 ();
 b15zdnd11an1n64x5 FILLER_26_1122 ();
 b15zdnd11an1n64x5 FILLER_26_1186 ();
 b15zdnd11an1n64x5 FILLER_26_1266 ();
 b15zdnd11an1n08x5 FILLER_26_1330 ();
 b15zdnd00an1n02x5 FILLER_26_1338 ();
 b15zdnd00an1n01x5 FILLER_26_1340 ();
 b15zdnd11an1n04x5 FILLER_26_1383 ();
 b15zdnd00an1n02x5 FILLER_26_1387 ();
 b15zdnd00an1n01x5 FILLER_26_1389 ();
 b15zdnd11an1n64x5 FILLER_26_1432 ();
 b15zdnd11an1n64x5 FILLER_26_1496 ();
 b15zdnd11an1n64x5 FILLER_26_1560 ();
 b15zdnd11an1n32x5 FILLER_26_1624 ();
 b15zdnd11an1n04x5 FILLER_26_1656 ();
 b15zdnd11an1n64x5 FILLER_26_1691 ();
 b15zdnd11an1n64x5 FILLER_26_1755 ();
 b15zdnd11an1n64x5 FILLER_26_1819 ();
 b15zdnd11an1n64x5 FILLER_26_1883 ();
 b15zdnd11an1n64x5 FILLER_26_1947 ();
 b15zdnd11an1n64x5 FILLER_26_2011 ();
 b15zdnd11an1n64x5 FILLER_26_2075 ();
 b15zdnd11an1n08x5 FILLER_26_2139 ();
 b15zdnd11an1n04x5 FILLER_26_2147 ();
 b15zdnd00an1n02x5 FILLER_26_2151 ();
 b15zdnd00an1n01x5 FILLER_26_2153 ();
 b15zdnd00an1n02x5 FILLER_26_2162 ();
 b15zdnd11an1n04x5 FILLER_26_2206 ();
 b15zdnd11an1n16x5 FILLER_26_2252 ();
 b15zdnd11an1n08x5 FILLER_26_2268 ();
 b15zdnd11an1n64x5 FILLER_27_0 ();
 b15zdnd11an1n64x5 FILLER_27_64 ();
 b15zdnd11an1n64x5 FILLER_27_128 ();
 b15zdnd11an1n64x5 FILLER_27_192 ();
 b15zdnd11an1n64x5 FILLER_27_256 ();
 b15zdnd11an1n64x5 FILLER_27_320 ();
 b15zdnd11an1n64x5 FILLER_27_384 ();
 b15zdnd11an1n64x5 FILLER_27_448 ();
 b15zdnd11an1n64x5 FILLER_27_512 ();
 b15zdnd11an1n64x5 FILLER_27_576 ();
 b15zdnd11an1n64x5 FILLER_27_640 ();
 b15zdnd11an1n64x5 FILLER_27_704 ();
 b15zdnd11an1n64x5 FILLER_27_768 ();
 b15zdnd11an1n64x5 FILLER_27_832 ();
 b15zdnd11an1n64x5 FILLER_27_896 ();
 b15zdnd11an1n64x5 FILLER_27_960 ();
 b15zdnd11an1n64x5 FILLER_27_1024 ();
 b15zdnd11an1n16x5 FILLER_27_1088 ();
 b15zdnd11an1n04x5 FILLER_27_1104 ();
 b15zdnd11an1n64x5 FILLER_27_1150 ();
 b15zdnd11an1n16x5 FILLER_27_1214 ();
 b15zdnd11an1n08x5 FILLER_27_1230 ();
 b15zdnd00an1n01x5 FILLER_27_1238 ();
 b15zdnd11an1n04x5 FILLER_27_1243 ();
 b15zdnd11an1n04x5 FILLER_27_1263 ();
 b15zdnd11an1n64x5 FILLER_27_1270 ();
 b15zdnd11an1n64x5 FILLER_27_1334 ();
 b15zdnd11an1n64x5 FILLER_27_1398 ();
 b15zdnd11an1n64x5 FILLER_27_1462 ();
 b15zdnd11an1n64x5 FILLER_27_1526 ();
 b15zdnd11an1n64x5 FILLER_27_1590 ();
 b15zdnd11an1n64x5 FILLER_27_1654 ();
 b15zdnd11an1n64x5 FILLER_27_1718 ();
 b15zdnd11an1n64x5 FILLER_27_1782 ();
 b15zdnd11an1n64x5 FILLER_27_1846 ();
 b15zdnd11an1n64x5 FILLER_27_1910 ();
 b15zdnd11an1n64x5 FILLER_27_1974 ();
 b15zdnd11an1n64x5 FILLER_27_2038 ();
 b15zdnd11an1n64x5 FILLER_27_2102 ();
 b15zdnd11an1n64x5 FILLER_27_2166 ();
 b15zdnd11an1n32x5 FILLER_27_2230 ();
 b15zdnd11an1n16x5 FILLER_27_2262 ();
 b15zdnd11an1n04x5 FILLER_27_2278 ();
 b15zdnd00an1n02x5 FILLER_27_2282 ();
 b15zdnd11an1n64x5 FILLER_28_8 ();
 b15zdnd11an1n64x5 FILLER_28_72 ();
 b15zdnd11an1n64x5 FILLER_28_136 ();
 b15zdnd11an1n64x5 FILLER_28_200 ();
 b15zdnd11an1n64x5 FILLER_28_264 ();
 b15zdnd11an1n64x5 FILLER_28_328 ();
 b15zdnd11an1n64x5 FILLER_28_392 ();
 b15zdnd11an1n64x5 FILLER_28_456 ();
 b15zdnd11an1n64x5 FILLER_28_520 ();
 b15zdnd11an1n64x5 FILLER_28_584 ();
 b15zdnd11an1n64x5 FILLER_28_648 ();
 b15zdnd11an1n04x5 FILLER_28_712 ();
 b15zdnd00an1n02x5 FILLER_28_716 ();
 b15zdnd11an1n64x5 FILLER_28_726 ();
 b15zdnd11an1n64x5 FILLER_28_790 ();
 b15zdnd11an1n64x5 FILLER_28_854 ();
 b15zdnd11an1n64x5 FILLER_28_918 ();
 b15zdnd11an1n64x5 FILLER_28_982 ();
 b15zdnd11an1n32x5 FILLER_28_1046 ();
 b15zdnd11an1n08x5 FILLER_28_1078 ();
 b15zdnd11an1n04x5 FILLER_28_1086 ();
 b15zdnd00an1n02x5 FILLER_28_1090 ();
 b15zdnd11an1n64x5 FILLER_28_1144 ();
 b15zdnd11an1n32x5 FILLER_28_1208 ();
 b15zdnd11an1n08x5 FILLER_28_1240 ();
 b15zdnd00an1n02x5 FILLER_28_1248 ();
 b15zdnd00an1n01x5 FILLER_28_1250 ();
 b15zdnd11an1n16x5 FILLER_28_1293 ();
 b15zdnd11an1n08x5 FILLER_28_1309 ();
 b15zdnd11an1n04x5 FILLER_28_1317 ();
 b15zdnd11an1n64x5 FILLER_28_1363 ();
 b15zdnd11an1n64x5 FILLER_28_1427 ();
 b15zdnd11an1n64x5 FILLER_28_1491 ();
 b15zdnd11an1n64x5 FILLER_28_1555 ();
 b15zdnd11an1n64x5 FILLER_28_1619 ();
 b15zdnd11an1n64x5 FILLER_28_1683 ();
 b15zdnd11an1n64x5 FILLER_28_1747 ();
 b15zdnd11an1n64x5 FILLER_28_1811 ();
 b15zdnd11an1n64x5 FILLER_28_1875 ();
 b15zdnd11an1n64x5 FILLER_28_1939 ();
 b15zdnd11an1n64x5 FILLER_28_2003 ();
 b15zdnd11an1n64x5 FILLER_28_2067 ();
 b15zdnd11an1n16x5 FILLER_28_2131 ();
 b15zdnd11an1n04x5 FILLER_28_2147 ();
 b15zdnd00an1n02x5 FILLER_28_2151 ();
 b15zdnd00an1n01x5 FILLER_28_2153 ();
 b15zdnd11an1n64x5 FILLER_28_2162 ();
 b15zdnd11an1n32x5 FILLER_28_2226 ();
 b15zdnd11an1n16x5 FILLER_28_2258 ();
 b15zdnd00an1n02x5 FILLER_28_2274 ();
 b15zdnd11an1n64x5 FILLER_29_0 ();
 b15zdnd11an1n64x5 FILLER_29_64 ();
 b15zdnd11an1n64x5 FILLER_29_128 ();
 b15zdnd11an1n64x5 FILLER_29_192 ();
 b15zdnd11an1n64x5 FILLER_29_256 ();
 b15zdnd11an1n64x5 FILLER_29_320 ();
 b15zdnd11an1n64x5 FILLER_29_384 ();
 b15zdnd11an1n64x5 FILLER_29_448 ();
 b15zdnd11an1n64x5 FILLER_29_512 ();
 b15zdnd11an1n64x5 FILLER_29_576 ();
 b15zdnd11an1n64x5 FILLER_29_640 ();
 b15zdnd11an1n64x5 FILLER_29_704 ();
 b15zdnd11an1n64x5 FILLER_29_768 ();
 b15zdnd11an1n64x5 FILLER_29_832 ();
 b15zdnd11an1n64x5 FILLER_29_896 ();
 b15zdnd11an1n16x5 FILLER_29_960 ();
 b15zdnd11an1n08x5 FILLER_29_976 ();
 b15zdnd00an1n01x5 FILLER_29_984 ();
 b15zdnd11an1n04x5 FILLER_29_1027 ();
 b15zdnd11an1n32x5 FILLER_29_1073 ();
 b15zdnd00an1n02x5 FILLER_29_1105 ();
 b15zdnd00an1n01x5 FILLER_29_1107 ();
 b15zdnd11an1n04x5 FILLER_29_1111 ();
 b15zdnd11an1n04x5 FILLER_29_1118 ();
 b15zdnd11an1n04x5 FILLER_29_1125 ();
 b15zdnd11an1n08x5 FILLER_29_1171 ();
 b15zdnd11an1n04x5 FILLER_29_1179 ();
 b15zdnd00an1n01x5 FILLER_29_1183 ();
 b15zdnd11an1n04x5 FILLER_29_1226 ();
 b15zdnd00an1n02x5 FILLER_29_1230 ();
 b15zdnd00an1n01x5 FILLER_29_1232 ();
 b15zdnd11an1n64x5 FILLER_29_1275 ();
 b15zdnd11an1n64x5 FILLER_29_1339 ();
 b15zdnd11an1n64x5 FILLER_29_1403 ();
 b15zdnd11an1n64x5 FILLER_29_1467 ();
 b15zdnd11an1n64x5 FILLER_29_1531 ();
 b15zdnd11an1n64x5 FILLER_29_1595 ();
 b15zdnd11an1n64x5 FILLER_29_1659 ();
 b15zdnd11an1n64x5 FILLER_29_1723 ();
 b15zdnd11an1n64x5 FILLER_29_1787 ();
 b15zdnd11an1n64x5 FILLER_29_1851 ();
 b15zdnd11an1n64x5 FILLER_29_1915 ();
 b15zdnd11an1n64x5 FILLER_29_1979 ();
 b15zdnd11an1n64x5 FILLER_29_2043 ();
 b15zdnd11an1n64x5 FILLER_29_2107 ();
 b15zdnd11an1n64x5 FILLER_29_2171 ();
 b15zdnd11an1n32x5 FILLER_29_2235 ();
 b15zdnd11an1n16x5 FILLER_29_2267 ();
 b15zdnd00an1n01x5 FILLER_29_2283 ();
 b15zdnd11an1n64x5 FILLER_30_8 ();
 b15zdnd11an1n64x5 FILLER_30_72 ();
 b15zdnd11an1n64x5 FILLER_30_136 ();
 b15zdnd11an1n64x5 FILLER_30_200 ();
 b15zdnd11an1n64x5 FILLER_30_264 ();
 b15zdnd11an1n64x5 FILLER_30_328 ();
 b15zdnd11an1n64x5 FILLER_30_392 ();
 b15zdnd11an1n32x5 FILLER_30_456 ();
 b15zdnd11an1n16x5 FILLER_30_488 ();
 b15zdnd11an1n08x5 FILLER_30_504 ();
 b15zdnd00an1n02x5 FILLER_30_512 ();
 b15zdnd00an1n01x5 FILLER_30_514 ();
 b15zdnd11an1n64x5 FILLER_30_532 ();
 b15zdnd11an1n64x5 FILLER_30_596 ();
 b15zdnd11an1n32x5 FILLER_30_660 ();
 b15zdnd11an1n16x5 FILLER_30_692 ();
 b15zdnd11an1n08x5 FILLER_30_708 ();
 b15zdnd00an1n02x5 FILLER_30_716 ();
 b15zdnd11an1n64x5 FILLER_30_726 ();
 b15zdnd11an1n64x5 FILLER_30_790 ();
 b15zdnd11an1n32x5 FILLER_30_854 ();
 b15zdnd11an1n16x5 FILLER_30_886 ();
 b15zdnd00an1n02x5 FILLER_30_902 ();
 b15zdnd00an1n01x5 FILLER_30_904 ();
 b15zdnd11an1n04x5 FILLER_30_914 ();
 b15zdnd00an1n02x5 FILLER_30_918 ();
 b15zdnd11an1n64x5 FILLER_30_929 ();
 b15zdnd11an1n64x5 FILLER_30_993 ();
 b15zdnd11an1n32x5 FILLER_30_1057 ();
 b15zdnd11an1n04x5 FILLER_30_1089 ();
 b15zdnd00an1n02x5 FILLER_30_1093 ();
 b15zdnd11an1n64x5 FILLER_30_1147 ();
 b15zdnd11an1n32x5 FILLER_30_1211 ();
 b15zdnd00an1n02x5 FILLER_30_1243 ();
 b15zdnd11an1n08x5 FILLER_30_1255 ();
 b15zdnd00an1n01x5 FILLER_30_1263 ();
 b15zdnd11an1n64x5 FILLER_30_1280 ();
 b15zdnd11an1n64x5 FILLER_30_1344 ();
 b15zdnd11an1n64x5 FILLER_30_1408 ();
 b15zdnd11an1n64x5 FILLER_30_1472 ();
 b15zdnd11an1n64x5 FILLER_30_1536 ();
 b15zdnd11an1n64x5 FILLER_30_1600 ();
 b15zdnd11an1n64x5 FILLER_30_1664 ();
 b15zdnd11an1n32x5 FILLER_30_1728 ();
 b15zdnd11an1n08x5 FILLER_30_1760 ();
 b15zdnd11an1n04x5 FILLER_30_1768 ();
 b15zdnd11an1n64x5 FILLER_30_1775 ();
 b15zdnd11an1n64x5 FILLER_30_1839 ();
 b15zdnd11an1n08x5 FILLER_30_1903 ();
 b15zdnd11an1n64x5 FILLER_30_1914 ();
 b15zdnd11an1n64x5 FILLER_30_1978 ();
 b15zdnd11an1n64x5 FILLER_30_2042 ();
 b15zdnd11an1n32x5 FILLER_30_2106 ();
 b15zdnd11an1n16x5 FILLER_30_2138 ();
 b15zdnd11an1n64x5 FILLER_30_2162 ();
 b15zdnd11an1n32x5 FILLER_30_2226 ();
 b15zdnd11an1n16x5 FILLER_30_2258 ();
 b15zdnd00an1n02x5 FILLER_30_2274 ();
 b15zdnd11an1n64x5 FILLER_31_0 ();
 b15zdnd11an1n64x5 FILLER_31_64 ();
 b15zdnd11an1n64x5 FILLER_31_128 ();
 b15zdnd11an1n64x5 FILLER_31_192 ();
 b15zdnd11an1n64x5 FILLER_31_256 ();
 b15zdnd11an1n64x5 FILLER_31_320 ();
 b15zdnd11an1n64x5 FILLER_31_384 ();
 b15zdnd11an1n64x5 FILLER_31_448 ();
 b15zdnd11an1n64x5 FILLER_31_512 ();
 b15zdnd11an1n04x5 FILLER_31_576 ();
 b15zdnd11an1n04x5 FILLER_31_583 ();
 b15zdnd00an1n01x5 FILLER_31_587 ();
 b15zdnd11an1n64x5 FILLER_31_591 ();
 b15zdnd11an1n64x5 FILLER_31_655 ();
 b15zdnd11an1n64x5 FILLER_31_719 ();
 b15zdnd11an1n64x5 FILLER_31_783 ();
 b15zdnd11an1n64x5 FILLER_31_847 ();
 b15zdnd11an1n64x5 FILLER_31_911 ();
 b15zdnd11an1n64x5 FILLER_31_975 ();
 b15zdnd11an1n64x5 FILLER_31_1039 ();
 b15zdnd11an1n16x5 FILLER_31_1103 ();
 b15zdnd11an1n04x5 FILLER_31_1119 ();
 b15zdnd00an1n02x5 FILLER_31_1123 ();
 b15zdnd00an1n01x5 FILLER_31_1125 ();
 b15zdnd11an1n08x5 FILLER_31_1129 ();
 b15zdnd11an1n04x5 FILLER_31_1137 ();
 b15zdnd00an1n02x5 FILLER_31_1141 ();
 b15zdnd00an1n01x5 FILLER_31_1143 ();
 b15zdnd11an1n16x5 FILLER_31_1151 ();
 b15zdnd11an1n04x5 FILLER_31_1167 ();
 b15zdnd00an1n02x5 FILLER_31_1171 ();
 b15zdnd11an1n64x5 FILLER_31_1180 ();
 b15zdnd11an1n08x5 FILLER_31_1244 ();
 b15zdnd00an1n01x5 FILLER_31_1252 ();
 b15zdnd11an1n04x5 FILLER_31_1263 ();
 b15zdnd11an1n64x5 FILLER_31_1274 ();
 b15zdnd11an1n64x5 FILLER_31_1338 ();
 b15zdnd11an1n64x5 FILLER_31_1402 ();
 b15zdnd11an1n08x5 FILLER_31_1466 ();
 b15zdnd11an1n04x5 FILLER_31_1474 ();
 b15zdnd11an1n32x5 FILLER_31_1481 ();
 b15zdnd11an1n16x5 FILLER_31_1513 ();
 b15zdnd11an1n04x5 FILLER_31_1529 ();
 b15zdnd00an1n02x5 FILLER_31_1533 ();
 b15zdnd00an1n01x5 FILLER_31_1535 ();
 b15zdnd11an1n16x5 FILLER_31_1578 ();
 b15zdnd00an1n01x5 FILLER_31_1594 ();
 b15zdnd11an1n32x5 FILLER_31_1598 ();
 b15zdnd11an1n16x5 FILLER_31_1630 ();
 b15zdnd11an1n08x5 FILLER_31_1646 ();
 b15zdnd11an1n04x5 FILLER_31_1654 ();
 b15zdnd00an1n01x5 FILLER_31_1658 ();
 b15zdnd11an1n64x5 FILLER_31_1683 ();
 b15zdnd11an1n16x5 FILLER_31_1747 ();
 b15zdnd11an1n08x5 FILLER_31_1763 ();
 b15zdnd00an1n01x5 FILLER_31_1771 ();
 b15zdnd11an1n64x5 FILLER_31_1775 ();
 b15zdnd11an1n64x5 FILLER_31_1839 ();
 b15zdnd11an1n04x5 FILLER_31_1903 ();
 b15zdnd00an1n02x5 FILLER_31_1907 ();
 b15zdnd11an1n04x5 FILLER_31_1912 ();
 b15zdnd11an1n64x5 FILLER_31_1919 ();
 b15zdnd11an1n32x5 FILLER_31_1983 ();
 b15zdnd11an1n08x5 FILLER_31_2015 ();
 b15zdnd00an1n02x5 FILLER_31_2023 ();
 b15zdnd00an1n01x5 FILLER_31_2025 ();
 b15zdnd11an1n64x5 FILLER_31_2078 ();
 b15zdnd11an1n64x5 FILLER_31_2142 ();
 b15zdnd11an1n64x5 FILLER_31_2206 ();
 b15zdnd11an1n08x5 FILLER_31_2270 ();
 b15zdnd11an1n04x5 FILLER_31_2278 ();
 b15zdnd00an1n02x5 FILLER_31_2282 ();
 b15zdnd11an1n64x5 FILLER_32_8 ();
 b15zdnd11an1n64x5 FILLER_32_72 ();
 b15zdnd11an1n64x5 FILLER_32_136 ();
 b15zdnd11an1n64x5 FILLER_32_200 ();
 b15zdnd11an1n64x5 FILLER_32_264 ();
 b15zdnd11an1n64x5 FILLER_32_328 ();
 b15zdnd11an1n64x5 FILLER_32_392 ();
 b15zdnd11an1n64x5 FILLER_32_456 ();
 b15zdnd11an1n32x5 FILLER_32_520 ();
 b15zdnd11an1n08x5 FILLER_32_552 ();
 b15zdnd00an1n01x5 FILLER_32_560 ();
 b15zdnd11an1n64x5 FILLER_32_603 ();
 b15zdnd11an1n32x5 FILLER_32_667 ();
 b15zdnd11an1n16x5 FILLER_32_699 ();
 b15zdnd00an1n02x5 FILLER_32_715 ();
 b15zdnd00an1n01x5 FILLER_32_717 ();
 b15zdnd11an1n64x5 FILLER_32_726 ();
 b15zdnd11an1n64x5 FILLER_32_790 ();
 b15zdnd11an1n64x5 FILLER_32_854 ();
 b15zdnd11an1n64x5 FILLER_32_918 ();
 b15zdnd00an1n02x5 FILLER_32_982 ();
 b15zdnd11an1n04x5 FILLER_32_987 ();
 b15zdnd11an1n64x5 FILLER_32_994 ();
 b15zdnd11an1n64x5 FILLER_32_1058 ();
 b15zdnd11an1n64x5 FILLER_32_1122 ();
 b15zdnd11an1n64x5 FILLER_32_1186 ();
 b15zdnd11an1n04x5 FILLER_32_1250 ();
 b15zdnd11an1n64x5 FILLER_32_1273 ();
 b15zdnd11an1n64x5 FILLER_32_1337 ();
 b15zdnd11an1n32x5 FILLER_32_1401 ();
 b15zdnd11an1n08x5 FILLER_32_1433 ();
 b15zdnd11an1n04x5 FILLER_32_1441 ();
 b15zdnd00an1n02x5 FILLER_32_1445 ();
 b15zdnd00an1n01x5 FILLER_32_1447 ();
 b15zdnd11an1n08x5 FILLER_32_1490 ();
 b15zdnd11an1n04x5 FILLER_32_1498 ();
 b15zdnd00an1n02x5 FILLER_32_1502 ();
 b15zdnd00an1n01x5 FILLER_32_1504 ();
 b15zdnd11an1n32x5 FILLER_32_1547 ();
 b15zdnd11an1n08x5 FILLER_32_1579 ();
 b15zdnd00an1n01x5 FILLER_32_1587 ();
 b15zdnd11an1n32x5 FILLER_32_1630 ();
 b15zdnd11an1n04x5 FILLER_32_1662 ();
 b15zdnd00an1n02x5 FILLER_32_1666 ();
 b15zdnd00an1n01x5 FILLER_32_1668 ();
 b15zdnd11an1n04x5 FILLER_32_1672 ();
 b15zdnd11an1n08x5 FILLER_32_1679 ();
 b15zdnd11an1n04x5 FILLER_32_1687 ();
 b15zdnd00an1n01x5 FILLER_32_1691 ();
 b15zdnd11an1n16x5 FILLER_32_1719 ();
 b15zdnd11an1n08x5 FILLER_32_1735 ();
 b15zdnd11an1n04x5 FILLER_32_1743 ();
 b15zdnd11an1n04x5 FILLER_32_1799 ();
 b15zdnd11an1n64x5 FILLER_32_1823 ();
 b15zdnd11an1n04x5 FILLER_32_1887 ();
 b15zdnd11an1n64x5 FILLER_32_1943 ();
 b15zdnd11an1n32x5 FILLER_32_2007 ();
 b15zdnd11an1n04x5 FILLER_32_2039 ();
 b15zdnd00an1n01x5 FILLER_32_2043 ();
 b15zdnd11an1n04x5 FILLER_32_2047 ();
 b15zdnd11an1n64x5 FILLER_32_2054 ();
 b15zdnd11an1n32x5 FILLER_32_2118 ();
 b15zdnd11an1n04x5 FILLER_32_2150 ();
 b15zdnd11an1n64x5 FILLER_32_2162 ();
 b15zdnd11an1n32x5 FILLER_32_2226 ();
 b15zdnd11an1n16x5 FILLER_32_2258 ();
 b15zdnd00an1n02x5 FILLER_32_2274 ();
 b15zdnd11an1n64x5 FILLER_33_0 ();
 b15zdnd11an1n64x5 FILLER_33_64 ();
 b15zdnd11an1n64x5 FILLER_33_128 ();
 b15zdnd11an1n64x5 FILLER_33_192 ();
 b15zdnd11an1n64x5 FILLER_33_256 ();
 b15zdnd11an1n32x5 FILLER_33_320 ();
 b15zdnd11an1n16x5 FILLER_33_352 ();
 b15zdnd11an1n04x5 FILLER_33_368 ();
 b15zdnd00an1n02x5 FILLER_33_372 ();
 b15zdnd11an1n64x5 FILLER_33_377 ();
 b15zdnd11an1n64x5 FILLER_33_441 ();
 b15zdnd11an1n32x5 FILLER_33_505 ();
 b15zdnd11an1n16x5 FILLER_33_537 ();
 b15zdnd11an1n04x5 FILLER_33_553 ();
 b15zdnd11an1n64x5 FILLER_33_609 ();
 b15zdnd11an1n16x5 FILLER_33_673 ();
 b15zdnd00an1n02x5 FILLER_33_689 ();
 b15zdnd00an1n01x5 FILLER_33_691 ();
 b15zdnd11an1n04x5 FILLER_33_695 ();
 b15zdnd00an1n02x5 FILLER_33_699 ();
 b15zdnd00an1n01x5 FILLER_33_701 ();
 b15zdnd11an1n64x5 FILLER_33_729 ();
 b15zdnd11an1n64x5 FILLER_33_793 ();
 b15zdnd11an1n64x5 FILLER_33_857 ();
 b15zdnd11an1n32x5 FILLER_33_921 ();
 b15zdnd11an1n08x5 FILLER_33_953 ();
 b15zdnd00an1n02x5 FILLER_33_961 ();
 b15zdnd00an1n01x5 FILLER_33_963 ();
 b15zdnd11an1n64x5 FILLER_33_1016 ();
 b15zdnd11an1n64x5 FILLER_33_1080 ();
 b15zdnd11an1n64x5 FILLER_33_1144 ();
 b15zdnd11an1n64x5 FILLER_33_1208 ();
 b15zdnd11an1n64x5 FILLER_33_1272 ();
 b15zdnd00an1n02x5 FILLER_33_1336 ();
 b15zdnd00an1n01x5 FILLER_33_1338 ();
 b15zdnd11an1n64x5 FILLER_33_1391 ();
 b15zdnd00an1n02x5 FILLER_33_1455 ();
 b15zdnd00an1n01x5 FILLER_33_1457 ();
 b15zdnd11an1n64x5 FILLER_33_1485 ();
 b15zdnd11an1n16x5 FILLER_33_1549 ();
 b15zdnd11an1n04x5 FILLER_33_1565 ();
 b15zdnd11an1n16x5 FILLER_33_1621 ();
 b15zdnd11an1n08x5 FILLER_33_1637 ();
 b15zdnd11an1n04x5 FILLER_33_1645 ();
 b15zdnd00an1n02x5 FILLER_33_1649 ();
 b15zdnd11an1n64x5 FILLER_33_1703 ();
 b15zdnd11an1n04x5 FILLER_33_1767 ();
 b15zdnd00an1n01x5 FILLER_33_1771 ();
 b15zdnd11an1n04x5 FILLER_33_1775 ();
 b15zdnd11an1n04x5 FILLER_33_1803 ();
 b15zdnd11an1n64x5 FILLER_33_1810 ();
 b15zdnd11an1n16x5 FILLER_33_1874 ();
 b15zdnd11an1n08x5 FILLER_33_1890 ();
 b15zdnd11an1n04x5 FILLER_33_1898 ();
 b15zdnd11an1n64x5 FILLER_33_1954 ();
 b15zdnd11an1n16x5 FILLER_33_2018 ();
 b15zdnd11an1n08x5 FILLER_33_2034 ();
 b15zdnd11an1n04x5 FILLER_33_2042 ();
 b15zdnd00an1n02x5 FILLER_33_2046 ();
 b15zdnd00an1n01x5 FILLER_33_2048 ();
 b15zdnd11an1n64x5 FILLER_33_2052 ();
 b15zdnd11an1n64x5 FILLER_33_2116 ();
 b15zdnd11an1n64x5 FILLER_33_2180 ();
 b15zdnd11an1n32x5 FILLER_33_2244 ();
 b15zdnd11an1n08x5 FILLER_33_2276 ();
 b15zdnd11an1n64x5 FILLER_34_8 ();
 b15zdnd11an1n64x5 FILLER_34_72 ();
 b15zdnd11an1n64x5 FILLER_34_136 ();
 b15zdnd11an1n64x5 FILLER_34_200 ();
 b15zdnd11an1n64x5 FILLER_34_264 ();
 b15zdnd11an1n32x5 FILLER_34_328 ();
 b15zdnd11an1n08x5 FILLER_34_360 ();
 b15zdnd11an1n04x5 FILLER_34_371 ();
 b15zdnd11an1n04x5 FILLER_34_378 ();
 b15zdnd11an1n64x5 FILLER_34_385 ();
 b15zdnd11an1n64x5 FILLER_34_449 ();
 b15zdnd11an1n64x5 FILLER_34_513 ();
 b15zdnd11an1n08x5 FILLER_34_577 ();
 b15zdnd00an1n01x5 FILLER_34_585 ();
 b15zdnd11an1n64x5 FILLER_34_589 ();
 b15zdnd11an1n64x5 FILLER_34_653 ();
 b15zdnd00an1n01x5 FILLER_34_717 ();
 b15zdnd11an1n08x5 FILLER_34_726 ();
 b15zdnd11an1n04x5 FILLER_34_734 ();
 b15zdnd11an1n04x5 FILLER_34_741 ();
 b15zdnd00an1n01x5 FILLER_34_745 ();
 b15zdnd11an1n64x5 FILLER_34_766 ();
 b15zdnd11an1n64x5 FILLER_34_830 ();
 b15zdnd11an1n32x5 FILLER_34_894 ();
 b15zdnd11an1n16x5 FILLER_34_926 ();
 b15zdnd11an1n08x5 FILLER_34_942 ();
 b15zdnd00an1n02x5 FILLER_34_950 ();
 b15zdnd00an1n01x5 FILLER_34_952 ();
 b15zdnd11an1n04x5 FILLER_34_956 ();
 b15zdnd11an1n04x5 FILLER_34_963 ();
 b15zdnd11an1n64x5 FILLER_34_970 ();
 b15zdnd11an1n64x5 FILLER_34_1034 ();
 b15zdnd11an1n64x5 FILLER_34_1098 ();
 b15zdnd11an1n64x5 FILLER_34_1162 ();
 b15zdnd11an1n64x5 FILLER_34_1226 ();
 b15zdnd11an1n64x5 FILLER_34_1290 ();
 b15zdnd11an1n04x5 FILLER_34_1354 ();
 b15zdnd11an1n04x5 FILLER_34_1361 ();
 b15zdnd11an1n64x5 FILLER_34_1368 ();
 b15zdnd11an1n16x5 FILLER_34_1432 ();
 b15zdnd00an1n02x5 FILLER_34_1448 ();
 b15zdnd00an1n01x5 FILLER_34_1450 ();
 b15zdnd11an1n64x5 FILLER_34_1503 ();
 b15zdnd11an1n16x5 FILLER_34_1567 ();
 b15zdnd11an1n04x5 FILLER_34_1583 ();
 b15zdnd11an1n04x5 FILLER_34_1590 ();
 b15zdnd11an1n64x5 FILLER_34_1597 ();
 b15zdnd11an1n08x5 FILLER_34_1661 ();
 b15zdnd11an1n04x5 FILLER_34_1669 ();
 b15zdnd00an1n02x5 FILLER_34_1673 ();
 b15zdnd00an1n01x5 FILLER_34_1675 ();
 b15zdnd11an1n08x5 FILLER_34_1679 ();
 b15zdnd11an1n04x5 FILLER_34_1687 ();
 b15zdnd00an1n02x5 FILLER_34_1691 ();
 b15zdnd00an1n01x5 FILLER_34_1693 ();
 b15zdnd11an1n64x5 FILLER_34_1697 ();
 b15zdnd00an1n02x5 FILLER_34_1761 ();
 b15zdnd11an1n64x5 FILLER_34_1815 ();
 b15zdnd11an1n16x5 FILLER_34_1879 ();
 b15zdnd11an1n04x5 FILLER_34_1895 ();
 b15zdnd00an1n01x5 FILLER_34_1899 ();
 b15zdnd11an1n64x5 FILLER_34_1952 ();
 b15zdnd11an1n64x5 FILLER_34_2016 ();
 b15zdnd11an1n64x5 FILLER_34_2080 ();
 b15zdnd11an1n08x5 FILLER_34_2144 ();
 b15zdnd00an1n02x5 FILLER_34_2152 ();
 b15zdnd11an1n64x5 FILLER_34_2162 ();
 b15zdnd11an1n32x5 FILLER_34_2226 ();
 b15zdnd11an1n16x5 FILLER_34_2258 ();
 b15zdnd00an1n02x5 FILLER_34_2274 ();
 b15zdnd11an1n64x5 FILLER_35_0 ();
 b15zdnd11an1n64x5 FILLER_35_64 ();
 b15zdnd11an1n64x5 FILLER_35_128 ();
 b15zdnd11an1n64x5 FILLER_35_192 ();
 b15zdnd11an1n64x5 FILLER_35_256 ();
 b15zdnd11an1n16x5 FILLER_35_320 ();
 b15zdnd11an1n08x5 FILLER_35_336 ();
 b15zdnd11an1n04x5 FILLER_35_344 ();
 b15zdnd00an1n01x5 FILLER_35_348 ();
 b15zdnd11an1n64x5 FILLER_35_401 ();
 b15zdnd11an1n04x5 FILLER_35_465 ();
 b15zdnd00an1n01x5 FILLER_35_469 ();
 b15zdnd11an1n64x5 FILLER_35_473 ();
 b15zdnd11an1n32x5 FILLER_35_537 ();
 b15zdnd00an1n01x5 FILLER_35_569 ();
 b15zdnd11an1n64x5 FILLER_35_590 ();
 b15zdnd11an1n32x5 FILLER_35_654 ();
 b15zdnd11an1n16x5 FILLER_35_686 ();
 b15zdnd11an1n08x5 FILLER_35_702 ();
 b15zdnd00an1n01x5 FILLER_35_710 ();
 b15zdnd11an1n64x5 FILLER_35_763 ();
 b15zdnd11an1n64x5 FILLER_35_827 ();
 b15zdnd11an1n32x5 FILLER_35_891 ();
 b15zdnd11an1n04x5 FILLER_35_923 ();
 b15zdnd00an1n02x5 FILLER_35_927 ();
 b15zdnd00an1n01x5 FILLER_35_929 ();
 b15zdnd11an1n04x5 FILLER_35_982 ();
 b15zdnd11an1n64x5 FILLER_35_989 ();
 b15zdnd11an1n64x5 FILLER_35_1053 ();
 b15zdnd11an1n64x5 FILLER_35_1117 ();
 b15zdnd11an1n64x5 FILLER_35_1181 ();
 b15zdnd11an1n64x5 FILLER_35_1245 ();
 b15zdnd11an1n32x5 FILLER_35_1309 ();
 b15zdnd11an1n16x5 FILLER_35_1341 ();
 b15zdnd11an1n04x5 FILLER_35_1357 ();
 b15zdnd00an1n02x5 FILLER_35_1361 ();
 b15zdnd00an1n01x5 FILLER_35_1363 ();
 b15zdnd11an1n64x5 FILLER_35_1367 ();
 b15zdnd11an1n16x5 FILLER_35_1431 ();
 b15zdnd11an1n08x5 FILLER_35_1447 ();
 b15zdnd11an1n04x5 FILLER_35_1455 ();
 b15zdnd00an1n01x5 FILLER_35_1459 ();
 b15zdnd11an1n04x5 FILLER_35_1463 ();
 b15zdnd00an1n02x5 FILLER_35_1467 ();
 b15zdnd00an1n01x5 FILLER_35_1469 ();
 b15zdnd11an1n04x5 FILLER_35_1473 ();
 b15zdnd11an1n64x5 FILLER_35_1480 ();
 b15zdnd11an1n32x5 FILLER_35_1544 ();
 b15zdnd11an1n16x5 FILLER_35_1576 ();
 b15zdnd11an1n08x5 FILLER_35_1592 ();
 b15zdnd00an1n02x5 FILLER_35_1600 ();
 b15zdnd11an1n64x5 FILLER_35_1605 ();
 b15zdnd11an1n64x5 FILLER_35_1669 ();
 b15zdnd11an1n32x5 FILLER_35_1733 ();
 b15zdnd11an1n16x5 FILLER_35_1765 ();
 b15zdnd11an1n04x5 FILLER_35_1784 ();
 b15zdnd11an1n64x5 FILLER_35_1791 ();
 b15zdnd11an1n32x5 FILLER_35_1855 ();
 b15zdnd11an1n16x5 FILLER_35_1887 ();
 b15zdnd11an1n08x5 FILLER_35_1903 ();
 b15zdnd11an1n04x5 FILLER_35_1911 ();
 b15zdnd00an1n02x5 FILLER_35_1915 ();
 b15zdnd00an1n01x5 FILLER_35_1917 ();
 b15zdnd11an1n04x5 FILLER_35_1921 ();
 b15zdnd11an1n04x5 FILLER_35_1928 ();
 b15zdnd11an1n04x5 FILLER_35_1935 ();
 b15zdnd11an1n64x5 FILLER_35_1942 ();
 b15zdnd11an1n64x5 FILLER_35_2006 ();
 b15zdnd11an1n64x5 FILLER_35_2070 ();
 b15zdnd11an1n64x5 FILLER_35_2134 ();
 b15zdnd11an1n64x5 FILLER_35_2198 ();
 b15zdnd11an1n16x5 FILLER_35_2262 ();
 b15zdnd11an1n04x5 FILLER_35_2278 ();
 b15zdnd00an1n02x5 FILLER_35_2282 ();
 b15zdnd11an1n64x5 FILLER_36_8 ();
 b15zdnd11an1n64x5 FILLER_36_72 ();
 b15zdnd11an1n64x5 FILLER_36_136 ();
 b15zdnd11an1n64x5 FILLER_36_200 ();
 b15zdnd11an1n64x5 FILLER_36_264 ();
 b15zdnd11an1n16x5 FILLER_36_328 ();
 b15zdnd11an1n04x5 FILLER_36_344 ();
 b15zdnd11an1n32x5 FILLER_36_400 ();
 b15zdnd11an1n16x5 FILLER_36_432 ();
 b15zdnd00an1n02x5 FILLER_36_448 ();
 b15zdnd11an1n64x5 FILLER_36_502 ();
 b15zdnd11an1n64x5 FILLER_36_566 ();
 b15zdnd11an1n64x5 FILLER_36_630 ();
 b15zdnd11an1n16x5 FILLER_36_694 ();
 b15zdnd11an1n08x5 FILLER_36_710 ();
 b15zdnd00an1n02x5 FILLER_36_726 ();
 b15zdnd00an1n01x5 FILLER_36_728 ();
 b15zdnd11an1n04x5 FILLER_36_732 ();
 b15zdnd11an1n64x5 FILLER_36_739 ();
 b15zdnd11an1n64x5 FILLER_36_803 ();
 b15zdnd11an1n64x5 FILLER_36_867 ();
 b15zdnd11an1n64x5 FILLER_36_931 ();
 b15zdnd11an1n64x5 FILLER_36_995 ();
 b15zdnd11an1n64x5 FILLER_36_1059 ();
 b15zdnd11an1n32x5 FILLER_36_1123 ();
 b15zdnd11an1n16x5 FILLER_36_1155 ();
 b15zdnd11an1n04x5 FILLER_36_1171 ();
 b15zdnd11an1n64x5 FILLER_36_1185 ();
 b15zdnd11an1n64x5 FILLER_36_1249 ();
 b15zdnd11an1n64x5 FILLER_36_1313 ();
 b15zdnd11an1n64x5 FILLER_36_1377 ();
 b15zdnd11an1n16x5 FILLER_36_1441 ();
 b15zdnd11an1n08x5 FILLER_36_1457 ();
 b15zdnd00an1n02x5 FILLER_36_1465 ();
 b15zdnd11an1n64x5 FILLER_36_1519 ();
 b15zdnd11an1n16x5 FILLER_36_1583 ();
 b15zdnd00an1n02x5 FILLER_36_1599 ();
 b15zdnd00an1n01x5 FILLER_36_1601 ();
 b15zdnd11an1n04x5 FILLER_36_1605 ();
 b15zdnd11an1n64x5 FILLER_36_1612 ();
 b15zdnd11an1n64x5 FILLER_36_1676 ();
 b15zdnd11an1n64x5 FILLER_36_1740 ();
 b15zdnd11an1n64x5 FILLER_36_1804 ();
 b15zdnd11an1n32x5 FILLER_36_1868 ();
 b15zdnd11an1n16x5 FILLER_36_1900 ();
 b15zdnd11an1n04x5 FILLER_36_1916 ();
 b15zdnd11an1n04x5 FILLER_36_1923 ();
 b15zdnd11an1n64x5 FILLER_36_1930 ();
 b15zdnd11an1n08x5 FILLER_36_1994 ();
 b15zdnd11an1n04x5 FILLER_36_2002 ();
 b15zdnd00an1n02x5 FILLER_36_2006 ();
 b15zdnd11an1n04x5 FILLER_36_2011 ();
 b15zdnd11an1n64x5 FILLER_36_2042 ();
 b15zdnd11an1n32x5 FILLER_36_2106 ();
 b15zdnd11an1n16x5 FILLER_36_2138 ();
 b15zdnd11an1n64x5 FILLER_36_2162 ();
 b15zdnd11an1n32x5 FILLER_36_2226 ();
 b15zdnd11an1n16x5 FILLER_36_2258 ();
 b15zdnd00an1n02x5 FILLER_36_2274 ();
 b15zdnd11an1n64x5 FILLER_37_0 ();
 b15zdnd11an1n64x5 FILLER_37_64 ();
 b15zdnd11an1n64x5 FILLER_37_128 ();
 b15zdnd11an1n64x5 FILLER_37_192 ();
 b15zdnd11an1n64x5 FILLER_37_256 ();
 b15zdnd11an1n32x5 FILLER_37_320 ();
 b15zdnd11an1n16x5 FILLER_37_352 ();
 b15zdnd00an1n01x5 FILLER_37_368 ();
 b15zdnd11an1n32x5 FILLER_37_421 ();
 b15zdnd11an1n64x5 FILLER_37_505 ();
 b15zdnd11an1n64x5 FILLER_37_569 ();
 b15zdnd11an1n32x5 FILLER_37_633 ();
 b15zdnd11an1n16x5 FILLER_37_665 ();
 b15zdnd11an1n04x5 FILLER_37_681 ();
 b15zdnd00an1n01x5 FILLER_37_685 ();
 b15zdnd11an1n64x5 FILLER_37_689 ();
 b15zdnd11an1n64x5 FILLER_37_770 ();
 b15zdnd11an1n32x5 FILLER_37_834 ();
 b15zdnd11an1n16x5 FILLER_37_866 ();
 b15zdnd11an1n64x5 FILLER_37_885 ();
 b15zdnd11an1n64x5 FILLER_37_949 ();
 b15zdnd11an1n64x5 FILLER_37_1013 ();
 b15zdnd11an1n64x5 FILLER_37_1077 ();
 b15zdnd11an1n64x5 FILLER_37_1141 ();
 b15zdnd11an1n64x5 FILLER_37_1205 ();
 b15zdnd11an1n64x5 FILLER_37_1269 ();
 b15zdnd11an1n64x5 FILLER_37_1333 ();
 b15zdnd11an1n64x5 FILLER_37_1397 ();
 b15zdnd11an1n16x5 FILLER_37_1461 ();
 b15zdnd11an1n08x5 FILLER_37_1477 ();
 b15zdnd11an1n04x5 FILLER_37_1488 ();
 b15zdnd11an1n64x5 FILLER_37_1495 ();
 b15zdnd11an1n16x5 FILLER_37_1559 ();
 b15zdnd11an1n04x5 FILLER_37_1575 ();
 b15zdnd11an1n64x5 FILLER_37_1631 ();
 b15zdnd11an1n64x5 FILLER_37_1695 ();
 b15zdnd11an1n64x5 FILLER_37_1759 ();
 b15zdnd11an1n64x5 FILLER_37_1823 ();
 b15zdnd11an1n64x5 FILLER_37_1887 ();
 b15zdnd11an1n64x5 FILLER_37_1951 ();
 b15zdnd11an1n64x5 FILLER_37_2015 ();
 b15zdnd11an1n64x5 FILLER_37_2079 ();
 b15zdnd11an1n64x5 FILLER_37_2143 ();
 b15zdnd11an1n16x5 FILLER_37_2207 ();
 b15zdnd11an1n16x5 FILLER_37_2265 ();
 b15zdnd00an1n02x5 FILLER_37_2281 ();
 b15zdnd00an1n01x5 FILLER_37_2283 ();
 b15zdnd11an1n64x5 FILLER_38_8 ();
 b15zdnd11an1n64x5 FILLER_38_72 ();
 b15zdnd11an1n64x5 FILLER_38_136 ();
 b15zdnd11an1n64x5 FILLER_38_200 ();
 b15zdnd11an1n64x5 FILLER_38_264 ();
 b15zdnd11an1n32x5 FILLER_38_328 ();
 b15zdnd11an1n04x5 FILLER_38_360 ();
 b15zdnd00an1n01x5 FILLER_38_364 ();
 b15zdnd11an1n04x5 FILLER_38_368 ();
 b15zdnd11an1n08x5 FILLER_38_375 ();
 b15zdnd00an1n02x5 FILLER_38_383 ();
 b15zdnd00an1n01x5 FILLER_38_385 ();
 b15zdnd11an1n04x5 FILLER_38_389 ();
 b15zdnd11an1n64x5 FILLER_38_396 ();
 b15zdnd11an1n04x5 FILLER_38_460 ();
 b15zdnd00an1n01x5 FILLER_38_464 ();
 b15zdnd11an1n04x5 FILLER_38_468 ();
 b15zdnd11an1n04x5 FILLER_38_475 ();
 b15zdnd11an1n04x5 FILLER_38_482 ();
 b15zdnd11an1n64x5 FILLER_38_489 ();
 b15zdnd11an1n32x5 FILLER_38_553 ();
 b15zdnd11an1n08x5 FILLER_38_585 ();
 b15zdnd00an1n02x5 FILLER_38_593 ();
 b15zdnd00an1n01x5 FILLER_38_595 ();
 b15zdnd11an1n64x5 FILLER_38_599 ();
 b15zdnd00an1n01x5 FILLER_38_663 ();
 b15zdnd00an1n02x5 FILLER_38_716 ();
 b15zdnd11an1n64x5 FILLER_38_726 ();
 b15zdnd11an1n32x5 FILLER_38_790 ();
 b15zdnd11an1n16x5 FILLER_38_822 ();
 b15zdnd11an1n08x5 FILLER_38_838 ();
 b15zdnd00an1n02x5 FILLER_38_846 ();
 b15zdnd00an1n01x5 FILLER_38_848 ();
 b15zdnd11an1n04x5 FILLER_38_876 ();
 b15zdnd11an1n04x5 FILLER_38_883 ();
 b15zdnd11an1n64x5 FILLER_38_890 ();
 b15zdnd11an1n64x5 FILLER_38_954 ();
 b15zdnd11an1n64x5 FILLER_38_1018 ();
 b15zdnd11an1n64x5 FILLER_38_1082 ();
 b15zdnd11an1n64x5 FILLER_38_1146 ();
 b15zdnd11an1n32x5 FILLER_38_1210 ();
 b15zdnd11an1n16x5 FILLER_38_1242 ();
 b15zdnd11an1n08x5 FILLER_38_1258 ();
 b15zdnd11an1n04x5 FILLER_38_1266 ();
 b15zdnd00an1n01x5 FILLER_38_1270 ();
 b15zdnd11an1n64x5 FILLER_38_1278 ();
 b15zdnd11an1n64x5 FILLER_38_1342 ();
 b15zdnd11an1n64x5 FILLER_38_1406 ();
 b15zdnd11an1n16x5 FILLER_38_1470 ();
 b15zdnd11an1n04x5 FILLER_38_1486 ();
 b15zdnd00an1n01x5 FILLER_38_1490 ();
 b15zdnd11an1n64x5 FILLER_38_1494 ();
 b15zdnd11an1n64x5 FILLER_38_1558 ();
 b15zdnd11an1n64x5 FILLER_38_1622 ();
 b15zdnd11an1n64x5 FILLER_38_1686 ();
 b15zdnd11an1n64x5 FILLER_38_1750 ();
 b15zdnd11an1n64x5 FILLER_38_1814 ();
 b15zdnd11an1n64x5 FILLER_38_1878 ();
 b15zdnd11an1n64x5 FILLER_38_1942 ();
 b15zdnd11an1n64x5 FILLER_38_2006 ();
 b15zdnd11an1n64x5 FILLER_38_2070 ();
 b15zdnd11an1n16x5 FILLER_38_2134 ();
 b15zdnd11an1n04x5 FILLER_38_2150 ();
 b15zdnd11an1n16x5 FILLER_38_2162 ();
 b15zdnd11an1n08x5 FILLER_38_2178 ();
 b15zdnd00an1n02x5 FILLER_38_2186 ();
 b15zdnd11an1n32x5 FILLER_38_2230 ();
 b15zdnd11an1n08x5 FILLER_38_2262 ();
 b15zdnd11an1n04x5 FILLER_38_2270 ();
 b15zdnd00an1n02x5 FILLER_38_2274 ();
 b15zdnd11an1n64x5 FILLER_39_0 ();
 b15zdnd11an1n64x5 FILLER_39_64 ();
 b15zdnd11an1n64x5 FILLER_39_128 ();
 b15zdnd11an1n64x5 FILLER_39_192 ();
 b15zdnd11an1n64x5 FILLER_39_256 ();
 b15zdnd11an1n64x5 FILLER_39_320 ();
 b15zdnd11an1n08x5 FILLER_39_384 ();
 b15zdnd00an1n02x5 FILLER_39_392 ();
 b15zdnd11an1n64x5 FILLER_39_397 ();
 b15zdnd11an1n08x5 FILLER_39_461 ();
 b15zdnd11an1n04x5 FILLER_39_469 ();
 b15zdnd00an1n02x5 FILLER_39_473 ();
 b15zdnd00an1n01x5 FILLER_39_475 ();
 b15zdnd11an1n64x5 FILLER_39_479 ();
 b15zdnd11an1n16x5 FILLER_39_543 ();
 b15zdnd11an1n08x5 FILLER_39_559 ();
 b15zdnd00an1n02x5 FILLER_39_567 ();
 b15zdnd11an1n64x5 FILLER_39_621 ();
 b15zdnd11an1n04x5 FILLER_39_688 ();
 b15zdnd00an1n01x5 FILLER_39_692 ();
 b15zdnd11an1n64x5 FILLER_39_696 ();
 b15zdnd11an1n64x5 FILLER_39_760 ();
 b15zdnd11an1n16x5 FILLER_39_824 ();
 b15zdnd11an1n08x5 FILLER_39_840 ();
 b15zdnd00an1n02x5 FILLER_39_848 ();
 b15zdnd11an1n04x5 FILLER_39_853 ();
 b15zdnd11an1n64x5 FILLER_39_909 ();
 b15zdnd11an1n64x5 FILLER_39_973 ();
 b15zdnd11an1n64x5 FILLER_39_1037 ();
 b15zdnd11an1n64x5 FILLER_39_1101 ();
 b15zdnd11an1n64x5 FILLER_39_1165 ();
 b15zdnd11an1n32x5 FILLER_39_1229 ();
 b15zdnd11an1n04x5 FILLER_39_1261 ();
 b15zdnd00an1n01x5 FILLER_39_1265 ();
 b15zdnd11an1n08x5 FILLER_39_1278 ();
 b15zdnd00an1n01x5 FILLER_39_1286 ();
 b15zdnd11an1n32x5 FILLER_39_1292 ();
 b15zdnd11an1n16x5 FILLER_39_1324 ();
 b15zdnd11an1n08x5 FILLER_39_1340 ();
 b15zdnd00an1n02x5 FILLER_39_1348 ();
 b15zdnd00an1n01x5 FILLER_39_1350 ();
 b15zdnd11an1n04x5 FILLER_39_1383 ();
 b15zdnd11an1n04x5 FILLER_39_1390 ();
 b15zdnd11an1n64x5 FILLER_39_1397 ();
 b15zdnd11an1n64x5 FILLER_39_1461 ();
 b15zdnd11an1n64x5 FILLER_39_1525 ();
 b15zdnd11an1n64x5 FILLER_39_1589 ();
 b15zdnd11an1n64x5 FILLER_39_1653 ();
 b15zdnd11an1n64x5 FILLER_39_1717 ();
 b15zdnd11an1n64x5 FILLER_39_1781 ();
 b15zdnd11an1n64x5 FILLER_39_1845 ();
 b15zdnd11an1n64x5 FILLER_39_1909 ();
 b15zdnd11an1n64x5 FILLER_39_1973 ();
 b15zdnd11an1n64x5 FILLER_39_2037 ();
 b15zdnd11an1n64x5 FILLER_39_2101 ();
 b15zdnd11an1n64x5 FILLER_39_2165 ();
 b15zdnd11an1n32x5 FILLER_39_2229 ();
 b15zdnd11an1n16x5 FILLER_39_2261 ();
 b15zdnd11an1n04x5 FILLER_39_2277 ();
 b15zdnd00an1n02x5 FILLER_39_2281 ();
 b15zdnd00an1n01x5 FILLER_39_2283 ();
 b15zdnd11an1n64x5 FILLER_40_8 ();
 b15zdnd11an1n64x5 FILLER_40_72 ();
 b15zdnd11an1n64x5 FILLER_40_136 ();
 b15zdnd11an1n64x5 FILLER_40_200 ();
 b15zdnd11an1n64x5 FILLER_40_264 ();
 b15zdnd11an1n64x5 FILLER_40_328 ();
 b15zdnd11an1n64x5 FILLER_40_392 ();
 b15zdnd11an1n64x5 FILLER_40_456 ();
 b15zdnd11an1n64x5 FILLER_40_520 ();
 b15zdnd11an1n04x5 FILLER_40_584 ();
 b15zdnd11an1n04x5 FILLER_40_591 ();
 b15zdnd11an1n64x5 FILLER_40_598 ();
 b15zdnd11an1n32x5 FILLER_40_662 ();
 b15zdnd11an1n16x5 FILLER_40_694 ();
 b15zdnd11an1n08x5 FILLER_40_710 ();
 b15zdnd11an1n64x5 FILLER_40_726 ();
 b15zdnd11an1n64x5 FILLER_40_790 ();
 b15zdnd11an1n04x5 FILLER_40_854 ();
 b15zdnd00an1n02x5 FILLER_40_858 ();
 b15zdnd00an1n01x5 FILLER_40_860 ();
 b15zdnd11an1n08x5 FILLER_40_864 ();
 b15zdnd00an1n02x5 FILLER_40_872 ();
 b15zdnd11an1n04x5 FILLER_40_877 ();
 b15zdnd00an1n02x5 FILLER_40_881 ();
 b15zdnd11an1n64x5 FILLER_40_886 ();
 b15zdnd11an1n64x5 FILLER_40_950 ();
 b15zdnd11an1n64x5 FILLER_40_1014 ();
 b15zdnd11an1n64x5 FILLER_40_1078 ();
 b15zdnd11an1n16x5 FILLER_40_1142 ();
 b15zdnd00an1n02x5 FILLER_40_1158 ();
 b15zdnd11an1n64x5 FILLER_40_1181 ();
 b15zdnd11an1n64x5 FILLER_40_1245 ();
 b15zdnd11an1n64x5 FILLER_40_1309 ();
 b15zdnd11an1n64x5 FILLER_40_1373 ();
 b15zdnd11an1n64x5 FILLER_40_1437 ();
 b15zdnd11an1n32x5 FILLER_40_1501 ();
 b15zdnd11an1n08x5 FILLER_40_1533 ();
 b15zdnd00an1n02x5 FILLER_40_1541 ();
 b15zdnd00an1n01x5 FILLER_40_1543 ();
 b15zdnd11an1n64x5 FILLER_40_1553 ();
 b15zdnd11an1n64x5 FILLER_40_1617 ();
 b15zdnd11an1n16x5 FILLER_40_1681 ();
 b15zdnd11an1n08x5 FILLER_40_1697 ();
 b15zdnd11an1n04x5 FILLER_40_1705 ();
 b15zdnd00an1n01x5 FILLER_40_1709 ();
 b15zdnd11an1n64x5 FILLER_40_1719 ();
 b15zdnd11an1n64x5 FILLER_40_1783 ();
 b15zdnd11an1n64x5 FILLER_40_1847 ();
 b15zdnd11an1n16x5 FILLER_40_1911 ();
 b15zdnd11an1n04x5 FILLER_40_1927 ();
 b15zdnd00an1n01x5 FILLER_40_1931 ();
 b15zdnd11an1n32x5 FILLER_40_1941 ();
 b15zdnd11an1n08x5 FILLER_40_1973 ();
 b15zdnd11an1n04x5 FILLER_40_1981 ();
 b15zdnd00an1n02x5 FILLER_40_1985 ();
 b15zdnd00an1n01x5 FILLER_40_1987 ();
 b15zdnd11an1n64x5 FILLER_40_1997 ();
 b15zdnd11an1n64x5 FILLER_40_2061 ();
 b15zdnd11an1n16x5 FILLER_40_2125 ();
 b15zdnd11an1n08x5 FILLER_40_2141 ();
 b15zdnd11an1n04x5 FILLER_40_2149 ();
 b15zdnd00an1n01x5 FILLER_40_2153 ();
 b15zdnd11an1n64x5 FILLER_40_2162 ();
 b15zdnd11an1n32x5 FILLER_40_2226 ();
 b15zdnd11an1n16x5 FILLER_40_2258 ();
 b15zdnd00an1n02x5 FILLER_40_2274 ();
 b15zdnd11an1n64x5 FILLER_41_0 ();
 b15zdnd11an1n64x5 FILLER_41_64 ();
 b15zdnd11an1n64x5 FILLER_41_128 ();
 b15zdnd11an1n64x5 FILLER_41_192 ();
 b15zdnd11an1n64x5 FILLER_41_256 ();
 b15zdnd11an1n64x5 FILLER_41_320 ();
 b15zdnd11an1n64x5 FILLER_41_384 ();
 b15zdnd11an1n64x5 FILLER_41_448 ();
 b15zdnd11an1n64x5 FILLER_41_512 ();
 b15zdnd11an1n64x5 FILLER_41_576 ();
 b15zdnd11an1n64x5 FILLER_41_640 ();
 b15zdnd11an1n64x5 FILLER_41_704 ();
 b15zdnd11an1n64x5 FILLER_41_768 ();
 b15zdnd11an1n04x5 FILLER_41_832 ();
 b15zdnd00an1n02x5 FILLER_41_836 ();
 b15zdnd00an1n01x5 FILLER_41_838 ();
 b15zdnd11an1n64x5 FILLER_41_891 ();
 b15zdnd11an1n64x5 FILLER_41_955 ();
 b15zdnd11an1n64x5 FILLER_41_1019 ();
 b15zdnd11an1n64x5 FILLER_41_1083 ();
 b15zdnd11an1n16x5 FILLER_41_1151 ();
 b15zdnd11an1n64x5 FILLER_41_1179 ();
 b15zdnd11an1n16x5 FILLER_41_1243 ();
 b15zdnd11an1n64x5 FILLER_41_1263 ();
 b15zdnd11an1n64x5 FILLER_41_1327 ();
 b15zdnd11an1n64x5 FILLER_41_1391 ();
 b15zdnd11an1n64x5 FILLER_41_1455 ();
 b15zdnd11an1n64x5 FILLER_41_1519 ();
 b15zdnd11an1n64x5 FILLER_41_1583 ();
 b15zdnd11an1n64x5 FILLER_41_1647 ();
 b15zdnd11an1n64x5 FILLER_41_1711 ();
 b15zdnd11an1n64x5 FILLER_41_1775 ();
 b15zdnd11an1n64x5 FILLER_41_1839 ();
 b15zdnd11an1n64x5 FILLER_41_1903 ();
 b15zdnd11an1n64x5 FILLER_41_1967 ();
 b15zdnd11an1n64x5 FILLER_41_2031 ();
 b15zdnd11an1n64x5 FILLER_41_2095 ();
 b15zdnd11an1n64x5 FILLER_41_2159 ();
 b15zdnd11an1n32x5 FILLER_41_2223 ();
 b15zdnd11an1n16x5 FILLER_41_2255 ();
 b15zdnd11an1n08x5 FILLER_41_2271 ();
 b15zdnd11an1n04x5 FILLER_41_2279 ();
 b15zdnd00an1n01x5 FILLER_41_2283 ();
 b15zdnd11an1n64x5 FILLER_42_8 ();
 b15zdnd11an1n64x5 FILLER_42_72 ();
 b15zdnd11an1n64x5 FILLER_42_136 ();
 b15zdnd11an1n64x5 FILLER_42_200 ();
 b15zdnd11an1n64x5 FILLER_42_264 ();
 b15zdnd11an1n64x5 FILLER_42_328 ();
 b15zdnd11an1n64x5 FILLER_42_392 ();
 b15zdnd11an1n64x5 FILLER_42_456 ();
 b15zdnd11an1n64x5 FILLER_42_520 ();
 b15zdnd11an1n64x5 FILLER_42_584 ();
 b15zdnd11an1n08x5 FILLER_42_648 ();
 b15zdnd11an1n32x5 FILLER_42_673 ();
 b15zdnd11an1n08x5 FILLER_42_705 ();
 b15zdnd11an1n04x5 FILLER_42_713 ();
 b15zdnd00an1n01x5 FILLER_42_717 ();
 b15zdnd11an1n64x5 FILLER_42_726 ();
 b15zdnd11an1n64x5 FILLER_42_790 ();
 b15zdnd11an1n64x5 FILLER_42_854 ();
 b15zdnd11an1n64x5 FILLER_42_918 ();
 b15zdnd11an1n64x5 FILLER_42_982 ();
 b15zdnd11an1n64x5 FILLER_42_1046 ();
 b15zdnd11an1n32x5 FILLER_42_1110 ();
 b15zdnd11an1n08x5 FILLER_42_1142 ();
 b15zdnd00an1n02x5 FILLER_42_1150 ();
 b15zdnd11an1n04x5 FILLER_42_1160 ();
 b15zdnd11an1n08x5 FILLER_42_1170 ();
 b15zdnd11an1n04x5 FILLER_42_1178 ();
 b15zdnd00an1n02x5 FILLER_42_1182 ();
 b15zdnd11an1n64x5 FILLER_42_1188 ();
 b15zdnd11an1n64x5 FILLER_42_1267 ();
 b15zdnd11an1n64x5 FILLER_42_1331 ();
 b15zdnd11an1n64x5 FILLER_42_1395 ();
 b15zdnd11an1n64x5 FILLER_42_1459 ();
 b15zdnd11an1n64x5 FILLER_42_1523 ();
 b15zdnd11an1n64x5 FILLER_42_1587 ();
 b15zdnd11an1n64x5 FILLER_42_1651 ();
 b15zdnd11an1n64x5 FILLER_42_1715 ();
 b15zdnd11an1n64x5 FILLER_42_1779 ();
 b15zdnd11an1n64x5 FILLER_42_1843 ();
 b15zdnd11an1n64x5 FILLER_42_1907 ();
 b15zdnd11an1n04x5 FILLER_42_1971 ();
 b15zdnd00an1n02x5 FILLER_42_1975 ();
 b15zdnd11an1n32x5 FILLER_42_1986 ();
 b15zdnd11an1n08x5 FILLER_42_2018 ();
 b15zdnd00an1n02x5 FILLER_42_2026 ();
 b15zdnd00an1n01x5 FILLER_42_2028 ();
 b15zdnd11an1n64x5 FILLER_42_2032 ();
 b15zdnd11an1n32x5 FILLER_42_2096 ();
 b15zdnd11an1n16x5 FILLER_42_2128 ();
 b15zdnd11an1n08x5 FILLER_42_2144 ();
 b15zdnd00an1n02x5 FILLER_42_2152 ();
 b15zdnd11an1n64x5 FILLER_42_2162 ();
 b15zdnd11an1n32x5 FILLER_42_2226 ();
 b15zdnd11an1n16x5 FILLER_42_2258 ();
 b15zdnd00an1n02x5 FILLER_42_2274 ();
 b15zdnd11an1n64x5 FILLER_43_0 ();
 b15zdnd11an1n64x5 FILLER_43_64 ();
 b15zdnd11an1n64x5 FILLER_43_128 ();
 b15zdnd11an1n64x5 FILLER_43_192 ();
 b15zdnd11an1n64x5 FILLER_43_256 ();
 b15zdnd11an1n64x5 FILLER_43_320 ();
 b15zdnd11an1n64x5 FILLER_43_384 ();
 b15zdnd11an1n64x5 FILLER_43_448 ();
 b15zdnd11an1n64x5 FILLER_43_512 ();
 b15zdnd11an1n64x5 FILLER_43_576 ();
 b15zdnd11an1n64x5 FILLER_43_640 ();
 b15zdnd11an1n64x5 FILLER_43_704 ();
 b15zdnd11an1n64x5 FILLER_43_768 ();
 b15zdnd11an1n64x5 FILLER_43_832 ();
 b15zdnd11an1n64x5 FILLER_43_896 ();
 b15zdnd11an1n64x5 FILLER_43_960 ();
 b15zdnd11an1n64x5 FILLER_43_1024 ();
 b15zdnd11an1n64x5 FILLER_43_1088 ();
 b15zdnd11an1n08x5 FILLER_43_1152 ();
 b15zdnd11an1n08x5 FILLER_43_1174 ();
 b15zdnd00an1n02x5 FILLER_43_1182 ();
 b15zdnd00an1n01x5 FILLER_43_1184 ();
 b15zdnd11an1n64x5 FILLER_43_1188 ();
 b15zdnd11an1n64x5 FILLER_43_1252 ();
 b15zdnd11an1n64x5 FILLER_43_1316 ();
 b15zdnd11an1n64x5 FILLER_43_1380 ();
 b15zdnd11an1n64x5 FILLER_43_1444 ();
 b15zdnd11an1n64x5 FILLER_43_1508 ();
 b15zdnd11an1n64x5 FILLER_43_1572 ();
 b15zdnd11an1n32x5 FILLER_43_1636 ();
 b15zdnd11an1n08x5 FILLER_43_1668 ();
 b15zdnd11an1n04x5 FILLER_43_1679 ();
 b15zdnd11an1n64x5 FILLER_43_1686 ();
 b15zdnd11an1n64x5 FILLER_43_1750 ();
 b15zdnd11an1n64x5 FILLER_43_1814 ();
 b15zdnd11an1n64x5 FILLER_43_1878 ();
 b15zdnd11an1n64x5 FILLER_43_1942 ();
 b15zdnd11an1n16x5 FILLER_43_2006 ();
 b15zdnd11an1n04x5 FILLER_43_2022 ();
 b15zdnd00an1n02x5 FILLER_43_2026 ();
 b15zdnd00an1n01x5 FILLER_43_2028 ();
 b15zdnd11an1n04x5 FILLER_43_2032 ();
 b15zdnd11an1n64x5 FILLER_43_2039 ();
 b15zdnd11an1n64x5 FILLER_43_2103 ();
 b15zdnd11an1n64x5 FILLER_43_2167 ();
 b15zdnd11an1n32x5 FILLER_43_2231 ();
 b15zdnd11an1n16x5 FILLER_43_2263 ();
 b15zdnd11an1n04x5 FILLER_43_2279 ();
 b15zdnd00an1n01x5 FILLER_43_2283 ();
 b15zdnd11an1n64x5 FILLER_44_8 ();
 b15zdnd11an1n64x5 FILLER_44_72 ();
 b15zdnd11an1n64x5 FILLER_44_136 ();
 b15zdnd11an1n64x5 FILLER_44_200 ();
 b15zdnd11an1n64x5 FILLER_44_264 ();
 b15zdnd11an1n64x5 FILLER_44_328 ();
 b15zdnd11an1n64x5 FILLER_44_392 ();
 b15zdnd11an1n64x5 FILLER_44_456 ();
 b15zdnd11an1n64x5 FILLER_44_520 ();
 b15zdnd11an1n64x5 FILLER_44_584 ();
 b15zdnd11an1n64x5 FILLER_44_648 ();
 b15zdnd11an1n04x5 FILLER_44_712 ();
 b15zdnd00an1n02x5 FILLER_44_716 ();
 b15zdnd11an1n64x5 FILLER_44_726 ();
 b15zdnd11an1n64x5 FILLER_44_790 ();
 b15zdnd11an1n64x5 FILLER_44_854 ();
 b15zdnd11an1n64x5 FILLER_44_918 ();
 b15zdnd11an1n64x5 FILLER_44_982 ();
 b15zdnd11an1n64x5 FILLER_44_1046 ();
 b15zdnd11an1n32x5 FILLER_44_1110 ();
 b15zdnd11an1n08x5 FILLER_44_1142 ();
 b15zdnd11an1n64x5 FILLER_44_1156 ();
 b15zdnd11an1n32x5 FILLER_44_1220 ();
 b15zdnd11an1n16x5 FILLER_44_1252 ();
 b15zdnd11an1n08x5 FILLER_44_1268 ();
 b15zdnd11an1n04x5 FILLER_44_1276 ();
 b15zdnd11an1n04x5 FILLER_44_1322 ();
 b15zdnd00an1n02x5 FILLER_44_1326 ();
 b15zdnd00an1n01x5 FILLER_44_1328 ();
 b15zdnd11an1n64x5 FILLER_44_1371 ();
 b15zdnd11an1n32x5 FILLER_44_1435 ();
 b15zdnd11an1n16x5 FILLER_44_1467 ();
 b15zdnd11an1n04x5 FILLER_44_1483 ();
 b15zdnd00an1n02x5 FILLER_44_1487 ();
 b15zdnd11an1n08x5 FILLER_44_1531 ();
 b15zdnd00an1n02x5 FILLER_44_1539 ();
 b15zdnd11an1n64x5 FILLER_44_1583 ();
 b15zdnd11an1n04x5 FILLER_44_1647 ();
 b15zdnd11an1n32x5 FILLER_44_1703 ();
 b15zdnd00an1n02x5 FILLER_44_1735 ();
 b15zdnd00an1n01x5 FILLER_44_1737 ();
 b15zdnd11an1n64x5 FILLER_44_1747 ();
 b15zdnd11an1n64x5 FILLER_44_1811 ();
 b15zdnd11an1n64x5 FILLER_44_1875 ();
 b15zdnd11an1n64x5 FILLER_44_1939 ();
 b15zdnd00an1n02x5 FILLER_44_2003 ();
 b15zdnd00an1n01x5 FILLER_44_2005 ();
 b15zdnd11an1n64x5 FILLER_44_2058 ();
 b15zdnd11an1n32x5 FILLER_44_2122 ();
 b15zdnd11an1n64x5 FILLER_44_2162 ();
 b15zdnd11an1n32x5 FILLER_44_2226 ();
 b15zdnd11an1n16x5 FILLER_44_2258 ();
 b15zdnd00an1n02x5 FILLER_44_2274 ();
 b15zdnd11an1n64x5 FILLER_45_0 ();
 b15zdnd11an1n64x5 FILLER_45_64 ();
 b15zdnd11an1n64x5 FILLER_45_128 ();
 b15zdnd11an1n64x5 FILLER_45_192 ();
 b15zdnd11an1n64x5 FILLER_45_256 ();
 b15zdnd11an1n64x5 FILLER_45_320 ();
 b15zdnd11an1n64x5 FILLER_45_384 ();
 b15zdnd11an1n64x5 FILLER_45_448 ();
 b15zdnd11an1n64x5 FILLER_45_512 ();
 b15zdnd11an1n32x5 FILLER_45_576 ();
 b15zdnd11an1n16x5 FILLER_45_608 ();
 b15zdnd00an1n02x5 FILLER_45_624 ();
 b15zdnd00an1n01x5 FILLER_45_626 ();
 b15zdnd11an1n32x5 FILLER_45_636 ();
 b15zdnd00an1n01x5 FILLER_45_668 ();
 b15zdnd11an1n04x5 FILLER_45_678 ();
 b15zdnd11an1n64x5 FILLER_45_691 ();
 b15zdnd11an1n64x5 FILLER_45_755 ();
 b15zdnd11an1n64x5 FILLER_45_819 ();
 b15zdnd11an1n64x5 FILLER_45_883 ();
 b15zdnd11an1n64x5 FILLER_45_947 ();
 b15zdnd11an1n64x5 FILLER_45_1011 ();
 b15zdnd11an1n64x5 FILLER_45_1075 ();
 b15zdnd11an1n64x5 FILLER_45_1139 ();
 b15zdnd11an1n64x5 FILLER_45_1203 ();
 b15zdnd00an1n02x5 FILLER_45_1267 ();
 b15zdnd11an1n16x5 FILLER_45_1273 ();
 b15zdnd11an1n64x5 FILLER_45_1292 ();
 b15zdnd11an1n64x5 FILLER_45_1356 ();
 b15zdnd11an1n64x5 FILLER_45_1420 ();
 b15zdnd11an1n64x5 FILLER_45_1484 ();
 b15zdnd11an1n64x5 FILLER_45_1548 ();
 b15zdnd11an1n64x5 FILLER_45_1612 ();
 b15zdnd11an1n32x5 FILLER_45_1679 ();
 b15zdnd11an1n16x5 FILLER_45_1711 ();
 b15zdnd11an1n08x5 FILLER_45_1727 ();
 b15zdnd11an1n04x5 FILLER_45_1735 ();
 b15zdnd11an1n64x5 FILLER_45_1748 ();
 b15zdnd11an1n64x5 FILLER_45_1812 ();
 b15zdnd11an1n64x5 FILLER_45_1876 ();
 b15zdnd11an1n64x5 FILLER_45_1940 ();
 b15zdnd11an1n64x5 FILLER_45_2004 ();
 b15zdnd11an1n64x5 FILLER_45_2068 ();
 b15zdnd11an1n64x5 FILLER_45_2132 ();
 b15zdnd11an1n64x5 FILLER_45_2196 ();
 b15zdnd11an1n16x5 FILLER_45_2260 ();
 b15zdnd11an1n08x5 FILLER_45_2276 ();
 b15zdnd11an1n64x5 FILLER_46_8 ();
 b15zdnd11an1n64x5 FILLER_46_72 ();
 b15zdnd11an1n64x5 FILLER_46_136 ();
 b15zdnd11an1n64x5 FILLER_46_200 ();
 b15zdnd11an1n64x5 FILLER_46_264 ();
 b15zdnd11an1n64x5 FILLER_46_328 ();
 b15zdnd11an1n64x5 FILLER_46_392 ();
 b15zdnd11an1n64x5 FILLER_46_456 ();
 b15zdnd11an1n64x5 FILLER_46_520 ();
 b15zdnd11an1n64x5 FILLER_46_584 ();
 b15zdnd11an1n64x5 FILLER_46_648 ();
 b15zdnd11an1n04x5 FILLER_46_712 ();
 b15zdnd00an1n02x5 FILLER_46_716 ();
 b15zdnd11an1n64x5 FILLER_46_726 ();
 b15zdnd11an1n64x5 FILLER_46_790 ();
 b15zdnd11an1n64x5 FILLER_46_854 ();
 b15zdnd11an1n64x5 FILLER_46_918 ();
 b15zdnd11an1n64x5 FILLER_46_982 ();
 b15zdnd11an1n64x5 FILLER_46_1046 ();
 b15zdnd11an1n64x5 FILLER_46_1110 ();
 b15zdnd11an1n64x5 FILLER_46_1174 ();
 b15zdnd11an1n04x5 FILLER_46_1238 ();
 b15zdnd00an1n02x5 FILLER_46_1242 ();
 b15zdnd11an1n04x5 FILLER_46_1256 ();
 b15zdnd11an1n64x5 FILLER_46_1268 ();
 b15zdnd11an1n64x5 FILLER_46_1332 ();
 b15zdnd11an1n64x5 FILLER_46_1396 ();
 b15zdnd11an1n64x5 FILLER_46_1460 ();
 b15zdnd11an1n64x5 FILLER_46_1524 ();
 b15zdnd11an1n64x5 FILLER_46_1588 ();
 b15zdnd11an1n64x5 FILLER_46_1652 ();
 b15zdnd11an1n64x5 FILLER_46_1716 ();
 b15zdnd11an1n64x5 FILLER_46_1780 ();
 b15zdnd11an1n64x5 FILLER_46_1844 ();
 b15zdnd11an1n64x5 FILLER_46_1908 ();
 b15zdnd11an1n64x5 FILLER_46_1972 ();
 b15zdnd11an1n64x5 FILLER_46_2036 ();
 b15zdnd11an1n32x5 FILLER_46_2100 ();
 b15zdnd11an1n16x5 FILLER_46_2132 ();
 b15zdnd11an1n04x5 FILLER_46_2148 ();
 b15zdnd00an1n02x5 FILLER_46_2152 ();
 b15zdnd11an1n64x5 FILLER_46_2162 ();
 b15zdnd11an1n32x5 FILLER_46_2226 ();
 b15zdnd11an1n16x5 FILLER_46_2258 ();
 b15zdnd00an1n02x5 FILLER_46_2274 ();
 b15zdnd11an1n64x5 FILLER_47_0 ();
 b15zdnd11an1n64x5 FILLER_47_64 ();
 b15zdnd11an1n64x5 FILLER_47_128 ();
 b15zdnd11an1n64x5 FILLER_47_192 ();
 b15zdnd11an1n64x5 FILLER_47_256 ();
 b15zdnd11an1n64x5 FILLER_47_320 ();
 b15zdnd11an1n64x5 FILLER_47_384 ();
 b15zdnd11an1n64x5 FILLER_47_448 ();
 b15zdnd11an1n64x5 FILLER_47_532 ();
 b15zdnd11an1n64x5 FILLER_47_596 ();
 b15zdnd11an1n64x5 FILLER_47_660 ();
 b15zdnd11an1n64x5 FILLER_47_724 ();
 b15zdnd11an1n64x5 FILLER_47_788 ();
 b15zdnd11an1n64x5 FILLER_47_852 ();
 b15zdnd11an1n64x5 FILLER_47_916 ();
 b15zdnd11an1n64x5 FILLER_47_980 ();
 b15zdnd11an1n64x5 FILLER_47_1044 ();
 b15zdnd11an1n64x5 FILLER_47_1108 ();
 b15zdnd11an1n64x5 FILLER_47_1172 ();
 b15zdnd11an1n16x5 FILLER_47_1236 ();
 b15zdnd11an1n08x5 FILLER_47_1252 ();
 b15zdnd11an1n04x5 FILLER_47_1260 ();
 b15zdnd00an1n02x5 FILLER_47_1264 ();
 b15zdnd00an1n01x5 FILLER_47_1266 ();
 b15zdnd11an1n64x5 FILLER_47_1273 ();
 b15zdnd11an1n64x5 FILLER_47_1337 ();
 b15zdnd11an1n64x5 FILLER_47_1401 ();
 b15zdnd11an1n64x5 FILLER_47_1465 ();
 b15zdnd11an1n16x5 FILLER_47_1529 ();
 b15zdnd11an1n64x5 FILLER_47_1554 ();
 b15zdnd11an1n64x5 FILLER_47_1618 ();
 b15zdnd11an1n64x5 FILLER_47_1682 ();
 b15zdnd11an1n64x5 FILLER_47_1746 ();
 b15zdnd11an1n64x5 FILLER_47_1810 ();
 b15zdnd11an1n64x5 FILLER_47_1874 ();
 b15zdnd11an1n64x5 FILLER_47_1938 ();
 b15zdnd11an1n64x5 FILLER_47_2002 ();
 b15zdnd11an1n64x5 FILLER_47_2066 ();
 b15zdnd11an1n64x5 FILLER_47_2130 ();
 b15zdnd11an1n64x5 FILLER_47_2194 ();
 b15zdnd11an1n16x5 FILLER_47_2258 ();
 b15zdnd11an1n08x5 FILLER_47_2274 ();
 b15zdnd00an1n02x5 FILLER_47_2282 ();
 b15zdnd11an1n64x5 FILLER_48_8 ();
 b15zdnd11an1n64x5 FILLER_48_72 ();
 b15zdnd11an1n64x5 FILLER_48_136 ();
 b15zdnd11an1n64x5 FILLER_48_200 ();
 b15zdnd11an1n64x5 FILLER_48_264 ();
 b15zdnd11an1n64x5 FILLER_48_328 ();
 b15zdnd11an1n64x5 FILLER_48_392 ();
 b15zdnd11an1n64x5 FILLER_48_456 ();
 b15zdnd11an1n64x5 FILLER_48_520 ();
 b15zdnd11an1n64x5 FILLER_48_584 ();
 b15zdnd11an1n64x5 FILLER_48_648 ();
 b15zdnd11an1n04x5 FILLER_48_712 ();
 b15zdnd00an1n02x5 FILLER_48_716 ();
 b15zdnd11an1n64x5 FILLER_48_726 ();
 b15zdnd11an1n64x5 FILLER_48_790 ();
 b15zdnd11an1n64x5 FILLER_48_854 ();
 b15zdnd11an1n64x5 FILLER_48_918 ();
 b15zdnd11an1n64x5 FILLER_48_982 ();
 b15zdnd11an1n16x5 FILLER_48_1046 ();
 b15zdnd11an1n64x5 FILLER_48_1104 ();
 b15zdnd11an1n64x5 FILLER_48_1168 ();
 b15zdnd11an1n16x5 FILLER_48_1232 ();
 b15zdnd11an1n04x5 FILLER_48_1248 ();
 b15zdnd00an1n02x5 FILLER_48_1252 ();
 b15zdnd11an1n04x5 FILLER_48_1261 ();
 b15zdnd11an1n64x5 FILLER_48_1283 ();
 b15zdnd11an1n64x5 FILLER_48_1347 ();
 b15zdnd11an1n64x5 FILLER_48_1411 ();
 b15zdnd11an1n64x5 FILLER_48_1475 ();
 b15zdnd11an1n64x5 FILLER_48_1539 ();
 b15zdnd11an1n64x5 FILLER_48_1603 ();
 b15zdnd11an1n64x5 FILLER_48_1667 ();
 b15zdnd11an1n64x5 FILLER_48_1731 ();
 b15zdnd11an1n64x5 FILLER_48_1795 ();
 b15zdnd11an1n64x5 FILLER_48_1859 ();
 b15zdnd11an1n64x5 FILLER_48_1923 ();
 b15zdnd11an1n64x5 FILLER_48_1987 ();
 b15zdnd11an1n64x5 FILLER_48_2051 ();
 b15zdnd11an1n32x5 FILLER_48_2115 ();
 b15zdnd11an1n04x5 FILLER_48_2147 ();
 b15zdnd00an1n02x5 FILLER_48_2151 ();
 b15zdnd00an1n01x5 FILLER_48_2153 ();
 b15zdnd11an1n64x5 FILLER_48_2162 ();
 b15zdnd11an1n32x5 FILLER_48_2226 ();
 b15zdnd11an1n16x5 FILLER_48_2258 ();
 b15zdnd00an1n02x5 FILLER_48_2274 ();
 b15zdnd11an1n64x5 FILLER_49_0 ();
 b15zdnd11an1n64x5 FILLER_49_64 ();
 b15zdnd11an1n64x5 FILLER_49_128 ();
 b15zdnd11an1n64x5 FILLER_49_192 ();
 b15zdnd11an1n64x5 FILLER_49_256 ();
 b15zdnd11an1n64x5 FILLER_49_320 ();
 b15zdnd11an1n64x5 FILLER_49_384 ();
 b15zdnd11an1n64x5 FILLER_49_448 ();
 b15zdnd11an1n64x5 FILLER_49_512 ();
 b15zdnd11an1n64x5 FILLER_49_576 ();
 b15zdnd11an1n64x5 FILLER_49_640 ();
 b15zdnd11an1n64x5 FILLER_49_704 ();
 b15zdnd11an1n64x5 FILLER_49_768 ();
 b15zdnd11an1n64x5 FILLER_49_832 ();
 b15zdnd11an1n64x5 FILLER_49_896 ();
 b15zdnd11an1n32x5 FILLER_49_960 ();
 b15zdnd11an1n16x5 FILLER_49_992 ();
 b15zdnd11an1n08x5 FILLER_49_1008 ();
 b15zdnd00an1n02x5 FILLER_49_1016 ();
 b15zdnd00an1n01x5 FILLER_49_1018 ();
 b15zdnd11an1n08x5 FILLER_49_1061 ();
 b15zdnd11an1n04x5 FILLER_49_1069 ();
 b15zdnd11an1n08x5 FILLER_49_1115 ();
 b15zdnd11an1n04x5 FILLER_49_1123 ();
 b15zdnd00an1n02x5 FILLER_49_1127 ();
 b15zdnd00an1n01x5 FILLER_49_1129 ();
 b15zdnd11an1n04x5 FILLER_49_1172 ();
 b15zdnd00an1n02x5 FILLER_49_1176 ();
 b15zdnd00an1n01x5 FILLER_49_1178 ();
 b15zdnd11an1n32x5 FILLER_49_1221 ();
 b15zdnd11an1n08x5 FILLER_49_1253 ();
 b15zdnd11an1n04x5 FILLER_49_1261 ();
 b15zdnd00an1n01x5 FILLER_49_1265 ();
 b15zdnd11an1n64x5 FILLER_49_1279 ();
 b15zdnd11an1n64x5 FILLER_49_1343 ();
 b15zdnd11an1n64x5 FILLER_49_1407 ();
 b15zdnd11an1n32x5 FILLER_49_1471 ();
 b15zdnd11an1n08x5 FILLER_49_1503 ();
 b15zdnd11an1n04x5 FILLER_49_1511 ();
 b15zdnd00an1n01x5 FILLER_49_1515 ();
 b15zdnd11an1n64x5 FILLER_49_1525 ();
 b15zdnd11an1n64x5 FILLER_49_1589 ();
 b15zdnd11an1n64x5 FILLER_49_1653 ();
 b15zdnd11an1n64x5 FILLER_49_1717 ();
 b15zdnd11an1n64x5 FILLER_49_1781 ();
 b15zdnd11an1n64x5 FILLER_49_1845 ();
 b15zdnd11an1n64x5 FILLER_49_1909 ();
 b15zdnd11an1n64x5 FILLER_49_1973 ();
 b15zdnd11an1n64x5 FILLER_49_2037 ();
 b15zdnd11an1n64x5 FILLER_49_2101 ();
 b15zdnd11an1n64x5 FILLER_49_2165 ();
 b15zdnd11an1n32x5 FILLER_49_2229 ();
 b15zdnd11an1n16x5 FILLER_49_2261 ();
 b15zdnd11an1n04x5 FILLER_49_2277 ();
 b15zdnd00an1n02x5 FILLER_49_2281 ();
 b15zdnd00an1n01x5 FILLER_49_2283 ();
 b15zdnd11an1n64x5 FILLER_50_8 ();
 b15zdnd11an1n64x5 FILLER_50_72 ();
 b15zdnd11an1n64x5 FILLER_50_136 ();
 b15zdnd11an1n64x5 FILLER_50_200 ();
 b15zdnd11an1n32x5 FILLER_50_264 ();
 b15zdnd11an1n16x5 FILLER_50_296 ();
 b15zdnd11an1n04x5 FILLER_50_312 ();
 b15zdnd00an1n01x5 FILLER_50_316 ();
 b15zdnd11an1n04x5 FILLER_50_320 ();
 b15zdnd11an1n64x5 FILLER_50_327 ();
 b15zdnd11an1n64x5 FILLER_50_391 ();
 b15zdnd11an1n64x5 FILLER_50_455 ();
 b15zdnd11an1n64x5 FILLER_50_519 ();
 b15zdnd11an1n64x5 FILLER_50_583 ();
 b15zdnd11an1n64x5 FILLER_50_647 ();
 b15zdnd11an1n04x5 FILLER_50_711 ();
 b15zdnd00an1n02x5 FILLER_50_715 ();
 b15zdnd00an1n01x5 FILLER_50_717 ();
 b15zdnd11an1n64x5 FILLER_50_726 ();
 b15zdnd11an1n64x5 FILLER_50_790 ();
 b15zdnd11an1n64x5 FILLER_50_854 ();
 b15zdnd11an1n64x5 FILLER_50_918 ();
 b15zdnd11an1n64x5 FILLER_50_982 ();
 b15zdnd11an1n64x5 FILLER_50_1046 ();
 b15zdnd11an1n64x5 FILLER_50_1110 ();
 b15zdnd11an1n64x5 FILLER_50_1174 ();
 b15zdnd00an1n02x5 FILLER_50_1238 ();
 b15zdnd00an1n01x5 FILLER_50_1240 ();
 b15zdnd11an1n64x5 FILLER_50_1250 ();
 b15zdnd11an1n64x5 FILLER_50_1314 ();
 b15zdnd11an1n64x5 FILLER_50_1378 ();
 b15zdnd11an1n64x5 FILLER_50_1442 ();
 b15zdnd11an1n64x5 FILLER_50_1506 ();
 b15zdnd11an1n64x5 FILLER_50_1570 ();
 b15zdnd11an1n64x5 FILLER_50_1634 ();
 b15zdnd11an1n64x5 FILLER_50_1698 ();
 b15zdnd11an1n64x5 FILLER_50_1762 ();
 b15zdnd11an1n64x5 FILLER_50_1826 ();
 b15zdnd11an1n04x5 FILLER_50_1890 ();
 b15zdnd11an1n04x5 FILLER_50_1897 ();
 b15zdnd11an1n16x5 FILLER_50_1904 ();
 b15zdnd11an1n32x5 FILLER_50_1972 ();
 b15zdnd11an1n16x5 FILLER_50_2004 ();
 b15zdnd11an1n04x5 FILLER_50_2020 ();
 b15zdnd11an1n64x5 FILLER_50_2027 ();
 b15zdnd11an1n32x5 FILLER_50_2091 ();
 b15zdnd11an1n16x5 FILLER_50_2123 ();
 b15zdnd11an1n08x5 FILLER_50_2139 ();
 b15zdnd11an1n04x5 FILLER_50_2147 ();
 b15zdnd00an1n02x5 FILLER_50_2151 ();
 b15zdnd00an1n01x5 FILLER_50_2153 ();
 b15zdnd11an1n64x5 FILLER_50_2162 ();
 b15zdnd11an1n04x5 FILLER_50_2226 ();
 b15zdnd00an1n02x5 FILLER_50_2230 ();
 b15zdnd00an1n02x5 FILLER_50_2274 ();
 b15zdnd11an1n64x5 FILLER_51_0 ();
 b15zdnd11an1n64x5 FILLER_51_64 ();
 b15zdnd11an1n64x5 FILLER_51_128 ();
 b15zdnd11an1n16x5 FILLER_51_192 ();
 b15zdnd11an1n08x5 FILLER_51_208 ();
 b15zdnd11an1n04x5 FILLER_51_216 ();
 b15zdnd00an1n02x5 FILLER_51_220 ();
 b15zdnd11an1n64x5 FILLER_51_225 ();
 b15zdnd11an1n08x5 FILLER_51_289 ();
 b15zdnd00an1n02x5 FILLER_51_297 ();
 b15zdnd11an1n64x5 FILLER_51_351 ();
 b15zdnd11an1n64x5 FILLER_51_415 ();
 b15zdnd11an1n64x5 FILLER_51_479 ();
 b15zdnd11an1n64x5 FILLER_51_543 ();
 b15zdnd11an1n64x5 FILLER_51_607 ();
 b15zdnd11an1n32x5 FILLER_51_671 ();
 b15zdnd11an1n08x5 FILLER_51_703 ();
 b15zdnd11an1n04x5 FILLER_51_711 ();
 b15zdnd00an1n02x5 FILLER_51_715 ();
 b15zdnd00an1n01x5 FILLER_51_717 ();
 b15zdnd11an1n64x5 FILLER_51_770 ();
 b15zdnd11an1n64x5 FILLER_51_834 ();
 b15zdnd11an1n64x5 FILLER_51_898 ();
 b15zdnd11an1n64x5 FILLER_51_962 ();
 b15zdnd11an1n04x5 FILLER_51_1026 ();
 b15zdnd00an1n01x5 FILLER_51_1030 ();
 b15zdnd11an1n64x5 FILLER_51_1034 ();
 b15zdnd11an1n64x5 FILLER_51_1098 ();
 b15zdnd11an1n64x5 FILLER_51_1162 ();
 b15zdnd11an1n64x5 FILLER_51_1226 ();
 b15zdnd11an1n64x5 FILLER_51_1290 ();
 b15zdnd11an1n16x5 FILLER_51_1354 ();
 b15zdnd11an1n08x5 FILLER_51_1370 ();
 b15zdnd00an1n01x5 FILLER_51_1378 ();
 b15zdnd11an1n64x5 FILLER_51_1421 ();
 b15zdnd11an1n64x5 FILLER_51_1485 ();
 b15zdnd11an1n64x5 FILLER_51_1549 ();
 b15zdnd11an1n64x5 FILLER_51_1613 ();
 b15zdnd11an1n64x5 FILLER_51_1677 ();
 b15zdnd11an1n64x5 FILLER_51_1741 ();
 b15zdnd11an1n64x5 FILLER_51_1805 ();
 b15zdnd11an1n04x5 FILLER_51_1869 ();
 b15zdnd00an1n02x5 FILLER_51_1873 ();
 b15zdnd00an1n01x5 FILLER_51_1875 ();
 b15zdnd11an1n08x5 FILLER_51_1928 ();
 b15zdnd00an1n02x5 FILLER_51_1936 ();
 b15zdnd11an1n04x5 FILLER_51_1941 ();
 b15zdnd11an1n64x5 FILLER_51_1948 ();
 b15zdnd11an1n08x5 FILLER_51_2012 ();
 b15zdnd00an1n02x5 FILLER_51_2020 ();
 b15zdnd00an1n01x5 FILLER_51_2022 ();
 b15zdnd11an1n04x5 FILLER_51_2026 ();
 b15zdnd00an1n02x5 FILLER_51_2030 ();
 b15zdnd11an1n64x5 FILLER_51_2035 ();
 b15zdnd11an1n64x5 FILLER_51_2099 ();
 b15zdnd11an1n64x5 FILLER_51_2163 ();
 b15zdnd11an1n04x5 FILLER_51_2227 ();
 b15zdnd00an1n02x5 FILLER_51_2231 ();
 b15zdnd11an1n08x5 FILLER_51_2275 ();
 b15zdnd00an1n01x5 FILLER_51_2283 ();
 b15zdnd11an1n08x5 FILLER_52_8 ();
 b15zdnd11an1n04x5 FILLER_52_16 ();
 b15zdnd00an1n02x5 FILLER_52_20 ();
 b15zdnd00an1n01x5 FILLER_52_22 ();
 b15zdnd11an1n64x5 FILLER_52_26 ();
 b15zdnd11an1n64x5 FILLER_52_90 ();
 b15zdnd11an1n32x5 FILLER_52_154 ();
 b15zdnd11an1n08x5 FILLER_52_186 ();
 b15zdnd11an1n04x5 FILLER_52_194 ();
 b15zdnd11an1n64x5 FILLER_52_250 ();
 b15zdnd11an1n08x5 FILLER_52_314 ();
 b15zdnd11an1n64x5 FILLER_52_325 ();
 b15zdnd11an1n64x5 FILLER_52_389 ();
 b15zdnd11an1n16x5 FILLER_52_453 ();
 b15zdnd11an1n08x5 FILLER_52_469 ();
 b15zdnd11an1n04x5 FILLER_52_477 ();
 b15zdnd11an1n04x5 FILLER_52_495 ();
 b15zdnd11an1n64x5 FILLER_52_519 ();
 b15zdnd11an1n64x5 FILLER_52_583 ();
 b15zdnd11an1n64x5 FILLER_52_647 ();
 b15zdnd11an1n04x5 FILLER_52_711 ();
 b15zdnd00an1n02x5 FILLER_52_715 ();
 b15zdnd00an1n01x5 FILLER_52_717 ();
 b15zdnd11an1n08x5 FILLER_52_726 ();
 b15zdnd11an1n04x5 FILLER_52_734 ();
 b15zdnd00an1n02x5 FILLER_52_738 ();
 b15zdnd11an1n04x5 FILLER_52_743 ();
 b15zdnd11an1n04x5 FILLER_52_750 ();
 b15zdnd11an1n64x5 FILLER_52_757 ();
 b15zdnd11an1n64x5 FILLER_52_821 ();
 b15zdnd11an1n64x5 FILLER_52_885 ();
 b15zdnd11an1n32x5 FILLER_52_949 ();
 b15zdnd00an1n01x5 FILLER_52_981 ();
 b15zdnd11an1n64x5 FILLER_52_1034 ();
 b15zdnd11an1n64x5 FILLER_52_1098 ();
 b15zdnd11an1n64x5 FILLER_52_1162 ();
 b15zdnd11an1n32x5 FILLER_52_1226 ();
 b15zdnd11an1n16x5 FILLER_52_1258 ();
 b15zdnd11an1n04x5 FILLER_52_1274 ();
 b15zdnd11an1n64x5 FILLER_52_1284 ();
 b15zdnd11an1n64x5 FILLER_52_1348 ();
 b15zdnd11an1n64x5 FILLER_52_1412 ();
 b15zdnd11an1n64x5 FILLER_52_1476 ();
 b15zdnd11an1n64x5 FILLER_52_1540 ();
 b15zdnd11an1n64x5 FILLER_52_1604 ();
 b15zdnd11an1n64x5 FILLER_52_1668 ();
 b15zdnd11an1n32x5 FILLER_52_1732 ();
 b15zdnd11an1n04x5 FILLER_52_1764 ();
 b15zdnd00an1n01x5 FILLER_52_1768 ();
 b15zdnd11an1n04x5 FILLER_52_1772 ();
 b15zdnd00an1n01x5 FILLER_52_1776 ();
 b15zdnd11an1n64x5 FILLER_52_1780 ();
 b15zdnd11an1n32x5 FILLER_52_1844 ();
 b15zdnd11an1n16x5 FILLER_52_1876 ();
 b15zdnd11an1n08x5 FILLER_52_1892 ();
 b15zdnd00an1n01x5 FILLER_52_1900 ();
 b15zdnd11an1n32x5 FILLER_52_1904 ();
 b15zdnd11an1n08x5 FILLER_52_1936 ();
 b15zdnd00an1n01x5 FILLER_52_1944 ();
 b15zdnd11an1n32x5 FILLER_52_1948 ();
 b15zdnd11an1n16x5 FILLER_52_1980 ();
 b15zdnd00an1n02x5 FILLER_52_1996 ();
 b15zdnd00an1n01x5 FILLER_52_1998 ();
 b15zdnd11an1n64x5 FILLER_52_2051 ();
 b15zdnd11an1n32x5 FILLER_52_2115 ();
 b15zdnd11an1n04x5 FILLER_52_2147 ();
 b15zdnd00an1n02x5 FILLER_52_2151 ();
 b15zdnd00an1n01x5 FILLER_52_2153 ();
 b15zdnd11an1n64x5 FILLER_52_2162 ();
 b15zdnd11an1n32x5 FILLER_52_2226 ();
 b15zdnd11an1n16x5 FILLER_52_2258 ();
 b15zdnd00an1n02x5 FILLER_52_2274 ();
 b15zdnd11an1n16x5 FILLER_53_0 ();
 b15zdnd11an1n04x5 FILLER_53_16 ();
 b15zdnd00an1n02x5 FILLER_53_20 ();
 b15zdnd00an1n01x5 FILLER_53_22 ();
 b15zdnd11an1n64x5 FILLER_53_26 ();
 b15zdnd11an1n64x5 FILLER_53_90 ();
 b15zdnd11an1n32x5 FILLER_53_154 ();
 b15zdnd11an1n16x5 FILLER_53_186 ();
 b15zdnd11an1n08x5 FILLER_53_202 ();
 b15zdnd11an1n04x5 FILLER_53_210 ();
 b15zdnd00an1n02x5 FILLER_53_214 ();
 b15zdnd11an1n04x5 FILLER_53_219 ();
 b15zdnd11an1n64x5 FILLER_53_226 ();
 b15zdnd11an1n64x5 FILLER_53_290 ();
 b15zdnd11an1n64x5 FILLER_53_354 ();
 b15zdnd11an1n64x5 FILLER_53_418 ();
 b15zdnd11an1n64x5 FILLER_53_482 ();
 b15zdnd11an1n64x5 FILLER_53_546 ();
 b15zdnd11an1n08x5 FILLER_53_610 ();
 b15zdnd00an1n01x5 FILLER_53_618 ();
 b15zdnd11an1n64x5 FILLER_53_622 ();
 b15zdnd11an1n32x5 FILLER_53_686 ();
 b15zdnd00an1n02x5 FILLER_53_718 ();
 b15zdnd11an1n64x5 FILLER_53_772 ();
 b15zdnd11an1n64x5 FILLER_53_836 ();
 b15zdnd11an1n16x5 FILLER_53_900 ();
 b15zdnd11an1n08x5 FILLER_53_916 ();
 b15zdnd11an1n04x5 FILLER_53_924 ();
 b15zdnd00an1n01x5 FILLER_53_928 ();
 b15zdnd11an1n64x5 FILLER_53_932 ();
 b15zdnd11an1n64x5 FILLER_53_996 ();
 b15zdnd11an1n64x5 FILLER_53_1060 ();
 b15zdnd11an1n64x5 FILLER_53_1124 ();
 b15zdnd11an1n64x5 FILLER_53_1188 ();
 b15zdnd11an1n64x5 FILLER_53_1252 ();
 b15zdnd11an1n64x5 FILLER_53_1316 ();
 b15zdnd11an1n64x5 FILLER_53_1380 ();
 b15zdnd11an1n64x5 FILLER_53_1444 ();
 b15zdnd11an1n64x5 FILLER_53_1508 ();
 b15zdnd11an1n64x5 FILLER_53_1572 ();
 b15zdnd11an1n64x5 FILLER_53_1636 ();
 b15zdnd11an1n32x5 FILLER_53_1700 ();
 b15zdnd11an1n04x5 FILLER_53_1732 ();
 b15zdnd11an1n04x5 FILLER_53_1778 ();
 b15zdnd11an1n04x5 FILLER_53_1785 ();
 b15zdnd11an1n64x5 FILLER_53_1792 ();
 b15zdnd11an1n64x5 FILLER_53_1856 ();
 b15zdnd11an1n64x5 FILLER_53_1920 ();
 b15zdnd11an1n64x5 FILLER_53_1984 ();
 b15zdnd11an1n64x5 FILLER_53_2048 ();
 b15zdnd11an1n64x5 FILLER_53_2112 ();
 b15zdnd11an1n64x5 FILLER_53_2176 ();
 b15zdnd11an1n32x5 FILLER_53_2240 ();
 b15zdnd11an1n08x5 FILLER_53_2272 ();
 b15zdnd11an1n04x5 FILLER_53_2280 ();
 b15zdnd11an1n64x5 FILLER_54_8 ();
 b15zdnd11an1n64x5 FILLER_54_72 ();
 b15zdnd11an1n64x5 FILLER_54_136 ();
 b15zdnd11an1n32x5 FILLER_54_200 ();
 b15zdnd00an1n02x5 FILLER_54_232 ();
 b15zdnd11an1n64x5 FILLER_54_261 ();
 b15zdnd11an1n64x5 FILLER_54_325 ();
 b15zdnd11an1n32x5 FILLER_54_389 ();
 b15zdnd11an1n08x5 FILLER_54_421 ();
 b15zdnd11an1n04x5 FILLER_54_429 ();
 b15zdnd00an1n01x5 FILLER_54_433 ();
 b15zdnd11an1n32x5 FILLER_54_454 ();
 b15zdnd11an1n16x5 FILLER_54_486 ();
 b15zdnd00an1n01x5 FILLER_54_502 ();
 b15zdnd11an1n04x5 FILLER_54_517 ();
 b15zdnd11an1n32x5 FILLER_54_533 ();
 b15zdnd11an1n16x5 FILLER_54_565 ();
 b15zdnd11an1n08x5 FILLER_54_581 ();
 b15zdnd11an1n04x5 FILLER_54_589 ();
 b15zdnd00an1n01x5 FILLER_54_593 ();
 b15zdnd11an1n64x5 FILLER_54_646 ();
 b15zdnd11an1n08x5 FILLER_54_710 ();
 b15zdnd11an1n08x5 FILLER_54_726 ();
 b15zdnd11an1n04x5 FILLER_54_734 ();
 b15zdnd11an1n04x5 FILLER_54_741 ();
 b15zdnd11an1n32x5 FILLER_54_748 ();
 b15zdnd11an1n16x5 FILLER_54_780 ();
 b15zdnd11an1n08x5 FILLER_54_796 ();
 b15zdnd11an1n04x5 FILLER_54_804 ();
 b15zdnd00an1n02x5 FILLER_54_808 ();
 b15zdnd11an1n64x5 FILLER_54_827 ();
 b15zdnd11an1n08x5 FILLER_54_891 ();
 b15zdnd00an1n02x5 FILLER_54_899 ();
 b15zdnd00an1n01x5 FILLER_54_901 ();
 b15zdnd11an1n32x5 FILLER_54_954 ();
 b15zdnd11an1n16x5 FILLER_54_986 ();
 b15zdnd00an1n01x5 FILLER_54_1002 ();
 b15zdnd11an1n32x5 FILLER_54_1006 ();
 b15zdnd00an1n01x5 FILLER_54_1038 ();
 b15zdnd11an1n64x5 FILLER_54_1042 ();
 b15zdnd11an1n64x5 FILLER_54_1106 ();
 b15zdnd11an1n64x5 FILLER_54_1170 ();
 b15zdnd00an1n01x5 FILLER_54_1234 ();
 b15zdnd11an1n04x5 FILLER_54_1255 ();
 b15zdnd11an1n64x5 FILLER_54_1263 ();
 b15zdnd11an1n64x5 FILLER_54_1327 ();
 b15zdnd11an1n64x5 FILLER_54_1391 ();
 b15zdnd11an1n64x5 FILLER_54_1455 ();
 b15zdnd11an1n64x5 FILLER_54_1519 ();
 b15zdnd11an1n64x5 FILLER_54_1583 ();
 b15zdnd11an1n64x5 FILLER_54_1647 ();
 b15zdnd11an1n32x5 FILLER_54_1711 ();
 b15zdnd11an1n08x5 FILLER_54_1743 ();
 b15zdnd00an1n01x5 FILLER_54_1751 ();
 b15zdnd11an1n64x5 FILLER_54_1804 ();
 b15zdnd11an1n64x5 FILLER_54_1868 ();
 b15zdnd11an1n64x5 FILLER_54_1932 ();
 b15zdnd11an1n64x5 FILLER_54_1996 ();
 b15zdnd11an1n64x5 FILLER_54_2060 ();
 b15zdnd11an1n16x5 FILLER_54_2124 ();
 b15zdnd11an1n08x5 FILLER_54_2140 ();
 b15zdnd11an1n04x5 FILLER_54_2148 ();
 b15zdnd00an1n02x5 FILLER_54_2152 ();
 b15zdnd11an1n64x5 FILLER_54_2162 ();
 b15zdnd11an1n32x5 FILLER_54_2226 ();
 b15zdnd11an1n16x5 FILLER_54_2258 ();
 b15zdnd00an1n02x5 FILLER_54_2274 ();
 b15zdnd11an1n64x5 FILLER_55_0 ();
 b15zdnd11an1n64x5 FILLER_55_64 ();
 b15zdnd11an1n64x5 FILLER_55_128 ();
 b15zdnd11an1n32x5 FILLER_55_192 ();
 b15zdnd11an1n08x5 FILLER_55_224 ();
 b15zdnd00an1n02x5 FILLER_55_232 ();
 b15zdnd11an1n64x5 FILLER_55_237 ();
 b15zdnd11an1n64x5 FILLER_55_301 ();
 b15zdnd11an1n64x5 FILLER_55_365 ();
 b15zdnd11an1n64x5 FILLER_55_429 ();
 b15zdnd11an1n08x5 FILLER_55_493 ();
 b15zdnd11an1n04x5 FILLER_55_501 ();
 b15zdnd00an1n02x5 FILLER_55_505 ();
 b15zdnd11an1n64x5 FILLER_55_527 ();
 b15zdnd11an1n08x5 FILLER_55_591 ();
 b15zdnd11an1n04x5 FILLER_55_599 ();
 b15zdnd00an1n02x5 FILLER_55_603 ();
 b15zdnd00an1n01x5 FILLER_55_605 ();
 b15zdnd11an1n64x5 FILLER_55_658 ();
 b15zdnd11an1n16x5 FILLER_55_722 ();
 b15zdnd11an1n04x5 FILLER_55_738 ();
 b15zdnd00an1n02x5 FILLER_55_742 ();
 b15zdnd11an1n64x5 FILLER_55_747 ();
 b15zdnd11an1n64x5 FILLER_55_811 ();
 b15zdnd11an1n32x5 FILLER_55_875 ();
 b15zdnd11an1n08x5 FILLER_55_907 ();
 b15zdnd11an1n04x5 FILLER_55_915 ();
 b15zdnd00an1n01x5 FILLER_55_919 ();
 b15zdnd11an1n04x5 FILLER_55_923 ();
 b15zdnd11an1n32x5 FILLER_55_930 ();
 b15zdnd11an1n16x5 FILLER_55_962 ();
 b15zdnd11an1n08x5 FILLER_55_978 ();
 b15zdnd00an1n02x5 FILLER_55_986 ();
 b15zdnd11an1n04x5 FILLER_55_1040 ();
 b15zdnd00an1n02x5 FILLER_55_1044 ();
 b15zdnd11an1n64x5 FILLER_55_1049 ();
 b15zdnd11an1n32x5 FILLER_55_1113 ();
 b15zdnd11an1n08x5 FILLER_55_1145 ();
 b15zdnd11an1n04x5 FILLER_55_1156 ();
 b15zdnd11an1n04x5 FILLER_55_1163 ();
 b15zdnd11an1n64x5 FILLER_55_1170 ();
 b15zdnd11an1n04x5 FILLER_55_1234 ();
 b15zdnd00an1n02x5 FILLER_55_1238 ();
 b15zdnd11an1n08x5 FILLER_55_1250 ();
 b15zdnd00an1n02x5 FILLER_55_1258 ();
 b15zdnd00an1n01x5 FILLER_55_1260 ();
 b15zdnd11an1n16x5 FILLER_55_1303 ();
 b15zdnd11an1n04x5 FILLER_55_1319 ();
 b15zdnd00an1n01x5 FILLER_55_1323 ();
 b15zdnd11an1n64x5 FILLER_55_1366 ();
 b15zdnd11an1n64x5 FILLER_55_1430 ();
 b15zdnd11an1n64x5 FILLER_55_1494 ();
 b15zdnd11an1n64x5 FILLER_55_1558 ();
 b15zdnd11an1n32x5 FILLER_55_1622 ();
 b15zdnd11an1n16x5 FILLER_55_1654 ();
 b15zdnd11an1n04x5 FILLER_55_1670 ();
 b15zdnd11an1n04x5 FILLER_55_1677 ();
 b15zdnd11an1n64x5 FILLER_55_1684 ();
 b15zdnd00an1n02x5 FILLER_55_1748 ();
 b15zdnd11an1n64x5 FILLER_55_1802 ();
 b15zdnd11an1n64x5 FILLER_55_1866 ();
 b15zdnd11an1n64x5 FILLER_55_1930 ();
 b15zdnd11an1n64x5 FILLER_55_1994 ();
 b15zdnd11an1n64x5 FILLER_55_2058 ();
 b15zdnd11an1n64x5 FILLER_55_2122 ();
 b15zdnd11an1n64x5 FILLER_55_2186 ();
 b15zdnd11an1n32x5 FILLER_55_2250 ();
 b15zdnd00an1n02x5 FILLER_55_2282 ();
 b15zdnd11an1n64x5 FILLER_56_8 ();
 b15zdnd11an1n64x5 FILLER_56_72 ();
 b15zdnd11an1n64x5 FILLER_56_136 ();
 b15zdnd11an1n64x5 FILLER_56_200 ();
 b15zdnd11an1n64x5 FILLER_56_264 ();
 b15zdnd11an1n64x5 FILLER_56_328 ();
 b15zdnd11an1n64x5 FILLER_56_392 ();
 b15zdnd11an1n32x5 FILLER_56_456 ();
 b15zdnd11an1n16x5 FILLER_56_488 ();
 b15zdnd11an1n08x5 FILLER_56_504 ();
 b15zdnd11an1n04x5 FILLER_56_512 ();
 b15zdnd00an1n02x5 FILLER_56_516 ();
 b15zdnd11an1n04x5 FILLER_56_538 ();
 b15zdnd11an1n32x5 FILLER_56_556 ();
 b15zdnd11an1n16x5 FILLER_56_588 ();
 b15zdnd11an1n08x5 FILLER_56_604 ();
 b15zdnd11an1n04x5 FILLER_56_615 ();
 b15zdnd11an1n04x5 FILLER_56_622 ();
 b15zdnd11an1n04x5 FILLER_56_629 ();
 b15zdnd11an1n64x5 FILLER_56_636 ();
 b15zdnd11an1n16x5 FILLER_56_700 ();
 b15zdnd00an1n02x5 FILLER_56_716 ();
 b15zdnd11an1n64x5 FILLER_56_726 ();
 b15zdnd11an1n64x5 FILLER_56_790 ();
 b15zdnd11an1n64x5 FILLER_56_854 ();
 b15zdnd11an1n64x5 FILLER_56_918 ();
 b15zdnd11an1n16x5 FILLER_56_982 ();
 b15zdnd11an1n08x5 FILLER_56_998 ();
 b15zdnd00an1n02x5 FILLER_56_1006 ();
 b15zdnd11an1n08x5 FILLER_56_1011 ();
 b15zdnd00an1n02x5 FILLER_56_1019 ();
 b15zdnd00an1n01x5 FILLER_56_1021 ();
 b15zdnd11an1n16x5 FILLER_56_1025 ();
 b15zdnd11an1n04x5 FILLER_56_1041 ();
 b15zdnd00an1n01x5 FILLER_56_1045 ();
 b15zdnd11an1n64x5 FILLER_56_1049 ();
 b15zdnd11an1n16x5 FILLER_56_1113 ();
 b15zdnd11an1n04x5 FILLER_56_1129 ();
 b15zdnd00an1n02x5 FILLER_56_1133 ();
 b15zdnd11an1n64x5 FILLER_56_1187 ();
 b15zdnd00an1n02x5 FILLER_56_1251 ();
 b15zdnd00an1n01x5 FILLER_56_1253 ();
 b15zdnd11an1n16x5 FILLER_56_1268 ();
 b15zdnd11an1n08x5 FILLER_56_1284 ();
 b15zdnd11an1n04x5 FILLER_56_1324 ();
 b15zdnd11an1n64x5 FILLER_56_1331 ();
 b15zdnd11an1n04x5 FILLER_56_1395 ();
 b15zdnd11an1n32x5 FILLER_56_1402 ();
 b15zdnd11an1n16x5 FILLER_56_1434 ();
 b15zdnd11an1n08x5 FILLER_56_1450 ();
 b15zdnd11an1n04x5 FILLER_56_1458 ();
 b15zdnd00an1n01x5 FILLER_56_1462 ();
 b15zdnd11an1n04x5 FILLER_56_1466 ();
 b15zdnd11an1n04x5 FILLER_56_1473 ();
 b15zdnd11an1n64x5 FILLER_56_1480 ();
 b15zdnd11an1n64x5 FILLER_56_1544 ();
 b15zdnd11an1n32x5 FILLER_56_1608 ();
 b15zdnd11an1n16x5 FILLER_56_1640 ();
 b15zdnd11an1n08x5 FILLER_56_1656 ();
 b15zdnd00an1n02x5 FILLER_56_1664 ();
 b15zdnd00an1n01x5 FILLER_56_1666 ();
 b15zdnd11an1n08x5 FILLER_56_1670 ();
 b15zdnd00an1n01x5 FILLER_56_1678 ();
 b15zdnd11an1n32x5 FILLER_56_1721 ();
 b15zdnd11an1n08x5 FILLER_56_1753 ();
 b15zdnd00an1n02x5 FILLER_56_1761 ();
 b15zdnd00an1n01x5 FILLER_56_1763 ();
 b15zdnd11an1n64x5 FILLER_56_1816 ();
 b15zdnd11an1n64x5 FILLER_56_1880 ();
 b15zdnd11an1n64x5 FILLER_56_1944 ();
 b15zdnd11an1n64x5 FILLER_56_2008 ();
 b15zdnd11an1n64x5 FILLER_56_2072 ();
 b15zdnd11an1n16x5 FILLER_56_2136 ();
 b15zdnd00an1n02x5 FILLER_56_2152 ();
 b15zdnd11an1n64x5 FILLER_56_2162 ();
 b15zdnd11an1n32x5 FILLER_56_2226 ();
 b15zdnd11an1n16x5 FILLER_56_2258 ();
 b15zdnd00an1n02x5 FILLER_56_2274 ();
 b15zdnd11an1n64x5 FILLER_57_0 ();
 b15zdnd11an1n64x5 FILLER_57_64 ();
 b15zdnd11an1n64x5 FILLER_57_128 ();
 b15zdnd11an1n64x5 FILLER_57_192 ();
 b15zdnd11an1n64x5 FILLER_57_256 ();
 b15zdnd11an1n64x5 FILLER_57_320 ();
 b15zdnd11an1n64x5 FILLER_57_384 ();
 b15zdnd11an1n64x5 FILLER_57_448 ();
 b15zdnd11an1n64x5 FILLER_57_512 ();
 b15zdnd11an1n32x5 FILLER_57_576 ();
 b15zdnd11an1n16x5 FILLER_57_608 ();
 b15zdnd11an1n08x5 FILLER_57_624 ();
 b15zdnd11an1n64x5 FILLER_57_635 ();
 b15zdnd11an1n64x5 FILLER_57_699 ();
 b15zdnd11an1n64x5 FILLER_57_763 ();
 b15zdnd11an1n64x5 FILLER_57_827 ();
 b15zdnd11an1n04x5 FILLER_57_891 ();
 b15zdnd11an1n64x5 FILLER_57_926 ();
 b15zdnd11an1n08x5 FILLER_57_990 ();
 b15zdnd11an1n04x5 FILLER_57_998 ();
 b15zdnd00an1n02x5 FILLER_57_1002 ();
 b15zdnd11an1n04x5 FILLER_57_1046 ();
 b15zdnd11an1n64x5 FILLER_57_1092 ();
 b15zdnd11an1n16x5 FILLER_57_1156 ();
 b15zdnd00an1n02x5 FILLER_57_1172 ();
 b15zdnd11an1n64x5 FILLER_57_1184 ();
 b15zdnd00an1n02x5 FILLER_57_1248 ();
 b15zdnd11an1n32x5 FILLER_57_1260 ();
 b15zdnd11an1n16x5 FILLER_57_1292 ();
 b15zdnd11an1n08x5 FILLER_57_1308 ();
 b15zdnd11an1n32x5 FILLER_57_1319 ();
 b15zdnd11an1n16x5 FILLER_57_1351 ();
 b15zdnd11an1n04x5 FILLER_57_1367 ();
 b15zdnd00an1n02x5 FILLER_57_1371 ();
 b15zdnd11an1n16x5 FILLER_57_1425 ();
 b15zdnd11an1n04x5 FILLER_57_1441 ();
 b15zdnd00an1n01x5 FILLER_57_1445 ();
 b15zdnd11an1n04x5 FILLER_57_1498 ();
 b15zdnd11an1n32x5 FILLER_57_1554 ();
 b15zdnd11an1n16x5 FILLER_57_1586 ();
 b15zdnd11an1n08x5 FILLER_57_1602 ();
 b15zdnd11an1n04x5 FILLER_57_1610 ();
 b15zdnd00an1n02x5 FILLER_57_1614 ();
 b15zdnd00an1n01x5 FILLER_57_1616 ();
 b15zdnd11an1n16x5 FILLER_57_1620 ();
 b15zdnd11an1n08x5 FILLER_57_1636 ();
 b15zdnd11an1n04x5 FILLER_57_1644 ();
 b15zdnd00an1n01x5 FILLER_57_1648 ();
 b15zdnd11an1n64x5 FILLER_57_1701 ();
 b15zdnd11an1n08x5 FILLER_57_1765 ();
 b15zdnd00an1n02x5 FILLER_57_1773 ();
 b15zdnd11an1n04x5 FILLER_57_1778 ();
 b15zdnd11an1n04x5 FILLER_57_1785 ();
 b15zdnd11an1n04x5 FILLER_57_1792 ();
 b15zdnd11an1n64x5 FILLER_57_1799 ();
 b15zdnd11an1n64x5 FILLER_57_1863 ();
 b15zdnd11an1n64x5 FILLER_57_1927 ();
 b15zdnd11an1n64x5 FILLER_57_1991 ();
 b15zdnd11an1n64x5 FILLER_57_2055 ();
 b15zdnd11an1n64x5 FILLER_57_2119 ();
 b15zdnd11an1n64x5 FILLER_57_2183 ();
 b15zdnd11an1n32x5 FILLER_57_2247 ();
 b15zdnd11an1n04x5 FILLER_57_2279 ();
 b15zdnd00an1n01x5 FILLER_57_2283 ();
 b15zdnd11an1n64x5 FILLER_58_8 ();
 b15zdnd11an1n64x5 FILLER_58_72 ();
 b15zdnd11an1n64x5 FILLER_58_136 ();
 b15zdnd11an1n64x5 FILLER_58_200 ();
 b15zdnd11an1n64x5 FILLER_58_264 ();
 b15zdnd11an1n64x5 FILLER_58_328 ();
 b15zdnd11an1n64x5 FILLER_58_392 ();
 b15zdnd11an1n64x5 FILLER_58_456 ();
 b15zdnd11an1n64x5 FILLER_58_520 ();
 b15zdnd11an1n64x5 FILLER_58_584 ();
 b15zdnd11an1n64x5 FILLER_58_648 ();
 b15zdnd11an1n04x5 FILLER_58_712 ();
 b15zdnd00an1n02x5 FILLER_58_716 ();
 b15zdnd11an1n64x5 FILLER_58_726 ();
 b15zdnd11an1n64x5 FILLER_58_790 ();
 b15zdnd11an1n64x5 FILLER_58_854 ();
 b15zdnd11an1n64x5 FILLER_58_918 ();
 b15zdnd11an1n32x5 FILLER_58_982 ();
 b15zdnd11an1n04x5 FILLER_58_1014 ();
 b15zdnd00an1n01x5 FILLER_58_1018 ();
 b15zdnd11an1n64x5 FILLER_58_1071 ();
 b15zdnd11an1n64x5 FILLER_58_1135 ();
 b15zdnd11an1n64x5 FILLER_58_1199 ();
 b15zdnd11an1n64x5 FILLER_58_1263 ();
 b15zdnd11an1n64x5 FILLER_58_1327 ();
 b15zdnd11an1n04x5 FILLER_58_1391 ();
 b15zdnd00an1n02x5 FILLER_58_1395 ();
 b15zdnd00an1n01x5 FILLER_58_1397 ();
 b15zdnd11an1n64x5 FILLER_58_1401 ();
 b15zdnd11an1n32x5 FILLER_58_1465 ();
 b15zdnd11an1n16x5 FILLER_58_1497 ();
 b15zdnd11an1n08x5 FILLER_58_1513 ();
 b15zdnd11an1n04x5 FILLER_58_1524 ();
 b15zdnd11an1n04x5 FILLER_58_1531 ();
 b15zdnd11an1n64x5 FILLER_58_1538 ();
 b15zdnd11an1n04x5 FILLER_58_1602 ();
 b15zdnd00an1n02x5 FILLER_58_1606 ();
 b15zdnd11an1n04x5 FILLER_58_1611 ();
 b15zdnd11an1n64x5 FILLER_58_1618 ();
 b15zdnd11an1n64x5 FILLER_58_1682 ();
 b15zdnd11an1n16x5 FILLER_58_1746 ();
 b15zdnd11an1n08x5 FILLER_58_1762 ();
 b15zdnd11an1n04x5 FILLER_58_1770 ();
 b15zdnd00an1n01x5 FILLER_58_1774 ();
 b15zdnd11an1n64x5 FILLER_58_1778 ();
 b15zdnd11an1n64x5 FILLER_58_1842 ();
 b15zdnd11an1n64x5 FILLER_58_1906 ();
 b15zdnd11an1n64x5 FILLER_58_1970 ();
 b15zdnd11an1n64x5 FILLER_58_2034 ();
 b15zdnd11an1n32x5 FILLER_58_2098 ();
 b15zdnd11an1n16x5 FILLER_58_2130 ();
 b15zdnd11an1n08x5 FILLER_58_2146 ();
 b15zdnd11an1n64x5 FILLER_58_2162 ();
 b15zdnd11an1n32x5 FILLER_58_2226 ();
 b15zdnd11an1n16x5 FILLER_58_2258 ();
 b15zdnd00an1n02x5 FILLER_58_2274 ();
 b15zdnd11an1n64x5 FILLER_59_0 ();
 b15zdnd11an1n64x5 FILLER_59_64 ();
 b15zdnd11an1n64x5 FILLER_59_128 ();
 b15zdnd11an1n64x5 FILLER_59_192 ();
 b15zdnd11an1n08x5 FILLER_59_256 ();
 b15zdnd00an1n02x5 FILLER_59_264 ();
 b15zdnd11an1n16x5 FILLER_59_275 ();
 b15zdnd00an1n02x5 FILLER_59_291 ();
 b15zdnd00an1n01x5 FILLER_59_293 ();
 b15zdnd11an1n64x5 FILLER_59_303 ();
 b15zdnd11an1n64x5 FILLER_59_367 ();
 b15zdnd11an1n32x5 FILLER_59_431 ();
 b15zdnd11an1n16x5 FILLER_59_463 ();
 b15zdnd11an1n08x5 FILLER_59_479 ();
 b15zdnd11an1n04x5 FILLER_59_487 ();
 b15zdnd11an1n64x5 FILLER_59_508 ();
 b15zdnd11an1n64x5 FILLER_59_572 ();
 b15zdnd11an1n64x5 FILLER_59_636 ();
 b15zdnd11an1n64x5 FILLER_59_700 ();
 b15zdnd11an1n64x5 FILLER_59_764 ();
 b15zdnd11an1n64x5 FILLER_59_828 ();
 b15zdnd11an1n64x5 FILLER_59_892 ();
 b15zdnd11an1n04x5 FILLER_59_956 ();
 b15zdnd11an1n64x5 FILLER_59_969 ();
 b15zdnd11an1n04x5 FILLER_59_1033 ();
 b15zdnd00an1n01x5 FILLER_59_1037 ();
 b15zdnd11an1n04x5 FILLER_59_1041 ();
 b15zdnd11an1n64x5 FILLER_59_1048 ();
 b15zdnd11an1n64x5 FILLER_59_1112 ();
 b15zdnd11an1n64x5 FILLER_59_1176 ();
 b15zdnd11an1n64x5 FILLER_59_1240 ();
 b15zdnd11an1n64x5 FILLER_59_1304 ();
 b15zdnd11an1n16x5 FILLER_59_1368 ();
 b15zdnd11an1n08x5 FILLER_59_1384 ();
 b15zdnd11an1n04x5 FILLER_59_1392 ();
 b15zdnd00an1n01x5 FILLER_59_1396 ();
 b15zdnd11an1n64x5 FILLER_59_1400 ();
 b15zdnd11an1n32x5 FILLER_59_1464 ();
 b15zdnd11an1n16x5 FILLER_59_1496 ();
 b15zdnd11an1n08x5 FILLER_59_1512 ();
 b15zdnd00an1n02x5 FILLER_59_1520 ();
 b15zdnd00an1n01x5 FILLER_59_1522 ();
 b15zdnd11an1n16x5 FILLER_59_1575 ();
 b15zdnd00an1n01x5 FILLER_59_1591 ();
 b15zdnd11an1n04x5 FILLER_59_1644 ();
 b15zdnd11an1n64x5 FILLER_59_1668 ();
 b15zdnd11an1n64x5 FILLER_59_1732 ();
 b15zdnd11an1n64x5 FILLER_59_1796 ();
 b15zdnd11an1n64x5 FILLER_59_1860 ();
 b15zdnd11an1n64x5 FILLER_59_1924 ();
 b15zdnd11an1n64x5 FILLER_59_1988 ();
 b15zdnd11an1n64x5 FILLER_59_2052 ();
 b15zdnd11an1n64x5 FILLER_59_2116 ();
 b15zdnd11an1n64x5 FILLER_59_2180 ();
 b15zdnd11an1n32x5 FILLER_59_2244 ();
 b15zdnd11an1n08x5 FILLER_59_2276 ();
 b15zdnd11an1n64x5 FILLER_60_8 ();
 b15zdnd11an1n64x5 FILLER_60_72 ();
 b15zdnd11an1n64x5 FILLER_60_136 ();
 b15zdnd11an1n32x5 FILLER_60_200 ();
 b15zdnd00an1n02x5 FILLER_60_232 ();
 b15zdnd00an1n01x5 FILLER_60_234 ();
 b15zdnd11an1n32x5 FILLER_60_238 ();
 b15zdnd11an1n16x5 FILLER_60_270 ();
 b15zdnd11an1n08x5 FILLER_60_286 ();
 b15zdnd00an1n02x5 FILLER_60_294 ();
 b15zdnd00an1n01x5 FILLER_60_296 ();
 b15zdnd11an1n64x5 FILLER_60_306 ();
 b15zdnd11an1n64x5 FILLER_60_370 ();
 b15zdnd11an1n64x5 FILLER_60_434 ();
 b15zdnd11an1n04x5 FILLER_60_498 ();
 b15zdnd00an1n01x5 FILLER_60_502 ();
 b15zdnd11an1n32x5 FILLER_60_517 ();
 b15zdnd11an1n64x5 FILLER_60_563 ();
 b15zdnd11an1n64x5 FILLER_60_627 ();
 b15zdnd11an1n16x5 FILLER_60_691 ();
 b15zdnd11an1n08x5 FILLER_60_707 ();
 b15zdnd00an1n02x5 FILLER_60_715 ();
 b15zdnd00an1n01x5 FILLER_60_717 ();
 b15zdnd11an1n64x5 FILLER_60_726 ();
 b15zdnd11an1n64x5 FILLER_60_790 ();
 b15zdnd11an1n32x5 FILLER_60_854 ();
 b15zdnd11an1n16x5 FILLER_60_886 ();
 b15zdnd00an1n02x5 FILLER_60_902 ();
 b15zdnd11an1n64x5 FILLER_60_907 ();
 b15zdnd11an1n64x5 FILLER_60_971 ();
 b15zdnd11an1n64x5 FILLER_60_1035 ();
 b15zdnd11an1n64x5 FILLER_60_1099 ();
 b15zdnd11an1n64x5 FILLER_60_1163 ();
 b15zdnd11an1n16x5 FILLER_60_1227 ();
 b15zdnd11an1n08x5 FILLER_60_1243 ();
 b15zdnd11an1n64x5 FILLER_60_1267 ();
 b15zdnd11an1n64x5 FILLER_60_1331 ();
 b15zdnd11an1n64x5 FILLER_60_1395 ();
 b15zdnd11an1n64x5 FILLER_60_1459 ();
 b15zdnd11an1n08x5 FILLER_60_1523 ();
 b15zdnd11an1n04x5 FILLER_60_1531 ();
 b15zdnd00an1n02x5 FILLER_60_1535 ();
 b15zdnd11an1n08x5 FILLER_60_1540 ();
 b15zdnd00an1n01x5 FILLER_60_1548 ();
 b15zdnd11an1n64x5 FILLER_60_1552 ();
 b15zdnd11an1n08x5 FILLER_60_1616 ();
 b15zdnd00an1n02x5 FILLER_60_1624 ();
 b15zdnd11an1n64x5 FILLER_60_1657 ();
 b15zdnd11an1n64x5 FILLER_60_1721 ();
 b15zdnd11an1n64x5 FILLER_60_1785 ();
 b15zdnd11an1n64x5 FILLER_60_1849 ();
 b15zdnd11an1n64x5 FILLER_60_1913 ();
 b15zdnd11an1n64x5 FILLER_60_1977 ();
 b15zdnd11an1n64x5 FILLER_60_2041 ();
 b15zdnd11an1n32x5 FILLER_60_2105 ();
 b15zdnd11an1n16x5 FILLER_60_2137 ();
 b15zdnd00an1n01x5 FILLER_60_2153 ();
 b15zdnd11an1n64x5 FILLER_60_2162 ();
 b15zdnd11an1n32x5 FILLER_60_2226 ();
 b15zdnd11an1n08x5 FILLER_60_2258 ();
 b15zdnd11an1n04x5 FILLER_60_2270 ();
 b15zdnd00an1n02x5 FILLER_60_2274 ();
 b15zdnd11an1n64x5 FILLER_61_0 ();
 b15zdnd11an1n64x5 FILLER_61_64 ();
 b15zdnd11an1n64x5 FILLER_61_128 ();
 b15zdnd11an1n08x5 FILLER_61_192 ();
 b15zdnd11an1n04x5 FILLER_61_200 ();
 b15zdnd00an1n02x5 FILLER_61_204 ();
 b15zdnd00an1n01x5 FILLER_61_206 ();
 b15zdnd11an1n64x5 FILLER_61_259 ();
 b15zdnd11an1n64x5 FILLER_61_323 ();
 b15zdnd11an1n64x5 FILLER_61_387 ();
 b15zdnd11an1n16x5 FILLER_61_451 ();
 b15zdnd11an1n08x5 FILLER_61_467 ();
 b15zdnd11an1n04x5 FILLER_61_475 ();
 b15zdnd11an1n16x5 FILLER_61_493 ();
 b15zdnd00an1n02x5 FILLER_61_509 ();
 b15zdnd00an1n01x5 FILLER_61_511 ();
 b15zdnd11an1n64x5 FILLER_61_532 ();
 b15zdnd11an1n64x5 FILLER_61_596 ();
 b15zdnd11an1n64x5 FILLER_61_660 ();
 b15zdnd11an1n64x5 FILLER_61_724 ();
 b15zdnd11an1n08x5 FILLER_61_788 ();
 b15zdnd11an1n04x5 FILLER_61_796 ();
 b15zdnd11an1n64x5 FILLER_61_820 ();
 b15zdnd11an1n16x5 FILLER_61_884 ();
 b15zdnd11an1n04x5 FILLER_61_900 ();
 b15zdnd11an1n64x5 FILLER_61_907 ();
 b15zdnd11an1n64x5 FILLER_61_971 ();
 b15zdnd11an1n64x5 FILLER_61_1035 ();
 b15zdnd11an1n64x5 FILLER_61_1099 ();
 b15zdnd11an1n64x5 FILLER_61_1163 ();
 b15zdnd11an1n08x5 FILLER_61_1227 ();
 b15zdnd00an1n02x5 FILLER_61_1235 ();
 b15zdnd11an1n16x5 FILLER_61_1245 ();
 b15zdnd11an1n04x5 FILLER_61_1261 ();
 b15zdnd00an1n01x5 FILLER_61_1265 ();
 b15zdnd11an1n64x5 FILLER_61_1270 ();
 b15zdnd11an1n64x5 FILLER_61_1334 ();
 b15zdnd11an1n64x5 FILLER_61_1398 ();
 b15zdnd11an1n64x5 FILLER_61_1462 ();
 b15zdnd11an1n16x5 FILLER_61_1526 ();
 b15zdnd11an1n04x5 FILLER_61_1542 ();
 b15zdnd11an1n64x5 FILLER_61_1549 ();
 b15zdnd11an1n64x5 FILLER_61_1613 ();
 b15zdnd11an1n64x5 FILLER_61_1677 ();
 b15zdnd11an1n64x5 FILLER_61_1741 ();
 b15zdnd11an1n64x5 FILLER_61_1805 ();
 b15zdnd11an1n64x5 FILLER_61_1869 ();
 b15zdnd11an1n64x5 FILLER_61_1933 ();
 b15zdnd11an1n64x5 FILLER_61_1997 ();
 b15zdnd11an1n64x5 FILLER_61_2061 ();
 b15zdnd11an1n64x5 FILLER_61_2125 ();
 b15zdnd11an1n32x5 FILLER_61_2189 ();
 b15zdnd11an1n16x5 FILLER_61_2221 ();
 b15zdnd00an1n02x5 FILLER_61_2237 ();
 b15zdnd00an1n01x5 FILLER_61_2239 ();
 b15zdnd00an1n02x5 FILLER_61_2282 ();
 b15zdnd11an1n64x5 FILLER_62_8 ();
 b15zdnd11an1n64x5 FILLER_62_72 ();
 b15zdnd11an1n64x5 FILLER_62_136 ();
 b15zdnd11an1n16x5 FILLER_62_200 ();
 b15zdnd11an1n08x5 FILLER_62_216 ();
 b15zdnd11an1n04x5 FILLER_62_224 ();
 b15zdnd00an1n02x5 FILLER_62_228 ();
 b15zdnd11an1n64x5 FILLER_62_233 ();
 b15zdnd11an1n64x5 FILLER_62_297 ();
 b15zdnd11an1n08x5 FILLER_62_361 ();
 b15zdnd11an1n04x5 FILLER_62_369 ();
 b15zdnd00an1n01x5 FILLER_62_373 ();
 b15zdnd11an1n64x5 FILLER_62_377 ();
 b15zdnd11an1n32x5 FILLER_62_441 ();
 b15zdnd11an1n08x5 FILLER_62_473 ();
 b15zdnd11an1n04x5 FILLER_62_481 ();
 b15zdnd11an1n64x5 FILLER_62_505 ();
 b15zdnd11an1n64x5 FILLER_62_569 ();
 b15zdnd11an1n64x5 FILLER_62_633 ();
 b15zdnd11an1n16x5 FILLER_62_697 ();
 b15zdnd11an1n04x5 FILLER_62_713 ();
 b15zdnd00an1n01x5 FILLER_62_717 ();
 b15zdnd11an1n64x5 FILLER_62_726 ();
 b15zdnd11an1n64x5 FILLER_62_790 ();
 b15zdnd11an1n16x5 FILLER_62_854 ();
 b15zdnd11an1n08x5 FILLER_62_870 ();
 b15zdnd00an1n02x5 FILLER_62_878 ();
 b15zdnd11an1n64x5 FILLER_62_932 ();
 b15zdnd11an1n64x5 FILLER_62_996 ();
 b15zdnd11an1n64x5 FILLER_62_1060 ();
 b15zdnd11an1n32x5 FILLER_62_1124 ();
 b15zdnd11an1n08x5 FILLER_62_1156 ();
 b15zdnd00an1n01x5 FILLER_62_1164 ();
 b15zdnd11an1n64x5 FILLER_62_1168 ();
 b15zdnd11an1n64x5 FILLER_62_1232 ();
 b15zdnd11an1n64x5 FILLER_62_1296 ();
 b15zdnd11an1n64x5 FILLER_62_1360 ();
 b15zdnd11an1n32x5 FILLER_62_1424 ();
 b15zdnd11an1n04x5 FILLER_62_1456 ();
 b15zdnd00an1n02x5 FILLER_62_1460 ();
 b15zdnd00an1n01x5 FILLER_62_1462 ();
 b15zdnd11an1n16x5 FILLER_62_1476 ();
 b15zdnd11an1n04x5 FILLER_62_1492 ();
 b15zdnd00an1n02x5 FILLER_62_1496 ();
 b15zdnd00an1n01x5 FILLER_62_1498 ();
 b15zdnd11an1n64x5 FILLER_62_1541 ();
 b15zdnd11an1n64x5 FILLER_62_1605 ();
 b15zdnd11an1n64x5 FILLER_62_1669 ();
 b15zdnd11an1n64x5 FILLER_62_1733 ();
 b15zdnd11an1n64x5 FILLER_62_1797 ();
 b15zdnd11an1n64x5 FILLER_62_1861 ();
 b15zdnd11an1n64x5 FILLER_62_1925 ();
 b15zdnd11an1n64x5 FILLER_62_1989 ();
 b15zdnd11an1n64x5 FILLER_62_2053 ();
 b15zdnd11an1n32x5 FILLER_62_2117 ();
 b15zdnd11an1n04x5 FILLER_62_2149 ();
 b15zdnd00an1n01x5 FILLER_62_2153 ();
 b15zdnd11an1n64x5 FILLER_62_2162 ();
 b15zdnd11an1n04x5 FILLER_62_2226 ();
 b15zdnd00an1n02x5 FILLER_62_2230 ();
 b15zdnd00an1n02x5 FILLER_62_2274 ();
 b15zdnd11an1n64x5 FILLER_63_0 ();
 b15zdnd11an1n64x5 FILLER_63_64 ();
 b15zdnd11an1n64x5 FILLER_63_128 ();
 b15zdnd11an1n32x5 FILLER_63_192 ();
 b15zdnd11an1n04x5 FILLER_63_224 ();
 b15zdnd00an1n02x5 FILLER_63_228 ();
 b15zdnd00an1n01x5 FILLER_63_230 ();
 b15zdnd11an1n64x5 FILLER_63_234 ();
 b15zdnd11an1n64x5 FILLER_63_298 ();
 b15zdnd11an1n08x5 FILLER_63_362 ();
 b15zdnd00an1n02x5 FILLER_63_370 ();
 b15zdnd11an1n04x5 FILLER_63_375 ();
 b15zdnd11an1n04x5 FILLER_63_382 ();
 b15zdnd11an1n64x5 FILLER_63_389 ();
 b15zdnd11an1n16x5 FILLER_63_453 ();
 b15zdnd11an1n08x5 FILLER_63_469 ();
 b15zdnd00an1n02x5 FILLER_63_477 ();
 b15zdnd00an1n01x5 FILLER_63_479 ();
 b15zdnd11an1n64x5 FILLER_63_492 ();
 b15zdnd11an1n64x5 FILLER_63_556 ();
 b15zdnd11an1n64x5 FILLER_63_620 ();
 b15zdnd11an1n64x5 FILLER_63_684 ();
 b15zdnd11an1n64x5 FILLER_63_748 ();
 b15zdnd11an1n64x5 FILLER_63_812 ();
 b15zdnd11an1n08x5 FILLER_63_876 ();
 b15zdnd11an1n04x5 FILLER_63_904 ();
 b15zdnd11an1n64x5 FILLER_63_911 ();
 b15zdnd11an1n64x5 FILLER_63_975 ();
 b15zdnd11an1n64x5 FILLER_63_1039 ();
 b15zdnd11an1n64x5 FILLER_63_1103 ();
 b15zdnd11an1n64x5 FILLER_63_1167 ();
 b15zdnd11an1n64x5 FILLER_63_1231 ();
 b15zdnd11an1n64x5 FILLER_63_1295 ();
 b15zdnd11an1n16x5 FILLER_63_1359 ();
 b15zdnd11an1n04x5 FILLER_63_1375 ();
 b15zdnd11an1n04x5 FILLER_63_1411 ();
 b15zdnd11an1n08x5 FILLER_63_1418 ();
 b15zdnd11an1n04x5 FILLER_63_1426 ();
 b15zdnd00an1n02x5 FILLER_63_1430 ();
 b15zdnd11an1n08x5 FILLER_63_1474 ();
 b15zdnd00an1n02x5 FILLER_63_1482 ();
 b15zdnd00an1n01x5 FILLER_63_1484 ();
 b15zdnd11an1n16x5 FILLER_63_1527 ();
 b15zdnd11an1n04x5 FILLER_63_1543 ();
 b15zdnd00an1n02x5 FILLER_63_1547 ();
 b15zdnd00an1n01x5 FILLER_63_1549 ();
 b15zdnd11an1n32x5 FILLER_63_1592 ();
 b15zdnd11an1n16x5 FILLER_63_1624 ();
 b15zdnd11an1n04x5 FILLER_63_1640 ();
 b15zdnd11an1n04x5 FILLER_63_1668 ();
 b15zdnd11an1n64x5 FILLER_63_1703 ();
 b15zdnd11an1n64x5 FILLER_63_1767 ();
 b15zdnd11an1n64x5 FILLER_63_1831 ();
 b15zdnd11an1n08x5 FILLER_63_1895 ();
 b15zdnd11an1n64x5 FILLER_63_1934 ();
 b15zdnd11an1n32x5 FILLER_63_1998 ();
 b15zdnd11an1n16x5 FILLER_63_2030 ();
 b15zdnd11an1n04x5 FILLER_63_2046 ();
 b15zdnd11an1n64x5 FILLER_63_2102 ();
 b15zdnd11an1n64x5 FILLER_63_2166 ();
 b15zdnd11an1n08x5 FILLER_63_2230 ();
 b15zdnd00an1n02x5 FILLER_63_2238 ();
 b15zdnd00an1n02x5 FILLER_63_2282 ();
 b15zdnd11an1n64x5 FILLER_64_8 ();
 b15zdnd11an1n64x5 FILLER_64_72 ();
 b15zdnd11an1n64x5 FILLER_64_136 ();
 b15zdnd11an1n64x5 FILLER_64_200 ();
 b15zdnd11an1n64x5 FILLER_64_264 ();
 b15zdnd11an1n16x5 FILLER_64_328 ();
 b15zdnd11an1n08x5 FILLER_64_344 ();
 b15zdnd11an1n64x5 FILLER_64_404 ();
 b15zdnd11an1n64x5 FILLER_64_468 ();
 b15zdnd11an1n64x5 FILLER_64_532 ();
 b15zdnd11an1n64x5 FILLER_64_596 ();
 b15zdnd11an1n32x5 FILLER_64_660 ();
 b15zdnd11an1n16x5 FILLER_64_692 ();
 b15zdnd11an1n08x5 FILLER_64_708 ();
 b15zdnd00an1n02x5 FILLER_64_716 ();
 b15zdnd11an1n64x5 FILLER_64_726 ();
 b15zdnd00an1n02x5 FILLER_64_790 ();
 b15zdnd00an1n01x5 FILLER_64_792 ();
 b15zdnd11an1n64x5 FILLER_64_807 ();
 b15zdnd11an1n64x5 FILLER_64_871 ();
 b15zdnd11an1n64x5 FILLER_64_935 ();
 b15zdnd11an1n64x5 FILLER_64_999 ();
 b15zdnd11an1n64x5 FILLER_64_1063 ();
 b15zdnd11an1n32x5 FILLER_64_1127 ();
 b15zdnd11an1n16x5 FILLER_64_1159 ();
 b15zdnd11an1n08x5 FILLER_64_1175 ();
 b15zdnd00an1n02x5 FILLER_64_1183 ();
 b15zdnd00an1n01x5 FILLER_64_1185 ();
 b15zdnd11an1n64x5 FILLER_64_1228 ();
 b15zdnd11an1n64x5 FILLER_64_1292 ();
 b15zdnd11an1n32x5 FILLER_64_1356 ();
 b15zdnd11an1n16x5 FILLER_64_1388 ();
 b15zdnd00an1n02x5 FILLER_64_1404 ();
 b15zdnd00an1n01x5 FILLER_64_1406 ();
 b15zdnd11an1n64x5 FILLER_64_1410 ();
 b15zdnd11an1n64x5 FILLER_64_1474 ();
 b15zdnd11an1n64x5 FILLER_64_1538 ();
 b15zdnd11an1n32x5 FILLER_64_1602 ();
 b15zdnd11an1n08x5 FILLER_64_1634 ();
 b15zdnd00an1n02x5 FILLER_64_1642 ();
 b15zdnd11an1n64x5 FILLER_64_1661 ();
 b15zdnd11an1n64x5 FILLER_64_1725 ();
 b15zdnd11an1n64x5 FILLER_64_1789 ();
 b15zdnd11an1n64x5 FILLER_64_1853 ();
 b15zdnd11an1n64x5 FILLER_64_1917 ();
 b15zdnd11an1n32x5 FILLER_64_1981 ();
 b15zdnd11an1n16x5 FILLER_64_2013 ();
 b15zdnd11an1n04x5 FILLER_64_2029 ();
 b15zdnd11an1n04x5 FILLER_64_2085 ();
 b15zdnd11an1n32x5 FILLER_64_2092 ();
 b15zdnd11an1n16x5 FILLER_64_2124 ();
 b15zdnd11an1n08x5 FILLER_64_2140 ();
 b15zdnd11an1n04x5 FILLER_64_2148 ();
 b15zdnd00an1n02x5 FILLER_64_2152 ();
 b15zdnd11an1n64x5 FILLER_64_2162 ();
 b15zdnd11an1n04x5 FILLER_64_2226 ();
 b15zdnd00an1n02x5 FILLER_64_2230 ();
 b15zdnd00an1n02x5 FILLER_64_2274 ();
 b15zdnd11an1n64x5 FILLER_65_0 ();
 b15zdnd11an1n64x5 FILLER_65_64 ();
 b15zdnd11an1n64x5 FILLER_65_128 ();
 b15zdnd11an1n64x5 FILLER_65_192 ();
 b15zdnd11an1n64x5 FILLER_65_256 ();
 b15zdnd11an1n32x5 FILLER_65_320 ();
 b15zdnd11an1n16x5 FILLER_65_352 ();
 b15zdnd11an1n04x5 FILLER_65_368 ();
 b15zdnd00an1n02x5 FILLER_65_372 ();
 b15zdnd11an1n08x5 FILLER_65_377 ();
 b15zdnd00an1n01x5 FILLER_65_385 ();
 b15zdnd11an1n64x5 FILLER_65_389 ();
 b15zdnd11an1n64x5 FILLER_65_453 ();
 b15zdnd11an1n08x5 FILLER_65_517 ();
 b15zdnd11an1n04x5 FILLER_65_525 ();
 b15zdnd00an1n02x5 FILLER_65_529 ();
 b15zdnd00an1n01x5 FILLER_65_531 ();
 b15zdnd11an1n64x5 FILLER_65_549 ();
 b15zdnd11an1n64x5 FILLER_65_613 ();
 b15zdnd11an1n64x5 FILLER_65_677 ();
 b15zdnd11an1n64x5 FILLER_65_741 ();
 b15zdnd11an1n32x5 FILLER_65_805 ();
 b15zdnd11an1n16x5 FILLER_65_837 ();
 b15zdnd11an1n08x5 FILLER_65_853 ();
 b15zdnd11an1n64x5 FILLER_65_878 ();
 b15zdnd11an1n32x5 FILLER_65_942 ();
 b15zdnd00an1n02x5 FILLER_65_974 ();
 b15zdnd00an1n01x5 FILLER_65_976 ();
 b15zdnd11an1n64x5 FILLER_65_986 ();
 b15zdnd11an1n64x5 FILLER_65_1050 ();
 b15zdnd11an1n32x5 FILLER_65_1114 ();
 b15zdnd11an1n08x5 FILLER_65_1146 ();
 b15zdnd00an1n02x5 FILLER_65_1154 ();
 b15zdnd00an1n01x5 FILLER_65_1156 ();
 b15zdnd11an1n64x5 FILLER_65_1199 ();
 b15zdnd11an1n64x5 FILLER_65_1263 ();
 b15zdnd11an1n64x5 FILLER_65_1327 ();
 b15zdnd11an1n64x5 FILLER_65_1391 ();
 b15zdnd11an1n64x5 FILLER_65_1455 ();
 b15zdnd11an1n32x5 FILLER_65_1519 ();
 b15zdnd11an1n16x5 FILLER_65_1551 ();
 b15zdnd11an1n08x5 FILLER_65_1567 ();
 b15zdnd00an1n02x5 FILLER_65_1575 ();
 b15zdnd11an1n32x5 FILLER_65_1586 ();
 b15zdnd11an1n16x5 FILLER_65_1618 ();
 b15zdnd11an1n08x5 FILLER_65_1634 ();
 b15zdnd00an1n02x5 FILLER_65_1642 ();
 b15zdnd11an1n64x5 FILLER_65_1668 ();
 b15zdnd11an1n64x5 FILLER_65_1732 ();
 b15zdnd11an1n64x5 FILLER_65_1796 ();
 b15zdnd11an1n32x5 FILLER_65_1860 ();
 b15zdnd11an1n16x5 FILLER_65_1892 ();
 b15zdnd11an1n64x5 FILLER_65_1928 ();
 b15zdnd11an1n32x5 FILLER_65_1992 ();
 b15zdnd11an1n16x5 FILLER_65_2024 ();
 b15zdnd11an1n08x5 FILLER_65_2040 ();
 b15zdnd00an1n02x5 FILLER_65_2048 ();
 b15zdnd00an1n01x5 FILLER_65_2050 ();
 b15zdnd11an1n04x5 FILLER_65_2054 ();
 b15zdnd11an1n04x5 FILLER_65_2061 ();
 b15zdnd00an1n02x5 FILLER_65_2065 ();
 b15zdnd00an1n01x5 FILLER_65_2067 ();
 b15zdnd11an1n04x5 FILLER_65_2071 ();
 b15zdnd11an1n64x5 FILLER_65_2078 ();
 b15zdnd11an1n64x5 FILLER_65_2142 ();
 b15zdnd11an1n32x5 FILLER_65_2206 ();
 b15zdnd11an1n04x5 FILLER_65_2238 ();
 b15zdnd00an1n02x5 FILLER_65_2242 ();
 b15zdnd11an1n32x5 FILLER_65_2248 ();
 b15zdnd11an1n04x5 FILLER_65_2280 ();
 b15zdnd11an1n64x5 FILLER_66_8 ();
 b15zdnd11an1n64x5 FILLER_66_72 ();
 b15zdnd11an1n64x5 FILLER_66_136 ();
 b15zdnd00an1n01x5 FILLER_66_200 ();
 b15zdnd11an1n04x5 FILLER_66_204 ();
 b15zdnd11an1n64x5 FILLER_66_211 ();
 b15zdnd11an1n64x5 FILLER_66_275 ();
 b15zdnd11an1n08x5 FILLER_66_339 ();
 b15zdnd11an1n04x5 FILLER_66_347 ();
 b15zdnd00an1n02x5 FILLER_66_351 ();
 b15zdnd11an1n04x5 FILLER_66_356 ();
 b15zdnd11an1n32x5 FILLER_66_412 ();
 b15zdnd11an1n16x5 FILLER_66_444 ();
 b15zdnd11an1n08x5 FILLER_66_460 ();
 b15zdnd11an1n04x5 FILLER_66_468 ();
 b15zdnd00an1n02x5 FILLER_66_472 ();
 b15zdnd11an1n32x5 FILLER_66_494 ();
 b15zdnd11an1n16x5 FILLER_66_526 ();
 b15zdnd00an1n02x5 FILLER_66_542 ();
 b15zdnd11an1n64x5 FILLER_66_586 ();
 b15zdnd11an1n64x5 FILLER_66_650 ();
 b15zdnd11an1n04x5 FILLER_66_714 ();
 b15zdnd11an1n16x5 FILLER_66_726 ();
 b15zdnd11an1n64x5 FILLER_66_759 ();
 b15zdnd11an1n64x5 FILLER_66_823 ();
 b15zdnd11an1n64x5 FILLER_66_887 ();
 b15zdnd11an1n64x5 FILLER_66_951 ();
 b15zdnd11an1n64x5 FILLER_66_1015 ();
 b15zdnd11an1n64x5 FILLER_66_1079 ();
 b15zdnd11an1n64x5 FILLER_66_1143 ();
 b15zdnd11an1n16x5 FILLER_66_1207 ();
 b15zdnd11an1n04x5 FILLER_66_1223 ();
 b15zdnd00an1n02x5 FILLER_66_1227 ();
 b15zdnd11an1n08x5 FILLER_66_1237 ();
 b15zdnd00an1n02x5 FILLER_66_1245 ();
 b15zdnd00an1n01x5 FILLER_66_1247 ();
 b15zdnd11an1n32x5 FILLER_66_1254 ();
 b15zdnd11an1n16x5 FILLER_66_1286 ();
 b15zdnd11an1n08x5 FILLER_66_1302 ();
 b15zdnd11an1n04x5 FILLER_66_1310 ();
 b15zdnd00an1n02x5 FILLER_66_1314 ();
 b15zdnd00an1n01x5 FILLER_66_1316 ();
 b15zdnd11an1n64x5 FILLER_66_1359 ();
 b15zdnd00an1n02x5 FILLER_66_1423 ();
 b15zdnd11an1n08x5 FILLER_66_1467 ();
 b15zdnd11an1n64x5 FILLER_66_1517 ();
 b15zdnd11an1n32x5 FILLER_66_1581 ();
 b15zdnd11an1n16x5 FILLER_66_1613 ();
 b15zdnd11an1n08x5 FILLER_66_1629 ();
 b15zdnd00an1n02x5 FILLER_66_1637 ();
 b15zdnd00an1n01x5 FILLER_66_1639 ();
 b15zdnd11an1n64x5 FILLER_66_1664 ();
 b15zdnd11an1n64x5 FILLER_66_1728 ();
 b15zdnd11an1n64x5 FILLER_66_1792 ();
 b15zdnd11an1n32x5 FILLER_66_1856 ();
 b15zdnd11an1n16x5 FILLER_66_1888 ();
 b15zdnd00an1n02x5 FILLER_66_1904 ();
 b15zdnd11an1n04x5 FILLER_66_1926 ();
 b15zdnd11an1n64x5 FILLER_66_1933 ();
 b15zdnd11an1n32x5 FILLER_66_1997 ();
 b15zdnd11an1n16x5 FILLER_66_2029 ();
 b15zdnd11an1n08x5 FILLER_66_2045 ();
 b15zdnd11an1n04x5 FILLER_66_2053 ();
 b15zdnd00an1n01x5 FILLER_66_2057 ();
 b15zdnd11an1n64x5 FILLER_66_2061 ();
 b15zdnd11an1n16x5 FILLER_66_2125 ();
 b15zdnd11an1n08x5 FILLER_66_2141 ();
 b15zdnd11an1n04x5 FILLER_66_2149 ();
 b15zdnd00an1n01x5 FILLER_66_2153 ();
 b15zdnd11an1n64x5 FILLER_66_2162 ();
 b15zdnd11an1n32x5 FILLER_66_2226 ();
 b15zdnd11an1n16x5 FILLER_66_2258 ();
 b15zdnd00an1n02x5 FILLER_66_2274 ();
 b15zdnd11an1n16x5 FILLER_67_0 ();
 b15zdnd11an1n04x5 FILLER_67_16 ();
 b15zdnd00an1n02x5 FILLER_67_20 ();
 b15zdnd00an1n01x5 FILLER_67_22 ();
 b15zdnd11an1n64x5 FILLER_67_26 ();
 b15zdnd11an1n64x5 FILLER_67_90 ();
 b15zdnd11an1n16x5 FILLER_67_154 ();
 b15zdnd11an1n08x5 FILLER_67_170 ();
 b15zdnd00an1n02x5 FILLER_67_178 ();
 b15zdnd00an1n01x5 FILLER_67_180 ();
 b15zdnd11an1n64x5 FILLER_67_233 ();
 b15zdnd11an1n16x5 FILLER_67_297 ();
 b15zdnd11an1n08x5 FILLER_67_313 ();
 b15zdnd11an1n04x5 FILLER_67_321 ();
 b15zdnd00an1n01x5 FILLER_67_325 ();
 b15zdnd11an1n64x5 FILLER_67_378 ();
 b15zdnd11an1n64x5 FILLER_67_442 ();
 b15zdnd11an1n64x5 FILLER_67_506 ();
 b15zdnd11an1n64x5 FILLER_67_570 ();
 b15zdnd11an1n64x5 FILLER_67_634 ();
 b15zdnd00an1n02x5 FILLER_67_698 ();
 b15zdnd11an1n32x5 FILLER_67_709 ();
 b15zdnd11an1n16x5 FILLER_67_741 ();
 b15zdnd00an1n02x5 FILLER_67_757 ();
 b15zdnd11an1n64x5 FILLER_67_779 ();
 b15zdnd00an1n02x5 FILLER_67_843 ();
 b15zdnd00an1n01x5 FILLER_67_845 ();
 b15zdnd11an1n16x5 FILLER_67_860 ();
 b15zdnd00an1n02x5 FILLER_67_876 ();
 b15zdnd11an1n64x5 FILLER_67_898 ();
 b15zdnd11an1n64x5 FILLER_67_962 ();
 b15zdnd11an1n64x5 FILLER_67_1026 ();
 b15zdnd11an1n64x5 FILLER_67_1090 ();
 b15zdnd11an1n64x5 FILLER_67_1154 ();
 b15zdnd11an1n64x5 FILLER_67_1218 ();
 b15zdnd11an1n64x5 FILLER_67_1282 ();
 b15zdnd11an1n64x5 FILLER_67_1346 ();
 b15zdnd11an1n64x5 FILLER_67_1410 ();
 b15zdnd11an1n64x5 FILLER_67_1474 ();
 b15zdnd11an1n64x5 FILLER_67_1538 ();
 b15zdnd11an1n64x5 FILLER_67_1602 ();
 b15zdnd11an1n64x5 FILLER_67_1666 ();
 b15zdnd11an1n64x5 FILLER_67_1730 ();
 b15zdnd11an1n64x5 FILLER_67_1794 ();
 b15zdnd11an1n64x5 FILLER_67_1858 ();
 b15zdnd11an1n04x5 FILLER_67_1922 ();
 b15zdnd00an1n01x5 FILLER_67_1926 ();
 b15zdnd11an1n64x5 FILLER_67_1954 ();
 b15zdnd11an1n64x5 FILLER_67_2018 ();
 b15zdnd11an1n64x5 FILLER_67_2082 ();
 b15zdnd11an1n64x5 FILLER_67_2146 ();
 b15zdnd11an1n64x5 FILLER_67_2210 ();
 b15zdnd11an1n08x5 FILLER_67_2274 ();
 b15zdnd00an1n02x5 FILLER_67_2282 ();
 b15zdnd11an1n08x5 FILLER_68_8 ();
 b15zdnd11an1n04x5 FILLER_68_16 ();
 b15zdnd00an1n02x5 FILLER_68_20 ();
 b15zdnd11an1n64x5 FILLER_68_25 ();
 b15zdnd11an1n64x5 FILLER_68_89 ();
 b15zdnd11an1n16x5 FILLER_68_153 ();
 b15zdnd11an1n08x5 FILLER_68_169 ();
 b15zdnd11an1n04x5 FILLER_68_177 ();
 b15zdnd11an1n64x5 FILLER_68_233 ();
 b15zdnd11an1n32x5 FILLER_68_297 ();
 b15zdnd11an1n16x5 FILLER_68_329 ();
 b15zdnd11an1n04x5 FILLER_68_345 ();
 b15zdnd00an1n02x5 FILLER_68_349 ();
 b15zdnd00an1n01x5 FILLER_68_351 ();
 b15zdnd11an1n64x5 FILLER_68_355 ();
 b15zdnd11an1n64x5 FILLER_68_419 ();
 b15zdnd11an1n32x5 FILLER_68_483 ();
 b15zdnd11an1n16x5 FILLER_68_515 ();
 b15zdnd11an1n08x5 FILLER_68_531 ();
 b15zdnd00an1n02x5 FILLER_68_539 ();
 b15zdnd11an1n64x5 FILLER_68_561 ();
 b15zdnd11an1n64x5 FILLER_68_625 ();
 b15zdnd11an1n16x5 FILLER_68_689 ();
 b15zdnd11an1n08x5 FILLER_68_705 ();
 b15zdnd11an1n04x5 FILLER_68_713 ();
 b15zdnd00an1n01x5 FILLER_68_717 ();
 b15zdnd11an1n64x5 FILLER_68_726 ();
 b15zdnd11an1n64x5 FILLER_68_790 ();
 b15zdnd11an1n64x5 FILLER_68_854 ();
 b15zdnd11an1n32x5 FILLER_68_918 ();
 b15zdnd11an1n08x5 FILLER_68_950 ();
 b15zdnd00an1n02x5 FILLER_68_958 ();
 b15zdnd11an1n64x5 FILLER_68_969 ();
 b15zdnd11an1n64x5 FILLER_68_1033 ();
 b15zdnd11an1n64x5 FILLER_68_1097 ();
 b15zdnd11an1n64x5 FILLER_68_1161 ();
 b15zdnd11an1n64x5 FILLER_68_1225 ();
 b15zdnd11an1n64x5 FILLER_68_1289 ();
 b15zdnd11an1n04x5 FILLER_68_1353 ();
 b15zdnd00an1n01x5 FILLER_68_1357 ();
 b15zdnd11an1n16x5 FILLER_68_1363 ();
 b15zdnd11an1n08x5 FILLER_68_1379 ();
 b15zdnd11an1n04x5 FILLER_68_1387 ();
 b15zdnd11an1n64x5 FILLER_68_1396 ();
 b15zdnd11an1n64x5 FILLER_68_1460 ();
 b15zdnd11an1n64x5 FILLER_68_1524 ();
 b15zdnd11an1n64x5 FILLER_68_1588 ();
 b15zdnd11an1n64x5 FILLER_68_1652 ();
 b15zdnd11an1n64x5 FILLER_68_1716 ();
 b15zdnd11an1n64x5 FILLER_68_1780 ();
 b15zdnd11an1n32x5 FILLER_68_1844 ();
 b15zdnd11an1n16x5 FILLER_68_1876 ();
 b15zdnd11an1n08x5 FILLER_68_1892 ();
 b15zdnd11an1n04x5 FILLER_68_1900 ();
 b15zdnd00an1n01x5 FILLER_68_1904 ();
 b15zdnd11an1n64x5 FILLER_68_1957 ();
 b15zdnd11an1n64x5 FILLER_68_2021 ();
 b15zdnd11an1n64x5 FILLER_68_2085 ();
 b15zdnd11an1n04x5 FILLER_68_2149 ();
 b15zdnd00an1n01x5 FILLER_68_2153 ();
 b15zdnd11an1n64x5 FILLER_68_2162 ();
 b15zdnd11an1n32x5 FILLER_68_2226 ();
 b15zdnd11an1n16x5 FILLER_68_2258 ();
 b15zdnd00an1n02x5 FILLER_68_2274 ();
 b15zdnd11an1n64x5 FILLER_69_0 ();
 b15zdnd11an1n64x5 FILLER_69_64 ();
 b15zdnd11an1n64x5 FILLER_69_128 ();
 b15zdnd11an1n08x5 FILLER_69_192 ();
 b15zdnd00an1n01x5 FILLER_69_200 ();
 b15zdnd11an1n04x5 FILLER_69_204 ();
 b15zdnd11an1n64x5 FILLER_69_211 ();
 b15zdnd11an1n64x5 FILLER_69_275 ();
 b15zdnd11an1n08x5 FILLER_69_339 ();
 b15zdnd00an1n02x5 FILLER_69_347 ();
 b15zdnd00an1n01x5 FILLER_69_349 ();
 b15zdnd11an1n64x5 FILLER_69_353 ();
 b15zdnd11an1n64x5 FILLER_69_417 ();
 b15zdnd11an1n32x5 FILLER_69_481 ();
 b15zdnd11an1n16x5 FILLER_69_513 ();
 b15zdnd00an1n01x5 FILLER_69_529 ();
 b15zdnd11an1n64x5 FILLER_69_547 ();
 b15zdnd11an1n16x5 FILLER_69_611 ();
 b15zdnd11an1n04x5 FILLER_69_627 ();
 b15zdnd00an1n02x5 FILLER_69_631 ();
 b15zdnd11an1n16x5 FILLER_69_645 ();
 b15zdnd00an1n02x5 FILLER_69_661 ();
 b15zdnd00an1n01x5 FILLER_69_663 ();
 b15zdnd11an1n04x5 FILLER_69_678 ();
 b15zdnd11an1n32x5 FILLER_69_702 ();
 b15zdnd00an1n01x5 FILLER_69_734 ();
 b15zdnd11an1n64x5 FILLER_69_755 ();
 b15zdnd11an1n64x5 FILLER_69_819 ();
 b15zdnd11an1n64x5 FILLER_69_883 ();
 b15zdnd11an1n64x5 FILLER_69_947 ();
 b15zdnd11an1n64x5 FILLER_69_1011 ();
 b15zdnd11an1n64x5 FILLER_69_1075 ();
 b15zdnd11an1n32x5 FILLER_69_1139 ();
 b15zdnd11an1n04x5 FILLER_69_1171 ();
 b15zdnd00an1n01x5 FILLER_69_1175 ();
 b15zdnd11an1n32x5 FILLER_69_1179 ();
 b15zdnd11an1n16x5 FILLER_69_1211 ();
 b15zdnd11an1n08x5 FILLER_69_1227 ();
 b15zdnd11an1n04x5 FILLER_69_1235 ();
 b15zdnd00an1n02x5 FILLER_69_1239 ();
 b15zdnd11an1n64x5 FILLER_69_1269 ();
 b15zdnd11an1n64x5 FILLER_69_1333 ();
 b15zdnd11an1n64x5 FILLER_69_1397 ();
 b15zdnd11an1n64x5 FILLER_69_1461 ();
 b15zdnd11an1n64x5 FILLER_69_1525 ();
 b15zdnd11an1n64x5 FILLER_69_1589 ();
 b15zdnd11an1n64x5 FILLER_69_1653 ();
 b15zdnd11an1n64x5 FILLER_69_1717 ();
 b15zdnd11an1n64x5 FILLER_69_1781 ();
 b15zdnd11an1n64x5 FILLER_69_1845 ();
 b15zdnd11an1n08x5 FILLER_69_1909 ();
 b15zdnd11an1n04x5 FILLER_69_1917 ();
 b15zdnd00an1n01x5 FILLER_69_1921 ();
 b15zdnd11an1n04x5 FILLER_69_1925 ();
 b15zdnd11an1n04x5 FILLER_69_1932 ();
 b15zdnd11an1n64x5 FILLER_69_1939 ();
 b15zdnd11an1n64x5 FILLER_69_2003 ();
 b15zdnd11an1n64x5 FILLER_69_2067 ();
 b15zdnd11an1n64x5 FILLER_69_2131 ();
 b15zdnd11an1n64x5 FILLER_69_2195 ();
 b15zdnd11an1n16x5 FILLER_69_2259 ();
 b15zdnd11an1n08x5 FILLER_69_2275 ();
 b15zdnd00an1n01x5 FILLER_69_2283 ();
 b15zdnd11an1n64x5 FILLER_70_8 ();
 b15zdnd11an1n64x5 FILLER_70_72 ();
 b15zdnd11an1n64x5 FILLER_70_136 ();
 b15zdnd11an1n04x5 FILLER_70_203 ();
 b15zdnd11an1n64x5 FILLER_70_210 ();
 b15zdnd11an1n64x5 FILLER_70_274 ();
 b15zdnd11an1n64x5 FILLER_70_338 ();
 b15zdnd11an1n64x5 FILLER_70_402 ();
 b15zdnd11an1n64x5 FILLER_70_466 ();
 b15zdnd11an1n64x5 FILLER_70_530 ();
 b15zdnd11an1n64x5 FILLER_70_594 ();
 b15zdnd11an1n32x5 FILLER_70_658 ();
 b15zdnd11an1n16x5 FILLER_70_690 ();
 b15zdnd11an1n08x5 FILLER_70_706 ();
 b15zdnd11an1n04x5 FILLER_70_714 ();
 b15zdnd11an1n64x5 FILLER_70_726 ();
 b15zdnd11an1n64x5 FILLER_70_790 ();
 b15zdnd11an1n64x5 FILLER_70_854 ();
 b15zdnd11an1n64x5 FILLER_70_918 ();
 b15zdnd11an1n64x5 FILLER_70_982 ();
 b15zdnd11an1n64x5 FILLER_70_1046 ();
 b15zdnd11an1n64x5 FILLER_70_1110 ();
 b15zdnd11an1n04x5 FILLER_70_1177 ();
 b15zdnd11an1n64x5 FILLER_70_1184 ();
 b15zdnd11an1n64x5 FILLER_70_1248 ();
 b15zdnd11an1n64x5 FILLER_70_1312 ();
 b15zdnd11an1n64x5 FILLER_70_1376 ();
 b15zdnd11an1n64x5 FILLER_70_1440 ();
 b15zdnd11an1n64x5 FILLER_70_1504 ();
 b15zdnd11an1n64x5 FILLER_70_1568 ();
 b15zdnd11an1n64x5 FILLER_70_1632 ();
 b15zdnd11an1n64x5 FILLER_70_1696 ();
 b15zdnd11an1n64x5 FILLER_70_1760 ();
 b15zdnd11an1n64x5 FILLER_70_1824 ();
 b15zdnd11an1n64x5 FILLER_70_1888 ();
 b15zdnd11an1n64x5 FILLER_70_1952 ();
 b15zdnd11an1n64x5 FILLER_70_2016 ();
 b15zdnd11an1n64x5 FILLER_70_2080 ();
 b15zdnd11an1n08x5 FILLER_70_2144 ();
 b15zdnd00an1n02x5 FILLER_70_2152 ();
 b15zdnd11an1n64x5 FILLER_70_2162 ();
 b15zdnd11an1n32x5 FILLER_70_2226 ();
 b15zdnd11an1n16x5 FILLER_70_2258 ();
 b15zdnd00an1n02x5 FILLER_70_2274 ();
 b15zdnd11an1n64x5 FILLER_71_0 ();
 b15zdnd11an1n64x5 FILLER_71_64 ();
 b15zdnd11an1n64x5 FILLER_71_128 ();
 b15zdnd11an1n64x5 FILLER_71_192 ();
 b15zdnd11an1n64x5 FILLER_71_256 ();
 b15zdnd11an1n64x5 FILLER_71_320 ();
 b15zdnd11an1n64x5 FILLER_71_384 ();
 b15zdnd11an1n64x5 FILLER_71_448 ();
 b15zdnd11an1n08x5 FILLER_71_512 ();
 b15zdnd00an1n01x5 FILLER_71_520 ();
 b15zdnd11an1n08x5 FILLER_71_541 ();
 b15zdnd00an1n02x5 FILLER_71_549 ();
 b15zdnd00an1n01x5 FILLER_71_551 ();
 b15zdnd11an1n64x5 FILLER_71_572 ();
 b15zdnd11an1n64x5 FILLER_71_636 ();
 b15zdnd11an1n64x5 FILLER_71_700 ();
 b15zdnd11an1n16x5 FILLER_71_764 ();
 b15zdnd11an1n04x5 FILLER_71_780 ();
 b15zdnd11an1n64x5 FILLER_71_808 ();
 b15zdnd11an1n64x5 FILLER_71_872 ();
 b15zdnd11an1n64x5 FILLER_71_936 ();
 b15zdnd11an1n64x5 FILLER_71_1000 ();
 b15zdnd11an1n64x5 FILLER_71_1064 ();
 b15zdnd11an1n32x5 FILLER_71_1128 ();
 b15zdnd11an1n08x5 FILLER_71_1160 ();
 b15zdnd00an1n01x5 FILLER_71_1168 ();
 b15zdnd11an1n64x5 FILLER_71_1189 ();
 b15zdnd11an1n64x5 FILLER_71_1253 ();
 b15zdnd11an1n64x5 FILLER_71_1317 ();
 b15zdnd11an1n64x5 FILLER_71_1381 ();
 b15zdnd11an1n64x5 FILLER_71_1445 ();
 b15zdnd11an1n64x5 FILLER_71_1509 ();
 b15zdnd11an1n64x5 FILLER_71_1573 ();
 b15zdnd11an1n64x5 FILLER_71_1637 ();
 b15zdnd11an1n64x5 FILLER_71_1701 ();
 b15zdnd11an1n64x5 FILLER_71_1765 ();
 b15zdnd11an1n64x5 FILLER_71_1829 ();
 b15zdnd11an1n64x5 FILLER_71_1893 ();
 b15zdnd11an1n64x5 FILLER_71_1957 ();
 b15zdnd11an1n64x5 FILLER_71_2021 ();
 b15zdnd11an1n64x5 FILLER_71_2085 ();
 b15zdnd11an1n64x5 FILLER_71_2149 ();
 b15zdnd11an1n64x5 FILLER_71_2213 ();
 b15zdnd11an1n04x5 FILLER_71_2277 ();
 b15zdnd00an1n02x5 FILLER_71_2281 ();
 b15zdnd00an1n01x5 FILLER_71_2283 ();
 b15zdnd11an1n16x5 FILLER_72_8 ();
 b15zdnd11an1n08x5 FILLER_72_24 ();
 b15zdnd11an1n04x5 FILLER_72_32 ();
 b15zdnd11an1n64x5 FILLER_72_39 ();
 b15zdnd11an1n64x5 FILLER_72_103 ();
 b15zdnd11an1n64x5 FILLER_72_167 ();
 b15zdnd11an1n64x5 FILLER_72_231 ();
 b15zdnd11an1n64x5 FILLER_72_295 ();
 b15zdnd11an1n64x5 FILLER_72_359 ();
 b15zdnd11an1n64x5 FILLER_72_423 ();
 b15zdnd11an1n32x5 FILLER_72_487 ();
 b15zdnd11an1n08x5 FILLER_72_519 ();
 b15zdnd00an1n02x5 FILLER_72_527 ();
 b15zdnd11an1n64x5 FILLER_72_546 ();
 b15zdnd11an1n64x5 FILLER_72_610 ();
 b15zdnd11an1n32x5 FILLER_72_674 ();
 b15zdnd11an1n08x5 FILLER_72_706 ();
 b15zdnd11an1n04x5 FILLER_72_714 ();
 b15zdnd11an1n16x5 FILLER_72_726 ();
 b15zdnd00an1n02x5 FILLER_72_742 ();
 b15zdnd00an1n01x5 FILLER_72_744 ();
 b15zdnd11an1n64x5 FILLER_72_768 ();
 b15zdnd11an1n32x5 FILLER_72_832 ();
 b15zdnd11an1n04x5 FILLER_72_864 ();
 b15zdnd00an1n02x5 FILLER_72_868 ();
 b15zdnd11an1n64x5 FILLER_72_890 ();
 b15zdnd11an1n64x5 FILLER_72_954 ();
 b15zdnd11an1n64x5 FILLER_72_1018 ();
 b15zdnd11an1n64x5 FILLER_72_1082 ();
 b15zdnd11an1n08x5 FILLER_72_1146 ();
 b15zdnd00an1n02x5 FILLER_72_1154 ();
 b15zdnd11an1n64x5 FILLER_72_1208 ();
 b15zdnd11an1n64x5 FILLER_72_1272 ();
 b15zdnd11an1n64x5 FILLER_72_1336 ();
 b15zdnd11an1n64x5 FILLER_72_1400 ();
 b15zdnd11an1n08x5 FILLER_72_1464 ();
 b15zdnd00an1n02x5 FILLER_72_1472 ();
 b15zdnd00an1n01x5 FILLER_72_1474 ();
 b15zdnd11an1n64x5 FILLER_72_1495 ();
 b15zdnd11an1n64x5 FILLER_72_1559 ();
 b15zdnd11an1n64x5 FILLER_72_1623 ();
 b15zdnd11an1n64x5 FILLER_72_1687 ();
 b15zdnd11an1n64x5 FILLER_72_1751 ();
 b15zdnd11an1n64x5 FILLER_72_1815 ();
 b15zdnd11an1n64x5 FILLER_72_1879 ();
 b15zdnd11an1n64x5 FILLER_72_1943 ();
 b15zdnd11an1n64x5 FILLER_72_2007 ();
 b15zdnd11an1n64x5 FILLER_72_2071 ();
 b15zdnd11an1n16x5 FILLER_72_2135 ();
 b15zdnd00an1n02x5 FILLER_72_2151 ();
 b15zdnd00an1n01x5 FILLER_72_2153 ();
 b15zdnd11an1n64x5 FILLER_72_2162 ();
 b15zdnd11an1n32x5 FILLER_72_2226 ();
 b15zdnd11an1n16x5 FILLER_72_2258 ();
 b15zdnd00an1n02x5 FILLER_72_2274 ();
 b15zdnd11an1n16x5 FILLER_73_0 ();
 b15zdnd00an1n01x5 FILLER_73_16 ();
 b15zdnd11an1n04x5 FILLER_73_20 ();
 b15zdnd11an1n04x5 FILLER_73_27 ();
 b15zdnd11an1n04x5 FILLER_73_34 ();
 b15zdnd11an1n64x5 FILLER_73_41 ();
 b15zdnd11an1n64x5 FILLER_73_105 ();
 b15zdnd11an1n64x5 FILLER_73_169 ();
 b15zdnd11an1n64x5 FILLER_73_233 ();
 b15zdnd11an1n64x5 FILLER_73_297 ();
 b15zdnd11an1n64x5 FILLER_73_361 ();
 b15zdnd11an1n08x5 FILLER_73_425 ();
 b15zdnd11an1n04x5 FILLER_73_433 ();
 b15zdnd00an1n02x5 FILLER_73_437 ();
 b15zdnd00an1n01x5 FILLER_73_439 ();
 b15zdnd11an1n64x5 FILLER_73_460 ();
 b15zdnd11an1n32x5 FILLER_73_524 ();
 b15zdnd11an1n16x5 FILLER_73_556 ();
 b15zdnd11an1n08x5 FILLER_73_572 ();
 b15zdnd00an1n01x5 FILLER_73_580 ();
 b15zdnd11an1n16x5 FILLER_73_598 ();
 b15zdnd11an1n04x5 FILLER_73_614 ();
 b15zdnd11an1n16x5 FILLER_73_638 ();
 b15zdnd11an1n04x5 FILLER_73_654 ();
 b15zdnd11an1n64x5 FILLER_73_678 ();
 b15zdnd11an1n64x5 FILLER_73_742 ();
 b15zdnd11an1n64x5 FILLER_73_806 ();
 b15zdnd11an1n32x5 FILLER_73_870 ();
 b15zdnd11an1n64x5 FILLER_73_905 ();
 b15zdnd11an1n64x5 FILLER_73_969 ();
 b15zdnd11an1n64x5 FILLER_73_1033 ();
 b15zdnd11an1n08x5 FILLER_73_1097 ();
 b15zdnd11an1n04x5 FILLER_73_1105 ();
 b15zdnd00an1n02x5 FILLER_73_1109 ();
 b15zdnd11an1n04x5 FILLER_73_1153 ();
 b15zdnd11an1n16x5 FILLER_73_1199 ();
 b15zdnd00an1n01x5 FILLER_73_1215 ();
 b15zdnd11an1n64x5 FILLER_73_1224 ();
 b15zdnd11an1n64x5 FILLER_73_1288 ();
 b15zdnd11an1n64x5 FILLER_73_1352 ();
 b15zdnd11an1n64x5 FILLER_73_1416 ();
 b15zdnd11an1n64x5 FILLER_73_1480 ();
 b15zdnd11an1n64x5 FILLER_73_1544 ();
 b15zdnd11an1n64x5 FILLER_73_1608 ();
 b15zdnd11an1n64x5 FILLER_73_1672 ();
 b15zdnd11an1n04x5 FILLER_73_1736 ();
 b15zdnd00an1n01x5 FILLER_73_1740 ();
 b15zdnd11an1n64x5 FILLER_73_1753 ();
 b15zdnd11an1n64x5 FILLER_73_1817 ();
 b15zdnd11an1n64x5 FILLER_73_1881 ();
 b15zdnd11an1n08x5 FILLER_73_1945 ();
 b15zdnd11an1n04x5 FILLER_73_1953 ();
 b15zdnd00an1n02x5 FILLER_73_1957 ();
 b15zdnd00an1n01x5 FILLER_73_1959 ();
 b15zdnd11an1n32x5 FILLER_73_1969 ();
 b15zdnd11an1n08x5 FILLER_73_2001 ();
 b15zdnd11an1n04x5 FILLER_73_2009 ();
 b15zdnd00an1n02x5 FILLER_73_2013 ();
 b15zdnd00an1n01x5 FILLER_73_2015 ();
 b15zdnd11an1n64x5 FILLER_73_2025 ();
 b15zdnd11an1n64x5 FILLER_73_2089 ();
 b15zdnd11an1n64x5 FILLER_73_2153 ();
 b15zdnd11an1n64x5 FILLER_73_2217 ();
 b15zdnd00an1n02x5 FILLER_73_2281 ();
 b15zdnd00an1n01x5 FILLER_73_2283 ();
 b15zdnd11an1n16x5 FILLER_74_8 ();
 b15zdnd00an1n02x5 FILLER_74_24 ();
 b15zdnd11an1n64x5 FILLER_74_29 ();
 b15zdnd11an1n64x5 FILLER_74_93 ();
 b15zdnd11an1n64x5 FILLER_74_157 ();
 b15zdnd11an1n64x5 FILLER_74_221 ();
 b15zdnd11an1n64x5 FILLER_74_285 ();
 b15zdnd11an1n64x5 FILLER_74_349 ();
 b15zdnd11an1n64x5 FILLER_74_413 ();
 b15zdnd11an1n64x5 FILLER_74_477 ();
 b15zdnd11an1n64x5 FILLER_74_541 ();
 b15zdnd11an1n16x5 FILLER_74_605 ();
 b15zdnd11an1n08x5 FILLER_74_621 ();
 b15zdnd00an1n02x5 FILLER_74_629 ();
 b15zdnd00an1n01x5 FILLER_74_631 ();
 b15zdnd11an1n04x5 FILLER_74_649 ();
 b15zdnd00an1n02x5 FILLER_74_653 ();
 b15zdnd11an1n32x5 FILLER_74_675 ();
 b15zdnd11an1n08x5 FILLER_74_707 ();
 b15zdnd00an1n02x5 FILLER_74_715 ();
 b15zdnd00an1n01x5 FILLER_74_717 ();
 b15zdnd11an1n64x5 FILLER_74_726 ();
 b15zdnd11an1n04x5 FILLER_74_790 ();
 b15zdnd00an1n02x5 FILLER_74_794 ();
 b15zdnd00an1n01x5 FILLER_74_796 ();
 b15zdnd11an1n16x5 FILLER_74_811 ();
 b15zdnd11an1n08x5 FILLER_74_827 ();
 b15zdnd00an1n01x5 FILLER_74_835 ();
 b15zdnd11an1n16x5 FILLER_74_850 ();
 b15zdnd11an1n08x5 FILLER_74_866 ();
 b15zdnd00an1n01x5 FILLER_74_874 ();
 b15zdnd11an1n64x5 FILLER_74_927 ();
 b15zdnd11an1n64x5 FILLER_74_991 ();
 b15zdnd11an1n32x5 FILLER_74_1055 ();
 b15zdnd11an1n08x5 FILLER_74_1087 ();
 b15zdnd00an1n01x5 FILLER_74_1095 ();
 b15zdnd11an1n08x5 FILLER_74_1138 ();
 b15zdnd00an1n02x5 FILLER_74_1146 ();
 b15zdnd00an1n01x5 FILLER_74_1148 ();
 b15zdnd11an1n64x5 FILLER_74_1191 ();
 b15zdnd11an1n64x5 FILLER_74_1255 ();
 b15zdnd11an1n64x5 FILLER_74_1319 ();
 b15zdnd11an1n32x5 FILLER_74_1383 ();
 b15zdnd11an1n16x5 FILLER_74_1415 ();
 b15zdnd00an1n01x5 FILLER_74_1431 ();
 b15zdnd11an1n64x5 FILLER_74_1452 ();
 b15zdnd11an1n64x5 FILLER_74_1516 ();
 b15zdnd11an1n64x5 FILLER_74_1580 ();
 b15zdnd11an1n64x5 FILLER_74_1644 ();
 b15zdnd11an1n32x5 FILLER_74_1708 ();
 b15zdnd11an1n04x5 FILLER_74_1740 ();
 b15zdnd00an1n01x5 FILLER_74_1744 ();
 b15zdnd11an1n64x5 FILLER_74_1765 ();
 b15zdnd11an1n64x5 FILLER_74_1829 ();
 b15zdnd11an1n64x5 FILLER_74_1893 ();
 b15zdnd11an1n32x5 FILLER_74_1957 ();
 b15zdnd11an1n08x5 FILLER_74_1989 ();
 b15zdnd11an1n04x5 FILLER_74_1997 ();
 b15zdnd00an1n01x5 FILLER_74_2001 ();
 b15zdnd11an1n64x5 FILLER_74_2011 ();
 b15zdnd11an1n64x5 FILLER_74_2075 ();
 b15zdnd11an1n08x5 FILLER_74_2139 ();
 b15zdnd11an1n04x5 FILLER_74_2147 ();
 b15zdnd00an1n02x5 FILLER_74_2151 ();
 b15zdnd00an1n01x5 FILLER_74_2153 ();
 b15zdnd11an1n64x5 FILLER_74_2162 ();
 b15zdnd11an1n32x5 FILLER_74_2226 ();
 b15zdnd11an1n16x5 FILLER_74_2258 ();
 b15zdnd00an1n02x5 FILLER_74_2274 ();
 b15zdnd11an1n16x5 FILLER_75_0 ();
 b15zdnd11an1n04x5 FILLER_75_16 ();
 b15zdnd00an1n01x5 FILLER_75_20 ();
 b15zdnd11an1n64x5 FILLER_75_24 ();
 b15zdnd11an1n64x5 FILLER_75_88 ();
 b15zdnd11an1n64x5 FILLER_75_152 ();
 b15zdnd11an1n64x5 FILLER_75_216 ();
 b15zdnd11an1n64x5 FILLER_75_280 ();
 b15zdnd11an1n64x5 FILLER_75_344 ();
 b15zdnd11an1n64x5 FILLER_75_408 ();
 b15zdnd11an1n64x5 FILLER_75_472 ();
 b15zdnd11an1n64x5 FILLER_75_536 ();
 b15zdnd11an1n16x5 FILLER_75_600 ();
 b15zdnd11an1n04x5 FILLER_75_616 ();
 b15zdnd00an1n02x5 FILLER_75_620 ();
 b15zdnd00an1n01x5 FILLER_75_622 ();
 b15zdnd11an1n32x5 FILLER_75_635 ();
 b15zdnd11an1n08x5 FILLER_75_667 ();
 b15zdnd11an1n04x5 FILLER_75_675 ();
 b15zdnd00an1n02x5 FILLER_75_679 ();
 b15zdnd11an1n04x5 FILLER_75_695 ();
 b15zdnd11an1n16x5 FILLER_75_711 ();
 b15zdnd11an1n08x5 FILLER_75_727 ();
 b15zdnd00an1n01x5 FILLER_75_735 ();
 b15zdnd11an1n64x5 FILLER_75_756 ();
 b15zdnd11an1n64x5 FILLER_75_820 ();
 b15zdnd11an1n16x5 FILLER_75_884 ();
 b15zdnd11an1n04x5 FILLER_75_900 ();
 b15zdnd00an1n02x5 FILLER_75_904 ();
 b15zdnd11an1n04x5 FILLER_75_909 ();
 b15zdnd11an1n32x5 FILLER_75_916 ();
 b15zdnd11an1n16x5 FILLER_75_948 ();
 b15zdnd11an1n08x5 FILLER_75_964 ();
 b15zdnd00an1n02x5 FILLER_75_972 ();
 b15zdnd11an1n32x5 FILLER_75_977 ();
 b15zdnd11an1n16x5 FILLER_75_1009 ();
 b15zdnd11an1n04x5 FILLER_75_1025 ();
 b15zdnd00an1n01x5 FILLER_75_1029 ();
 b15zdnd11an1n08x5 FILLER_75_1041 ();
 b15zdnd00an1n01x5 FILLER_75_1049 ();
 b15zdnd11an1n64x5 FILLER_75_1053 ();
 b15zdnd11an1n32x5 FILLER_75_1117 ();
 b15zdnd11an1n08x5 FILLER_75_1149 ();
 b15zdnd00an1n01x5 FILLER_75_1157 ();
 b15zdnd11an1n64x5 FILLER_75_1178 ();
 b15zdnd11an1n64x5 FILLER_75_1242 ();
 b15zdnd11an1n08x5 FILLER_75_1306 ();
 b15zdnd11an1n04x5 FILLER_75_1346 ();
 b15zdnd11an1n64x5 FILLER_75_1353 ();
 b15zdnd11an1n08x5 FILLER_75_1417 ();
 b15zdnd11an1n64x5 FILLER_75_1451 ();
 b15zdnd11an1n64x5 FILLER_75_1515 ();
 b15zdnd11an1n64x5 FILLER_75_1579 ();
 b15zdnd11an1n64x5 FILLER_75_1643 ();
 b15zdnd11an1n32x5 FILLER_75_1707 ();
 b15zdnd11an1n16x5 FILLER_75_1739 ();
 b15zdnd11an1n08x5 FILLER_75_1755 ();
 b15zdnd11an1n04x5 FILLER_75_1763 ();
 b15zdnd11an1n64x5 FILLER_75_1787 ();
 b15zdnd11an1n08x5 FILLER_75_1851 ();
 b15zdnd11an1n04x5 FILLER_75_1859 ();
 b15zdnd00an1n02x5 FILLER_75_1863 ();
 b15zdnd00an1n01x5 FILLER_75_1865 ();
 b15zdnd11an1n64x5 FILLER_75_1883 ();
 b15zdnd11an1n64x5 FILLER_75_1947 ();
 b15zdnd11an1n64x5 FILLER_75_2011 ();
 b15zdnd11an1n64x5 FILLER_75_2075 ();
 b15zdnd11an1n64x5 FILLER_75_2139 ();
 b15zdnd11an1n64x5 FILLER_75_2203 ();
 b15zdnd11an1n16x5 FILLER_75_2267 ();
 b15zdnd00an1n01x5 FILLER_75_2283 ();
 b15zdnd11an1n16x5 FILLER_76_8 ();
 b15zdnd00an1n02x5 FILLER_76_24 ();
 b15zdnd00an1n01x5 FILLER_76_26 ();
 b15zdnd11an1n64x5 FILLER_76_30 ();
 b15zdnd11an1n64x5 FILLER_76_94 ();
 b15zdnd11an1n64x5 FILLER_76_158 ();
 b15zdnd11an1n64x5 FILLER_76_222 ();
 b15zdnd11an1n64x5 FILLER_76_286 ();
 b15zdnd11an1n32x5 FILLER_76_350 ();
 b15zdnd11an1n64x5 FILLER_76_402 ();
 b15zdnd11an1n64x5 FILLER_76_466 ();
 b15zdnd11an1n64x5 FILLER_76_530 ();
 b15zdnd11an1n64x5 FILLER_76_594 ();
 b15zdnd11an1n16x5 FILLER_76_658 ();
 b15zdnd11an1n04x5 FILLER_76_674 ();
 b15zdnd11an1n16x5 FILLER_76_698 ();
 b15zdnd11an1n04x5 FILLER_76_714 ();
 b15zdnd11an1n64x5 FILLER_76_726 ();
 b15zdnd11an1n64x5 FILLER_76_790 ();
 b15zdnd11an1n64x5 FILLER_76_854 ();
 b15zdnd11an1n32x5 FILLER_76_918 ();
 b15zdnd11an1n08x5 FILLER_76_950 ();
 b15zdnd11an1n04x5 FILLER_76_969 ();
 b15zdnd11an1n16x5 FILLER_76_976 ();
 b15zdnd11an1n04x5 FILLER_76_992 ();
 b15zdnd00an1n01x5 FILLER_76_996 ();
 b15zdnd11an1n04x5 FILLER_76_1000 ();
 b15zdnd11an1n16x5 FILLER_76_1031 ();
 b15zdnd00an1n02x5 FILLER_76_1047 ();
 b15zdnd00an1n01x5 FILLER_76_1049 ();
 b15zdnd11an1n16x5 FILLER_76_1053 ();
 b15zdnd11an1n04x5 FILLER_76_1069 ();
 b15zdnd11an1n64x5 FILLER_76_1097 ();
 b15zdnd11an1n64x5 FILLER_76_1161 ();
 b15zdnd11an1n64x5 FILLER_76_1225 ();
 b15zdnd11an1n32x5 FILLER_76_1289 ();
 b15zdnd11an1n16x5 FILLER_76_1321 ();
 b15zdnd11an1n04x5 FILLER_76_1337 ();
 b15zdnd11an1n64x5 FILLER_76_1344 ();
 b15zdnd11an1n64x5 FILLER_76_1408 ();
 b15zdnd11an1n64x5 FILLER_76_1472 ();
 b15zdnd11an1n64x5 FILLER_76_1536 ();
 b15zdnd11an1n64x5 FILLER_76_1600 ();
 b15zdnd11an1n04x5 FILLER_76_1664 ();
 b15zdnd00an1n02x5 FILLER_76_1668 ();
 b15zdnd00an1n01x5 FILLER_76_1670 ();
 b15zdnd11an1n64x5 FILLER_76_1688 ();
 b15zdnd11an1n16x5 FILLER_76_1752 ();
 b15zdnd11an1n08x5 FILLER_76_1768 ();
 b15zdnd00an1n02x5 FILLER_76_1776 ();
 b15zdnd11an1n16x5 FILLER_76_1790 ();
 b15zdnd11an1n04x5 FILLER_76_1806 ();
 b15zdnd00an1n02x5 FILLER_76_1810 ();
 b15zdnd11an1n64x5 FILLER_76_1829 ();
 b15zdnd11an1n64x5 FILLER_76_1893 ();
 b15zdnd11an1n64x5 FILLER_76_1957 ();
 b15zdnd11an1n64x5 FILLER_76_2021 ();
 b15zdnd11an1n64x5 FILLER_76_2085 ();
 b15zdnd11an1n04x5 FILLER_76_2149 ();
 b15zdnd00an1n01x5 FILLER_76_2153 ();
 b15zdnd11an1n64x5 FILLER_76_2162 ();
 b15zdnd11an1n32x5 FILLER_76_2226 ();
 b15zdnd11an1n16x5 FILLER_76_2258 ();
 b15zdnd00an1n02x5 FILLER_76_2274 ();
 b15zdnd11an1n64x5 FILLER_77_0 ();
 b15zdnd11an1n64x5 FILLER_77_64 ();
 b15zdnd11an1n64x5 FILLER_77_128 ();
 b15zdnd11an1n64x5 FILLER_77_192 ();
 b15zdnd11an1n64x5 FILLER_77_256 ();
 b15zdnd11an1n64x5 FILLER_77_320 ();
 b15zdnd11an1n64x5 FILLER_77_384 ();
 b15zdnd11an1n64x5 FILLER_77_448 ();
 b15zdnd11an1n08x5 FILLER_77_512 ();
 b15zdnd11an1n64x5 FILLER_77_537 ();
 b15zdnd11an1n64x5 FILLER_77_601 ();
 b15zdnd11an1n64x5 FILLER_77_665 ();
 b15zdnd11an1n64x5 FILLER_77_729 ();
 b15zdnd11an1n64x5 FILLER_77_793 ();
 b15zdnd11an1n64x5 FILLER_77_857 ();
 b15zdnd11an1n16x5 FILLER_77_921 ();
 b15zdnd11an1n08x5 FILLER_77_937 ();
 b15zdnd11an1n04x5 FILLER_77_945 ();
 b15zdnd00an1n01x5 FILLER_77_949 ();
 b15zdnd11an1n16x5 FILLER_77_1002 ();
 b15zdnd11an1n08x5 FILLER_77_1018 ();
 b15zdnd00an1n01x5 FILLER_77_1026 ();
 b15zdnd11an1n32x5 FILLER_77_1079 ();
 b15zdnd11an1n08x5 FILLER_77_1111 ();
 b15zdnd11an1n04x5 FILLER_77_1119 ();
 b15zdnd00an1n02x5 FILLER_77_1123 ();
 b15zdnd11an1n64x5 FILLER_77_1141 ();
 b15zdnd11an1n64x5 FILLER_77_1205 ();
 b15zdnd11an1n64x5 FILLER_77_1269 ();
 b15zdnd11an1n64x5 FILLER_77_1333 ();
 b15zdnd11an1n64x5 FILLER_77_1397 ();
 b15zdnd11an1n64x5 FILLER_77_1461 ();
 b15zdnd11an1n64x5 FILLER_77_1525 ();
 b15zdnd11an1n64x5 FILLER_77_1589 ();
 b15zdnd11an1n16x5 FILLER_77_1653 ();
 b15zdnd00an1n02x5 FILLER_77_1669 ();
 b15zdnd00an1n01x5 FILLER_77_1671 ();
 b15zdnd11an1n64x5 FILLER_77_1686 ();
 b15zdnd11an1n08x5 FILLER_77_1750 ();
 b15zdnd11an1n04x5 FILLER_77_1758 ();
 b15zdnd00an1n01x5 FILLER_77_1762 ();
 b15zdnd11an1n08x5 FILLER_77_1775 ();
 b15zdnd11an1n04x5 FILLER_77_1783 ();
 b15zdnd00an1n01x5 FILLER_77_1787 ();
 b15zdnd11an1n64x5 FILLER_77_1802 ();
 b15zdnd11an1n64x5 FILLER_77_1866 ();
 b15zdnd11an1n64x5 FILLER_77_1930 ();
 b15zdnd11an1n64x5 FILLER_77_1994 ();
 b15zdnd00an1n02x5 FILLER_77_2058 ();
 b15zdnd00an1n01x5 FILLER_77_2060 ();
 b15zdnd11an1n04x5 FILLER_77_2064 ();
 b15zdnd11an1n64x5 FILLER_77_2071 ();
 b15zdnd11an1n64x5 FILLER_77_2135 ();
 b15zdnd11an1n64x5 FILLER_77_2199 ();
 b15zdnd11an1n16x5 FILLER_77_2263 ();
 b15zdnd11an1n04x5 FILLER_77_2279 ();
 b15zdnd00an1n01x5 FILLER_77_2283 ();
 b15zdnd11an1n08x5 FILLER_78_8 ();
 b15zdnd11an1n04x5 FILLER_78_16 ();
 b15zdnd00an1n02x5 FILLER_78_20 ();
 b15zdnd11an1n04x5 FILLER_78_25 ();
 b15zdnd11an1n04x5 FILLER_78_32 ();
 b15zdnd11an1n64x5 FILLER_78_39 ();
 b15zdnd11an1n64x5 FILLER_78_103 ();
 b15zdnd11an1n64x5 FILLER_78_167 ();
 b15zdnd11an1n64x5 FILLER_78_231 ();
 b15zdnd11an1n64x5 FILLER_78_295 ();
 b15zdnd11an1n32x5 FILLER_78_359 ();
 b15zdnd11an1n04x5 FILLER_78_391 ();
 b15zdnd11an1n64x5 FILLER_78_415 ();
 b15zdnd11an1n64x5 FILLER_78_479 ();
 b15zdnd11an1n64x5 FILLER_78_543 ();
 b15zdnd11an1n64x5 FILLER_78_607 ();
 b15zdnd11an1n32x5 FILLER_78_671 ();
 b15zdnd11an1n08x5 FILLER_78_703 ();
 b15zdnd11an1n04x5 FILLER_78_711 ();
 b15zdnd00an1n02x5 FILLER_78_715 ();
 b15zdnd00an1n01x5 FILLER_78_717 ();
 b15zdnd11an1n64x5 FILLER_78_726 ();
 b15zdnd11an1n64x5 FILLER_78_790 ();
 b15zdnd11an1n64x5 FILLER_78_854 ();
 b15zdnd11an1n32x5 FILLER_78_918 ();
 b15zdnd00an1n02x5 FILLER_78_950 ();
 b15zdnd11an1n08x5 FILLER_78_963 ();
 b15zdnd11an1n04x5 FILLER_78_971 ();
 b15zdnd00an1n01x5 FILLER_78_975 ();
 b15zdnd11an1n32x5 FILLER_78_979 ();
 b15zdnd11an1n16x5 FILLER_78_1011 ();
 b15zdnd11an1n04x5 FILLER_78_1027 ();
 b15zdnd00an1n01x5 FILLER_78_1031 ();
 b15zdnd11an1n08x5 FILLER_78_1043 ();
 b15zdnd11an1n04x5 FILLER_78_1051 ();
 b15zdnd11an1n64x5 FILLER_78_1058 ();
 b15zdnd11an1n64x5 FILLER_78_1122 ();
 b15zdnd11an1n64x5 FILLER_78_1186 ();
 b15zdnd11an1n64x5 FILLER_78_1250 ();
 b15zdnd11an1n64x5 FILLER_78_1314 ();
 b15zdnd11an1n64x5 FILLER_78_1378 ();
 b15zdnd11an1n32x5 FILLER_78_1442 ();
 b15zdnd11an1n16x5 FILLER_78_1474 ();
 b15zdnd11an1n04x5 FILLER_78_1490 ();
 b15zdnd00an1n01x5 FILLER_78_1494 ();
 b15zdnd11an1n64x5 FILLER_78_1498 ();
 b15zdnd11an1n64x5 FILLER_78_1562 ();
 b15zdnd11an1n32x5 FILLER_78_1626 ();
 b15zdnd11an1n08x5 FILLER_78_1658 ();
 b15zdnd11an1n64x5 FILLER_78_1686 ();
 b15zdnd11an1n64x5 FILLER_78_1750 ();
 b15zdnd11an1n08x5 FILLER_78_1814 ();
 b15zdnd11an1n04x5 FILLER_78_1822 ();
 b15zdnd00an1n02x5 FILLER_78_1826 ();
 b15zdnd00an1n01x5 FILLER_78_1828 ();
 b15zdnd11an1n64x5 FILLER_78_1849 ();
 b15zdnd11an1n08x5 FILLER_78_1913 ();
 b15zdnd00an1n02x5 FILLER_78_1921 ();
 b15zdnd11an1n64x5 FILLER_78_1926 ();
 b15zdnd11an1n32x5 FILLER_78_1990 ();
 b15zdnd11an1n16x5 FILLER_78_2022 ();
 b15zdnd11an1n04x5 FILLER_78_2038 ();
 b15zdnd00an1n01x5 FILLER_78_2042 ();
 b15zdnd11an1n32x5 FILLER_78_2095 ();
 b15zdnd11an1n16x5 FILLER_78_2127 ();
 b15zdnd11an1n08x5 FILLER_78_2143 ();
 b15zdnd00an1n02x5 FILLER_78_2151 ();
 b15zdnd00an1n01x5 FILLER_78_2153 ();
 b15zdnd11an1n64x5 FILLER_78_2162 ();
 b15zdnd11an1n32x5 FILLER_78_2226 ();
 b15zdnd11an1n16x5 FILLER_78_2258 ();
 b15zdnd00an1n02x5 FILLER_78_2274 ();
 b15zdnd11an1n32x5 FILLER_79_0 ();
 b15zdnd11an1n04x5 FILLER_79_32 ();
 b15zdnd11an1n64x5 FILLER_79_39 ();
 b15zdnd11an1n64x5 FILLER_79_103 ();
 b15zdnd11an1n64x5 FILLER_79_167 ();
 b15zdnd11an1n64x5 FILLER_79_231 ();
 b15zdnd11an1n64x5 FILLER_79_295 ();
 b15zdnd11an1n64x5 FILLER_79_359 ();
 b15zdnd11an1n64x5 FILLER_79_423 ();
 b15zdnd11an1n64x5 FILLER_79_487 ();
 b15zdnd11an1n64x5 FILLER_79_551 ();
 b15zdnd11an1n64x5 FILLER_79_615 ();
 b15zdnd11an1n32x5 FILLER_79_702 ();
 b15zdnd11an1n04x5 FILLER_79_734 ();
 b15zdnd11an1n32x5 FILLER_79_752 ();
 b15zdnd11an1n08x5 FILLER_79_784 ();
 b15zdnd00an1n02x5 FILLER_79_792 ();
 b15zdnd00an1n01x5 FILLER_79_794 ();
 b15zdnd11an1n64x5 FILLER_79_809 ();
 b15zdnd11an1n64x5 FILLER_79_873 ();
 b15zdnd11an1n64x5 FILLER_79_937 ();
 b15zdnd11an1n64x5 FILLER_79_1001 ();
 b15zdnd11an1n64x5 FILLER_79_1065 ();
 b15zdnd11an1n64x5 FILLER_79_1129 ();
 b15zdnd11an1n64x5 FILLER_79_1193 ();
 b15zdnd11an1n64x5 FILLER_79_1257 ();
 b15zdnd11an1n64x5 FILLER_79_1321 ();
 b15zdnd11an1n64x5 FILLER_79_1385 ();
 b15zdnd11an1n16x5 FILLER_79_1449 ();
 b15zdnd11an1n04x5 FILLER_79_1465 ();
 b15zdnd11an1n64x5 FILLER_79_1521 ();
 b15zdnd11an1n64x5 FILLER_79_1585 ();
 b15zdnd11an1n08x5 FILLER_79_1649 ();
 b15zdnd11an1n04x5 FILLER_79_1657 ();
 b15zdnd00an1n02x5 FILLER_79_1661 ();
 b15zdnd11an1n08x5 FILLER_79_1675 ();
 b15zdnd00an1n02x5 FILLER_79_1683 ();
 b15zdnd00an1n01x5 FILLER_79_1685 ();
 b15zdnd11an1n64x5 FILLER_79_1706 ();
 b15zdnd11an1n64x5 FILLER_79_1770 ();
 b15zdnd11an1n32x5 FILLER_79_1834 ();
 b15zdnd11an1n16x5 FILLER_79_1866 ();
 b15zdnd11an1n08x5 FILLER_79_1882 ();
 b15zdnd11an1n04x5 FILLER_79_1890 ();
 b15zdnd00an1n02x5 FILLER_79_1894 ();
 b15zdnd00an1n01x5 FILLER_79_1896 ();
 b15zdnd11an1n64x5 FILLER_79_1949 ();
 b15zdnd11an1n32x5 FILLER_79_2013 ();
 b15zdnd11an1n16x5 FILLER_79_2045 ();
 b15zdnd11an1n04x5 FILLER_79_2061 ();
 b15zdnd00an1n02x5 FILLER_79_2065 ();
 b15zdnd00an1n01x5 FILLER_79_2067 ();
 b15zdnd11an1n64x5 FILLER_79_2071 ();
 b15zdnd11an1n64x5 FILLER_79_2135 ();
 b15zdnd11an1n64x5 FILLER_79_2199 ();
 b15zdnd11an1n16x5 FILLER_79_2263 ();
 b15zdnd11an1n04x5 FILLER_79_2279 ();
 b15zdnd00an1n01x5 FILLER_79_2283 ();
 b15zdnd11an1n04x5 FILLER_80_8 ();
 b15zdnd00an1n02x5 FILLER_80_12 ();
 b15zdnd00an1n01x5 FILLER_80_14 ();
 b15zdnd11an1n04x5 FILLER_80_18 ();
 b15zdnd11an1n64x5 FILLER_80_25 ();
 b15zdnd11an1n64x5 FILLER_80_89 ();
 b15zdnd11an1n64x5 FILLER_80_153 ();
 b15zdnd11an1n64x5 FILLER_80_217 ();
 b15zdnd11an1n64x5 FILLER_80_281 ();
 b15zdnd11an1n64x5 FILLER_80_345 ();
 b15zdnd11an1n64x5 FILLER_80_409 ();
 b15zdnd11an1n64x5 FILLER_80_473 ();
 b15zdnd11an1n32x5 FILLER_80_537 ();
 b15zdnd11an1n04x5 FILLER_80_569 ();
 b15zdnd00an1n02x5 FILLER_80_573 ();
 b15zdnd11an1n64x5 FILLER_80_595 ();
 b15zdnd11an1n32x5 FILLER_80_659 ();
 b15zdnd11an1n16x5 FILLER_80_691 ();
 b15zdnd11an1n08x5 FILLER_80_707 ();
 b15zdnd00an1n02x5 FILLER_80_715 ();
 b15zdnd00an1n01x5 FILLER_80_717 ();
 b15zdnd11an1n64x5 FILLER_80_726 ();
 b15zdnd11an1n64x5 FILLER_80_790 ();
 b15zdnd11an1n64x5 FILLER_80_854 ();
 b15zdnd11an1n64x5 FILLER_80_918 ();
 b15zdnd11an1n64x5 FILLER_80_982 ();
 b15zdnd11an1n32x5 FILLER_80_1046 ();
 b15zdnd11an1n08x5 FILLER_80_1078 ();
 b15zdnd11an1n04x5 FILLER_80_1086 ();
 b15zdnd00an1n02x5 FILLER_80_1090 ();
 b15zdnd00an1n01x5 FILLER_80_1092 ();
 b15zdnd11an1n04x5 FILLER_80_1096 ();
 b15zdnd11an1n04x5 FILLER_80_1103 ();
 b15zdnd11an1n64x5 FILLER_80_1110 ();
 b15zdnd11an1n64x5 FILLER_80_1174 ();
 b15zdnd11an1n64x5 FILLER_80_1238 ();
 b15zdnd11an1n64x5 FILLER_80_1302 ();
 b15zdnd11an1n64x5 FILLER_80_1366 ();
 b15zdnd11an1n32x5 FILLER_80_1430 ();
 b15zdnd11an1n16x5 FILLER_80_1462 ();
 b15zdnd11an1n08x5 FILLER_80_1478 ();
 b15zdnd00an1n02x5 FILLER_80_1486 ();
 b15zdnd00an1n01x5 FILLER_80_1488 ();
 b15zdnd11an1n04x5 FILLER_80_1492 ();
 b15zdnd11an1n64x5 FILLER_80_1499 ();
 b15zdnd11an1n16x5 FILLER_80_1563 ();
 b15zdnd00an1n01x5 FILLER_80_1579 ();
 b15zdnd11an1n64x5 FILLER_80_1583 ();
 b15zdnd11an1n64x5 FILLER_80_1647 ();
 b15zdnd11an1n64x5 FILLER_80_1711 ();
 b15zdnd11an1n64x5 FILLER_80_1775 ();
 b15zdnd11an1n64x5 FILLER_80_1839 ();
 b15zdnd11an1n16x5 FILLER_80_1903 ();
 b15zdnd00an1n02x5 FILLER_80_1919 ();
 b15zdnd00an1n01x5 FILLER_80_1921 ();
 b15zdnd11an1n04x5 FILLER_80_1925 ();
 b15zdnd11an1n04x5 FILLER_80_1932 ();
 b15zdnd11an1n04x5 FILLER_80_1939 ();
 b15zdnd00an1n01x5 FILLER_80_1943 ();
 b15zdnd11an1n64x5 FILLER_80_1947 ();
 b15zdnd11an1n32x5 FILLER_80_2011 ();
 b15zdnd11an1n16x5 FILLER_80_2043 ();
 b15zdnd00an1n02x5 FILLER_80_2059 ();
 b15zdnd11an1n04x5 FILLER_80_2064 ();
 b15zdnd11an1n64x5 FILLER_80_2071 ();
 b15zdnd11an1n16x5 FILLER_80_2135 ();
 b15zdnd00an1n02x5 FILLER_80_2151 ();
 b15zdnd00an1n01x5 FILLER_80_2153 ();
 b15zdnd11an1n64x5 FILLER_80_2162 ();
 b15zdnd11an1n32x5 FILLER_80_2226 ();
 b15zdnd11an1n16x5 FILLER_80_2258 ();
 b15zdnd00an1n02x5 FILLER_80_2274 ();
 b15zdnd11an1n16x5 FILLER_81_0 ();
 b15zdnd11an1n04x5 FILLER_81_16 ();
 b15zdnd11an1n04x5 FILLER_81_23 ();
 b15zdnd11an1n04x5 FILLER_81_30 ();
 b15zdnd11an1n64x5 FILLER_81_37 ();
 b15zdnd11an1n64x5 FILLER_81_101 ();
 b15zdnd11an1n64x5 FILLER_81_165 ();
 b15zdnd11an1n64x5 FILLER_81_229 ();
 b15zdnd11an1n64x5 FILLER_81_293 ();
 b15zdnd11an1n64x5 FILLER_81_357 ();
 b15zdnd11an1n64x5 FILLER_81_421 ();
 b15zdnd11an1n64x5 FILLER_81_485 ();
 b15zdnd11an1n64x5 FILLER_81_549 ();
 b15zdnd11an1n64x5 FILLER_81_613 ();
 b15zdnd11an1n64x5 FILLER_81_677 ();
 b15zdnd11an1n64x5 FILLER_81_741 ();
 b15zdnd11an1n64x5 FILLER_81_805 ();
 b15zdnd11an1n64x5 FILLER_81_869 ();
 b15zdnd11an1n64x5 FILLER_81_933 ();
 b15zdnd11an1n32x5 FILLER_81_997 ();
 b15zdnd11an1n16x5 FILLER_81_1029 ();
 b15zdnd11an1n08x5 FILLER_81_1045 ();
 b15zdnd11an1n04x5 FILLER_81_1053 ();
 b15zdnd00an1n01x5 FILLER_81_1057 ();
 b15zdnd11an1n04x5 FILLER_81_1081 ();
 b15zdnd00an1n01x5 FILLER_81_1085 ();
 b15zdnd11an1n64x5 FILLER_81_1128 ();
 b15zdnd11an1n64x5 FILLER_81_1192 ();
 b15zdnd11an1n64x5 FILLER_81_1256 ();
 b15zdnd11an1n64x5 FILLER_81_1320 ();
 b15zdnd11an1n64x5 FILLER_81_1384 ();
 b15zdnd11an1n64x5 FILLER_81_1448 ();
 b15zdnd11an1n32x5 FILLER_81_1512 ();
 b15zdnd11an1n08x5 FILLER_81_1544 ();
 b15zdnd11an1n04x5 FILLER_81_1552 ();
 b15zdnd00an1n02x5 FILLER_81_1556 ();
 b15zdnd11an1n16x5 FILLER_81_1561 ();
 b15zdnd00an1n02x5 FILLER_81_1577 ();
 b15zdnd11an1n64x5 FILLER_81_1582 ();
 b15zdnd11an1n64x5 FILLER_81_1646 ();
 b15zdnd11an1n64x5 FILLER_81_1710 ();
 b15zdnd00an1n02x5 FILLER_81_1774 ();
 b15zdnd11an1n64x5 FILLER_81_1796 ();
 b15zdnd11an1n32x5 FILLER_81_1860 ();
 b15zdnd11an1n16x5 FILLER_81_1892 ();
 b15zdnd11an1n04x5 FILLER_81_1908 ();
 b15zdnd11an1n64x5 FILLER_81_1964 ();
 b15zdnd11an1n08x5 FILLER_81_2028 ();
 b15zdnd11an1n04x5 FILLER_81_2036 ();
 b15zdnd00an1n02x5 FILLER_81_2040 ();
 b15zdnd00an1n01x5 FILLER_81_2042 ();
 b15zdnd11an1n64x5 FILLER_81_2095 ();
 b15zdnd11an1n64x5 FILLER_81_2159 ();
 b15zdnd11an1n32x5 FILLER_81_2223 ();
 b15zdnd11an1n16x5 FILLER_81_2255 ();
 b15zdnd11an1n08x5 FILLER_81_2271 ();
 b15zdnd11an1n04x5 FILLER_81_2279 ();
 b15zdnd00an1n01x5 FILLER_81_2283 ();
 b15zdnd11an1n16x5 FILLER_82_8 ();
 b15zdnd00an1n01x5 FILLER_82_24 ();
 b15zdnd11an1n04x5 FILLER_82_28 ();
 b15zdnd11an1n04x5 FILLER_82_35 ();
 b15zdnd11an1n64x5 FILLER_82_42 ();
 b15zdnd11an1n64x5 FILLER_82_106 ();
 b15zdnd11an1n08x5 FILLER_82_170 ();
 b15zdnd11an1n04x5 FILLER_82_178 ();
 b15zdnd00an1n02x5 FILLER_82_182 ();
 b15zdnd11an1n64x5 FILLER_82_215 ();
 b15zdnd11an1n64x5 FILLER_82_279 ();
 b15zdnd11an1n64x5 FILLER_82_343 ();
 b15zdnd11an1n16x5 FILLER_82_407 ();
 b15zdnd11an1n08x5 FILLER_82_423 ();
 b15zdnd11an1n04x5 FILLER_82_431 ();
 b15zdnd00an1n01x5 FILLER_82_435 ();
 b15zdnd11an1n64x5 FILLER_82_450 ();
 b15zdnd11an1n64x5 FILLER_82_514 ();
 b15zdnd11an1n64x5 FILLER_82_578 ();
 b15zdnd11an1n64x5 FILLER_82_642 ();
 b15zdnd11an1n08x5 FILLER_82_706 ();
 b15zdnd11an1n04x5 FILLER_82_714 ();
 b15zdnd11an1n64x5 FILLER_82_726 ();
 b15zdnd11an1n16x5 FILLER_82_790 ();
 b15zdnd11an1n08x5 FILLER_82_806 ();
 b15zdnd00an1n01x5 FILLER_82_814 ();
 b15zdnd11an1n64x5 FILLER_82_839 ();
 b15zdnd11an1n64x5 FILLER_82_903 ();
 b15zdnd11an1n64x5 FILLER_82_967 ();
 b15zdnd11an1n32x5 FILLER_82_1031 ();
 b15zdnd11an1n04x5 FILLER_82_1063 ();
 b15zdnd00an1n02x5 FILLER_82_1067 ();
 b15zdnd00an1n01x5 FILLER_82_1069 ();
 b15zdnd11an1n64x5 FILLER_82_1122 ();
 b15zdnd11an1n64x5 FILLER_82_1186 ();
 b15zdnd11an1n08x5 FILLER_82_1250 ();
 b15zdnd00an1n02x5 FILLER_82_1258 ();
 b15zdnd00an1n01x5 FILLER_82_1260 ();
 b15zdnd11an1n04x5 FILLER_82_1264 ();
 b15zdnd00an1n02x5 FILLER_82_1268 ();
 b15zdnd00an1n01x5 FILLER_82_1270 ();
 b15zdnd11an1n08x5 FILLER_82_1274 ();
 b15zdnd11an1n04x5 FILLER_82_1282 ();
 b15zdnd00an1n02x5 FILLER_82_1286 ();
 b15zdnd11an1n64x5 FILLER_82_1330 ();
 b15zdnd11an1n64x5 FILLER_82_1394 ();
 b15zdnd11an1n64x5 FILLER_82_1458 ();
 b15zdnd11an1n08x5 FILLER_82_1522 ();
 b15zdnd00an1n02x5 FILLER_82_1530 ();
 b15zdnd00an1n01x5 FILLER_82_1532 ();
 b15zdnd11an1n04x5 FILLER_82_1585 ();
 b15zdnd11an1n64x5 FILLER_82_1592 ();
 b15zdnd11an1n64x5 FILLER_82_1656 ();
 b15zdnd11an1n64x5 FILLER_82_1720 ();
 b15zdnd11an1n16x5 FILLER_82_1784 ();
 b15zdnd11an1n04x5 FILLER_82_1800 ();
 b15zdnd00an1n02x5 FILLER_82_1804 ();
 b15zdnd00an1n01x5 FILLER_82_1806 ();
 b15zdnd11an1n64x5 FILLER_82_1819 ();
 b15zdnd11an1n32x5 FILLER_82_1883 ();
 b15zdnd11an1n16x5 FILLER_82_1915 ();
 b15zdnd11an1n04x5 FILLER_82_1931 ();
 b15zdnd00an1n02x5 FILLER_82_1935 ();
 b15zdnd00an1n01x5 FILLER_82_1937 ();
 b15zdnd11an1n16x5 FILLER_82_1941 ();
 b15zdnd11an1n08x5 FILLER_82_1957 ();
 b15zdnd00an1n01x5 FILLER_82_1965 ();
 b15zdnd11an1n64x5 FILLER_82_1986 ();
 b15zdnd11an1n16x5 FILLER_82_2050 ();
 b15zdnd00an1n02x5 FILLER_82_2066 ();
 b15zdnd11an1n64x5 FILLER_82_2071 ();
 b15zdnd11an1n16x5 FILLER_82_2135 ();
 b15zdnd00an1n02x5 FILLER_82_2151 ();
 b15zdnd00an1n01x5 FILLER_82_2153 ();
 b15zdnd11an1n64x5 FILLER_82_2162 ();
 b15zdnd11an1n32x5 FILLER_82_2226 ();
 b15zdnd11an1n16x5 FILLER_82_2258 ();
 b15zdnd00an1n02x5 FILLER_82_2274 ();
 b15zdnd11an1n64x5 FILLER_83_0 ();
 b15zdnd11an1n64x5 FILLER_83_64 ();
 b15zdnd11an1n32x5 FILLER_83_128 ();
 b15zdnd11an1n16x5 FILLER_83_160 ();
 b15zdnd11an1n08x5 FILLER_83_176 ();
 b15zdnd00an1n02x5 FILLER_83_184 ();
 b15zdnd00an1n01x5 FILLER_83_186 ();
 b15zdnd11an1n64x5 FILLER_83_218 ();
 b15zdnd11an1n64x5 FILLER_83_282 ();
 b15zdnd11an1n64x5 FILLER_83_346 ();
 b15zdnd11an1n16x5 FILLER_83_410 ();
 b15zdnd11an1n04x5 FILLER_83_426 ();
 b15zdnd00an1n02x5 FILLER_83_430 ();
 b15zdnd00an1n01x5 FILLER_83_432 ();
 b15zdnd11an1n04x5 FILLER_83_453 ();
 b15zdnd11an1n64x5 FILLER_83_477 ();
 b15zdnd11an1n64x5 FILLER_83_541 ();
 b15zdnd11an1n64x5 FILLER_83_605 ();
 b15zdnd11an1n64x5 FILLER_83_669 ();
 b15zdnd11an1n64x5 FILLER_83_733 ();
 b15zdnd11an1n64x5 FILLER_83_797 ();
 b15zdnd11an1n64x5 FILLER_83_861 ();
 b15zdnd11an1n64x5 FILLER_83_925 ();
 b15zdnd11an1n64x5 FILLER_83_989 ();
 b15zdnd11an1n64x5 FILLER_83_1053 ();
 b15zdnd11an1n32x5 FILLER_83_1117 ();
 b15zdnd11an1n16x5 FILLER_83_1149 ();
 b15zdnd00an1n02x5 FILLER_83_1165 ();
 b15zdnd00an1n01x5 FILLER_83_1167 ();
 b15zdnd11an1n32x5 FILLER_83_1184 ();
 b15zdnd11an1n16x5 FILLER_83_1216 ();
 b15zdnd11an1n08x5 FILLER_83_1232 ();
 b15zdnd11an1n04x5 FILLER_83_1240 ();
 b15zdnd00an1n02x5 FILLER_83_1244 ();
 b15zdnd11an1n32x5 FILLER_83_1298 ();
 b15zdnd11an1n08x5 FILLER_83_1330 ();
 b15zdnd11an1n04x5 FILLER_83_1338 ();
 b15zdnd00an1n01x5 FILLER_83_1342 ();
 b15zdnd11an1n64x5 FILLER_83_1385 ();
 b15zdnd11an1n64x5 FILLER_83_1449 ();
 b15zdnd11an1n32x5 FILLER_83_1513 ();
 b15zdnd11an1n04x5 FILLER_83_1545 ();
 b15zdnd00an1n01x5 FILLER_83_1549 ();
 b15zdnd11an1n04x5 FILLER_83_1553 ();
 b15zdnd11an1n64x5 FILLER_83_1609 ();
 b15zdnd11an1n32x5 FILLER_83_1673 ();
 b15zdnd11an1n08x5 FILLER_83_1705 ();
 b15zdnd00an1n02x5 FILLER_83_1713 ();
 b15zdnd11an1n64x5 FILLER_83_1732 ();
 b15zdnd11an1n16x5 FILLER_83_1796 ();
 b15zdnd00an1n02x5 FILLER_83_1812 ();
 b15zdnd11an1n64x5 FILLER_83_1828 ();
 b15zdnd11an1n64x5 FILLER_83_1892 ();
 b15zdnd11an1n64x5 FILLER_83_1956 ();
 b15zdnd11an1n16x5 FILLER_83_2020 ();
 b15zdnd11an1n04x5 FILLER_83_2036 ();
 b15zdnd00an1n02x5 FILLER_83_2040 ();
 b15zdnd11an1n04x5 FILLER_83_2045 ();
 b15zdnd00an1n02x5 FILLER_83_2049 ();
 b15zdnd11an1n64x5 FILLER_83_2054 ();
 b15zdnd11an1n64x5 FILLER_83_2118 ();
 b15zdnd11an1n64x5 FILLER_83_2182 ();
 b15zdnd11an1n32x5 FILLER_83_2246 ();
 b15zdnd11an1n04x5 FILLER_83_2278 ();
 b15zdnd00an1n02x5 FILLER_83_2282 ();
 b15zdnd11an1n16x5 FILLER_84_8 ();
 b15zdnd11an1n08x5 FILLER_84_24 ();
 b15zdnd11an1n64x5 FILLER_84_35 ();
 b15zdnd11an1n64x5 FILLER_84_99 ();
 b15zdnd11an1n64x5 FILLER_84_163 ();
 b15zdnd11an1n64x5 FILLER_84_227 ();
 b15zdnd11an1n64x5 FILLER_84_291 ();
 b15zdnd11an1n64x5 FILLER_84_355 ();
 b15zdnd11an1n64x5 FILLER_84_419 ();
 b15zdnd11an1n16x5 FILLER_84_483 ();
 b15zdnd11an1n04x5 FILLER_84_499 ();
 b15zdnd11an1n64x5 FILLER_84_506 ();
 b15zdnd11an1n64x5 FILLER_84_570 ();
 b15zdnd11an1n64x5 FILLER_84_634 ();
 b15zdnd11an1n16x5 FILLER_84_698 ();
 b15zdnd11an1n04x5 FILLER_84_714 ();
 b15zdnd11an1n64x5 FILLER_84_726 ();
 b15zdnd11an1n64x5 FILLER_84_790 ();
 b15zdnd11an1n64x5 FILLER_84_854 ();
 b15zdnd11an1n64x5 FILLER_84_918 ();
 b15zdnd11an1n64x5 FILLER_84_982 ();
 b15zdnd11an1n64x5 FILLER_84_1046 ();
 b15zdnd00an1n02x5 FILLER_84_1110 ();
 b15zdnd11an1n64x5 FILLER_84_1128 ();
 b15zdnd11an1n32x5 FILLER_84_1192 ();
 b15zdnd11an1n08x5 FILLER_84_1224 ();
 b15zdnd11an1n04x5 FILLER_84_1232 ();
 b15zdnd11an1n04x5 FILLER_84_1288 ();
 b15zdnd11an1n64x5 FILLER_84_1334 ();
 b15zdnd11an1n64x5 FILLER_84_1398 ();
 b15zdnd11an1n64x5 FILLER_84_1462 ();
 b15zdnd11an1n16x5 FILLER_84_1526 ();
 b15zdnd11an1n08x5 FILLER_84_1542 ();
 b15zdnd11an1n04x5 FILLER_84_1550 ();
 b15zdnd00an1n02x5 FILLER_84_1554 ();
 b15zdnd00an1n01x5 FILLER_84_1556 ();
 b15zdnd11an1n64x5 FILLER_84_1560 ();
 b15zdnd11an1n64x5 FILLER_84_1624 ();
 b15zdnd00an1n01x5 FILLER_84_1688 ();
 b15zdnd11an1n32x5 FILLER_84_1706 ();
 b15zdnd11an1n16x5 FILLER_84_1738 ();
 b15zdnd11an1n08x5 FILLER_84_1754 ();
 b15zdnd11an1n04x5 FILLER_84_1762 ();
 b15zdnd00an1n02x5 FILLER_84_1766 ();
 b15zdnd00an1n01x5 FILLER_84_1768 ();
 b15zdnd11an1n08x5 FILLER_84_1786 ();
 b15zdnd00an1n01x5 FILLER_84_1794 ();
 b15zdnd11an1n04x5 FILLER_84_1809 ();
 b15zdnd00an1n01x5 FILLER_84_1813 ();
 b15zdnd11an1n64x5 FILLER_84_1834 ();
 b15zdnd11an1n64x5 FILLER_84_1898 ();
 b15zdnd11an1n32x5 FILLER_84_1962 ();
 b15zdnd11an1n16x5 FILLER_84_1994 ();
 b15zdnd11an1n08x5 FILLER_84_2010 ();
 b15zdnd00an1n01x5 FILLER_84_2018 ();
 b15zdnd11an1n64x5 FILLER_84_2071 ();
 b15zdnd11an1n16x5 FILLER_84_2135 ();
 b15zdnd00an1n02x5 FILLER_84_2151 ();
 b15zdnd00an1n01x5 FILLER_84_2153 ();
 b15zdnd11an1n64x5 FILLER_84_2162 ();
 b15zdnd11an1n32x5 FILLER_84_2226 ();
 b15zdnd11an1n16x5 FILLER_84_2258 ();
 b15zdnd00an1n02x5 FILLER_84_2274 ();
 b15zdnd11an1n32x5 FILLER_85_0 ();
 b15zdnd00an1n01x5 FILLER_85_32 ();
 b15zdnd11an1n64x5 FILLER_85_36 ();
 b15zdnd11an1n64x5 FILLER_85_100 ();
 b15zdnd11an1n32x5 FILLER_85_164 ();
 b15zdnd11an1n16x5 FILLER_85_196 ();
 b15zdnd00an1n01x5 FILLER_85_212 ();
 b15zdnd11an1n64x5 FILLER_85_216 ();
 b15zdnd11an1n32x5 FILLER_85_280 ();
 b15zdnd11an1n08x5 FILLER_85_312 ();
 b15zdnd11an1n64x5 FILLER_85_372 ();
 b15zdnd11an1n08x5 FILLER_85_436 ();
 b15zdnd00an1n02x5 FILLER_85_444 ();
 b15zdnd00an1n01x5 FILLER_85_446 ();
 b15zdnd11an1n04x5 FILLER_85_473 ();
 b15zdnd11an1n64x5 FILLER_85_529 ();
 b15zdnd11an1n64x5 FILLER_85_593 ();
 b15zdnd11an1n64x5 FILLER_85_657 ();
 b15zdnd11an1n32x5 FILLER_85_721 ();
 b15zdnd11an1n64x5 FILLER_85_773 ();
 b15zdnd11an1n64x5 FILLER_85_837 ();
 b15zdnd11an1n64x5 FILLER_85_901 ();
 b15zdnd11an1n64x5 FILLER_85_965 ();
 b15zdnd11an1n08x5 FILLER_85_1029 ();
 b15zdnd00an1n02x5 FILLER_85_1037 ();
 b15zdnd11an1n04x5 FILLER_85_1081 ();
 b15zdnd11an1n64x5 FILLER_85_1127 ();
 b15zdnd11an1n32x5 FILLER_85_1191 ();
 b15zdnd11an1n16x5 FILLER_85_1223 ();
 b15zdnd11an1n04x5 FILLER_85_1245 ();
 b15zdnd00an1n02x5 FILLER_85_1249 ();
 b15zdnd00an1n01x5 FILLER_85_1251 ();
 b15zdnd11an1n64x5 FILLER_85_1294 ();
 b15zdnd11an1n64x5 FILLER_85_1358 ();
 b15zdnd11an1n64x5 FILLER_85_1422 ();
 b15zdnd11an1n64x5 FILLER_85_1486 ();
 b15zdnd11an1n64x5 FILLER_85_1550 ();
 b15zdnd11an1n64x5 FILLER_85_1614 ();
 b15zdnd11an1n64x5 FILLER_85_1678 ();
 b15zdnd11an1n08x5 FILLER_85_1742 ();
 b15zdnd11an1n04x5 FILLER_85_1750 ();
 b15zdnd00an1n01x5 FILLER_85_1754 ();
 b15zdnd11an1n16x5 FILLER_85_1769 ();
 b15zdnd11an1n04x5 FILLER_85_1785 ();
 b15zdnd00an1n02x5 FILLER_85_1789 ();
 b15zdnd11an1n64x5 FILLER_85_1811 ();
 b15zdnd11an1n32x5 FILLER_85_1875 ();
 b15zdnd11an1n04x5 FILLER_85_1907 ();
 b15zdnd00an1n01x5 FILLER_85_1911 ();
 b15zdnd11an1n64x5 FILLER_85_1932 ();
 b15zdnd11an1n32x5 FILLER_85_1996 ();
 b15zdnd11an1n08x5 FILLER_85_2028 ();
 b15zdnd11an1n04x5 FILLER_85_2036 ();
 b15zdnd00an1n02x5 FILLER_85_2040 ();
 b15zdnd00an1n01x5 FILLER_85_2042 ();
 b15zdnd11an1n64x5 FILLER_85_2046 ();
 b15zdnd11an1n64x5 FILLER_85_2110 ();
 b15zdnd11an1n64x5 FILLER_85_2174 ();
 b15zdnd11an1n32x5 FILLER_85_2238 ();
 b15zdnd11an1n08x5 FILLER_85_2270 ();
 b15zdnd11an1n04x5 FILLER_85_2278 ();
 b15zdnd00an1n02x5 FILLER_85_2282 ();
 b15zdnd11an1n16x5 FILLER_86_8 ();
 b15zdnd11an1n64x5 FILLER_86_27 ();
 b15zdnd11an1n64x5 FILLER_86_91 ();
 b15zdnd11an1n16x5 FILLER_86_155 ();
 b15zdnd11an1n08x5 FILLER_86_171 ();
 b15zdnd11an1n04x5 FILLER_86_179 ();
 b15zdnd00an1n02x5 FILLER_86_183 ();
 b15zdnd00an1n01x5 FILLER_86_185 ();
 b15zdnd11an1n64x5 FILLER_86_238 ();
 b15zdnd11an1n32x5 FILLER_86_302 ();
 b15zdnd11an1n04x5 FILLER_86_334 ();
 b15zdnd00an1n02x5 FILLER_86_338 ();
 b15zdnd11an1n04x5 FILLER_86_343 ();
 b15zdnd11an1n64x5 FILLER_86_350 ();
 b15zdnd11an1n64x5 FILLER_86_414 ();
 b15zdnd11an1n08x5 FILLER_86_478 ();
 b15zdnd11an1n64x5 FILLER_86_538 ();
 b15zdnd11an1n64x5 FILLER_86_602 ();
 b15zdnd11an1n32x5 FILLER_86_666 ();
 b15zdnd11an1n16x5 FILLER_86_698 ();
 b15zdnd11an1n04x5 FILLER_86_714 ();
 b15zdnd11an1n16x5 FILLER_86_726 ();
 b15zdnd11an1n08x5 FILLER_86_742 ();
 b15zdnd11an1n04x5 FILLER_86_750 ();
 b15zdnd11an1n64x5 FILLER_86_761 ();
 b15zdnd11an1n64x5 FILLER_86_825 ();
 b15zdnd11an1n64x5 FILLER_86_889 ();
 b15zdnd11an1n64x5 FILLER_86_953 ();
 b15zdnd11an1n64x5 FILLER_86_1017 ();
 b15zdnd11an1n32x5 FILLER_86_1081 ();
 b15zdnd11an1n16x5 FILLER_86_1113 ();
 b15zdnd11an1n08x5 FILLER_86_1129 ();
 b15zdnd11an1n04x5 FILLER_86_1137 ();
 b15zdnd00an1n01x5 FILLER_86_1141 ();
 b15zdnd11an1n64x5 FILLER_86_1158 ();
 b15zdnd11an1n32x5 FILLER_86_1222 ();
 b15zdnd00an1n02x5 FILLER_86_1254 ();
 b15zdnd11an1n04x5 FILLER_86_1259 ();
 b15zdnd11an1n04x5 FILLER_86_1266 ();
 b15zdnd11an1n04x5 FILLER_86_1273 ();
 b15zdnd11an1n64x5 FILLER_86_1280 ();
 b15zdnd11an1n32x5 FILLER_86_1344 ();
 b15zdnd11an1n04x5 FILLER_86_1376 ();
 b15zdnd00an1n02x5 FILLER_86_1380 ();
 b15zdnd00an1n01x5 FILLER_86_1382 ();
 b15zdnd11an1n64x5 FILLER_86_1386 ();
 b15zdnd11an1n64x5 FILLER_86_1450 ();
 b15zdnd11an1n64x5 FILLER_86_1514 ();
 b15zdnd11an1n64x5 FILLER_86_1578 ();
 b15zdnd11an1n64x5 FILLER_86_1642 ();
 b15zdnd11an1n64x5 FILLER_86_1706 ();
 b15zdnd11an1n64x5 FILLER_86_1770 ();
 b15zdnd11an1n64x5 FILLER_86_1834 ();
 b15zdnd11an1n64x5 FILLER_86_1898 ();
 b15zdnd11an1n64x5 FILLER_86_1962 ();
 b15zdnd11an1n64x5 FILLER_86_2026 ();
 b15zdnd11an1n64x5 FILLER_86_2090 ();
 b15zdnd11an1n64x5 FILLER_86_2162 ();
 b15zdnd11an1n32x5 FILLER_86_2226 ();
 b15zdnd11an1n16x5 FILLER_86_2258 ();
 b15zdnd00an1n02x5 FILLER_86_2274 ();
 b15zdnd11an1n16x5 FILLER_87_0 ();
 b15zdnd11an1n08x5 FILLER_87_16 ();
 b15zdnd11an1n04x5 FILLER_87_27 ();
 b15zdnd00an1n02x5 FILLER_87_31 ();
 b15zdnd00an1n01x5 FILLER_87_33 ();
 b15zdnd11an1n04x5 FILLER_87_37 ();
 b15zdnd11an1n64x5 FILLER_87_44 ();
 b15zdnd11an1n64x5 FILLER_87_108 ();
 b15zdnd11an1n16x5 FILLER_87_172 ();
 b15zdnd00an1n01x5 FILLER_87_188 ();
 b15zdnd11an1n64x5 FILLER_87_241 ();
 b15zdnd11an1n32x5 FILLER_87_305 ();
 b15zdnd11an1n08x5 FILLER_87_337 ();
 b15zdnd00an1n01x5 FILLER_87_345 ();
 b15zdnd11an1n32x5 FILLER_87_349 ();
 b15zdnd11an1n64x5 FILLER_87_401 ();
 b15zdnd11an1n32x5 FILLER_87_465 ();
 b15zdnd00an1n02x5 FILLER_87_497 ();
 b15zdnd11an1n04x5 FILLER_87_502 ();
 b15zdnd11an1n04x5 FILLER_87_509 ();
 b15zdnd11an1n64x5 FILLER_87_516 ();
 b15zdnd11an1n64x5 FILLER_87_580 ();
 b15zdnd11an1n64x5 FILLER_87_644 ();
 b15zdnd11an1n64x5 FILLER_87_708 ();
 b15zdnd11an1n32x5 FILLER_87_772 ();
 b15zdnd11an1n16x5 FILLER_87_804 ();
 b15zdnd00an1n02x5 FILLER_87_820 ();
 b15zdnd11an1n04x5 FILLER_87_833 ();
 b15zdnd11an1n64x5 FILLER_87_840 ();
 b15zdnd11an1n64x5 FILLER_87_904 ();
 b15zdnd11an1n64x5 FILLER_87_968 ();
 b15zdnd11an1n64x5 FILLER_87_1032 ();
 b15zdnd11an1n64x5 FILLER_87_1096 ();
 b15zdnd11an1n64x5 FILLER_87_1160 ();
 b15zdnd11an1n08x5 FILLER_87_1224 ();
 b15zdnd11an1n04x5 FILLER_87_1232 ();
 b15zdnd00an1n02x5 FILLER_87_1236 ();
 b15zdnd00an1n01x5 FILLER_87_1238 ();
 b15zdnd11an1n64x5 FILLER_87_1278 ();
 b15zdnd11an1n08x5 FILLER_87_1342 ();
 b15zdnd11an1n04x5 FILLER_87_1350 ();
 b15zdnd00an1n02x5 FILLER_87_1354 ();
 b15zdnd00an1n01x5 FILLER_87_1356 ();
 b15zdnd11an1n64x5 FILLER_87_1409 ();
 b15zdnd11an1n32x5 FILLER_87_1473 ();
 b15zdnd11an1n08x5 FILLER_87_1505 ();
 b15zdnd00an1n02x5 FILLER_87_1513 ();
 b15zdnd00an1n01x5 FILLER_87_1515 ();
 b15zdnd11an1n64x5 FILLER_87_1525 ();
 b15zdnd11an1n64x5 FILLER_87_1589 ();
 b15zdnd11an1n08x5 FILLER_87_1653 ();
 b15zdnd11an1n04x5 FILLER_87_1661 ();
 b15zdnd00an1n02x5 FILLER_87_1665 ();
 b15zdnd00an1n01x5 FILLER_87_1667 ();
 b15zdnd11an1n64x5 FILLER_87_1680 ();
 b15zdnd11an1n64x5 FILLER_87_1744 ();
 b15zdnd11an1n64x5 FILLER_87_1808 ();
 b15zdnd11an1n64x5 FILLER_87_1872 ();
 b15zdnd11an1n64x5 FILLER_87_1936 ();
 b15zdnd11an1n64x5 FILLER_87_2000 ();
 b15zdnd11an1n64x5 FILLER_87_2064 ();
 b15zdnd11an1n64x5 FILLER_87_2128 ();
 b15zdnd11an1n64x5 FILLER_87_2192 ();
 b15zdnd11an1n16x5 FILLER_87_2256 ();
 b15zdnd11an1n08x5 FILLER_87_2272 ();
 b15zdnd11an1n04x5 FILLER_87_2280 ();
 b15zdnd11an1n64x5 FILLER_88_8 ();
 b15zdnd11an1n64x5 FILLER_88_72 ();
 b15zdnd11an1n64x5 FILLER_88_136 ();
 b15zdnd00an1n02x5 FILLER_88_200 ();
 b15zdnd11an1n04x5 FILLER_88_205 ();
 b15zdnd11an1n04x5 FILLER_88_212 ();
 b15zdnd11an1n04x5 FILLER_88_219 ();
 b15zdnd11an1n64x5 FILLER_88_226 ();
 b15zdnd11an1n32x5 FILLER_88_290 ();
 b15zdnd11an1n08x5 FILLER_88_322 ();
 b15zdnd00an1n02x5 FILLER_88_330 ();
 b15zdnd00an1n01x5 FILLER_88_332 ();
 b15zdnd11an1n64x5 FILLER_88_385 ();
 b15zdnd11an1n32x5 FILLER_88_449 ();
 b15zdnd11an1n16x5 FILLER_88_481 ();
 b15zdnd11an1n04x5 FILLER_88_497 ();
 b15zdnd00an1n01x5 FILLER_88_501 ();
 b15zdnd11an1n04x5 FILLER_88_505 ();
 b15zdnd00an1n02x5 FILLER_88_509 ();
 b15zdnd00an1n01x5 FILLER_88_511 ();
 b15zdnd11an1n32x5 FILLER_88_515 ();
 b15zdnd11an1n08x5 FILLER_88_547 ();
 b15zdnd00an1n01x5 FILLER_88_555 ();
 b15zdnd11an1n64x5 FILLER_88_567 ();
 b15zdnd11an1n16x5 FILLER_88_631 ();
 b15zdnd11an1n04x5 FILLER_88_647 ();
 b15zdnd00an1n02x5 FILLER_88_651 ();
 b15zdnd11an1n32x5 FILLER_88_656 ();
 b15zdnd11an1n16x5 FILLER_88_688 ();
 b15zdnd11an1n08x5 FILLER_88_704 ();
 b15zdnd11an1n04x5 FILLER_88_712 ();
 b15zdnd00an1n02x5 FILLER_88_716 ();
 b15zdnd11an1n32x5 FILLER_88_726 ();
 b15zdnd11an1n16x5 FILLER_88_758 ();
 b15zdnd11an1n08x5 FILLER_88_774 ();
 b15zdnd11an1n04x5 FILLER_88_782 ();
 b15zdnd00an1n01x5 FILLER_88_786 ();
 b15zdnd11an1n64x5 FILLER_88_839 ();
 b15zdnd11an1n64x5 FILLER_88_903 ();
 b15zdnd11an1n64x5 FILLER_88_967 ();
 b15zdnd11an1n64x5 FILLER_88_1031 ();
 b15zdnd11an1n64x5 FILLER_88_1095 ();
 b15zdnd11an1n08x5 FILLER_88_1159 ();
 b15zdnd00an1n02x5 FILLER_88_1167 ();
 b15zdnd00an1n01x5 FILLER_88_1169 ();
 b15zdnd11an1n64x5 FILLER_88_1179 ();
 b15zdnd00an1n02x5 FILLER_88_1243 ();
 b15zdnd11an1n04x5 FILLER_88_1252 ();
 b15zdnd00an1n02x5 FILLER_88_1256 ();
 b15zdnd00an1n01x5 FILLER_88_1258 ();
 b15zdnd11an1n04x5 FILLER_88_1267 ();
 b15zdnd00an1n02x5 FILLER_88_1271 ();
 b15zdnd00an1n01x5 FILLER_88_1273 ();
 b15zdnd11an1n64x5 FILLER_88_1281 ();
 b15zdnd11an1n32x5 FILLER_88_1345 ();
 b15zdnd11an1n04x5 FILLER_88_1377 ();
 b15zdnd00an1n01x5 FILLER_88_1381 ();
 b15zdnd11an1n04x5 FILLER_88_1385 ();
 b15zdnd11an1n64x5 FILLER_88_1392 ();
 b15zdnd11an1n64x5 FILLER_88_1456 ();
 b15zdnd11an1n32x5 FILLER_88_1520 ();
 b15zdnd11an1n16x5 FILLER_88_1552 ();
 b15zdnd11an1n08x5 FILLER_88_1568 ();
 b15zdnd11an1n64x5 FILLER_88_1579 ();
 b15zdnd11an1n64x5 FILLER_88_1643 ();
 b15zdnd11an1n64x5 FILLER_88_1707 ();
 b15zdnd11an1n64x5 FILLER_88_1771 ();
 b15zdnd11an1n64x5 FILLER_88_1835 ();
 b15zdnd11an1n64x5 FILLER_88_1899 ();
 b15zdnd11an1n64x5 FILLER_88_1963 ();
 b15zdnd11an1n64x5 FILLER_88_2027 ();
 b15zdnd11an1n32x5 FILLER_88_2091 ();
 b15zdnd11an1n16x5 FILLER_88_2123 ();
 b15zdnd11an1n08x5 FILLER_88_2139 ();
 b15zdnd11an1n04x5 FILLER_88_2147 ();
 b15zdnd00an1n02x5 FILLER_88_2151 ();
 b15zdnd00an1n01x5 FILLER_88_2153 ();
 b15zdnd11an1n64x5 FILLER_88_2162 ();
 b15zdnd11an1n32x5 FILLER_88_2226 ();
 b15zdnd11an1n16x5 FILLER_88_2258 ();
 b15zdnd00an1n02x5 FILLER_88_2274 ();
 b15zdnd11an1n64x5 FILLER_89_0 ();
 b15zdnd11an1n64x5 FILLER_89_64 ();
 b15zdnd11an1n64x5 FILLER_89_128 ();
 b15zdnd11an1n16x5 FILLER_89_192 ();
 b15zdnd11an1n04x5 FILLER_89_208 ();
 b15zdnd11an1n16x5 FILLER_89_215 ();
 b15zdnd11an1n08x5 FILLER_89_231 ();
 b15zdnd11an1n04x5 FILLER_89_239 ();
 b15zdnd00an1n02x5 FILLER_89_243 ();
 b15zdnd00an1n01x5 FILLER_89_245 ();
 b15zdnd11an1n04x5 FILLER_89_249 ();
 b15zdnd11an1n64x5 FILLER_89_280 ();
 b15zdnd11an1n08x5 FILLER_89_344 ();
 b15zdnd00an1n01x5 FILLER_89_352 ();
 b15zdnd11an1n04x5 FILLER_89_356 ();
 b15zdnd11an1n64x5 FILLER_89_363 ();
 b15zdnd11an1n16x5 FILLER_89_427 ();
 b15zdnd00an1n02x5 FILLER_89_443 ();
 b15zdnd11an1n64x5 FILLER_89_465 ();
 b15zdnd11an1n64x5 FILLER_89_529 ();
 b15zdnd00an1n02x5 FILLER_89_593 ();
 b15zdnd11an1n04x5 FILLER_89_622 ();
 b15zdnd11an1n32x5 FILLER_89_678 ();
 b15zdnd11an1n04x5 FILLER_89_710 ();
 b15zdnd11an1n64x5 FILLER_89_734 ();
 b15zdnd11an1n08x5 FILLER_89_798 ();
 b15zdnd00an1n01x5 FILLER_89_806 ();
 b15zdnd11an1n04x5 FILLER_89_810 ();
 b15zdnd11an1n64x5 FILLER_89_866 ();
 b15zdnd11an1n64x5 FILLER_89_930 ();
 b15zdnd11an1n64x5 FILLER_89_994 ();
 b15zdnd11an1n64x5 FILLER_89_1058 ();
 b15zdnd11an1n64x5 FILLER_89_1122 ();
 b15zdnd11an1n64x5 FILLER_89_1186 ();
 b15zdnd11an1n64x5 FILLER_89_1250 ();
 b15zdnd11an1n64x5 FILLER_89_1314 ();
 b15zdnd11an1n04x5 FILLER_89_1378 ();
 b15zdnd00an1n01x5 FILLER_89_1382 ();
 b15zdnd11an1n64x5 FILLER_89_1388 ();
 b15zdnd00an1n02x5 FILLER_89_1452 ();
 b15zdnd11an1n04x5 FILLER_89_1457 ();
 b15zdnd11an1n64x5 FILLER_89_1464 ();
 b15zdnd11an1n32x5 FILLER_89_1528 ();
 b15zdnd11an1n08x5 FILLER_89_1560 ();
 b15zdnd11an1n04x5 FILLER_89_1568 ();
 b15zdnd00an1n02x5 FILLER_89_1572 ();
 b15zdnd11an1n04x5 FILLER_89_1577 ();
 b15zdnd11an1n64x5 FILLER_89_1584 ();
 b15zdnd11an1n64x5 FILLER_89_1648 ();
 b15zdnd11an1n64x5 FILLER_89_1712 ();
 b15zdnd11an1n64x5 FILLER_89_1776 ();
 b15zdnd11an1n64x5 FILLER_89_1840 ();
 b15zdnd11an1n64x5 FILLER_89_1904 ();
 b15zdnd11an1n64x5 FILLER_89_1968 ();
 b15zdnd11an1n64x5 FILLER_89_2032 ();
 b15zdnd11an1n64x5 FILLER_89_2096 ();
 b15zdnd11an1n64x5 FILLER_89_2160 ();
 b15zdnd11an1n32x5 FILLER_89_2224 ();
 b15zdnd11an1n16x5 FILLER_89_2256 ();
 b15zdnd11an1n08x5 FILLER_89_2272 ();
 b15zdnd11an1n04x5 FILLER_89_2280 ();
 b15zdnd11an1n64x5 FILLER_90_8 ();
 b15zdnd11an1n64x5 FILLER_90_72 ();
 b15zdnd11an1n64x5 FILLER_90_136 ();
 b15zdnd11an1n64x5 FILLER_90_200 ();
 b15zdnd11an1n64x5 FILLER_90_264 ();
 b15zdnd11an1n32x5 FILLER_90_328 ();
 b15zdnd00an1n01x5 FILLER_90_360 ();
 b15zdnd11an1n64x5 FILLER_90_364 ();
 b15zdnd11an1n64x5 FILLER_90_428 ();
 b15zdnd11an1n64x5 FILLER_90_492 ();
 b15zdnd11an1n32x5 FILLER_90_556 ();
 b15zdnd11an1n04x5 FILLER_90_588 ();
 b15zdnd00an1n02x5 FILLER_90_592 ();
 b15zdnd00an1n01x5 FILLER_90_594 ();
 b15zdnd11an1n32x5 FILLER_90_598 ();
 b15zdnd11an1n08x5 FILLER_90_630 ();
 b15zdnd11an1n04x5 FILLER_90_638 ();
 b15zdnd00an1n02x5 FILLER_90_642 ();
 b15zdnd00an1n01x5 FILLER_90_644 ();
 b15zdnd11an1n04x5 FILLER_90_648 ();
 b15zdnd11an1n32x5 FILLER_90_655 ();
 b15zdnd11an1n04x5 FILLER_90_711 ();
 b15zdnd00an1n02x5 FILLER_90_715 ();
 b15zdnd00an1n01x5 FILLER_90_717 ();
 b15zdnd11an1n64x5 FILLER_90_726 ();
 b15zdnd11an1n16x5 FILLER_90_790 ();
 b15zdnd00an1n01x5 FILLER_90_806 ();
 b15zdnd11an1n04x5 FILLER_90_810 ();
 b15zdnd11an1n16x5 FILLER_90_817 ();
 b15zdnd11an1n04x5 FILLER_90_833 ();
 b15zdnd11an1n08x5 FILLER_90_840 ();
 b15zdnd00an1n01x5 FILLER_90_848 ();
 b15zdnd11an1n64x5 FILLER_90_852 ();
 b15zdnd11an1n64x5 FILLER_90_916 ();
 b15zdnd11an1n64x5 FILLER_90_980 ();
 b15zdnd11an1n64x5 FILLER_90_1044 ();
 b15zdnd11an1n64x5 FILLER_90_1108 ();
 b15zdnd11an1n64x5 FILLER_90_1172 ();
 b15zdnd11an1n64x5 FILLER_90_1236 ();
 b15zdnd11an1n64x5 FILLER_90_1300 ();
 b15zdnd11an1n64x5 FILLER_90_1364 ();
 b15zdnd11an1n08x5 FILLER_90_1428 ();
 b15zdnd11an1n64x5 FILLER_90_1488 ();
 b15zdnd11an1n04x5 FILLER_90_1552 ();
 b15zdnd11an1n32x5 FILLER_90_1608 ();
 b15zdnd11an1n08x5 FILLER_90_1640 ();
 b15zdnd00an1n01x5 FILLER_90_1648 ();
 b15zdnd11an1n04x5 FILLER_90_1663 ();
 b15zdnd11an1n64x5 FILLER_90_1687 ();
 b15zdnd11an1n64x5 FILLER_90_1751 ();
 b15zdnd11an1n64x5 FILLER_90_1815 ();
 b15zdnd11an1n64x5 FILLER_90_1879 ();
 b15zdnd11an1n64x5 FILLER_90_1943 ();
 b15zdnd11an1n64x5 FILLER_90_2007 ();
 b15zdnd11an1n64x5 FILLER_90_2071 ();
 b15zdnd11an1n16x5 FILLER_90_2135 ();
 b15zdnd00an1n02x5 FILLER_90_2151 ();
 b15zdnd00an1n01x5 FILLER_90_2153 ();
 b15zdnd11an1n64x5 FILLER_90_2162 ();
 b15zdnd11an1n32x5 FILLER_90_2226 ();
 b15zdnd11an1n16x5 FILLER_90_2258 ();
 b15zdnd00an1n02x5 FILLER_90_2274 ();
 b15zdnd11an1n64x5 FILLER_91_0 ();
 b15zdnd11an1n64x5 FILLER_91_64 ();
 b15zdnd11an1n64x5 FILLER_91_128 ();
 b15zdnd11an1n64x5 FILLER_91_192 ();
 b15zdnd11an1n64x5 FILLER_91_256 ();
 b15zdnd11an1n64x5 FILLER_91_320 ();
 b15zdnd11an1n64x5 FILLER_91_384 ();
 b15zdnd11an1n64x5 FILLER_91_448 ();
 b15zdnd11an1n64x5 FILLER_91_512 ();
 b15zdnd11an1n64x5 FILLER_91_576 ();
 b15zdnd11an1n64x5 FILLER_91_640 ();
 b15zdnd11an1n64x5 FILLER_91_704 ();
 b15zdnd11an1n32x5 FILLER_91_768 ();
 b15zdnd11an1n16x5 FILLER_91_800 ();
 b15zdnd11an1n04x5 FILLER_91_816 ();
 b15zdnd00an1n02x5 FILLER_91_820 ();
 b15zdnd00an1n01x5 FILLER_91_822 ();
 b15zdnd11an1n64x5 FILLER_91_834 ();
 b15zdnd00an1n02x5 FILLER_91_898 ();
 b15zdnd11an1n32x5 FILLER_91_903 ();
 b15zdnd11an1n16x5 FILLER_91_935 ();
 b15zdnd11an1n04x5 FILLER_91_951 ();
 b15zdnd00an1n02x5 FILLER_91_955 ();
 b15zdnd11an1n64x5 FILLER_91_960 ();
 b15zdnd11an1n64x5 FILLER_91_1024 ();
 b15zdnd11an1n64x5 FILLER_91_1088 ();
 b15zdnd11an1n64x5 FILLER_91_1152 ();
 b15zdnd11an1n64x5 FILLER_91_1216 ();
 b15zdnd11an1n64x5 FILLER_91_1280 ();
 b15zdnd11an1n64x5 FILLER_91_1344 ();
 b15zdnd11an1n32x5 FILLER_91_1408 ();
 b15zdnd11an1n16x5 FILLER_91_1440 ();
 b15zdnd11an1n04x5 FILLER_91_1456 ();
 b15zdnd00an1n01x5 FILLER_91_1460 ();
 b15zdnd11an1n64x5 FILLER_91_1464 ();
 b15zdnd11an1n64x5 FILLER_91_1528 ();
 b15zdnd11an1n08x5 FILLER_91_1592 ();
 b15zdnd11an1n04x5 FILLER_91_1600 ();
 b15zdnd00an1n02x5 FILLER_91_1604 ();
 b15zdnd00an1n01x5 FILLER_91_1606 ();
 b15zdnd11an1n64x5 FILLER_91_1621 ();
 b15zdnd11an1n64x5 FILLER_91_1685 ();
 b15zdnd11an1n64x5 FILLER_91_1749 ();
 b15zdnd11an1n64x5 FILLER_91_1813 ();
 b15zdnd11an1n64x5 FILLER_91_1877 ();
 b15zdnd11an1n64x5 FILLER_91_1941 ();
 b15zdnd11an1n64x5 FILLER_91_2005 ();
 b15zdnd11an1n64x5 FILLER_91_2069 ();
 b15zdnd11an1n64x5 FILLER_91_2133 ();
 b15zdnd11an1n64x5 FILLER_91_2197 ();
 b15zdnd11an1n16x5 FILLER_91_2261 ();
 b15zdnd11an1n04x5 FILLER_91_2277 ();
 b15zdnd00an1n02x5 FILLER_91_2281 ();
 b15zdnd00an1n01x5 FILLER_91_2283 ();
 b15zdnd11an1n64x5 FILLER_92_8 ();
 b15zdnd11an1n64x5 FILLER_92_72 ();
 b15zdnd11an1n64x5 FILLER_92_136 ();
 b15zdnd11an1n32x5 FILLER_92_200 ();
 b15zdnd11an1n04x5 FILLER_92_232 ();
 b15zdnd00an1n02x5 FILLER_92_236 ();
 b15zdnd11an1n32x5 FILLER_92_247 ();
 b15zdnd11an1n08x5 FILLER_92_279 ();
 b15zdnd11an1n04x5 FILLER_92_287 ();
 b15zdnd00an1n02x5 FILLER_92_291 ();
 b15zdnd00an1n01x5 FILLER_92_293 ();
 b15zdnd11an1n64x5 FILLER_92_303 ();
 b15zdnd11an1n64x5 FILLER_92_367 ();
 b15zdnd11an1n64x5 FILLER_92_431 ();
 b15zdnd11an1n32x5 FILLER_92_495 ();
 b15zdnd11an1n16x5 FILLER_92_527 ();
 b15zdnd00an1n01x5 FILLER_92_543 ();
 b15zdnd11an1n32x5 FILLER_92_553 ();
 b15zdnd11an1n08x5 FILLER_92_585 ();
 b15zdnd11an1n04x5 FILLER_92_593 ();
 b15zdnd00an1n02x5 FILLER_92_597 ();
 b15zdnd11an1n64x5 FILLER_92_608 ();
 b15zdnd11an1n32x5 FILLER_92_672 ();
 b15zdnd11an1n08x5 FILLER_92_704 ();
 b15zdnd11an1n04x5 FILLER_92_712 ();
 b15zdnd00an1n02x5 FILLER_92_716 ();
 b15zdnd11an1n64x5 FILLER_92_726 ();
 b15zdnd11an1n64x5 FILLER_92_790 ();
 b15zdnd11an1n16x5 FILLER_92_854 ();
 b15zdnd11an1n04x5 FILLER_92_870 ();
 b15zdnd00an1n02x5 FILLER_92_874 ();
 b15zdnd00an1n01x5 FILLER_92_876 ();
 b15zdnd11an1n08x5 FILLER_92_886 ();
 b15zdnd11an1n04x5 FILLER_92_894 ();
 b15zdnd00an1n01x5 FILLER_92_898 ();
 b15zdnd11an1n04x5 FILLER_92_926 ();
 b15zdnd11an1n64x5 FILLER_92_982 ();
 b15zdnd11an1n64x5 FILLER_92_1046 ();
 b15zdnd11an1n64x5 FILLER_92_1110 ();
 b15zdnd11an1n64x5 FILLER_92_1174 ();
 b15zdnd11an1n64x5 FILLER_92_1238 ();
 b15zdnd11an1n64x5 FILLER_92_1302 ();
 b15zdnd11an1n64x5 FILLER_92_1366 ();
 b15zdnd11an1n64x5 FILLER_92_1430 ();
 b15zdnd11an1n16x5 FILLER_92_1494 ();
 b15zdnd11an1n04x5 FILLER_92_1510 ();
 b15zdnd00an1n02x5 FILLER_92_1514 ();
 b15zdnd11an1n64x5 FILLER_92_1525 ();
 b15zdnd11an1n64x5 FILLER_92_1589 ();
 b15zdnd11an1n64x5 FILLER_92_1653 ();
 b15zdnd11an1n64x5 FILLER_92_1717 ();
 b15zdnd11an1n64x5 FILLER_92_1781 ();
 b15zdnd11an1n64x5 FILLER_92_1845 ();
 b15zdnd11an1n64x5 FILLER_92_1909 ();
 b15zdnd11an1n64x5 FILLER_92_1973 ();
 b15zdnd11an1n64x5 FILLER_92_2037 ();
 b15zdnd11an1n32x5 FILLER_92_2101 ();
 b15zdnd11an1n16x5 FILLER_92_2133 ();
 b15zdnd11an1n04x5 FILLER_92_2149 ();
 b15zdnd00an1n01x5 FILLER_92_2153 ();
 b15zdnd11an1n64x5 FILLER_92_2162 ();
 b15zdnd11an1n32x5 FILLER_92_2226 ();
 b15zdnd11an1n16x5 FILLER_92_2258 ();
 b15zdnd00an1n02x5 FILLER_92_2274 ();
 b15zdnd11an1n64x5 FILLER_93_0 ();
 b15zdnd11an1n64x5 FILLER_93_64 ();
 b15zdnd11an1n64x5 FILLER_93_128 ();
 b15zdnd11an1n64x5 FILLER_93_192 ();
 b15zdnd11an1n64x5 FILLER_93_256 ();
 b15zdnd11an1n64x5 FILLER_93_320 ();
 b15zdnd11an1n64x5 FILLER_93_384 ();
 b15zdnd11an1n64x5 FILLER_93_448 ();
 b15zdnd11an1n64x5 FILLER_93_512 ();
 b15zdnd11an1n32x5 FILLER_93_576 ();
 b15zdnd11an1n16x5 FILLER_93_608 ();
 b15zdnd11an1n04x5 FILLER_93_624 ();
 b15zdnd00an1n02x5 FILLER_93_628 ();
 b15zdnd00an1n01x5 FILLER_93_630 ();
 b15zdnd11an1n64x5 FILLER_93_645 ();
 b15zdnd11an1n64x5 FILLER_93_709 ();
 b15zdnd11an1n64x5 FILLER_93_773 ();
 b15zdnd11an1n64x5 FILLER_93_837 ();
 b15zdnd11an1n32x5 FILLER_93_901 ();
 b15zdnd11an1n08x5 FILLER_93_933 ();
 b15zdnd11an1n04x5 FILLER_93_941 ();
 b15zdnd00an1n02x5 FILLER_93_945 ();
 b15zdnd00an1n01x5 FILLER_93_947 ();
 b15zdnd11an1n04x5 FILLER_93_951 ();
 b15zdnd11an1n64x5 FILLER_93_958 ();
 b15zdnd11an1n64x5 FILLER_93_1022 ();
 b15zdnd11an1n64x5 FILLER_93_1086 ();
 b15zdnd11an1n64x5 FILLER_93_1150 ();
 b15zdnd11an1n64x5 FILLER_93_1214 ();
 b15zdnd11an1n64x5 FILLER_93_1278 ();
 b15zdnd11an1n32x5 FILLER_93_1342 ();
 b15zdnd00an1n02x5 FILLER_93_1374 ();
 b15zdnd00an1n01x5 FILLER_93_1376 ();
 b15zdnd11an1n64x5 FILLER_93_1382 ();
 b15zdnd11an1n64x5 FILLER_93_1446 ();
 b15zdnd11an1n16x5 FILLER_93_1510 ();
 b15zdnd11an1n04x5 FILLER_93_1526 ();
 b15zdnd00an1n02x5 FILLER_93_1530 ();
 b15zdnd00an1n01x5 FILLER_93_1532 ();
 b15zdnd11an1n64x5 FILLER_93_1542 ();
 b15zdnd11an1n32x5 FILLER_93_1606 ();
 b15zdnd11an1n04x5 FILLER_93_1638 ();
 b15zdnd11an1n04x5 FILLER_93_1662 ();
 b15zdnd11an1n64x5 FILLER_93_1692 ();
 b15zdnd11an1n64x5 FILLER_93_1756 ();
 b15zdnd11an1n64x5 FILLER_93_1820 ();
 b15zdnd11an1n08x5 FILLER_93_1884 ();
 b15zdnd00an1n01x5 FILLER_93_1892 ();
 b15zdnd11an1n64x5 FILLER_93_1913 ();
 b15zdnd11an1n64x5 FILLER_93_1977 ();
 b15zdnd11an1n64x5 FILLER_93_2041 ();
 b15zdnd11an1n64x5 FILLER_93_2105 ();
 b15zdnd11an1n64x5 FILLER_93_2169 ();
 b15zdnd11an1n32x5 FILLER_93_2233 ();
 b15zdnd11an1n16x5 FILLER_93_2265 ();
 b15zdnd00an1n02x5 FILLER_93_2281 ();
 b15zdnd00an1n01x5 FILLER_93_2283 ();
 b15zdnd11an1n64x5 FILLER_94_8 ();
 b15zdnd11an1n64x5 FILLER_94_72 ();
 b15zdnd11an1n32x5 FILLER_94_136 ();
 b15zdnd11an1n16x5 FILLER_94_168 ();
 b15zdnd11an1n08x5 FILLER_94_184 ();
 b15zdnd00an1n01x5 FILLER_94_192 ();
 b15zdnd11an1n64x5 FILLER_94_224 ();
 b15zdnd11an1n64x5 FILLER_94_288 ();
 b15zdnd11an1n64x5 FILLER_94_352 ();
 b15zdnd11an1n64x5 FILLER_94_416 ();
 b15zdnd11an1n64x5 FILLER_94_480 ();
 b15zdnd11an1n64x5 FILLER_94_544 ();
 b15zdnd11an1n16x5 FILLER_94_608 ();
 b15zdnd11an1n04x5 FILLER_94_624 ();
 b15zdnd00an1n02x5 FILLER_94_628 ();
 b15zdnd11an1n32x5 FILLER_94_682 ();
 b15zdnd11an1n04x5 FILLER_94_714 ();
 b15zdnd11an1n64x5 FILLER_94_726 ();
 b15zdnd11an1n64x5 FILLER_94_790 ();
 b15zdnd11an1n64x5 FILLER_94_854 ();
 b15zdnd11an1n64x5 FILLER_94_918 ();
 b15zdnd11an1n64x5 FILLER_94_982 ();
 b15zdnd11an1n08x5 FILLER_94_1046 ();
 b15zdnd11an1n04x5 FILLER_94_1054 ();
 b15zdnd00an1n02x5 FILLER_94_1058 ();
 b15zdnd00an1n01x5 FILLER_94_1060 ();
 b15zdnd11an1n16x5 FILLER_94_1077 ();
 b15zdnd11an1n04x5 FILLER_94_1093 ();
 b15zdnd11an1n64x5 FILLER_94_1113 ();
 b15zdnd11an1n64x5 FILLER_94_1177 ();
 b15zdnd11an1n64x5 FILLER_94_1241 ();
 b15zdnd11an1n64x5 FILLER_94_1305 ();
 b15zdnd11an1n64x5 FILLER_94_1369 ();
 b15zdnd11an1n32x5 FILLER_94_1433 ();
 b15zdnd11an1n08x5 FILLER_94_1465 ();
 b15zdnd11an1n04x5 FILLER_94_1473 ();
 b15zdnd00an1n02x5 FILLER_94_1477 ();
 b15zdnd00an1n01x5 FILLER_94_1479 ();
 b15zdnd11an1n04x5 FILLER_94_1522 ();
 b15zdnd00an1n02x5 FILLER_94_1526 ();
 b15zdnd00an1n01x5 FILLER_94_1528 ();
 b15zdnd11an1n64x5 FILLER_94_1571 ();
 b15zdnd11an1n16x5 FILLER_94_1635 ();
 b15zdnd11an1n04x5 FILLER_94_1668 ();
 b15zdnd11an1n16x5 FILLER_94_1686 ();
 b15zdnd11an1n04x5 FILLER_94_1702 ();
 b15zdnd00an1n02x5 FILLER_94_1706 ();
 b15zdnd11an1n64x5 FILLER_94_1728 ();
 b15zdnd11an1n64x5 FILLER_94_1792 ();
 b15zdnd11an1n64x5 FILLER_94_1856 ();
 b15zdnd11an1n64x5 FILLER_94_1920 ();
 b15zdnd11an1n64x5 FILLER_94_1984 ();
 b15zdnd11an1n64x5 FILLER_94_2048 ();
 b15zdnd11an1n32x5 FILLER_94_2112 ();
 b15zdnd11an1n08x5 FILLER_94_2144 ();
 b15zdnd00an1n02x5 FILLER_94_2152 ();
 b15zdnd11an1n64x5 FILLER_94_2162 ();
 b15zdnd11an1n32x5 FILLER_94_2226 ();
 b15zdnd11an1n16x5 FILLER_94_2258 ();
 b15zdnd00an1n02x5 FILLER_94_2274 ();
 b15zdnd11an1n64x5 FILLER_95_0 ();
 b15zdnd11an1n64x5 FILLER_95_64 ();
 b15zdnd11an1n64x5 FILLER_95_128 ();
 b15zdnd11an1n08x5 FILLER_95_192 ();
 b15zdnd11an1n04x5 FILLER_95_200 ();
 b15zdnd11an1n32x5 FILLER_95_230 ();
 b15zdnd11an1n16x5 FILLER_95_262 ();
 b15zdnd11an1n08x5 FILLER_95_278 ();
 b15zdnd11an1n64x5 FILLER_95_295 ();
 b15zdnd11an1n64x5 FILLER_95_359 ();
 b15zdnd11an1n64x5 FILLER_95_423 ();
 b15zdnd11an1n64x5 FILLER_95_487 ();
 b15zdnd11an1n64x5 FILLER_95_551 ();
 b15zdnd11an1n32x5 FILLER_95_615 ();
 b15zdnd00an1n01x5 FILLER_95_647 ();
 b15zdnd11an1n04x5 FILLER_95_651 ();
 b15zdnd11an1n04x5 FILLER_95_658 ();
 b15zdnd11an1n64x5 FILLER_95_665 ();
 b15zdnd11an1n64x5 FILLER_95_729 ();
 b15zdnd11an1n64x5 FILLER_95_793 ();
 b15zdnd11an1n64x5 FILLER_95_857 ();
 b15zdnd11an1n64x5 FILLER_95_921 ();
 b15zdnd11an1n64x5 FILLER_95_985 ();
 b15zdnd11an1n32x5 FILLER_95_1049 ();
 b15zdnd11an1n08x5 FILLER_95_1081 ();
 b15zdnd11an1n04x5 FILLER_95_1089 ();
 b15zdnd11an1n64x5 FILLER_95_1109 ();
 b15zdnd11an1n32x5 FILLER_95_1173 ();
 b15zdnd11an1n16x5 FILLER_95_1205 ();
 b15zdnd11an1n04x5 FILLER_95_1221 ();
 b15zdnd00an1n02x5 FILLER_95_1225 ();
 b15zdnd11an1n64x5 FILLER_95_1230 ();
 b15zdnd11an1n64x5 FILLER_95_1294 ();
 b15zdnd11an1n64x5 FILLER_95_1358 ();
 b15zdnd11an1n08x5 FILLER_95_1422 ();
 b15zdnd00an1n02x5 FILLER_95_1430 ();
 b15zdnd11an1n08x5 FILLER_95_1474 ();
 b15zdnd00an1n01x5 FILLER_95_1482 ();
 b15zdnd11an1n64x5 FILLER_95_1525 ();
 b15zdnd11an1n64x5 FILLER_95_1589 ();
 b15zdnd11an1n64x5 FILLER_95_1653 ();
 b15zdnd11an1n64x5 FILLER_95_1717 ();
 b15zdnd11an1n16x5 FILLER_95_1781 ();
 b15zdnd11an1n08x5 FILLER_95_1797 ();
 b15zdnd00an1n01x5 FILLER_95_1805 ();
 b15zdnd11an1n64x5 FILLER_95_1823 ();
 b15zdnd11an1n64x5 FILLER_95_1887 ();
 b15zdnd11an1n64x5 FILLER_95_1951 ();
 b15zdnd11an1n64x5 FILLER_95_2015 ();
 b15zdnd11an1n64x5 FILLER_95_2079 ();
 b15zdnd11an1n64x5 FILLER_95_2143 ();
 b15zdnd11an1n64x5 FILLER_95_2207 ();
 b15zdnd11an1n08x5 FILLER_95_2271 ();
 b15zdnd11an1n04x5 FILLER_95_2279 ();
 b15zdnd00an1n01x5 FILLER_95_2283 ();
 b15zdnd11an1n08x5 FILLER_96_8 ();
 b15zdnd11an1n04x5 FILLER_96_16 ();
 b15zdnd00an1n02x5 FILLER_96_20 ();
 b15zdnd00an1n01x5 FILLER_96_22 ();
 b15zdnd11an1n64x5 FILLER_96_26 ();
 b15zdnd11an1n64x5 FILLER_96_90 ();
 b15zdnd11an1n32x5 FILLER_96_154 ();
 b15zdnd11an1n16x5 FILLER_96_186 ();
 b15zdnd11an1n08x5 FILLER_96_202 ();
 b15zdnd11an1n04x5 FILLER_96_210 ();
 b15zdnd11an1n64x5 FILLER_96_234 ();
 b15zdnd11an1n64x5 FILLER_96_298 ();
 b15zdnd11an1n64x5 FILLER_96_362 ();
 b15zdnd11an1n64x5 FILLER_96_426 ();
 b15zdnd11an1n64x5 FILLER_96_490 ();
 b15zdnd11an1n16x5 FILLER_96_554 ();
 b15zdnd11an1n08x5 FILLER_96_570 ();
 b15zdnd00an1n01x5 FILLER_96_578 ();
 b15zdnd11an1n64x5 FILLER_96_588 ();
 b15zdnd11an1n64x5 FILLER_96_652 ();
 b15zdnd00an1n02x5 FILLER_96_716 ();
 b15zdnd11an1n64x5 FILLER_96_726 ();
 b15zdnd11an1n64x5 FILLER_96_790 ();
 b15zdnd11an1n64x5 FILLER_96_854 ();
 b15zdnd11an1n64x5 FILLER_96_918 ();
 b15zdnd11an1n64x5 FILLER_96_982 ();
 b15zdnd11an1n32x5 FILLER_96_1046 ();
 b15zdnd11an1n08x5 FILLER_96_1078 ();
 b15zdnd11an1n32x5 FILLER_96_1102 ();
 b15zdnd11an1n08x5 FILLER_96_1134 ();
 b15zdnd00an1n01x5 FILLER_96_1142 ();
 b15zdnd11an1n32x5 FILLER_96_1146 ();
 b15zdnd11an1n16x5 FILLER_96_1178 ();
 b15zdnd11an1n04x5 FILLER_96_1194 ();
 b15zdnd00an1n02x5 FILLER_96_1198 ();
 b15zdnd00an1n01x5 FILLER_96_1200 ();
 b15zdnd11an1n64x5 FILLER_96_1253 ();
 b15zdnd11an1n64x5 FILLER_96_1317 ();
 b15zdnd11an1n64x5 FILLER_96_1381 ();
 b15zdnd11an1n64x5 FILLER_96_1445 ();
 b15zdnd11an1n64x5 FILLER_96_1509 ();
 b15zdnd11an1n64x5 FILLER_96_1573 ();
 b15zdnd11an1n64x5 FILLER_96_1637 ();
 b15zdnd11an1n64x5 FILLER_96_1701 ();
 b15zdnd11an1n16x5 FILLER_96_1765 ();
 b15zdnd11an1n08x5 FILLER_96_1781 ();
 b15zdnd11an1n32x5 FILLER_96_1809 ();
 b15zdnd11an1n16x5 FILLER_96_1841 ();
 b15zdnd11an1n08x5 FILLER_96_1857 ();
 b15zdnd11an1n04x5 FILLER_96_1865 ();
 b15zdnd00an1n02x5 FILLER_96_1869 ();
 b15zdnd11an1n64x5 FILLER_96_1888 ();
 b15zdnd11an1n64x5 FILLER_96_1952 ();
 b15zdnd11an1n64x5 FILLER_96_2016 ();
 b15zdnd11an1n64x5 FILLER_96_2080 ();
 b15zdnd11an1n08x5 FILLER_96_2144 ();
 b15zdnd00an1n02x5 FILLER_96_2152 ();
 b15zdnd11an1n64x5 FILLER_96_2162 ();
 b15zdnd11an1n32x5 FILLER_96_2226 ();
 b15zdnd11an1n16x5 FILLER_96_2258 ();
 b15zdnd00an1n02x5 FILLER_96_2274 ();
 b15zdnd11an1n16x5 FILLER_97_0 ();
 b15zdnd11an1n04x5 FILLER_97_16 ();
 b15zdnd00an1n01x5 FILLER_97_20 ();
 b15zdnd11an1n64x5 FILLER_97_24 ();
 b15zdnd11an1n64x5 FILLER_97_88 ();
 b15zdnd11an1n64x5 FILLER_97_152 ();
 b15zdnd11an1n64x5 FILLER_97_216 ();
 b15zdnd11an1n64x5 FILLER_97_280 ();
 b15zdnd11an1n64x5 FILLER_97_344 ();
 b15zdnd11an1n64x5 FILLER_97_408 ();
 b15zdnd11an1n64x5 FILLER_97_472 ();
 b15zdnd11an1n64x5 FILLER_97_536 ();
 b15zdnd11an1n64x5 FILLER_97_600 ();
 b15zdnd11an1n64x5 FILLER_97_664 ();
 b15zdnd11an1n64x5 FILLER_97_728 ();
 b15zdnd11an1n64x5 FILLER_97_792 ();
 b15zdnd11an1n64x5 FILLER_97_856 ();
 b15zdnd11an1n64x5 FILLER_97_920 ();
 b15zdnd11an1n64x5 FILLER_97_984 ();
 b15zdnd11an1n32x5 FILLER_97_1048 ();
 b15zdnd11an1n08x5 FILLER_97_1080 ();
 b15zdnd00an1n02x5 FILLER_97_1088 ();
 b15zdnd00an1n01x5 FILLER_97_1090 ();
 b15zdnd11an1n08x5 FILLER_97_1107 ();
 b15zdnd00an1n01x5 FILLER_97_1115 ();
 b15zdnd11an1n32x5 FILLER_97_1168 ();
 b15zdnd11an1n16x5 FILLER_97_1200 ();
 b15zdnd00an1n02x5 FILLER_97_1216 ();
 b15zdnd00an1n01x5 FILLER_97_1218 ();
 b15zdnd11an1n04x5 FILLER_97_1222 ();
 b15zdnd11an1n64x5 FILLER_97_1229 ();
 b15zdnd11an1n64x5 FILLER_97_1293 ();
 b15zdnd11an1n64x5 FILLER_97_1357 ();
 b15zdnd11an1n64x5 FILLER_97_1421 ();
 b15zdnd11an1n64x5 FILLER_97_1485 ();
 b15zdnd11an1n64x5 FILLER_97_1549 ();
 b15zdnd11an1n64x5 FILLER_97_1613 ();
 b15zdnd11an1n64x5 FILLER_97_1677 ();
 b15zdnd11an1n32x5 FILLER_97_1741 ();
 b15zdnd11an1n08x5 FILLER_97_1773 ();
 b15zdnd11an1n04x5 FILLER_97_1781 ();
 b15zdnd00an1n01x5 FILLER_97_1785 ();
 b15zdnd11an1n64x5 FILLER_97_1806 ();
 b15zdnd11an1n32x5 FILLER_97_1870 ();
 b15zdnd11an1n08x5 FILLER_97_1902 ();
 b15zdnd00an1n02x5 FILLER_97_1910 ();
 b15zdnd11an1n64x5 FILLER_97_1926 ();
 b15zdnd11an1n64x5 FILLER_97_1990 ();
 b15zdnd11an1n64x5 FILLER_97_2054 ();
 b15zdnd11an1n64x5 FILLER_97_2118 ();
 b15zdnd11an1n64x5 FILLER_97_2182 ();
 b15zdnd11an1n32x5 FILLER_97_2246 ();
 b15zdnd11an1n04x5 FILLER_97_2278 ();
 b15zdnd00an1n02x5 FILLER_97_2282 ();
 b15zdnd11an1n64x5 FILLER_98_8 ();
 b15zdnd11an1n64x5 FILLER_98_72 ();
 b15zdnd11an1n64x5 FILLER_98_136 ();
 b15zdnd11an1n64x5 FILLER_98_200 ();
 b15zdnd11an1n64x5 FILLER_98_264 ();
 b15zdnd11an1n64x5 FILLER_98_328 ();
 b15zdnd11an1n64x5 FILLER_98_392 ();
 b15zdnd11an1n64x5 FILLER_98_456 ();
 b15zdnd11an1n16x5 FILLER_98_520 ();
 b15zdnd11an1n08x5 FILLER_98_536 ();
 b15zdnd00an1n01x5 FILLER_98_544 ();
 b15zdnd11an1n64x5 FILLER_98_587 ();
 b15zdnd11an1n64x5 FILLER_98_651 ();
 b15zdnd00an1n02x5 FILLER_98_715 ();
 b15zdnd00an1n01x5 FILLER_98_717 ();
 b15zdnd11an1n64x5 FILLER_98_726 ();
 b15zdnd11an1n64x5 FILLER_98_790 ();
 b15zdnd11an1n64x5 FILLER_98_854 ();
 b15zdnd11an1n64x5 FILLER_98_918 ();
 b15zdnd11an1n64x5 FILLER_98_982 ();
 b15zdnd11an1n64x5 FILLER_98_1046 ();
 b15zdnd11an1n16x5 FILLER_98_1110 ();
 b15zdnd11an1n08x5 FILLER_98_1126 ();
 b15zdnd00an1n01x5 FILLER_98_1134 ();
 b15zdnd11an1n04x5 FILLER_98_1138 ();
 b15zdnd11an1n64x5 FILLER_98_1145 ();
 b15zdnd11an1n64x5 FILLER_98_1209 ();
 b15zdnd11an1n64x5 FILLER_98_1273 ();
 b15zdnd11an1n64x5 FILLER_98_1337 ();
 b15zdnd11an1n04x5 FILLER_98_1401 ();
 b15zdnd00an1n02x5 FILLER_98_1405 ();
 b15zdnd00an1n01x5 FILLER_98_1407 ();
 b15zdnd11an1n64x5 FILLER_98_1421 ();
 b15zdnd11an1n64x5 FILLER_98_1485 ();
 b15zdnd11an1n64x5 FILLER_98_1549 ();
 b15zdnd11an1n64x5 FILLER_98_1613 ();
 b15zdnd11an1n64x5 FILLER_98_1677 ();
 b15zdnd11an1n32x5 FILLER_98_1741 ();
 b15zdnd11an1n08x5 FILLER_98_1773 ();
 b15zdnd00an1n02x5 FILLER_98_1781 ();
 b15zdnd00an1n01x5 FILLER_98_1783 ();
 b15zdnd11an1n64x5 FILLER_98_1798 ();
 b15zdnd11an1n32x5 FILLER_98_1862 ();
 b15zdnd11an1n16x5 FILLER_98_1894 ();
 b15zdnd11an1n08x5 FILLER_98_1910 ();
 b15zdnd00an1n02x5 FILLER_98_1918 ();
 b15zdnd00an1n01x5 FILLER_98_1920 ();
 b15zdnd11an1n64x5 FILLER_98_1924 ();
 b15zdnd11an1n32x5 FILLER_98_1988 ();
 b15zdnd11an1n04x5 FILLER_98_2020 ();
 b15zdnd00an1n01x5 FILLER_98_2024 ();
 b15zdnd11an1n64x5 FILLER_98_2028 ();
 b15zdnd11an1n32x5 FILLER_98_2092 ();
 b15zdnd11an1n16x5 FILLER_98_2124 ();
 b15zdnd11an1n08x5 FILLER_98_2140 ();
 b15zdnd11an1n04x5 FILLER_98_2148 ();
 b15zdnd00an1n02x5 FILLER_98_2152 ();
 b15zdnd11an1n64x5 FILLER_98_2162 ();
 b15zdnd11an1n32x5 FILLER_98_2226 ();
 b15zdnd11an1n16x5 FILLER_98_2258 ();
 b15zdnd00an1n02x5 FILLER_98_2274 ();
 b15zdnd11an1n64x5 FILLER_99_0 ();
 b15zdnd11an1n64x5 FILLER_99_64 ();
 b15zdnd11an1n64x5 FILLER_99_128 ();
 b15zdnd11an1n64x5 FILLER_99_192 ();
 b15zdnd11an1n64x5 FILLER_99_256 ();
 b15zdnd11an1n64x5 FILLER_99_320 ();
 b15zdnd11an1n64x5 FILLER_99_384 ();
 b15zdnd11an1n64x5 FILLER_99_448 ();
 b15zdnd11an1n64x5 FILLER_99_512 ();
 b15zdnd11an1n64x5 FILLER_99_576 ();
 b15zdnd11an1n64x5 FILLER_99_640 ();
 b15zdnd11an1n64x5 FILLER_99_704 ();
 b15zdnd11an1n64x5 FILLER_99_768 ();
 b15zdnd11an1n64x5 FILLER_99_832 ();
 b15zdnd11an1n64x5 FILLER_99_896 ();
 b15zdnd11an1n64x5 FILLER_99_960 ();
 b15zdnd11an1n64x5 FILLER_99_1024 ();
 b15zdnd11an1n04x5 FILLER_99_1088 ();
 b15zdnd00an1n01x5 FILLER_99_1092 ();
 b15zdnd11an1n64x5 FILLER_99_1109 ();
 b15zdnd11an1n64x5 FILLER_99_1173 ();
 b15zdnd11an1n64x5 FILLER_99_1237 ();
 b15zdnd11an1n64x5 FILLER_99_1301 ();
 b15zdnd11an1n64x5 FILLER_99_1365 ();
 b15zdnd11an1n64x5 FILLER_99_1429 ();
 b15zdnd11an1n64x5 FILLER_99_1493 ();
 b15zdnd11an1n64x5 FILLER_99_1557 ();
 b15zdnd11an1n64x5 FILLER_99_1621 ();
 b15zdnd11an1n64x5 FILLER_99_1685 ();
 b15zdnd11an1n32x5 FILLER_99_1749 ();
 b15zdnd11an1n08x5 FILLER_99_1781 ();
 b15zdnd11an1n04x5 FILLER_99_1803 ();
 b15zdnd11an1n64x5 FILLER_99_1821 ();
 b15zdnd11an1n08x5 FILLER_99_1885 ();
 b15zdnd00an1n02x5 FILLER_99_1893 ();
 b15zdnd11an1n64x5 FILLER_99_1947 ();
 b15zdnd11an1n04x5 FILLER_99_2011 ();
 b15zdnd00an1n01x5 FILLER_99_2015 ();
 b15zdnd11an1n04x5 FILLER_99_2019 ();
 b15zdnd11an1n08x5 FILLER_99_2026 ();
 b15zdnd11an1n04x5 FILLER_99_2034 ();
 b15zdnd00an1n02x5 FILLER_99_2038 ();
 b15zdnd11an1n64x5 FILLER_99_2043 ();
 b15zdnd11an1n64x5 FILLER_99_2107 ();
 b15zdnd11an1n64x5 FILLER_99_2171 ();
 b15zdnd11an1n32x5 FILLER_99_2235 ();
 b15zdnd11an1n16x5 FILLER_99_2267 ();
 b15zdnd00an1n01x5 FILLER_99_2283 ();
 b15zdnd11an1n64x5 FILLER_100_8 ();
 b15zdnd11an1n64x5 FILLER_100_72 ();
 b15zdnd11an1n64x5 FILLER_100_136 ();
 b15zdnd11an1n64x5 FILLER_100_200 ();
 b15zdnd11an1n64x5 FILLER_100_264 ();
 b15zdnd11an1n16x5 FILLER_100_328 ();
 b15zdnd11an1n08x5 FILLER_100_344 ();
 b15zdnd11an1n64x5 FILLER_100_355 ();
 b15zdnd11an1n64x5 FILLER_100_419 ();
 b15zdnd11an1n64x5 FILLER_100_483 ();
 b15zdnd11an1n64x5 FILLER_100_547 ();
 b15zdnd11an1n64x5 FILLER_100_611 ();
 b15zdnd11an1n32x5 FILLER_100_675 ();
 b15zdnd11an1n08x5 FILLER_100_707 ();
 b15zdnd00an1n02x5 FILLER_100_715 ();
 b15zdnd00an1n01x5 FILLER_100_717 ();
 b15zdnd11an1n64x5 FILLER_100_726 ();
 b15zdnd11an1n64x5 FILLER_100_790 ();
 b15zdnd11an1n16x5 FILLER_100_854 ();
 b15zdnd11an1n08x5 FILLER_100_870 ();
 b15zdnd11an1n04x5 FILLER_100_878 ();
 b15zdnd00an1n02x5 FILLER_100_882 ();
 b15zdnd00an1n01x5 FILLER_100_884 ();
 b15zdnd11an1n64x5 FILLER_100_894 ();
 b15zdnd11an1n64x5 FILLER_100_958 ();
 b15zdnd11an1n64x5 FILLER_100_1022 ();
 b15zdnd11an1n64x5 FILLER_100_1086 ();
 b15zdnd11an1n64x5 FILLER_100_1150 ();
 b15zdnd11an1n64x5 FILLER_100_1214 ();
 b15zdnd11an1n64x5 FILLER_100_1278 ();
 b15zdnd11an1n32x5 FILLER_100_1342 ();
 b15zdnd11an1n16x5 FILLER_100_1374 ();
 b15zdnd11an1n04x5 FILLER_100_1390 ();
 b15zdnd11an1n64x5 FILLER_100_1399 ();
 b15zdnd11an1n64x5 FILLER_100_1463 ();
 b15zdnd11an1n32x5 FILLER_100_1527 ();
 b15zdnd11an1n08x5 FILLER_100_1559 ();
 b15zdnd11an1n04x5 FILLER_100_1567 ();
 b15zdnd00an1n01x5 FILLER_100_1571 ();
 b15zdnd11an1n32x5 FILLER_100_1581 ();
 b15zdnd11an1n16x5 FILLER_100_1613 ();
 b15zdnd11an1n08x5 FILLER_100_1629 ();
 b15zdnd11an1n04x5 FILLER_100_1637 ();
 b15zdnd00an1n01x5 FILLER_100_1641 ();
 b15zdnd11an1n64x5 FILLER_100_1662 ();
 b15zdnd11an1n64x5 FILLER_100_1726 ();
 b15zdnd00an1n02x5 FILLER_100_1790 ();
 b15zdnd11an1n64x5 FILLER_100_1804 ();
 b15zdnd11an1n32x5 FILLER_100_1868 ();
 b15zdnd11an1n16x5 FILLER_100_1900 ();
 b15zdnd11an1n04x5 FILLER_100_1916 ();
 b15zdnd11an1n04x5 FILLER_100_1923 ();
 b15zdnd11an1n64x5 FILLER_100_1930 ();
 b15zdnd11an1n04x5 FILLER_100_1994 ();
 b15zdnd11an1n64x5 FILLER_100_2050 ();
 b15zdnd11an1n32x5 FILLER_100_2114 ();
 b15zdnd11an1n08x5 FILLER_100_2146 ();
 b15zdnd11an1n64x5 FILLER_100_2162 ();
 b15zdnd11an1n32x5 FILLER_100_2226 ();
 b15zdnd11an1n16x5 FILLER_100_2258 ();
 b15zdnd00an1n02x5 FILLER_100_2274 ();
 b15zdnd11an1n32x5 FILLER_101_0 ();
 b15zdnd00an1n01x5 FILLER_101_32 ();
 b15zdnd11an1n64x5 FILLER_101_36 ();
 b15zdnd11an1n64x5 FILLER_101_100 ();
 b15zdnd11an1n64x5 FILLER_101_164 ();
 b15zdnd11an1n64x5 FILLER_101_228 ();
 b15zdnd11an1n32x5 FILLER_101_292 ();
 b15zdnd11an1n16x5 FILLER_101_324 ();
 b15zdnd11an1n04x5 FILLER_101_340 ();
 b15zdnd00an1n02x5 FILLER_101_344 ();
 b15zdnd00an1n01x5 FILLER_101_346 ();
 b15zdnd11an1n04x5 FILLER_101_350 ();
 b15zdnd11an1n64x5 FILLER_101_357 ();
 b15zdnd11an1n16x5 FILLER_101_421 ();
 b15zdnd11an1n08x5 FILLER_101_437 ();
 b15zdnd11an1n04x5 FILLER_101_445 ();
 b15zdnd00an1n01x5 FILLER_101_449 ();
 b15zdnd11an1n64x5 FILLER_101_464 ();
 b15zdnd11an1n64x5 FILLER_101_528 ();
 b15zdnd11an1n32x5 FILLER_101_592 ();
 b15zdnd11an1n16x5 FILLER_101_624 ();
 b15zdnd11an1n08x5 FILLER_101_640 ();
 b15zdnd00an1n02x5 FILLER_101_648 ();
 b15zdnd11an1n64x5 FILLER_101_653 ();
 b15zdnd11an1n64x5 FILLER_101_717 ();
 b15zdnd11an1n64x5 FILLER_101_781 ();
 b15zdnd11an1n64x5 FILLER_101_845 ();
 b15zdnd11an1n64x5 FILLER_101_909 ();
 b15zdnd11an1n64x5 FILLER_101_973 ();
 b15zdnd11an1n64x5 FILLER_101_1037 ();
 b15zdnd11an1n64x5 FILLER_101_1101 ();
 b15zdnd11an1n64x5 FILLER_101_1165 ();
 b15zdnd11an1n64x5 FILLER_101_1229 ();
 b15zdnd11an1n32x5 FILLER_101_1293 ();
 b15zdnd11an1n08x5 FILLER_101_1325 ();
 b15zdnd11an1n04x5 FILLER_101_1333 ();
 b15zdnd00an1n02x5 FILLER_101_1337 ();
 b15zdnd00an1n01x5 FILLER_101_1339 ();
 b15zdnd11an1n64x5 FILLER_101_1356 ();
 b15zdnd11an1n64x5 FILLER_101_1420 ();
 b15zdnd11an1n64x5 FILLER_101_1484 ();
 b15zdnd11an1n64x5 FILLER_101_1548 ();
 b15zdnd11an1n16x5 FILLER_101_1612 ();
 b15zdnd00an1n01x5 FILLER_101_1628 ();
 b15zdnd11an1n16x5 FILLER_101_1649 ();
 b15zdnd11an1n04x5 FILLER_101_1665 ();
 b15zdnd00an1n02x5 FILLER_101_1669 ();
 b15zdnd11an1n64x5 FILLER_101_1691 ();
 b15zdnd11an1n64x5 FILLER_101_1755 ();
 b15zdnd11an1n64x5 FILLER_101_1819 ();
 b15zdnd11an1n64x5 FILLER_101_1883 ();
 b15zdnd11an1n64x5 FILLER_101_1947 ();
 b15zdnd00an1n02x5 FILLER_101_2011 ();
 b15zdnd11an1n64x5 FILLER_101_2065 ();
 b15zdnd11an1n64x5 FILLER_101_2129 ();
 b15zdnd11an1n64x5 FILLER_101_2193 ();
 b15zdnd11an1n16x5 FILLER_101_2257 ();
 b15zdnd11an1n08x5 FILLER_101_2273 ();
 b15zdnd00an1n02x5 FILLER_101_2281 ();
 b15zdnd00an1n01x5 FILLER_101_2283 ();
 b15zdnd11an1n16x5 FILLER_102_8 ();
 b15zdnd00an1n02x5 FILLER_102_24 ();
 b15zdnd00an1n01x5 FILLER_102_26 ();
 b15zdnd11an1n04x5 FILLER_102_30 ();
 b15zdnd11an1n64x5 FILLER_102_37 ();
 b15zdnd11an1n64x5 FILLER_102_101 ();
 b15zdnd11an1n32x5 FILLER_102_165 ();
 b15zdnd00an1n02x5 FILLER_102_197 ();
 b15zdnd00an1n01x5 FILLER_102_199 ();
 b15zdnd11an1n04x5 FILLER_102_203 ();
 b15zdnd11an1n32x5 FILLER_102_210 ();
 b15zdnd11an1n04x5 FILLER_102_242 ();
 b15zdnd00an1n01x5 FILLER_102_246 ();
 b15zdnd11an1n64x5 FILLER_102_250 ();
 b15zdnd11an1n08x5 FILLER_102_314 ();
 b15zdnd11an1n04x5 FILLER_102_322 ();
 b15zdnd00an1n01x5 FILLER_102_326 ();
 b15zdnd11an1n64x5 FILLER_102_379 ();
 b15zdnd11an1n08x5 FILLER_102_443 ();
 b15zdnd11an1n04x5 FILLER_102_451 ();
 b15zdnd00an1n02x5 FILLER_102_455 ();
 b15zdnd00an1n01x5 FILLER_102_457 ();
 b15zdnd11an1n64x5 FILLER_102_478 ();
 b15zdnd11an1n64x5 FILLER_102_542 ();
 b15zdnd11an1n16x5 FILLER_102_606 ();
 b15zdnd00an1n01x5 FILLER_102_622 ();
 b15zdnd11an1n32x5 FILLER_102_675 ();
 b15zdnd11an1n08x5 FILLER_102_707 ();
 b15zdnd00an1n02x5 FILLER_102_715 ();
 b15zdnd00an1n01x5 FILLER_102_717 ();
 b15zdnd11an1n64x5 FILLER_102_726 ();
 b15zdnd11an1n32x5 FILLER_102_790 ();
 b15zdnd11an1n16x5 FILLER_102_822 ();
 b15zdnd11an1n08x5 FILLER_102_838 ();
 b15zdnd00an1n02x5 FILLER_102_846 ();
 b15zdnd00an1n01x5 FILLER_102_848 ();
 b15zdnd11an1n64x5 FILLER_102_858 ();
 b15zdnd11an1n64x5 FILLER_102_922 ();
 b15zdnd11an1n32x5 FILLER_102_986 ();
 b15zdnd11an1n04x5 FILLER_102_1018 ();
 b15zdnd00an1n01x5 FILLER_102_1022 ();
 b15zdnd11an1n16x5 FILLER_102_1037 ();
 b15zdnd11an1n04x5 FILLER_102_1053 ();
 b15zdnd00an1n02x5 FILLER_102_1057 ();
 b15zdnd11an1n64x5 FILLER_102_1062 ();
 b15zdnd11an1n64x5 FILLER_102_1126 ();
 b15zdnd11an1n64x5 FILLER_102_1190 ();
 b15zdnd11an1n08x5 FILLER_102_1254 ();
 b15zdnd11an1n04x5 FILLER_102_1262 ();
 b15zdnd00an1n02x5 FILLER_102_1266 ();
 b15zdnd00an1n01x5 FILLER_102_1268 ();
 b15zdnd11an1n64x5 FILLER_102_1278 ();
 b15zdnd11an1n64x5 FILLER_102_1342 ();
 b15zdnd11an1n32x5 FILLER_102_1406 ();
 b15zdnd11an1n04x5 FILLER_102_1438 ();
 b15zdnd11an1n08x5 FILLER_102_1469 ();
 b15zdnd00an1n02x5 FILLER_102_1477 ();
 b15zdnd00an1n01x5 FILLER_102_1479 ();
 b15zdnd11an1n64x5 FILLER_102_1483 ();
 b15zdnd11an1n64x5 FILLER_102_1547 ();
 b15zdnd11an1n16x5 FILLER_102_1611 ();
 b15zdnd11an1n08x5 FILLER_102_1627 ();
 b15zdnd00an1n02x5 FILLER_102_1635 ();
 b15zdnd11an1n64x5 FILLER_102_1657 ();
 b15zdnd11an1n32x5 FILLER_102_1721 ();
 b15zdnd11an1n16x5 FILLER_102_1753 ();
 b15zdnd11an1n16x5 FILLER_102_1789 ();
 b15zdnd11an1n08x5 FILLER_102_1805 ();
 b15zdnd00an1n02x5 FILLER_102_1813 ();
 b15zdnd00an1n01x5 FILLER_102_1815 ();
 b15zdnd11an1n64x5 FILLER_102_1833 ();
 b15zdnd11an1n64x5 FILLER_102_1897 ();
 b15zdnd11an1n64x5 FILLER_102_1961 ();
 b15zdnd11an1n04x5 FILLER_102_2025 ();
 b15zdnd00an1n02x5 FILLER_102_2029 ();
 b15zdnd00an1n01x5 FILLER_102_2031 ();
 b15zdnd11an1n04x5 FILLER_102_2035 ();
 b15zdnd11an1n64x5 FILLER_102_2042 ();
 b15zdnd11an1n32x5 FILLER_102_2106 ();
 b15zdnd11an1n16x5 FILLER_102_2138 ();
 b15zdnd11an1n64x5 FILLER_102_2162 ();
 b15zdnd11an1n32x5 FILLER_102_2226 ();
 b15zdnd11an1n16x5 FILLER_102_2258 ();
 b15zdnd00an1n02x5 FILLER_102_2274 ();
 b15zdnd11an1n16x5 FILLER_103_0 ();
 b15zdnd11an1n08x5 FILLER_103_16 ();
 b15zdnd00an1n02x5 FILLER_103_24 ();
 b15zdnd11an1n64x5 FILLER_103_29 ();
 b15zdnd11an1n64x5 FILLER_103_93 ();
 b15zdnd11an1n16x5 FILLER_103_157 ();
 b15zdnd11an1n04x5 FILLER_103_173 ();
 b15zdnd00an1n02x5 FILLER_103_177 ();
 b15zdnd00an1n01x5 FILLER_103_179 ();
 b15zdnd11an1n08x5 FILLER_103_232 ();
 b15zdnd11an1n16x5 FILLER_103_292 ();
 b15zdnd11an1n04x5 FILLER_103_308 ();
 b15zdnd00an1n02x5 FILLER_103_312 ();
 b15zdnd11an1n64x5 FILLER_103_366 ();
 b15zdnd11an1n64x5 FILLER_103_430 ();
 b15zdnd00an1n02x5 FILLER_103_494 ();
 b15zdnd11an1n64x5 FILLER_103_499 ();
 b15zdnd11an1n64x5 FILLER_103_563 ();
 b15zdnd11an1n08x5 FILLER_103_627 ();
 b15zdnd11an1n04x5 FILLER_103_635 ();
 b15zdnd00an1n02x5 FILLER_103_639 ();
 b15zdnd11an1n04x5 FILLER_103_644 ();
 b15zdnd00an1n01x5 FILLER_103_648 ();
 b15zdnd11an1n16x5 FILLER_103_652 ();
 b15zdnd11an1n08x5 FILLER_103_668 ();
 b15zdnd11an1n64x5 FILLER_103_696 ();
 b15zdnd11an1n64x5 FILLER_103_760 ();
 b15zdnd11an1n64x5 FILLER_103_824 ();
 b15zdnd11an1n32x5 FILLER_103_888 ();
 b15zdnd11an1n16x5 FILLER_103_920 ();
 b15zdnd00an1n02x5 FILLER_103_936 ();
 b15zdnd11an1n64x5 FILLER_103_941 ();
 b15zdnd11an1n32x5 FILLER_103_1005 ();
 b15zdnd11an1n08x5 FILLER_103_1037 ();
 b15zdnd00an1n02x5 FILLER_103_1045 ();
 b15zdnd00an1n01x5 FILLER_103_1047 ();
 b15zdnd11an1n64x5 FILLER_103_1090 ();
 b15zdnd11an1n64x5 FILLER_103_1154 ();
 b15zdnd11an1n64x5 FILLER_103_1218 ();
 b15zdnd11an1n64x5 FILLER_103_1282 ();
 b15zdnd11an1n64x5 FILLER_103_1346 ();
 b15zdnd11an1n32x5 FILLER_103_1410 ();
 b15zdnd11an1n08x5 FILLER_103_1442 ();
 b15zdnd00an1n02x5 FILLER_103_1450 ();
 b15zdnd00an1n01x5 FILLER_103_1452 ();
 b15zdnd11an1n64x5 FILLER_103_1505 ();
 b15zdnd11an1n64x5 FILLER_103_1569 ();
 b15zdnd11an1n64x5 FILLER_103_1633 ();
 b15zdnd11an1n64x5 FILLER_103_1697 ();
 b15zdnd11an1n04x5 FILLER_103_1761 ();
 b15zdnd00an1n02x5 FILLER_103_1765 ();
 b15zdnd11an1n64x5 FILLER_103_1781 ();
 b15zdnd11an1n64x5 FILLER_103_1845 ();
 b15zdnd11an1n64x5 FILLER_103_1909 ();
 b15zdnd11an1n64x5 FILLER_103_1973 ();
 b15zdnd11an1n64x5 FILLER_103_2037 ();
 b15zdnd11an1n64x5 FILLER_103_2101 ();
 b15zdnd11an1n64x5 FILLER_103_2165 ();
 b15zdnd11an1n32x5 FILLER_103_2229 ();
 b15zdnd11an1n16x5 FILLER_103_2261 ();
 b15zdnd11an1n04x5 FILLER_103_2277 ();
 b15zdnd00an1n02x5 FILLER_103_2281 ();
 b15zdnd00an1n01x5 FILLER_103_2283 ();
 b15zdnd11an1n64x5 FILLER_104_8 ();
 b15zdnd11an1n64x5 FILLER_104_72 ();
 b15zdnd11an1n64x5 FILLER_104_136 ();
 b15zdnd11an1n04x5 FILLER_104_200 ();
 b15zdnd00an1n02x5 FILLER_104_204 ();
 b15zdnd11an1n32x5 FILLER_104_209 ();
 b15zdnd11an1n16x5 FILLER_104_241 ();
 b15zdnd11an1n04x5 FILLER_104_257 ();
 b15zdnd00an1n02x5 FILLER_104_261 ();
 b15zdnd11an1n04x5 FILLER_104_266 ();
 b15zdnd11an1n32x5 FILLER_104_273 ();
 b15zdnd11an1n16x5 FILLER_104_305 ();
 b15zdnd11an1n08x5 FILLER_104_321 ();
 b15zdnd11an1n04x5 FILLER_104_329 ();
 b15zdnd00an1n01x5 FILLER_104_333 ();
 b15zdnd11an1n04x5 FILLER_104_337 ();
 b15zdnd11an1n64x5 FILLER_104_344 ();
 b15zdnd11an1n32x5 FILLER_104_408 ();
 b15zdnd11an1n16x5 FILLER_104_440 ();
 b15zdnd11an1n08x5 FILLER_104_456 ();
 b15zdnd11an1n04x5 FILLER_104_464 ();
 b15zdnd00an1n01x5 FILLER_104_468 ();
 b15zdnd11an1n16x5 FILLER_104_521 ();
 b15zdnd11an1n04x5 FILLER_104_537 ();
 b15zdnd00an1n02x5 FILLER_104_541 ();
 b15zdnd11an1n64x5 FILLER_104_567 ();
 b15zdnd11an1n64x5 FILLER_104_631 ();
 b15zdnd11an1n16x5 FILLER_104_695 ();
 b15zdnd11an1n04x5 FILLER_104_711 ();
 b15zdnd00an1n02x5 FILLER_104_715 ();
 b15zdnd00an1n01x5 FILLER_104_717 ();
 b15zdnd11an1n64x5 FILLER_104_726 ();
 b15zdnd11an1n64x5 FILLER_104_790 ();
 b15zdnd11an1n32x5 FILLER_104_854 ();
 b15zdnd11an1n16x5 FILLER_104_886 ();
 b15zdnd11an1n08x5 FILLER_104_902 ();
 b15zdnd11an1n04x5 FILLER_104_910 ();
 b15zdnd00an1n01x5 FILLER_104_914 ();
 b15zdnd11an1n64x5 FILLER_104_967 ();
 b15zdnd00an1n01x5 FILLER_104_1031 ();
 b15zdnd11an1n64x5 FILLER_104_1084 ();
 b15zdnd11an1n64x5 FILLER_104_1148 ();
 b15zdnd11an1n32x5 FILLER_104_1212 ();
 b15zdnd11an1n08x5 FILLER_104_1244 ();
 b15zdnd00an1n01x5 FILLER_104_1252 ();
 b15zdnd11an1n64x5 FILLER_104_1258 ();
 b15zdnd11an1n64x5 FILLER_104_1322 ();
 b15zdnd11an1n32x5 FILLER_104_1386 ();
 b15zdnd11an1n16x5 FILLER_104_1418 ();
 b15zdnd00an1n02x5 FILLER_104_1434 ();
 b15zdnd00an1n01x5 FILLER_104_1436 ();
 b15zdnd11an1n16x5 FILLER_104_1440 ();
 b15zdnd11an1n08x5 FILLER_104_1456 ();
 b15zdnd11an1n04x5 FILLER_104_1464 ();
 b15zdnd00an1n02x5 FILLER_104_1468 ();
 b15zdnd11an1n08x5 FILLER_104_1473 ();
 b15zdnd00an1n01x5 FILLER_104_1481 ();
 b15zdnd11an1n64x5 FILLER_104_1485 ();
 b15zdnd11an1n16x5 FILLER_104_1549 ();
 b15zdnd11an1n64x5 FILLER_104_1617 ();
 b15zdnd11an1n64x5 FILLER_104_1681 ();
 b15zdnd11an1n64x5 FILLER_104_1745 ();
 b15zdnd11an1n64x5 FILLER_104_1809 ();
 b15zdnd11an1n32x5 FILLER_104_1873 ();
 b15zdnd11an1n04x5 FILLER_104_1905 ();
 b15zdnd11an1n04x5 FILLER_104_1912 ();
 b15zdnd11an1n64x5 FILLER_104_1919 ();
 b15zdnd11an1n64x5 FILLER_104_1983 ();
 b15zdnd11an1n64x5 FILLER_104_2047 ();
 b15zdnd11an1n32x5 FILLER_104_2111 ();
 b15zdnd11an1n08x5 FILLER_104_2143 ();
 b15zdnd00an1n02x5 FILLER_104_2151 ();
 b15zdnd00an1n01x5 FILLER_104_2153 ();
 b15zdnd11an1n64x5 FILLER_104_2162 ();
 b15zdnd11an1n32x5 FILLER_104_2226 ();
 b15zdnd11an1n16x5 FILLER_104_2258 ();
 b15zdnd00an1n02x5 FILLER_104_2274 ();
 b15zdnd11an1n64x5 FILLER_105_0 ();
 b15zdnd11an1n64x5 FILLER_105_64 ();
 b15zdnd11an1n64x5 FILLER_105_128 ();
 b15zdnd11an1n64x5 FILLER_105_192 ();
 b15zdnd11an1n64x5 FILLER_105_256 ();
 b15zdnd11an1n16x5 FILLER_105_320 ();
 b15zdnd11an1n04x5 FILLER_105_336 ();
 b15zdnd00an1n01x5 FILLER_105_340 ();
 b15zdnd11an1n64x5 FILLER_105_344 ();
 b15zdnd11an1n64x5 FILLER_105_408 ();
 b15zdnd00an1n02x5 FILLER_105_472 ();
 b15zdnd00an1n01x5 FILLER_105_474 ();
 b15zdnd11an1n32x5 FILLER_105_527 ();
 b15zdnd11an1n04x5 FILLER_105_559 ();
 b15zdnd11an1n64x5 FILLER_105_566 ();
 b15zdnd11an1n64x5 FILLER_105_630 ();
 b15zdnd11an1n64x5 FILLER_105_694 ();
 b15zdnd11an1n32x5 FILLER_105_758 ();
 b15zdnd11an1n04x5 FILLER_105_790 ();
 b15zdnd00an1n01x5 FILLER_105_794 ();
 b15zdnd11an1n04x5 FILLER_105_847 ();
 b15zdnd11an1n64x5 FILLER_105_862 ();
 b15zdnd11an1n04x5 FILLER_105_926 ();
 b15zdnd00an1n02x5 FILLER_105_930 ();
 b15zdnd00an1n01x5 FILLER_105_932 ();
 b15zdnd11an1n04x5 FILLER_105_936 ();
 b15zdnd11an1n08x5 FILLER_105_943 ();
 b15zdnd11an1n04x5 FILLER_105_951 ();
 b15zdnd00an1n02x5 FILLER_105_955 ();
 b15zdnd00an1n01x5 FILLER_105_957 ();
 b15zdnd11an1n64x5 FILLER_105_972 ();
 b15zdnd11an1n16x5 FILLER_105_1036 ();
 b15zdnd11an1n04x5 FILLER_105_1052 ();
 b15zdnd00an1n02x5 FILLER_105_1056 ();
 b15zdnd11an1n04x5 FILLER_105_1061 ();
 b15zdnd11an1n64x5 FILLER_105_1068 ();
 b15zdnd11an1n64x5 FILLER_105_1132 ();
 b15zdnd11an1n64x5 FILLER_105_1196 ();
 b15zdnd11an1n32x5 FILLER_105_1260 ();
 b15zdnd00an1n02x5 FILLER_105_1292 ();
 b15zdnd11an1n64x5 FILLER_105_1310 ();
 b15zdnd11an1n64x5 FILLER_105_1374 ();
 b15zdnd11an1n64x5 FILLER_105_1438 ();
 b15zdnd11an1n32x5 FILLER_105_1502 ();
 b15zdnd00an1n02x5 FILLER_105_1534 ();
 b15zdnd11an1n32x5 FILLER_105_1539 ();
 b15zdnd11an1n16x5 FILLER_105_1571 ();
 b15zdnd11an1n04x5 FILLER_105_1587 ();
 b15zdnd00an1n02x5 FILLER_105_1591 ();
 b15zdnd11an1n64x5 FILLER_105_1596 ();
 b15zdnd11an1n32x5 FILLER_105_1660 ();
 b15zdnd11an1n08x5 FILLER_105_1692 ();
 b15zdnd11an1n04x5 FILLER_105_1700 ();
 b15zdnd00an1n02x5 FILLER_105_1704 ();
 b15zdnd00an1n01x5 FILLER_105_1706 ();
 b15zdnd11an1n04x5 FILLER_105_1721 ();
 b15zdnd11an1n04x5 FILLER_105_1745 ();
 b15zdnd00an1n02x5 FILLER_105_1749 ();
 b15zdnd11an1n64x5 FILLER_105_1768 ();
 b15zdnd11an1n32x5 FILLER_105_1832 ();
 b15zdnd11an1n16x5 FILLER_105_1864 ();
 b15zdnd11an1n08x5 FILLER_105_1880 ();
 b15zdnd00an1n02x5 FILLER_105_1888 ();
 b15zdnd00an1n01x5 FILLER_105_1890 ();
 b15zdnd11an1n64x5 FILLER_105_1943 ();
 b15zdnd11an1n64x5 FILLER_105_2007 ();
 b15zdnd11an1n64x5 FILLER_105_2071 ();
 b15zdnd11an1n64x5 FILLER_105_2135 ();
 b15zdnd11an1n64x5 FILLER_105_2199 ();
 b15zdnd11an1n16x5 FILLER_105_2263 ();
 b15zdnd11an1n04x5 FILLER_105_2279 ();
 b15zdnd00an1n01x5 FILLER_105_2283 ();
 b15zdnd11an1n64x5 FILLER_106_8 ();
 b15zdnd11an1n64x5 FILLER_106_72 ();
 b15zdnd11an1n64x5 FILLER_106_136 ();
 b15zdnd11an1n64x5 FILLER_106_200 ();
 b15zdnd11an1n64x5 FILLER_106_264 ();
 b15zdnd11an1n64x5 FILLER_106_328 ();
 b15zdnd11an1n64x5 FILLER_106_392 ();
 b15zdnd11an1n32x5 FILLER_106_456 ();
 b15zdnd11an1n04x5 FILLER_106_491 ();
 b15zdnd11an1n04x5 FILLER_106_498 ();
 b15zdnd11an1n04x5 FILLER_106_505 ();
 b15zdnd11an1n16x5 FILLER_106_512 ();
 b15zdnd11an1n08x5 FILLER_106_528 ();
 b15zdnd11an1n64x5 FILLER_106_588 ();
 b15zdnd11an1n64x5 FILLER_106_652 ();
 b15zdnd00an1n02x5 FILLER_106_716 ();
 b15zdnd11an1n64x5 FILLER_106_726 ();
 b15zdnd11an1n04x5 FILLER_106_790 ();
 b15zdnd00an1n01x5 FILLER_106_794 ();
 b15zdnd11an1n08x5 FILLER_106_806 ();
 b15zdnd00an1n02x5 FILLER_106_814 ();
 b15zdnd11an1n04x5 FILLER_106_819 ();
 b15zdnd11an1n64x5 FILLER_106_826 ();
 b15zdnd11an1n32x5 FILLER_106_890 ();
 b15zdnd11an1n64x5 FILLER_106_936 ();
 b15zdnd11an1n64x5 FILLER_106_1000 ();
 b15zdnd11an1n64x5 FILLER_106_1064 ();
 b15zdnd11an1n64x5 FILLER_106_1128 ();
 b15zdnd11an1n64x5 FILLER_106_1192 ();
 b15zdnd11an1n16x5 FILLER_106_1256 ();
 b15zdnd11an1n08x5 FILLER_106_1272 ();
 b15zdnd00an1n01x5 FILLER_106_1280 ();
 b15zdnd11an1n64x5 FILLER_106_1286 ();
 b15zdnd11an1n64x5 FILLER_106_1350 ();
 b15zdnd11an1n64x5 FILLER_106_1414 ();
 b15zdnd11an1n32x5 FILLER_106_1478 ();
 b15zdnd11an1n04x5 FILLER_106_1510 ();
 b15zdnd00an1n01x5 FILLER_106_1514 ();
 b15zdnd11an1n08x5 FILLER_106_1567 ();
 b15zdnd00an1n02x5 FILLER_106_1575 ();
 b15zdnd00an1n01x5 FILLER_106_1577 ();
 b15zdnd11an1n08x5 FILLER_106_1581 ();
 b15zdnd11an1n04x5 FILLER_106_1589 ();
 b15zdnd00an1n01x5 FILLER_106_1593 ();
 b15zdnd11an1n64x5 FILLER_106_1597 ();
 b15zdnd11an1n16x5 FILLER_106_1661 ();
 b15zdnd00an1n01x5 FILLER_106_1677 ();
 b15zdnd11an1n32x5 FILLER_106_1698 ();
 b15zdnd00an1n02x5 FILLER_106_1730 ();
 b15zdnd11an1n08x5 FILLER_106_1746 ();
 b15zdnd11an1n04x5 FILLER_106_1754 ();
 b15zdnd00an1n02x5 FILLER_106_1758 ();
 b15zdnd11an1n64x5 FILLER_106_1777 ();
 b15zdnd11an1n64x5 FILLER_106_1841 ();
 b15zdnd11an1n08x5 FILLER_106_1905 ();
 b15zdnd00an1n02x5 FILLER_106_1913 ();
 b15zdnd00an1n01x5 FILLER_106_1915 ();
 b15zdnd11an1n64x5 FILLER_106_1919 ();
 b15zdnd11an1n64x5 FILLER_106_1983 ();
 b15zdnd11an1n64x5 FILLER_106_2047 ();
 b15zdnd11an1n32x5 FILLER_106_2111 ();
 b15zdnd11an1n08x5 FILLER_106_2143 ();
 b15zdnd00an1n02x5 FILLER_106_2151 ();
 b15zdnd00an1n01x5 FILLER_106_2153 ();
 b15zdnd11an1n64x5 FILLER_106_2162 ();
 b15zdnd11an1n32x5 FILLER_106_2226 ();
 b15zdnd11an1n16x5 FILLER_106_2258 ();
 b15zdnd00an1n02x5 FILLER_106_2274 ();
 b15zdnd11an1n64x5 FILLER_107_0 ();
 b15zdnd11an1n64x5 FILLER_107_64 ();
 b15zdnd11an1n64x5 FILLER_107_128 ();
 b15zdnd11an1n64x5 FILLER_107_192 ();
 b15zdnd11an1n64x5 FILLER_107_256 ();
 b15zdnd11an1n64x5 FILLER_107_320 ();
 b15zdnd11an1n64x5 FILLER_107_384 ();
 b15zdnd11an1n32x5 FILLER_107_448 ();
 b15zdnd11an1n08x5 FILLER_107_480 ();
 b15zdnd11an1n04x5 FILLER_107_488 ();
 b15zdnd00an1n02x5 FILLER_107_492 ();
 b15zdnd11an1n32x5 FILLER_107_497 ();
 b15zdnd11an1n16x5 FILLER_107_529 ();
 b15zdnd11an1n08x5 FILLER_107_545 ();
 b15zdnd00an1n01x5 FILLER_107_553 ();
 b15zdnd11an1n04x5 FILLER_107_557 ();
 b15zdnd11an1n64x5 FILLER_107_564 ();
 b15zdnd11an1n64x5 FILLER_107_628 ();
 b15zdnd11an1n64x5 FILLER_107_692 ();
 b15zdnd11an1n32x5 FILLER_107_756 ();
 b15zdnd11an1n16x5 FILLER_107_788 ();
 b15zdnd11an1n08x5 FILLER_107_804 ();
 b15zdnd11an1n04x5 FILLER_107_812 ();
 b15zdnd00an1n02x5 FILLER_107_816 ();
 b15zdnd11an1n04x5 FILLER_107_821 ();
 b15zdnd11an1n64x5 FILLER_107_833 ();
 b15zdnd11an1n64x5 FILLER_107_897 ();
 b15zdnd11an1n64x5 FILLER_107_961 ();
 b15zdnd11an1n64x5 FILLER_107_1025 ();
 b15zdnd11an1n64x5 FILLER_107_1089 ();
 b15zdnd11an1n64x5 FILLER_107_1153 ();
 b15zdnd11an1n64x5 FILLER_107_1217 ();
 b15zdnd11an1n64x5 FILLER_107_1281 ();
 b15zdnd11an1n64x5 FILLER_107_1345 ();
 b15zdnd11an1n64x5 FILLER_107_1409 ();
 b15zdnd11an1n32x5 FILLER_107_1473 ();
 b15zdnd11an1n16x5 FILLER_107_1505 ();
 b15zdnd11an1n08x5 FILLER_107_1521 ();
 b15zdnd11an1n04x5 FILLER_107_1529 ();
 b15zdnd11an1n04x5 FILLER_107_1536 ();
 b15zdnd11an1n32x5 FILLER_107_1543 ();
 b15zdnd11an1n04x5 FILLER_107_1575 ();
 b15zdnd00an1n02x5 FILLER_107_1579 ();
 b15zdnd11an1n64x5 FILLER_107_1595 ();
 b15zdnd11an1n04x5 FILLER_107_1659 ();
 b15zdnd00an1n02x5 FILLER_107_1663 ();
 b15zdnd11an1n64x5 FILLER_107_1679 ();
 b15zdnd11an1n64x5 FILLER_107_1743 ();
 b15zdnd11an1n64x5 FILLER_107_1807 ();
 b15zdnd11an1n64x5 FILLER_107_1871 ();
 b15zdnd11an1n16x5 FILLER_107_1935 ();
 b15zdnd11an1n08x5 FILLER_107_1951 ();
 b15zdnd00an1n01x5 FILLER_107_1959 ();
 b15zdnd11an1n16x5 FILLER_107_1969 ();
 b15zdnd00an1n02x5 FILLER_107_1985 ();
 b15zdnd00an1n01x5 FILLER_107_1987 ();
 b15zdnd11an1n64x5 FILLER_107_1997 ();
 b15zdnd11an1n64x5 FILLER_107_2061 ();
 b15zdnd11an1n64x5 FILLER_107_2125 ();
 b15zdnd11an1n64x5 FILLER_107_2189 ();
 b15zdnd11an1n16x5 FILLER_107_2253 ();
 b15zdnd11an1n08x5 FILLER_107_2269 ();
 b15zdnd11an1n04x5 FILLER_107_2277 ();
 b15zdnd00an1n02x5 FILLER_107_2281 ();
 b15zdnd00an1n01x5 FILLER_107_2283 ();
 b15zdnd11an1n16x5 FILLER_108_8 ();
 b15zdnd11an1n04x5 FILLER_108_24 ();
 b15zdnd11an1n64x5 FILLER_108_38 ();
 b15zdnd11an1n64x5 FILLER_108_102 ();
 b15zdnd11an1n64x5 FILLER_108_166 ();
 b15zdnd11an1n64x5 FILLER_108_230 ();
 b15zdnd11an1n64x5 FILLER_108_294 ();
 b15zdnd11an1n64x5 FILLER_108_358 ();
 b15zdnd11an1n64x5 FILLER_108_422 ();
 b15zdnd11an1n64x5 FILLER_108_486 ();
 b15zdnd11an1n64x5 FILLER_108_550 ();
 b15zdnd11an1n64x5 FILLER_108_614 ();
 b15zdnd11an1n32x5 FILLER_108_678 ();
 b15zdnd11an1n08x5 FILLER_108_710 ();
 b15zdnd11an1n08x5 FILLER_108_726 ();
 b15zdnd11an1n04x5 FILLER_108_734 ();
 b15zdnd00an1n01x5 FILLER_108_738 ();
 b15zdnd11an1n32x5 FILLER_108_763 ();
 b15zdnd11an1n16x5 FILLER_108_795 ();
 b15zdnd11an1n08x5 FILLER_108_811 ();
 b15zdnd00an1n02x5 FILLER_108_819 ();
 b15zdnd00an1n01x5 FILLER_108_821 ();
 b15zdnd11an1n08x5 FILLER_108_825 ();
 b15zdnd11an1n64x5 FILLER_108_836 ();
 b15zdnd11an1n16x5 FILLER_108_900 ();
 b15zdnd11an1n04x5 FILLER_108_916 ();
 b15zdnd00an1n02x5 FILLER_108_920 ();
 b15zdnd11an1n04x5 FILLER_108_925 ();
 b15zdnd00an1n02x5 FILLER_108_929 ();
 b15zdnd00an1n01x5 FILLER_108_931 ();
 b15zdnd11an1n64x5 FILLER_108_935 ();
 b15zdnd11an1n64x5 FILLER_108_999 ();
 b15zdnd11an1n64x5 FILLER_108_1063 ();
 b15zdnd11an1n64x5 FILLER_108_1127 ();
 b15zdnd11an1n64x5 FILLER_108_1191 ();
 b15zdnd11an1n64x5 FILLER_108_1255 ();
 b15zdnd11an1n16x5 FILLER_108_1319 ();
 b15zdnd00an1n02x5 FILLER_108_1335 ();
 b15zdnd11an1n64x5 FILLER_108_1340 ();
 b15zdnd11an1n64x5 FILLER_108_1404 ();
 b15zdnd11an1n64x5 FILLER_108_1468 ();
 b15zdnd11an1n64x5 FILLER_108_1532 ();
 b15zdnd11an1n16x5 FILLER_108_1596 ();
 b15zdnd11an1n04x5 FILLER_108_1612 ();
 b15zdnd00an1n02x5 FILLER_108_1616 ();
 b15zdnd11an1n04x5 FILLER_108_1635 ();
 b15zdnd11an1n64x5 FILLER_108_1653 ();
 b15zdnd11an1n64x5 FILLER_108_1717 ();
 b15zdnd11an1n64x5 FILLER_108_1781 ();
 b15zdnd11an1n64x5 FILLER_108_1845 ();
 b15zdnd11an1n64x5 FILLER_108_1909 ();
 b15zdnd11an1n64x5 FILLER_108_1973 ();
 b15zdnd11an1n64x5 FILLER_108_2037 ();
 b15zdnd11an1n32x5 FILLER_108_2101 ();
 b15zdnd11an1n16x5 FILLER_108_2133 ();
 b15zdnd11an1n04x5 FILLER_108_2149 ();
 b15zdnd00an1n01x5 FILLER_108_2153 ();
 b15zdnd11an1n64x5 FILLER_108_2162 ();
 b15zdnd11an1n32x5 FILLER_108_2226 ();
 b15zdnd11an1n16x5 FILLER_108_2258 ();
 b15zdnd00an1n02x5 FILLER_108_2274 ();
 b15zdnd11an1n32x5 FILLER_109_0 ();
 b15zdnd11an1n08x5 FILLER_109_32 ();
 b15zdnd11an1n04x5 FILLER_109_40 ();
 b15zdnd00an1n02x5 FILLER_109_44 ();
 b15zdnd00an1n01x5 FILLER_109_46 ();
 b15zdnd11an1n04x5 FILLER_109_53 ();
 b15zdnd11an1n64x5 FILLER_109_63 ();
 b15zdnd11an1n64x5 FILLER_109_127 ();
 b15zdnd11an1n64x5 FILLER_109_191 ();
 b15zdnd11an1n64x5 FILLER_109_255 ();
 b15zdnd11an1n64x5 FILLER_109_319 ();
 b15zdnd11an1n64x5 FILLER_109_383 ();
 b15zdnd11an1n64x5 FILLER_109_447 ();
 b15zdnd11an1n64x5 FILLER_109_511 ();
 b15zdnd11an1n64x5 FILLER_109_575 ();
 b15zdnd11an1n64x5 FILLER_109_639 ();
 b15zdnd11an1n32x5 FILLER_109_703 ();
 b15zdnd11an1n04x5 FILLER_109_735 ();
 b15zdnd00an1n02x5 FILLER_109_739 ();
 b15zdnd00an1n01x5 FILLER_109_741 ();
 b15zdnd11an1n32x5 FILLER_109_762 ();
 b15zdnd11an1n04x5 FILLER_109_794 ();
 b15zdnd00an1n01x5 FILLER_109_798 ();
 b15zdnd11an1n32x5 FILLER_109_851 ();
 b15zdnd00an1n02x5 FILLER_109_883 ();
 b15zdnd11an1n64x5 FILLER_109_937 ();
 b15zdnd11an1n64x5 FILLER_109_1001 ();
 b15zdnd11an1n64x5 FILLER_109_1065 ();
 b15zdnd11an1n64x5 FILLER_109_1129 ();
 b15zdnd11an1n32x5 FILLER_109_1193 ();
 b15zdnd11an1n16x5 FILLER_109_1225 ();
 b15zdnd11an1n08x5 FILLER_109_1241 ();
 b15zdnd11an1n04x5 FILLER_109_1249 ();
 b15zdnd00an1n02x5 FILLER_109_1253 ();
 b15zdnd11an1n32x5 FILLER_109_1264 ();
 b15zdnd11an1n08x5 FILLER_109_1296 ();
 b15zdnd11an1n04x5 FILLER_109_1304 ();
 b15zdnd00an1n02x5 FILLER_109_1308 ();
 b15zdnd00an1n01x5 FILLER_109_1310 ();
 b15zdnd11an1n64x5 FILLER_109_1363 ();
 b15zdnd11an1n64x5 FILLER_109_1427 ();
 b15zdnd11an1n64x5 FILLER_109_1491 ();
 b15zdnd11an1n08x5 FILLER_109_1555 ();
 b15zdnd11an1n64x5 FILLER_109_1571 ();
 b15zdnd11an1n64x5 FILLER_109_1635 ();
 b15zdnd11an1n64x5 FILLER_109_1699 ();
 b15zdnd11an1n16x5 FILLER_109_1763 ();
 b15zdnd11an1n04x5 FILLER_109_1779 ();
 b15zdnd00an1n02x5 FILLER_109_1783 ();
 b15zdnd11an1n64x5 FILLER_109_1799 ();
 b15zdnd11an1n64x5 FILLER_109_1863 ();
 b15zdnd11an1n64x5 FILLER_109_1927 ();
 b15zdnd11an1n64x5 FILLER_109_1991 ();
 b15zdnd11an1n64x5 FILLER_109_2055 ();
 b15zdnd11an1n64x5 FILLER_109_2119 ();
 b15zdnd11an1n64x5 FILLER_109_2183 ();
 b15zdnd11an1n32x5 FILLER_109_2247 ();
 b15zdnd11an1n04x5 FILLER_109_2279 ();
 b15zdnd00an1n01x5 FILLER_109_2283 ();
 b15zdnd11an1n32x5 FILLER_110_8 ();
 b15zdnd11an1n08x5 FILLER_110_40 ();
 b15zdnd11an1n04x5 FILLER_110_48 ();
 b15zdnd11an1n04x5 FILLER_110_61 ();
 b15zdnd11an1n64x5 FILLER_110_71 ();
 b15zdnd11an1n64x5 FILLER_110_135 ();
 b15zdnd11an1n64x5 FILLER_110_199 ();
 b15zdnd11an1n64x5 FILLER_110_263 ();
 b15zdnd11an1n64x5 FILLER_110_327 ();
 b15zdnd11an1n64x5 FILLER_110_391 ();
 b15zdnd11an1n64x5 FILLER_110_455 ();
 b15zdnd11an1n32x5 FILLER_110_519 ();
 b15zdnd11an1n16x5 FILLER_110_551 ();
 b15zdnd11an1n04x5 FILLER_110_567 ();
 b15zdnd11an1n64x5 FILLER_110_591 ();
 b15zdnd11an1n32x5 FILLER_110_655 ();
 b15zdnd11an1n16x5 FILLER_110_687 ();
 b15zdnd11an1n08x5 FILLER_110_703 ();
 b15zdnd11an1n04x5 FILLER_110_711 ();
 b15zdnd00an1n02x5 FILLER_110_715 ();
 b15zdnd00an1n01x5 FILLER_110_717 ();
 b15zdnd11an1n64x5 FILLER_110_726 ();
 b15zdnd11an1n32x5 FILLER_110_790 ();
 b15zdnd00an1n02x5 FILLER_110_822 ();
 b15zdnd11an1n04x5 FILLER_110_827 ();
 b15zdnd11an1n08x5 FILLER_110_839 ();
 b15zdnd11an1n64x5 FILLER_110_850 ();
 b15zdnd11an1n16x5 FILLER_110_914 ();
 b15zdnd11an1n04x5 FILLER_110_930 ();
 b15zdnd00an1n02x5 FILLER_110_934 ();
 b15zdnd11an1n04x5 FILLER_110_939 ();
 b15zdnd00an1n02x5 FILLER_110_943 ();
 b15zdnd11an1n64x5 FILLER_110_956 ();
 b15zdnd11an1n64x5 FILLER_110_1020 ();
 b15zdnd11an1n64x5 FILLER_110_1084 ();
 b15zdnd11an1n64x5 FILLER_110_1148 ();
 b15zdnd11an1n64x5 FILLER_110_1212 ();
 b15zdnd11an1n32x5 FILLER_110_1276 ();
 b15zdnd11an1n16x5 FILLER_110_1308 ();
 b15zdnd11an1n04x5 FILLER_110_1324 ();
 b15zdnd00an1n01x5 FILLER_110_1328 ();
 b15zdnd11an1n04x5 FILLER_110_1332 ();
 b15zdnd11an1n64x5 FILLER_110_1339 ();
 b15zdnd11an1n64x5 FILLER_110_1403 ();
 b15zdnd11an1n16x5 FILLER_110_1467 ();
 b15zdnd11an1n08x5 FILLER_110_1483 ();
 b15zdnd00an1n02x5 FILLER_110_1491 ();
 b15zdnd11an1n64x5 FILLER_110_1501 ();
 b15zdnd11an1n64x5 FILLER_110_1565 ();
 b15zdnd11an1n32x5 FILLER_110_1629 ();
 b15zdnd11an1n08x5 FILLER_110_1661 ();
 b15zdnd00an1n02x5 FILLER_110_1669 ();
 b15zdnd11an1n64x5 FILLER_110_1685 ();
 b15zdnd11an1n32x5 FILLER_110_1749 ();
 b15zdnd11an1n16x5 FILLER_110_1781 ();
 b15zdnd11an1n64x5 FILLER_110_1811 ();
 b15zdnd11an1n64x5 FILLER_110_1875 ();
 b15zdnd11an1n32x5 FILLER_110_1939 ();
 b15zdnd11an1n08x5 FILLER_110_1971 ();
 b15zdnd11an1n04x5 FILLER_110_1979 ();
 b15zdnd00an1n02x5 FILLER_110_1983 ();
 b15zdnd00an1n01x5 FILLER_110_1985 ();
 b15zdnd11an1n64x5 FILLER_110_1995 ();
 b15zdnd11an1n64x5 FILLER_110_2059 ();
 b15zdnd11an1n16x5 FILLER_110_2123 ();
 b15zdnd11an1n08x5 FILLER_110_2139 ();
 b15zdnd11an1n04x5 FILLER_110_2147 ();
 b15zdnd00an1n02x5 FILLER_110_2151 ();
 b15zdnd00an1n01x5 FILLER_110_2153 ();
 b15zdnd11an1n64x5 FILLER_110_2162 ();
 b15zdnd11an1n32x5 FILLER_110_2226 ();
 b15zdnd11an1n16x5 FILLER_110_2258 ();
 b15zdnd00an1n02x5 FILLER_110_2274 ();
 b15zdnd11an1n16x5 FILLER_111_0 ();
 b15zdnd00an1n02x5 FILLER_111_16 ();
 b15zdnd00an1n01x5 FILLER_111_18 ();
 b15zdnd11an1n64x5 FILLER_111_22 ();
 b15zdnd11an1n64x5 FILLER_111_86 ();
 b15zdnd11an1n64x5 FILLER_111_150 ();
 b15zdnd11an1n64x5 FILLER_111_214 ();
 b15zdnd11an1n64x5 FILLER_111_278 ();
 b15zdnd11an1n64x5 FILLER_111_342 ();
 b15zdnd11an1n64x5 FILLER_111_406 ();
 b15zdnd11an1n64x5 FILLER_111_470 ();
 b15zdnd11an1n64x5 FILLER_111_534 ();
 b15zdnd11an1n64x5 FILLER_111_598 ();
 b15zdnd11an1n64x5 FILLER_111_662 ();
 b15zdnd11an1n64x5 FILLER_111_726 ();
 b15zdnd11an1n32x5 FILLER_111_790 ();
 b15zdnd11an1n32x5 FILLER_111_874 ();
 b15zdnd11an1n08x5 FILLER_111_906 ();
 b15zdnd11an1n64x5 FILLER_111_925 ();
 b15zdnd11an1n64x5 FILLER_111_989 ();
 b15zdnd11an1n64x5 FILLER_111_1053 ();
 b15zdnd11an1n64x5 FILLER_111_1117 ();
 b15zdnd11an1n64x5 FILLER_111_1181 ();
 b15zdnd11an1n32x5 FILLER_111_1245 ();
 b15zdnd11an1n08x5 FILLER_111_1277 ();
 b15zdnd00an1n02x5 FILLER_111_1285 ();
 b15zdnd11an1n64x5 FILLER_111_1297 ();
 b15zdnd11an1n64x5 FILLER_111_1361 ();
 b15zdnd11an1n64x5 FILLER_111_1425 ();
 b15zdnd11an1n64x5 FILLER_111_1489 ();
 b15zdnd11an1n64x5 FILLER_111_1553 ();
 b15zdnd11an1n64x5 FILLER_111_1617 ();
 b15zdnd11an1n64x5 FILLER_111_1681 ();
 b15zdnd11an1n64x5 FILLER_111_1745 ();
 b15zdnd11an1n64x5 FILLER_111_1809 ();
 b15zdnd11an1n64x5 FILLER_111_1873 ();
 b15zdnd11an1n64x5 FILLER_111_1937 ();
 b15zdnd11an1n64x5 FILLER_111_2001 ();
 b15zdnd11an1n64x5 FILLER_111_2065 ();
 b15zdnd11an1n64x5 FILLER_111_2129 ();
 b15zdnd11an1n32x5 FILLER_111_2193 ();
 b15zdnd11an1n08x5 FILLER_111_2225 ();
 b15zdnd11an1n04x5 FILLER_111_2233 ();
 b15zdnd00an1n02x5 FILLER_111_2237 ();
 b15zdnd00an1n01x5 FILLER_111_2239 ();
 b15zdnd00an1n02x5 FILLER_111_2282 ();
 b15zdnd11an1n08x5 FILLER_112_8 ();
 b15zdnd11an1n04x5 FILLER_112_16 ();
 b15zdnd11an1n16x5 FILLER_112_23 ();
 b15zdnd11an1n08x5 FILLER_112_39 ();
 b15zdnd11an1n64x5 FILLER_112_58 ();
 b15zdnd11an1n64x5 FILLER_112_122 ();
 b15zdnd11an1n64x5 FILLER_112_186 ();
 b15zdnd11an1n32x5 FILLER_112_250 ();
 b15zdnd11an1n16x5 FILLER_112_282 ();
 b15zdnd11an1n04x5 FILLER_112_298 ();
 b15zdnd00an1n02x5 FILLER_112_302 ();
 b15zdnd00an1n01x5 FILLER_112_304 ();
 b15zdnd11an1n64x5 FILLER_112_316 ();
 b15zdnd11an1n64x5 FILLER_112_380 ();
 b15zdnd11an1n16x5 FILLER_112_444 ();
 b15zdnd00an1n02x5 FILLER_112_460 ();
 b15zdnd00an1n01x5 FILLER_112_462 ();
 b15zdnd11an1n64x5 FILLER_112_486 ();
 b15zdnd11an1n64x5 FILLER_112_550 ();
 b15zdnd11an1n64x5 FILLER_112_614 ();
 b15zdnd11an1n32x5 FILLER_112_678 ();
 b15zdnd11an1n08x5 FILLER_112_710 ();
 b15zdnd11an1n32x5 FILLER_112_726 ();
 b15zdnd11an1n08x5 FILLER_112_758 ();
 b15zdnd11an1n04x5 FILLER_112_766 ();
 b15zdnd00an1n01x5 FILLER_112_770 ();
 b15zdnd11an1n32x5 FILLER_112_780 ();
 b15zdnd11an1n08x5 FILLER_112_812 ();
 b15zdnd11an1n04x5 FILLER_112_820 ();
 b15zdnd00an1n01x5 FILLER_112_824 ();
 b15zdnd11an1n04x5 FILLER_112_839 ();
 b15zdnd00an1n02x5 FILLER_112_843 ();
 b15zdnd11an1n04x5 FILLER_112_848 ();
 b15zdnd11an1n64x5 FILLER_112_866 ();
 b15zdnd11an1n64x5 FILLER_112_930 ();
 b15zdnd11an1n64x5 FILLER_112_994 ();
 b15zdnd11an1n08x5 FILLER_112_1058 ();
 b15zdnd00an1n02x5 FILLER_112_1066 ();
 b15zdnd00an1n01x5 FILLER_112_1068 ();
 b15zdnd11an1n64x5 FILLER_112_1121 ();
 b15zdnd11an1n64x5 FILLER_112_1185 ();
 b15zdnd11an1n64x5 FILLER_112_1249 ();
 b15zdnd11an1n64x5 FILLER_112_1313 ();
 b15zdnd11an1n64x5 FILLER_112_1377 ();
 b15zdnd11an1n64x5 FILLER_112_1441 ();
 b15zdnd11an1n32x5 FILLER_112_1505 ();
 b15zdnd11an1n16x5 FILLER_112_1537 ();
 b15zdnd11an1n08x5 FILLER_112_1553 ();
 b15zdnd00an1n02x5 FILLER_112_1561 ();
 b15zdnd00an1n01x5 FILLER_112_1563 ();
 b15zdnd11an1n64x5 FILLER_112_1581 ();
 b15zdnd11an1n64x5 FILLER_112_1645 ();
 b15zdnd11an1n64x5 FILLER_112_1709 ();
 b15zdnd11an1n64x5 FILLER_112_1773 ();
 b15zdnd11an1n64x5 FILLER_112_1837 ();
 b15zdnd11an1n64x5 FILLER_112_1901 ();
 b15zdnd11an1n64x5 FILLER_112_1965 ();
 b15zdnd11an1n64x5 FILLER_112_2029 ();
 b15zdnd11an1n32x5 FILLER_112_2093 ();
 b15zdnd11an1n16x5 FILLER_112_2125 ();
 b15zdnd11an1n08x5 FILLER_112_2141 ();
 b15zdnd11an1n04x5 FILLER_112_2149 ();
 b15zdnd00an1n01x5 FILLER_112_2153 ();
 b15zdnd11an1n64x5 FILLER_112_2162 ();
 b15zdnd11an1n04x5 FILLER_112_2226 ();
 b15zdnd00an1n02x5 FILLER_112_2230 ();
 b15zdnd00an1n02x5 FILLER_112_2274 ();
 b15zdnd11an1n64x5 FILLER_113_0 ();
 b15zdnd11an1n64x5 FILLER_113_64 ();
 b15zdnd11an1n64x5 FILLER_113_128 ();
 b15zdnd11an1n64x5 FILLER_113_192 ();
 b15zdnd11an1n64x5 FILLER_113_256 ();
 b15zdnd11an1n64x5 FILLER_113_320 ();
 b15zdnd11an1n64x5 FILLER_113_384 ();
 b15zdnd11an1n64x5 FILLER_113_448 ();
 b15zdnd11an1n64x5 FILLER_113_512 ();
 b15zdnd11an1n16x5 FILLER_113_576 ();
 b15zdnd11an1n08x5 FILLER_113_592 ();
 b15zdnd11an1n04x5 FILLER_113_600 ();
 b15zdnd00an1n02x5 FILLER_113_604 ();
 b15zdnd00an1n01x5 FILLER_113_606 ();
 b15zdnd11an1n64x5 FILLER_113_633 ();
 b15zdnd11an1n16x5 FILLER_113_697 ();
 b15zdnd11an1n04x5 FILLER_113_713 ();
 b15zdnd00an1n02x5 FILLER_113_717 ();
 b15zdnd00an1n01x5 FILLER_113_719 ();
 b15zdnd11an1n64x5 FILLER_113_740 ();
 b15zdnd11an1n32x5 FILLER_113_804 ();
 b15zdnd11an1n08x5 FILLER_113_836 ();
 b15zdnd00an1n02x5 FILLER_113_844 ();
 b15zdnd11an1n64x5 FILLER_113_849 ();
 b15zdnd11an1n64x5 FILLER_113_913 ();
 b15zdnd11an1n64x5 FILLER_113_977 ();
 b15zdnd11an1n32x5 FILLER_113_1041 ();
 b15zdnd11an1n16x5 FILLER_113_1073 ();
 b15zdnd11an1n04x5 FILLER_113_1092 ();
 b15zdnd11an1n16x5 FILLER_113_1099 ();
 b15zdnd11an1n08x5 FILLER_113_1115 ();
 b15zdnd11an1n32x5 FILLER_113_1165 ();
 b15zdnd11an1n08x5 FILLER_113_1197 ();
 b15zdnd00an1n01x5 FILLER_113_1205 ();
 b15zdnd11an1n64x5 FILLER_113_1237 ();
 b15zdnd11an1n64x5 FILLER_113_1301 ();
 b15zdnd11an1n64x5 FILLER_113_1365 ();
 b15zdnd11an1n64x5 FILLER_113_1429 ();
 b15zdnd11an1n64x5 FILLER_113_1493 ();
 b15zdnd11an1n64x5 FILLER_113_1557 ();
 b15zdnd11an1n64x5 FILLER_113_1621 ();
 b15zdnd11an1n64x5 FILLER_113_1685 ();
 b15zdnd11an1n64x5 FILLER_113_1749 ();
 b15zdnd11an1n64x5 FILLER_113_1813 ();
 b15zdnd11an1n64x5 FILLER_113_1877 ();
 b15zdnd11an1n64x5 FILLER_113_1941 ();
 b15zdnd11an1n64x5 FILLER_113_2005 ();
 b15zdnd11an1n64x5 FILLER_113_2069 ();
 b15zdnd11an1n64x5 FILLER_113_2133 ();
 b15zdnd11an1n32x5 FILLER_113_2197 ();
 b15zdnd11an1n08x5 FILLER_113_2229 ();
 b15zdnd00an1n02x5 FILLER_113_2237 ();
 b15zdnd00an1n01x5 FILLER_113_2239 ();
 b15zdnd00an1n02x5 FILLER_113_2282 ();
 b15zdnd11an1n64x5 FILLER_114_8 ();
 b15zdnd11an1n64x5 FILLER_114_72 ();
 b15zdnd11an1n64x5 FILLER_114_136 ();
 b15zdnd11an1n64x5 FILLER_114_200 ();
 b15zdnd11an1n64x5 FILLER_114_264 ();
 b15zdnd11an1n64x5 FILLER_114_328 ();
 b15zdnd11an1n64x5 FILLER_114_392 ();
 b15zdnd11an1n64x5 FILLER_114_456 ();
 b15zdnd11an1n64x5 FILLER_114_520 ();
 b15zdnd11an1n64x5 FILLER_114_584 ();
 b15zdnd11an1n16x5 FILLER_114_648 ();
 b15zdnd11an1n08x5 FILLER_114_664 ();
 b15zdnd00an1n02x5 FILLER_114_672 ();
 b15zdnd00an1n01x5 FILLER_114_674 ();
 b15zdnd11an1n04x5 FILLER_114_693 ();
 b15zdnd11an1n16x5 FILLER_114_702 ();
 b15zdnd11an1n64x5 FILLER_114_726 ();
 b15zdnd11an1n64x5 FILLER_114_790 ();
 b15zdnd11an1n64x5 FILLER_114_854 ();
 b15zdnd11an1n64x5 FILLER_114_918 ();
 b15zdnd11an1n64x5 FILLER_114_982 ();
 b15zdnd11an1n32x5 FILLER_114_1046 ();
 b15zdnd11an1n16x5 FILLER_114_1078 ();
 b15zdnd00an1n02x5 FILLER_114_1094 ();
 b15zdnd00an1n01x5 FILLER_114_1096 ();
 b15zdnd11an1n64x5 FILLER_114_1100 ();
 b15zdnd11an1n32x5 FILLER_114_1164 ();
 b15zdnd11an1n08x5 FILLER_114_1196 ();
 b15zdnd11an1n04x5 FILLER_114_1204 ();
 b15zdnd00an1n02x5 FILLER_114_1208 ();
 b15zdnd00an1n01x5 FILLER_114_1210 ();
 b15zdnd11an1n64x5 FILLER_114_1216 ();
 b15zdnd11an1n64x5 FILLER_114_1280 ();
 b15zdnd11an1n64x5 FILLER_114_1344 ();
 b15zdnd11an1n64x5 FILLER_114_1408 ();
 b15zdnd11an1n32x5 FILLER_114_1472 ();
 b15zdnd11an1n16x5 FILLER_114_1504 ();
 b15zdnd11an1n08x5 FILLER_114_1520 ();
 b15zdnd11an1n04x5 FILLER_114_1528 ();
 b15zdnd00an1n02x5 FILLER_114_1532 ();
 b15zdnd11an1n08x5 FILLER_114_1551 ();
 b15zdnd11an1n04x5 FILLER_114_1559 ();
 b15zdnd11an1n64x5 FILLER_114_1583 ();
 b15zdnd11an1n64x5 FILLER_114_1647 ();
 b15zdnd11an1n32x5 FILLER_114_1711 ();
 b15zdnd11an1n08x5 FILLER_114_1743 ();
 b15zdnd00an1n02x5 FILLER_114_1751 ();
 b15zdnd00an1n01x5 FILLER_114_1753 ();
 b15zdnd11an1n32x5 FILLER_114_1771 ();
 b15zdnd11an1n08x5 FILLER_114_1803 ();
 b15zdnd11an1n04x5 FILLER_114_1811 ();
 b15zdnd11an1n64x5 FILLER_114_1857 ();
 b15zdnd11an1n64x5 FILLER_114_1921 ();
 b15zdnd11an1n64x5 FILLER_114_1985 ();
 b15zdnd11an1n08x5 FILLER_114_2049 ();
 b15zdnd11an1n32x5 FILLER_114_2099 ();
 b15zdnd11an1n16x5 FILLER_114_2131 ();
 b15zdnd11an1n04x5 FILLER_114_2147 ();
 b15zdnd00an1n02x5 FILLER_114_2151 ();
 b15zdnd00an1n01x5 FILLER_114_2153 ();
 b15zdnd11an1n64x5 FILLER_114_2162 ();
 b15zdnd11an1n04x5 FILLER_114_2226 ();
 b15zdnd00an1n02x5 FILLER_114_2230 ();
 b15zdnd00an1n02x5 FILLER_114_2274 ();
 b15zdnd11an1n64x5 FILLER_115_0 ();
 b15zdnd11an1n64x5 FILLER_115_64 ();
 b15zdnd11an1n64x5 FILLER_115_128 ();
 b15zdnd11an1n64x5 FILLER_115_192 ();
 b15zdnd11an1n04x5 FILLER_115_256 ();
 b15zdnd00an1n01x5 FILLER_115_260 ();
 b15zdnd11an1n64x5 FILLER_115_273 ();
 b15zdnd11an1n64x5 FILLER_115_337 ();
 b15zdnd11an1n64x5 FILLER_115_401 ();
 b15zdnd11an1n64x5 FILLER_115_465 ();
 b15zdnd11an1n64x5 FILLER_115_529 ();
 b15zdnd11an1n64x5 FILLER_115_593 ();
 b15zdnd11an1n32x5 FILLER_115_657 ();
 b15zdnd00an1n02x5 FILLER_115_689 ();
 b15zdnd11an1n16x5 FILLER_115_709 ();
 b15zdnd11an1n04x5 FILLER_115_725 ();
 b15zdnd11an1n64x5 FILLER_115_745 ();
 b15zdnd11an1n64x5 FILLER_115_809 ();
 b15zdnd11an1n32x5 FILLER_115_873 ();
 b15zdnd11an1n64x5 FILLER_115_928 ();
 b15zdnd11an1n64x5 FILLER_115_992 ();
 b15zdnd11an1n64x5 FILLER_115_1056 ();
 b15zdnd11an1n64x5 FILLER_115_1120 ();
 b15zdnd11an1n16x5 FILLER_115_1184 ();
 b15zdnd11an1n08x5 FILLER_115_1200 ();
 b15zdnd11an1n64x5 FILLER_115_1216 ();
 b15zdnd11an1n64x5 FILLER_115_1280 ();
 b15zdnd11an1n64x5 FILLER_115_1344 ();
 b15zdnd11an1n64x5 FILLER_115_1408 ();
 b15zdnd11an1n64x5 FILLER_115_1472 ();
 b15zdnd11an1n64x5 FILLER_115_1536 ();
 b15zdnd11an1n64x5 FILLER_115_1600 ();
 b15zdnd11an1n32x5 FILLER_115_1664 ();
 b15zdnd11an1n16x5 FILLER_115_1696 ();
 b15zdnd11an1n04x5 FILLER_115_1712 ();
 b15zdnd00an1n02x5 FILLER_115_1716 ();
 b15zdnd11an1n32x5 FILLER_115_1738 ();
 b15zdnd11an1n16x5 FILLER_115_1770 ();
 b15zdnd11an1n08x5 FILLER_115_1786 ();
 b15zdnd11an1n04x5 FILLER_115_1794 ();
 b15zdnd00an1n02x5 FILLER_115_1798 ();
 b15zdnd11an1n64x5 FILLER_115_1842 ();
 b15zdnd11an1n64x5 FILLER_115_1906 ();
 b15zdnd11an1n64x5 FILLER_115_1970 ();
 b15zdnd11an1n16x5 FILLER_115_2034 ();
 b15zdnd11an1n04x5 FILLER_115_2050 ();
 b15zdnd11an1n64x5 FILLER_115_2096 ();
 b15zdnd11an1n64x5 FILLER_115_2160 ();
 b15zdnd11an1n32x5 FILLER_115_2224 ();
 b15zdnd00an1n02x5 FILLER_115_2256 ();
 b15zdnd00an1n01x5 FILLER_115_2258 ();
 b15zdnd11an1n08x5 FILLER_115_2263 ();
 b15zdnd11an1n04x5 FILLER_115_2271 ();
 b15zdnd00an1n02x5 FILLER_115_2275 ();
 b15zdnd00an1n01x5 FILLER_115_2277 ();
 b15zdnd00an1n02x5 FILLER_115_2282 ();
 b15zdnd11an1n64x5 FILLER_116_8 ();
 b15zdnd11an1n32x5 FILLER_116_72 ();
 b15zdnd11an1n08x5 FILLER_116_104 ();
 b15zdnd11an1n64x5 FILLER_116_127 ();
 b15zdnd11an1n32x5 FILLER_116_191 ();
 b15zdnd11an1n16x5 FILLER_116_223 ();
 b15zdnd11an1n08x5 FILLER_116_239 ();
 b15zdnd00an1n02x5 FILLER_116_247 ();
 b15zdnd11an1n64x5 FILLER_116_272 ();
 b15zdnd11an1n64x5 FILLER_116_336 ();
 b15zdnd11an1n64x5 FILLER_116_400 ();
 b15zdnd11an1n64x5 FILLER_116_464 ();
 b15zdnd11an1n64x5 FILLER_116_528 ();
 b15zdnd11an1n64x5 FILLER_116_592 ();
 b15zdnd11an1n32x5 FILLER_116_656 ();
 b15zdnd11an1n08x5 FILLER_116_688 ();
 b15zdnd11an1n04x5 FILLER_116_696 ();
 b15zdnd00an1n02x5 FILLER_116_716 ();
 b15zdnd11an1n64x5 FILLER_116_726 ();
 b15zdnd11an1n64x5 FILLER_116_790 ();
 b15zdnd11an1n64x5 FILLER_116_854 ();
 b15zdnd11an1n64x5 FILLER_116_918 ();
 b15zdnd11an1n32x5 FILLER_116_982 ();
 b15zdnd11an1n16x5 FILLER_116_1028 ();
 b15zdnd11an1n04x5 FILLER_116_1044 ();
 b15zdnd00an1n02x5 FILLER_116_1048 ();
 b15zdnd00an1n01x5 FILLER_116_1050 ();
 b15zdnd11an1n64x5 FILLER_116_1067 ();
 b15zdnd11an1n64x5 FILLER_116_1131 ();
 b15zdnd11an1n16x5 FILLER_116_1195 ();
 b15zdnd00an1n02x5 FILLER_116_1211 ();
 b15zdnd00an1n01x5 FILLER_116_1213 ();
 b15zdnd11an1n64x5 FILLER_116_1230 ();
 b15zdnd11an1n32x5 FILLER_116_1294 ();
 b15zdnd11an1n08x5 FILLER_116_1326 ();
 b15zdnd00an1n02x5 FILLER_116_1334 ();
 b15zdnd00an1n01x5 FILLER_116_1336 ();
 b15zdnd11an1n04x5 FILLER_116_1340 ();
 b15zdnd11an1n64x5 FILLER_116_1347 ();
 b15zdnd11an1n64x5 FILLER_116_1411 ();
 b15zdnd11an1n64x5 FILLER_116_1475 ();
 b15zdnd11an1n32x5 FILLER_116_1539 ();
 b15zdnd11an1n16x5 FILLER_116_1571 ();
 b15zdnd11an1n04x5 FILLER_116_1587 ();
 b15zdnd00an1n01x5 FILLER_116_1591 ();
 b15zdnd11an1n64x5 FILLER_116_1634 ();
 b15zdnd11an1n64x5 FILLER_116_1698 ();
 b15zdnd11an1n64x5 FILLER_116_1762 ();
 b15zdnd11an1n64x5 FILLER_116_1826 ();
 b15zdnd11an1n64x5 FILLER_116_1890 ();
 b15zdnd11an1n64x5 FILLER_116_1954 ();
 b15zdnd11an1n16x5 FILLER_116_2018 ();
 b15zdnd00an1n02x5 FILLER_116_2034 ();
 b15zdnd11an1n04x5 FILLER_116_2039 ();
 b15zdnd11an1n64x5 FILLER_116_2046 ();
 b15zdnd11an1n32x5 FILLER_116_2110 ();
 b15zdnd11an1n08x5 FILLER_116_2142 ();
 b15zdnd11an1n04x5 FILLER_116_2150 ();
 b15zdnd11an1n64x5 FILLER_116_2162 ();
 b15zdnd11an1n32x5 FILLER_116_2226 ();
 b15zdnd11an1n16x5 FILLER_116_2258 ();
 b15zdnd00an1n02x5 FILLER_116_2274 ();
 b15zdnd11an1n64x5 FILLER_117_0 ();
 b15zdnd11an1n64x5 FILLER_117_64 ();
 b15zdnd11an1n64x5 FILLER_117_128 ();
 b15zdnd11an1n64x5 FILLER_117_192 ();
 b15zdnd11an1n16x5 FILLER_117_256 ();
 b15zdnd11an1n04x5 FILLER_117_278 ();
 b15zdnd11an1n64x5 FILLER_117_298 ();
 b15zdnd11an1n64x5 FILLER_117_362 ();
 b15zdnd11an1n64x5 FILLER_117_426 ();
 b15zdnd11an1n64x5 FILLER_117_490 ();
 b15zdnd11an1n64x5 FILLER_117_554 ();
 b15zdnd11an1n64x5 FILLER_117_618 ();
 b15zdnd00an1n02x5 FILLER_117_682 ();
 b15zdnd11an1n16x5 FILLER_117_693 ();
 b15zdnd11an1n04x5 FILLER_117_709 ();
 b15zdnd11an1n64x5 FILLER_117_729 ();
 b15zdnd11an1n64x5 FILLER_117_793 ();
 b15zdnd11an1n64x5 FILLER_117_857 ();
 b15zdnd11an1n64x5 FILLER_117_921 ();
 b15zdnd11an1n64x5 FILLER_117_985 ();
 b15zdnd11an1n64x5 FILLER_117_1049 ();
 b15zdnd11an1n64x5 FILLER_117_1113 ();
 b15zdnd11an1n04x5 FILLER_117_1177 ();
 b15zdnd00an1n01x5 FILLER_117_1181 ();
 b15zdnd11an1n16x5 FILLER_117_1194 ();
 b15zdnd11an1n04x5 FILLER_117_1210 ();
 b15zdnd11an1n64x5 FILLER_117_1253 ();
 b15zdnd00an1n01x5 FILLER_117_1317 ();
 b15zdnd11an1n04x5 FILLER_117_1370 ();
 b15zdnd11an1n16x5 FILLER_117_1379 ();
 b15zdnd11an1n04x5 FILLER_117_1395 ();
 b15zdnd00an1n02x5 FILLER_117_1399 ();
 b15zdnd00an1n01x5 FILLER_117_1401 ();
 b15zdnd11an1n64x5 FILLER_117_1410 ();
 b15zdnd11an1n64x5 FILLER_117_1474 ();
 b15zdnd11an1n16x5 FILLER_117_1538 ();
 b15zdnd11an1n04x5 FILLER_117_1554 ();
 b15zdnd00an1n02x5 FILLER_117_1558 ();
 b15zdnd00an1n01x5 FILLER_117_1560 ();
 b15zdnd11an1n64x5 FILLER_117_1603 ();
 b15zdnd11an1n64x5 FILLER_117_1667 ();
 b15zdnd11an1n64x5 FILLER_117_1731 ();
 b15zdnd11an1n64x5 FILLER_117_1795 ();
 b15zdnd11an1n32x5 FILLER_117_1859 ();
 b15zdnd00an1n01x5 FILLER_117_1891 ();
 b15zdnd11an1n04x5 FILLER_117_1895 ();
 b15zdnd11an1n04x5 FILLER_117_1926 ();
 b15zdnd11an1n64x5 FILLER_117_1933 ();
 b15zdnd11an1n16x5 FILLER_117_1997 ();
 b15zdnd11an1n64x5 FILLER_117_2065 ();
 b15zdnd11an1n64x5 FILLER_117_2129 ();
 b15zdnd11an1n64x5 FILLER_117_2193 ();
 b15zdnd11an1n16x5 FILLER_117_2257 ();
 b15zdnd11an1n08x5 FILLER_117_2273 ();
 b15zdnd00an1n02x5 FILLER_117_2281 ();
 b15zdnd00an1n01x5 FILLER_117_2283 ();
 b15zdnd11an1n04x5 FILLER_118_8 ();
 b15zdnd00an1n02x5 FILLER_118_12 ();
 b15zdnd11an1n64x5 FILLER_118_18 ();
 b15zdnd11an1n64x5 FILLER_118_82 ();
 b15zdnd11an1n64x5 FILLER_118_146 ();
 b15zdnd11an1n64x5 FILLER_118_210 ();
 b15zdnd11an1n64x5 FILLER_118_274 ();
 b15zdnd11an1n64x5 FILLER_118_338 ();
 b15zdnd11an1n64x5 FILLER_118_402 ();
 b15zdnd11an1n64x5 FILLER_118_466 ();
 b15zdnd11an1n64x5 FILLER_118_530 ();
 b15zdnd11an1n64x5 FILLER_118_594 ();
 b15zdnd11an1n32x5 FILLER_118_658 ();
 b15zdnd11an1n16x5 FILLER_118_690 ();
 b15zdnd11an1n08x5 FILLER_118_706 ();
 b15zdnd11an1n04x5 FILLER_118_714 ();
 b15zdnd11an1n64x5 FILLER_118_726 ();
 b15zdnd11an1n64x5 FILLER_118_790 ();
 b15zdnd11an1n64x5 FILLER_118_854 ();
 b15zdnd11an1n64x5 FILLER_118_918 ();
 b15zdnd11an1n64x5 FILLER_118_982 ();
 b15zdnd11an1n32x5 FILLER_118_1046 ();
 b15zdnd11an1n08x5 FILLER_118_1078 ();
 b15zdnd11an1n04x5 FILLER_118_1086 ();
 b15zdnd11an1n64x5 FILLER_118_1095 ();
 b15zdnd11an1n32x5 FILLER_118_1159 ();
 b15zdnd11an1n16x5 FILLER_118_1191 ();
 b15zdnd11an1n04x5 FILLER_118_1207 ();
 b15zdnd11an1n64x5 FILLER_118_1222 ();
 b15zdnd11an1n32x5 FILLER_118_1286 ();
 b15zdnd11an1n16x5 FILLER_118_1318 ();
 b15zdnd11an1n04x5 FILLER_118_1334 ();
 b15zdnd00an1n02x5 FILLER_118_1338 ();
 b15zdnd00an1n01x5 FILLER_118_1340 ();
 b15zdnd11an1n64x5 FILLER_118_1344 ();
 b15zdnd11an1n64x5 FILLER_118_1408 ();
 b15zdnd11an1n64x5 FILLER_118_1472 ();
 b15zdnd11an1n64x5 FILLER_118_1536 ();
 b15zdnd11an1n64x5 FILLER_118_1600 ();
 b15zdnd11an1n64x5 FILLER_118_1664 ();
 b15zdnd11an1n64x5 FILLER_118_1728 ();
 b15zdnd11an1n64x5 FILLER_118_1792 ();
 b15zdnd11an1n32x5 FILLER_118_1856 ();
 b15zdnd11an1n08x5 FILLER_118_1888 ();
 b15zdnd11an1n04x5 FILLER_118_1896 ();
 b15zdnd00an1n02x5 FILLER_118_1900 ();
 b15zdnd00an1n01x5 FILLER_118_1902 ();
 b15zdnd11an1n32x5 FILLER_118_1955 ();
 b15zdnd11an1n16x5 FILLER_118_1987 ();
 b15zdnd11an1n08x5 FILLER_118_2003 ();
 b15zdnd11an1n04x5 FILLER_118_2011 ();
 b15zdnd00an1n02x5 FILLER_118_2015 ();
 b15zdnd11an1n64x5 FILLER_118_2069 ();
 b15zdnd11an1n16x5 FILLER_118_2133 ();
 b15zdnd11an1n04x5 FILLER_118_2149 ();
 b15zdnd00an1n01x5 FILLER_118_2153 ();
 b15zdnd11an1n64x5 FILLER_118_2162 ();
 b15zdnd11an1n32x5 FILLER_118_2226 ();
 b15zdnd11an1n16x5 FILLER_118_2258 ();
 b15zdnd00an1n02x5 FILLER_118_2274 ();
 b15zdnd11an1n08x5 FILLER_119_0 ();
 b15zdnd00an1n02x5 FILLER_119_8 ();
 b15zdnd00an1n01x5 FILLER_119_10 ();
 b15zdnd11an1n64x5 FILLER_119_17 ();
 b15zdnd11an1n64x5 FILLER_119_81 ();
 b15zdnd11an1n64x5 FILLER_119_145 ();
 b15zdnd11an1n64x5 FILLER_119_209 ();
 b15zdnd11an1n64x5 FILLER_119_273 ();
 b15zdnd11an1n64x5 FILLER_119_337 ();
 b15zdnd11an1n64x5 FILLER_119_401 ();
 b15zdnd11an1n64x5 FILLER_119_465 ();
 b15zdnd11an1n64x5 FILLER_119_529 ();
 b15zdnd11an1n64x5 FILLER_119_593 ();
 b15zdnd11an1n08x5 FILLER_119_657 ();
 b15zdnd11an1n04x5 FILLER_119_665 ();
 b15zdnd00an1n02x5 FILLER_119_669 ();
 b15zdnd00an1n01x5 FILLER_119_671 ();
 b15zdnd11an1n64x5 FILLER_119_675 ();
 b15zdnd11an1n64x5 FILLER_119_739 ();
 b15zdnd11an1n64x5 FILLER_119_803 ();
 b15zdnd11an1n64x5 FILLER_119_867 ();
 b15zdnd11an1n64x5 FILLER_119_931 ();
 b15zdnd11an1n64x5 FILLER_119_995 ();
 b15zdnd11an1n64x5 FILLER_119_1059 ();
 b15zdnd11an1n64x5 FILLER_119_1123 ();
 b15zdnd11an1n32x5 FILLER_119_1187 ();
 b15zdnd00an1n02x5 FILLER_119_1219 ();
 b15zdnd00an1n01x5 FILLER_119_1221 ();
 b15zdnd11an1n04x5 FILLER_119_1238 ();
 b15zdnd11an1n04x5 FILLER_119_1249 ();
 b15zdnd00an1n01x5 FILLER_119_1253 ();
 b15zdnd11an1n64x5 FILLER_119_1261 ();
 b15zdnd11an1n08x5 FILLER_119_1325 ();
 b15zdnd11an1n04x5 FILLER_119_1333 ();
 b15zdnd00an1n01x5 FILLER_119_1337 ();
 b15zdnd11an1n64x5 FILLER_119_1343 ();
 b15zdnd11an1n64x5 FILLER_119_1407 ();
 b15zdnd11an1n64x5 FILLER_119_1471 ();
 b15zdnd11an1n64x5 FILLER_119_1535 ();
 b15zdnd11an1n64x5 FILLER_119_1599 ();
 b15zdnd11an1n64x5 FILLER_119_1663 ();
 b15zdnd11an1n64x5 FILLER_119_1727 ();
 b15zdnd11an1n64x5 FILLER_119_1791 ();
 b15zdnd11an1n32x5 FILLER_119_1855 ();
 b15zdnd11an1n08x5 FILLER_119_1887 ();
 b15zdnd11an1n04x5 FILLER_119_1895 ();
 b15zdnd00an1n02x5 FILLER_119_1899 ();
 b15zdnd11an1n04x5 FILLER_119_1953 ();
 b15zdnd11an1n64x5 FILLER_119_1965 ();
 b15zdnd11an1n04x5 FILLER_119_2029 ();
 b15zdnd00an1n01x5 FILLER_119_2033 ();
 b15zdnd11an1n04x5 FILLER_119_2037 ();
 b15zdnd11an1n04x5 FILLER_119_2044 ();
 b15zdnd11an1n04x5 FILLER_119_2051 ();
 b15zdnd11an1n64x5 FILLER_119_2066 ();
 b15zdnd11an1n64x5 FILLER_119_2130 ();
 b15zdnd11an1n64x5 FILLER_119_2194 ();
 b15zdnd11an1n16x5 FILLER_119_2258 ();
 b15zdnd11an1n08x5 FILLER_119_2274 ();
 b15zdnd00an1n02x5 FILLER_119_2282 ();
 b15zdnd00an1n02x5 FILLER_120_8 ();
 b15zdnd11an1n04x5 FILLER_120_15 ();
 b15zdnd11an1n04x5 FILLER_120_23 ();
 b15zdnd00an1n02x5 FILLER_120_27 ();
 b15zdnd00an1n01x5 FILLER_120_29 ();
 b15zdnd11an1n08x5 FILLER_120_34 ();
 b15zdnd11an1n04x5 FILLER_120_42 ();
 b15zdnd11an1n16x5 FILLER_120_58 ();
 b15zdnd11an1n08x5 FILLER_120_74 ();
 b15zdnd11an1n04x5 FILLER_120_82 ();
 b15zdnd11an1n64x5 FILLER_120_110 ();
 b15zdnd11an1n64x5 FILLER_120_174 ();
 b15zdnd11an1n64x5 FILLER_120_238 ();
 b15zdnd11an1n64x5 FILLER_120_302 ();
 b15zdnd11an1n64x5 FILLER_120_366 ();
 b15zdnd11an1n64x5 FILLER_120_430 ();
 b15zdnd11an1n64x5 FILLER_120_494 ();
 b15zdnd11an1n64x5 FILLER_120_558 ();
 b15zdnd11an1n32x5 FILLER_120_622 ();
 b15zdnd11an1n16x5 FILLER_120_654 ();
 b15zdnd00an1n02x5 FILLER_120_670 ();
 b15zdnd00an1n01x5 FILLER_120_672 ();
 b15zdnd11an1n08x5 FILLER_120_676 ();
 b15zdnd11an1n16x5 FILLER_120_687 ();
 b15zdnd11an1n04x5 FILLER_120_703 ();
 b15zdnd00an1n01x5 FILLER_120_707 ();
 b15zdnd00an1n02x5 FILLER_120_715 ();
 b15zdnd00an1n01x5 FILLER_120_717 ();
 b15zdnd00an1n02x5 FILLER_120_726 ();
 b15zdnd11an1n64x5 FILLER_120_738 ();
 b15zdnd11an1n64x5 FILLER_120_802 ();
 b15zdnd11an1n64x5 FILLER_120_866 ();
 b15zdnd11an1n64x5 FILLER_120_930 ();
 b15zdnd11an1n64x5 FILLER_120_994 ();
 b15zdnd11an1n16x5 FILLER_120_1058 ();
 b15zdnd11an1n64x5 FILLER_120_1085 ();
 b15zdnd11an1n64x5 FILLER_120_1149 ();
 b15zdnd11an1n08x5 FILLER_120_1213 ();
 b15zdnd11an1n16x5 FILLER_120_1227 ();
 b15zdnd11an1n08x5 FILLER_120_1243 ();
 b15zdnd00an1n02x5 FILLER_120_1251 ();
 b15zdnd00an1n01x5 FILLER_120_1253 ();
 b15zdnd11an1n64x5 FILLER_120_1261 ();
 b15zdnd11an1n64x5 FILLER_120_1325 ();
 b15zdnd11an1n64x5 FILLER_120_1389 ();
 b15zdnd11an1n64x5 FILLER_120_1453 ();
 b15zdnd11an1n64x5 FILLER_120_1517 ();
 b15zdnd11an1n64x5 FILLER_120_1581 ();
 b15zdnd11an1n64x5 FILLER_120_1645 ();
 b15zdnd11an1n64x5 FILLER_120_1709 ();
 b15zdnd11an1n64x5 FILLER_120_1773 ();
 b15zdnd11an1n32x5 FILLER_120_1837 ();
 b15zdnd11an1n16x5 FILLER_120_1869 ();
 b15zdnd11an1n08x5 FILLER_120_1885 ();
 b15zdnd11an1n04x5 FILLER_120_1893 ();
 b15zdnd11an1n08x5 FILLER_120_1905 ();
 b15zdnd11an1n04x5 FILLER_120_1913 ();
 b15zdnd00an1n02x5 FILLER_120_1917 ();
 b15zdnd11an1n04x5 FILLER_120_1922 ();
 b15zdnd11an1n04x5 FILLER_120_1929 ();
 b15zdnd11an1n04x5 FILLER_120_1936 ();
 b15zdnd11an1n64x5 FILLER_120_1943 ();
 b15zdnd11an1n32x5 FILLER_120_2007 ();
 b15zdnd00an1n02x5 FILLER_120_2039 ();
 b15zdnd00an1n01x5 FILLER_120_2041 ();
 b15zdnd11an1n08x5 FILLER_120_2045 ();
 b15zdnd11an1n64x5 FILLER_120_2064 ();
 b15zdnd11an1n16x5 FILLER_120_2128 ();
 b15zdnd11an1n08x5 FILLER_120_2144 ();
 b15zdnd00an1n02x5 FILLER_120_2152 ();
 b15zdnd11an1n64x5 FILLER_120_2162 ();
 b15zdnd11an1n32x5 FILLER_120_2226 ();
 b15zdnd11an1n16x5 FILLER_120_2258 ();
 b15zdnd00an1n02x5 FILLER_120_2274 ();
 b15zdnd11an1n08x5 FILLER_121_0 ();
 b15zdnd11an1n04x5 FILLER_121_8 ();
 b15zdnd00an1n02x5 FILLER_121_12 ();
 b15zdnd00an1n01x5 FILLER_121_14 ();
 b15zdnd11an1n64x5 FILLER_121_23 ();
 b15zdnd11an1n32x5 FILLER_121_87 ();
 b15zdnd11an1n64x5 FILLER_121_122 ();
 b15zdnd11an1n64x5 FILLER_121_186 ();
 b15zdnd11an1n64x5 FILLER_121_250 ();
 b15zdnd11an1n64x5 FILLER_121_314 ();
 b15zdnd11an1n64x5 FILLER_121_378 ();
 b15zdnd11an1n64x5 FILLER_121_442 ();
 b15zdnd11an1n64x5 FILLER_121_506 ();
 b15zdnd11an1n64x5 FILLER_121_570 ();
 b15zdnd11an1n16x5 FILLER_121_634 ();
 b15zdnd00an1n02x5 FILLER_121_650 ();
 b15zdnd11an1n04x5 FILLER_121_704 ();
 b15zdnd11an1n64x5 FILLER_121_750 ();
 b15zdnd11an1n64x5 FILLER_121_814 ();
 b15zdnd11an1n64x5 FILLER_121_878 ();
 b15zdnd11an1n64x5 FILLER_121_942 ();
 b15zdnd11an1n64x5 FILLER_121_1006 ();
 b15zdnd11an1n64x5 FILLER_121_1070 ();
 b15zdnd11an1n08x5 FILLER_121_1134 ();
 b15zdnd11an1n64x5 FILLER_121_1170 ();
 b15zdnd11an1n64x5 FILLER_121_1234 ();
 b15zdnd11an1n64x5 FILLER_121_1298 ();
 b15zdnd11an1n64x5 FILLER_121_1362 ();
 b15zdnd11an1n64x5 FILLER_121_1426 ();
 b15zdnd11an1n64x5 FILLER_121_1490 ();
 b15zdnd11an1n64x5 FILLER_121_1554 ();
 b15zdnd11an1n64x5 FILLER_121_1618 ();
 b15zdnd11an1n32x5 FILLER_121_1682 ();
 b15zdnd11an1n04x5 FILLER_121_1714 ();
 b15zdnd00an1n01x5 FILLER_121_1718 ();
 b15zdnd11an1n08x5 FILLER_121_1722 ();
 b15zdnd11an1n04x5 FILLER_121_1730 ();
 b15zdnd00an1n01x5 FILLER_121_1734 ();
 b15zdnd11an1n04x5 FILLER_121_1738 ();
 b15zdnd11an1n32x5 FILLER_121_1745 ();
 b15zdnd11an1n16x5 FILLER_121_1777 ();
 b15zdnd11an1n64x5 FILLER_121_1824 ();
 b15zdnd11an1n32x5 FILLER_121_1888 ();
 b15zdnd11an1n08x5 FILLER_121_1920 ();
 b15zdnd00an1n01x5 FILLER_121_1928 ();
 b15zdnd11an1n64x5 FILLER_121_1932 ();
 b15zdnd11an1n64x5 FILLER_121_1996 ();
 b15zdnd11an1n64x5 FILLER_121_2060 ();
 b15zdnd11an1n64x5 FILLER_121_2124 ();
 b15zdnd11an1n64x5 FILLER_121_2188 ();
 b15zdnd11an1n32x5 FILLER_121_2252 ();
 b15zdnd11an1n16x5 FILLER_122_8 ();
 b15zdnd11an1n04x5 FILLER_122_24 ();
 b15zdnd00an1n02x5 FILLER_122_28 ();
 b15zdnd11an1n04x5 FILLER_122_33 ();
 b15zdnd11an1n64x5 FILLER_122_41 ();
 b15zdnd11an1n08x5 FILLER_122_105 ();
 b15zdnd00an1n02x5 FILLER_122_113 ();
 b15zdnd11an1n64x5 FILLER_122_135 ();
 b15zdnd11an1n64x5 FILLER_122_199 ();
 b15zdnd11an1n64x5 FILLER_122_263 ();
 b15zdnd11an1n64x5 FILLER_122_327 ();
 b15zdnd11an1n64x5 FILLER_122_391 ();
 b15zdnd11an1n64x5 FILLER_122_455 ();
 b15zdnd11an1n32x5 FILLER_122_519 ();
 b15zdnd11an1n16x5 FILLER_122_551 ();
 b15zdnd11an1n08x5 FILLER_122_567 ();
 b15zdnd00an1n02x5 FILLER_122_575 ();
 b15zdnd11an1n64x5 FILLER_122_587 ();
 b15zdnd11an1n04x5 FILLER_122_651 ();
 b15zdnd11an1n16x5 FILLER_122_697 ();
 b15zdnd11an1n04x5 FILLER_122_713 ();
 b15zdnd00an1n01x5 FILLER_122_717 ();
 b15zdnd11an1n64x5 FILLER_122_726 ();
 b15zdnd11an1n64x5 FILLER_122_790 ();
 b15zdnd11an1n64x5 FILLER_122_854 ();
 b15zdnd11an1n64x5 FILLER_122_918 ();
 b15zdnd11an1n64x5 FILLER_122_982 ();
 b15zdnd11an1n64x5 FILLER_122_1046 ();
 b15zdnd11an1n32x5 FILLER_122_1110 ();
 b15zdnd11an1n04x5 FILLER_122_1142 ();
 b15zdnd00an1n01x5 FILLER_122_1146 ();
 b15zdnd11an1n16x5 FILLER_122_1161 ();
 b15zdnd11an1n08x5 FILLER_122_1177 ();
 b15zdnd00an1n01x5 FILLER_122_1185 ();
 b15zdnd11an1n64x5 FILLER_122_1189 ();
 b15zdnd11an1n64x5 FILLER_122_1253 ();
 b15zdnd11an1n64x5 FILLER_122_1317 ();
 b15zdnd11an1n64x5 FILLER_122_1381 ();
 b15zdnd11an1n64x5 FILLER_122_1445 ();
 b15zdnd11an1n64x5 FILLER_122_1509 ();
 b15zdnd11an1n64x5 FILLER_122_1573 ();
 b15zdnd11an1n64x5 FILLER_122_1637 ();
 b15zdnd11an1n08x5 FILLER_122_1701 ();
 b15zdnd11an1n04x5 FILLER_122_1709 ();
 b15zdnd00an1n02x5 FILLER_122_1713 ();
 b15zdnd00an1n01x5 FILLER_122_1715 ();
 b15zdnd11an1n64x5 FILLER_122_1768 ();
 b15zdnd11an1n64x5 FILLER_122_1832 ();
 b15zdnd11an1n64x5 FILLER_122_1896 ();
 b15zdnd11an1n64x5 FILLER_122_1960 ();
 b15zdnd11an1n64x5 FILLER_122_2024 ();
 b15zdnd11an1n64x5 FILLER_122_2088 ();
 b15zdnd00an1n02x5 FILLER_122_2152 ();
 b15zdnd11an1n64x5 FILLER_122_2162 ();
 b15zdnd11an1n32x5 FILLER_122_2226 ();
 b15zdnd11an1n16x5 FILLER_122_2258 ();
 b15zdnd00an1n02x5 FILLER_122_2274 ();
 b15zdnd11an1n16x5 FILLER_123_0 ();
 b15zdnd00an1n02x5 FILLER_123_16 ();
 b15zdnd11an1n04x5 FILLER_123_23 ();
 b15zdnd00an1n01x5 FILLER_123_27 ();
 b15zdnd11an1n04x5 FILLER_123_31 ();
 b15zdnd11an1n64x5 FILLER_123_38 ();
 b15zdnd11an1n64x5 FILLER_123_102 ();
 b15zdnd11an1n64x5 FILLER_123_166 ();
 b15zdnd11an1n32x5 FILLER_123_230 ();
 b15zdnd11an1n08x5 FILLER_123_262 ();
 b15zdnd11an1n04x5 FILLER_123_270 ();
 b15zdnd00an1n02x5 FILLER_123_274 ();
 b15zdnd00an1n01x5 FILLER_123_276 ();
 b15zdnd11an1n32x5 FILLER_123_300 ();
 b15zdnd11an1n08x5 FILLER_123_332 ();
 b15zdnd00an1n02x5 FILLER_123_340 ();
 b15zdnd00an1n01x5 FILLER_123_342 ();
 b15zdnd11an1n64x5 FILLER_123_346 ();
 b15zdnd11an1n16x5 FILLER_123_410 ();
 b15zdnd11an1n08x5 FILLER_123_426 ();
 b15zdnd00an1n01x5 FILLER_123_434 ();
 b15zdnd11an1n64x5 FILLER_123_438 ();
 b15zdnd11an1n64x5 FILLER_123_502 ();
 b15zdnd11an1n64x5 FILLER_123_566 ();
 b15zdnd11an1n04x5 FILLER_123_630 ();
 b15zdnd00an1n02x5 FILLER_123_634 ();
 b15zdnd11an1n04x5 FILLER_123_661 ();
 b15zdnd11an1n16x5 FILLER_123_670 ();
 b15zdnd11an1n04x5 FILLER_123_686 ();
 b15zdnd00an1n01x5 FILLER_123_690 ();
 b15zdnd11an1n64x5 FILLER_123_714 ();
 b15zdnd11an1n64x5 FILLER_123_778 ();
 b15zdnd11an1n64x5 FILLER_123_842 ();
 b15zdnd11an1n64x5 FILLER_123_906 ();
 b15zdnd11an1n64x5 FILLER_123_970 ();
 b15zdnd11an1n64x5 FILLER_123_1034 ();
 b15zdnd11an1n64x5 FILLER_123_1098 ();
 b15zdnd11an1n08x5 FILLER_123_1162 ();
 b15zdnd00an1n02x5 FILLER_123_1170 ();
 b15zdnd11an1n64x5 FILLER_123_1175 ();
 b15zdnd11an1n64x5 FILLER_123_1239 ();
 b15zdnd11an1n32x5 FILLER_123_1303 ();
 b15zdnd11an1n08x5 FILLER_123_1335 ();
 b15zdnd00an1n02x5 FILLER_123_1343 ();
 b15zdnd00an1n01x5 FILLER_123_1345 ();
 b15zdnd11an1n64x5 FILLER_123_1351 ();
 b15zdnd11an1n64x5 FILLER_123_1415 ();
 b15zdnd11an1n64x5 FILLER_123_1479 ();
 b15zdnd11an1n64x5 FILLER_123_1543 ();
 b15zdnd11an1n64x5 FILLER_123_1607 ();
 b15zdnd11an1n16x5 FILLER_123_1671 ();
 b15zdnd11an1n04x5 FILLER_123_1687 ();
 b15zdnd00an1n01x5 FILLER_123_1691 ();
 b15zdnd11an1n64x5 FILLER_123_1744 ();
 b15zdnd11an1n04x5 FILLER_123_1808 ();
 b15zdnd11an1n64x5 FILLER_123_1836 ();
 b15zdnd11an1n64x5 FILLER_123_1900 ();
 b15zdnd11an1n64x5 FILLER_123_1964 ();
 b15zdnd11an1n64x5 FILLER_123_2028 ();
 b15zdnd11an1n64x5 FILLER_123_2092 ();
 b15zdnd11an1n64x5 FILLER_123_2156 ();
 b15zdnd11an1n64x5 FILLER_123_2220 ();
 b15zdnd00an1n02x5 FILLER_124_8 ();
 b15zdnd11an1n16x5 FILLER_124_52 ();
 b15zdnd11an1n08x5 FILLER_124_68 ();
 b15zdnd00an1n01x5 FILLER_124_76 ();
 b15zdnd11an1n64x5 FILLER_124_80 ();
 b15zdnd11an1n64x5 FILLER_124_144 ();
 b15zdnd11an1n64x5 FILLER_124_208 ();
 b15zdnd11an1n64x5 FILLER_124_272 ();
 b15zdnd00an1n02x5 FILLER_124_336 ();
 b15zdnd00an1n01x5 FILLER_124_338 ();
 b15zdnd11an1n08x5 FILLER_124_366 ();
 b15zdnd11an1n08x5 FILLER_124_381 ();
 b15zdnd11an1n04x5 FILLER_124_389 ();
 b15zdnd00an1n01x5 FILLER_124_393 ();
 b15zdnd11an1n04x5 FILLER_124_397 ();
 b15zdnd11an1n64x5 FILLER_124_443 ();
 b15zdnd11an1n64x5 FILLER_124_507 ();
 b15zdnd11an1n64x5 FILLER_124_571 ();
 b15zdnd00an1n02x5 FILLER_124_635 ();
 b15zdnd00an1n01x5 FILLER_124_637 ();
 b15zdnd11an1n32x5 FILLER_124_658 ();
 b15zdnd11an1n16x5 FILLER_124_690 ();
 b15zdnd11an1n08x5 FILLER_124_706 ();
 b15zdnd11an1n04x5 FILLER_124_714 ();
 b15zdnd11an1n64x5 FILLER_124_726 ();
 b15zdnd11an1n64x5 FILLER_124_790 ();
 b15zdnd11an1n64x5 FILLER_124_854 ();
 b15zdnd11an1n64x5 FILLER_124_918 ();
 b15zdnd11an1n64x5 FILLER_124_982 ();
 b15zdnd11an1n64x5 FILLER_124_1046 ();
 b15zdnd11an1n64x5 FILLER_124_1110 ();
 b15zdnd11an1n64x5 FILLER_124_1174 ();
 b15zdnd11an1n64x5 FILLER_124_1238 ();
 b15zdnd11an1n32x5 FILLER_124_1302 ();
 b15zdnd11an1n08x5 FILLER_124_1334 ();
 b15zdnd00an1n02x5 FILLER_124_1342 ();
 b15zdnd11an1n64x5 FILLER_124_1349 ();
 b15zdnd11an1n04x5 FILLER_124_1413 ();
 b15zdnd11an1n32x5 FILLER_124_1422 ();
 b15zdnd00an1n02x5 FILLER_124_1454 ();
 b15zdnd11an1n64x5 FILLER_124_1508 ();
 b15zdnd11an1n16x5 FILLER_124_1572 ();
 b15zdnd11an1n08x5 FILLER_124_1588 ();
 b15zdnd11an1n04x5 FILLER_124_1596 ();
 b15zdnd00an1n02x5 FILLER_124_1600 ();
 b15zdnd00an1n01x5 FILLER_124_1602 ();
 b15zdnd11an1n64x5 FILLER_124_1614 ();
 b15zdnd11an1n32x5 FILLER_124_1678 ();
 b15zdnd00an1n01x5 FILLER_124_1710 ();
 b15zdnd11an1n04x5 FILLER_124_1714 ();
 b15zdnd11an1n16x5 FILLER_124_1721 ();
 b15zdnd00an1n02x5 FILLER_124_1737 ();
 b15zdnd00an1n01x5 FILLER_124_1739 ();
 b15zdnd11an1n64x5 FILLER_124_1743 ();
 b15zdnd11an1n64x5 FILLER_124_1807 ();
 b15zdnd11an1n64x5 FILLER_124_1871 ();
 b15zdnd11an1n64x5 FILLER_124_1935 ();
 b15zdnd11an1n64x5 FILLER_124_1999 ();
 b15zdnd11an1n64x5 FILLER_124_2063 ();
 b15zdnd11an1n16x5 FILLER_124_2127 ();
 b15zdnd11an1n08x5 FILLER_124_2143 ();
 b15zdnd00an1n02x5 FILLER_124_2151 ();
 b15zdnd00an1n01x5 FILLER_124_2153 ();
 b15zdnd11an1n64x5 FILLER_124_2162 ();
 b15zdnd11an1n32x5 FILLER_124_2226 ();
 b15zdnd11an1n16x5 FILLER_124_2258 ();
 b15zdnd00an1n02x5 FILLER_124_2274 ();
 b15zdnd00an1n02x5 FILLER_125_0 ();
 b15zdnd11an1n04x5 FILLER_125_7 ();
 b15zdnd11an1n04x5 FILLER_125_53 ();
 b15zdnd11an1n64x5 FILLER_125_60 ();
 b15zdnd11an1n64x5 FILLER_125_124 ();
 b15zdnd11an1n64x5 FILLER_125_188 ();
 b15zdnd11an1n64x5 FILLER_125_252 ();
 b15zdnd11an1n04x5 FILLER_125_316 ();
 b15zdnd11an1n04x5 FILLER_125_372 ();
 b15zdnd11an1n04x5 FILLER_125_408 ();
 b15zdnd11an1n04x5 FILLER_125_464 ();
 b15zdnd11an1n32x5 FILLER_125_474 ();
 b15zdnd11an1n16x5 FILLER_125_506 ();
 b15zdnd00an1n01x5 FILLER_125_522 ();
 b15zdnd11an1n64x5 FILLER_125_542 ();
 b15zdnd11an1n64x5 FILLER_125_606 ();
 b15zdnd11an1n64x5 FILLER_125_670 ();
 b15zdnd11an1n64x5 FILLER_125_734 ();
 b15zdnd11an1n64x5 FILLER_125_798 ();
 b15zdnd11an1n64x5 FILLER_125_862 ();
 b15zdnd11an1n32x5 FILLER_125_926 ();
 b15zdnd11an1n16x5 FILLER_125_958 ();
 b15zdnd11an1n08x5 FILLER_125_974 ();
 b15zdnd00an1n02x5 FILLER_125_982 ();
 b15zdnd00an1n01x5 FILLER_125_984 ();
 b15zdnd11an1n64x5 FILLER_125_991 ();
 b15zdnd11an1n64x5 FILLER_125_1055 ();
 b15zdnd11an1n64x5 FILLER_125_1119 ();
 b15zdnd11an1n64x5 FILLER_125_1183 ();
 b15zdnd11an1n64x5 FILLER_125_1247 ();
 b15zdnd11an1n64x5 FILLER_125_1311 ();
 b15zdnd11an1n32x5 FILLER_125_1375 ();
 b15zdnd11an1n16x5 FILLER_125_1407 ();
 b15zdnd11an1n04x5 FILLER_125_1423 ();
 b15zdnd00an1n02x5 FILLER_125_1427 ();
 b15zdnd11an1n04x5 FILLER_125_1481 ();
 b15zdnd11an1n08x5 FILLER_125_1488 ();
 b15zdnd00an1n02x5 FILLER_125_1496 ();
 b15zdnd00an1n01x5 FILLER_125_1498 ();
 b15zdnd11an1n64x5 FILLER_125_1502 ();
 b15zdnd11an1n32x5 FILLER_125_1566 ();
 b15zdnd11an1n08x5 FILLER_125_1598 ();
 b15zdnd00an1n02x5 FILLER_125_1606 ();
 b15zdnd00an1n01x5 FILLER_125_1608 ();
 b15zdnd11an1n04x5 FILLER_125_1612 ();
 b15zdnd11an1n64x5 FILLER_125_1619 ();
 b15zdnd11an1n64x5 FILLER_125_1683 ();
 b15zdnd11an1n64x5 FILLER_125_1747 ();
 b15zdnd11an1n64x5 FILLER_125_1811 ();
 b15zdnd11an1n64x5 FILLER_125_1875 ();
 b15zdnd11an1n64x5 FILLER_125_1939 ();
 b15zdnd11an1n64x5 FILLER_125_2003 ();
 b15zdnd11an1n64x5 FILLER_125_2067 ();
 b15zdnd11an1n64x5 FILLER_125_2131 ();
 b15zdnd11an1n64x5 FILLER_125_2195 ();
 b15zdnd11an1n16x5 FILLER_125_2259 ();
 b15zdnd11an1n08x5 FILLER_125_2275 ();
 b15zdnd00an1n01x5 FILLER_125_2283 ();
 b15zdnd11an1n08x5 FILLER_126_8 ();
 b15zdnd00an1n02x5 FILLER_126_16 ();
 b15zdnd11an1n64x5 FILLER_126_60 ();
 b15zdnd11an1n64x5 FILLER_126_124 ();
 b15zdnd11an1n64x5 FILLER_126_188 ();
 b15zdnd11an1n64x5 FILLER_126_252 ();
 b15zdnd11an1n16x5 FILLER_126_316 ();
 b15zdnd11an1n04x5 FILLER_126_332 ();
 b15zdnd11an1n16x5 FILLER_126_378 ();
 b15zdnd11an1n08x5 FILLER_126_403 ();
 b15zdnd11an1n04x5 FILLER_126_411 ();
 b15zdnd11an1n04x5 FILLER_126_467 ();
 b15zdnd11an1n64x5 FILLER_126_478 ();
 b15zdnd11an1n16x5 FILLER_126_542 ();
 b15zdnd11an1n08x5 FILLER_126_558 ();
 b15zdnd11an1n04x5 FILLER_126_566 ();
 b15zdnd00an1n02x5 FILLER_126_570 ();
 b15zdnd00an1n01x5 FILLER_126_572 ();
 b15zdnd11an1n64x5 FILLER_126_615 ();
 b15zdnd11an1n32x5 FILLER_126_679 ();
 b15zdnd11an1n04x5 FILLER_126_711 ();
 b15zdnd00an1n02x5 FILLER_126_715 ();
 b15zdnd00an1n01x5 FILLER_126_717 ();
 b15zdnd11an1n64x5 FILLER_126_726 ();
 b15zdnd11an1n64x5 FILLER_126_790 ();
 b15zdnd11an1n64x5 FILLER_126_854 ();
 b15zdnd11an1n32x5 FILLER_126_918 ();
 b15zdnd11an1n04x5 FILLER_126_950 ();
 b15zdnd00an1n02x5 FILLER_126_954 ();
 b15zdnd00an1n01x5 FILLER_126_956 ();
 b15zdnd11an1n64x5 FILLER_126_960 ();
 b15zdnd11an1n64x5 FILLER_126_1024 ();
 b15zdnd11an1n64x5 FILLER_126_1088 ();
 b15zdnd11an1n64x5 FILLER_126_1152 ();
 b15zdnd11an1n64x5 FILLER_126_1216 ();
 b15zdnd11an1n64x5 FILLER_126_1280 ();
 b15zdnd11an1n64x5 FILLER_126_1344 ();
 b15zdnd11an1n32x5 FILLER_126_1408 ();
 b15zdnd11an1n08x5 FILLER_126_1440 ();
 b15zdnd11an1n04x5 FILLER_126_1451 ();
 b15zdnd11an1n04x5 FILLER_126_1458 ();
 b15zdnd11an1n16x5 FILLER_126_1465 ();
 b15zdnd11an1n04x5 FILLER_126_1481 ();
 b15zdnd00an1n01x5 FILLER_126_1485 ();
 b15zdnd11an1n64x5 FILLER_126_1489 ();
 b15zdnd11an1n32x5 FILLER_126_1553 ();
 b15zdnd11an1n04x5 FILLER_126_1585 ();
 b15zdnd00an1n02x5 FILLER_126_1589 ();
 b15zdnd11an1n04x5 FILLER_126_1643 ();
 b15zdnd11an1n64x5 FILLER_126_1658 ();
 b15zdnd11an1n64x5 FILLER_126_1722 ();
 b15zdnd11an1n64x5 FILLER_126_1786 ();
 b15zdnd11an1n64x5 FILLER_126_1850 ();
 b15zdnd11an1n64x5 FILLER_126_1914 ();
 b15zdnd11an1n64x5 FILLER_126_1978 ();
 b15zdnd11an1n64x5 FILLER_126_2042 ();
 b15zdnd11an1n32x5 FILLER_126_2106 ();
 b15zdnd11an1n16x5 FILLER_126_2138 ();
 b15zdnd11an1n64x5 FILLER_126_2162 ();
 b15zdnd11an1n32x5 FILLER_126_2226 ();
 b15zdnd11an1n16x5 FILLER_126_2258 ();
 b15zdnd00an1n02x5 FILLER_126_2274 ();
 b15zdnd11an1n08x5 FILLER_127_0 ();
 b15zdnd00an1n01x5 FILLER_127_8 ();
 b15zdnd11an1n04x5 FILLER_127_12 ();
 b15zdnd11an1n04x5 FILLER_127_20 ();
 b15zdnd11an1n64x5 FILLER_127_66 ();
 b15zdnd11an1n64x5 FILLER_127_130 ();
 b15zdnd11an1n64x5 FILLER_127_194 ();
 b15zdnd11an1n64x5 FILLER_127_258 ();
 b15zdnd11an1n04x5 FILLER_127_322 ();
 b15zdnd00an1n02x5 FILLER_127_326 ();
 b15zdnd00an1n01x5 FILLER_127_328 ();
 b15zdnd11an1n04x5 FILLER_127_361 ();
 b15zdnd11an1n04x5 FILLER_127_407 ();
 b15zdnd11an1n04x5 FILLER_127_420 ();
 b15zdnd11an1n04x5 FILLER_127_427 ();
 b15zdnd11an1n16x5 FILLER_127_473 ();
 b15zdnd11an1n08x5 FILLER_127_489 ();
 b15zdnd00an1n02x5 FILLER_127_497 ();
 b15zdnd00an1n01x5 FILLER_127_499 ();
 b15zdnd11an1n64x5 FILLER_127_507 ();
 b15zdnd11an1n64x5 FILLER_127_571 ();
 b15zdnd11an1n64x5 FILLER_127_635 ();
 b15zdnd11an1n64x5 FILLER_127_699 ();
 b15zdnd11an1n64x5 FILLER_127_763 ();
 b15zdnd11an1n64x5 FILLER_127_827 ();
 b15zdnd11an1n32x5 FILLER_127_891 ();
 b15zdnd11an1n16x5 FILLER_127_923 ();
 b15zdnd11an1n04x5 FILLER_127_939 ();
 b15zdnd00an1n02x5 FILLER_127_943 ();
 b15zdnd00an1n01x5 FILLER_127_945 ();
 b15zdnd11an1n64x5 FILLER_127_988 ();
 b15zdnd11an1n04x5 FILLER_127_1052 ();
 b15zdnd00an1n01x5 FILLER_127_1056 ();
 b15zdnd11an1n08x5 FILLER_127_1073 ();
 b15zdnd00an1n02x5 FILLER_127_1081 ();
 b15zdnd00an1n01x5 FILLER_127_1083 ();
 b15zdnd11an1n32x5 FILLER_127_1095 ();
 b15zdnd11an1n16x5 FILLER_127_1127 ();
 b15zdnd11an1n04x5 FILLER_127_1143 ();
 b15zdnd00an1n02x5 FILLER_127_1147 ();
 b15zdnd00an1n01x5 FILLER_127_1149 ();
 b15zdnd11an1n64x5 FILLER_127_1155 ();
 b15zdnd11an1n64x5 FILLER_127_1219 ();
 b15zdnd11an1n64x5 FILLER_127_1283 ();
 b15zdnd11an1n64x5 FILLER_127_1347 ();
 b15zdnd11an1n32x5 FILLER_127_1411 ();
 b15zdnd11an1n16x5 FILLER_127_1443 ();
 b15zdnd11an1n08x5 FILLER_127_1459 ();
 b15zdnd11an1n04x5 FILLER_127_1467 ();
 b15zdnd00an1n01x5 FILLER_127_1471 ();
 b15zdnd11an1n64x5 FILLER_127_1488 ();
 b15zdnd11an1n32x5 FILLER_127_1552 ();
 b15zdnd11an1n16x5 FILLER_127_1584 ();
 b15zdnd11an1n08x5 FILLER_127_1600 ();
 b15zdnd11an1n04x5 FILLER_127_1608 ();
 b15zdnd00an1n02x5 FILLER_127_1612 ();
 b15zdnd11an1n64x5 FILLER_127_1617 ();
 b15zdnd11an1n64x5 FILLER_127_1681 ();
 b15zdnd11an1n64x5 FILLER_127_1745 ();
 b15zdnd11an1n64x5 FILLER_127_1809 ();
 b15zdnd11an1n64x5 FILLER_127_1873 ();
 b15zdnd11an1n64x5 FILLER_127_1937 ();
 b15zdnd11an1n64x5 FILLER_127_2001 ();
 b15zdnd11an1n64x5 FILLER_127_2065 ();
 b15zdnd11an1n64x5 FILLER_127_2129 ();
 b15zdnd11an1n64x5 FILLER_127_2193 ();
 b15zdnd11an1n16x5 FILLER_127_2257 ();
 b15zdnd11an1n08x5 FILLER_127_2273 ();
 b15zdnd00an1n02x5 FILLER_127_2281 ();
 b15zdnd00an1n01x5 FILLER_127_2283 ();
 b15zdnd00an1n02x5 FILLER_128_8 ();
 b15zdnd11an1n08x5 FILLER_128_14 ();
 b15zdnd00an1n01x5 FILLER_128_22 ();
 b15zdnd11an1n04x5 FILLER_128_27 ();
 b15zdnd11an1n08x5 FILLER_128_35 ();
 b15zdnd11an1n04x5 FILLER_128_46 ();
 b15zdnd11an1n16x5 FILLER_128_53 ();
 b15zdnd11an1n08x5 FILLER_128_69 ();
 b15zdnd11an1n04x5 FILLER_128_77 ();
 b15zdnd11an1n08x5 FILLER_128_123 ();
 b15zdnd11an1n04x5 FILLER_128_131 ();
 b15zdnd00an1n02x5 FILLER_128_135 ();
 b15zdnd00an1n01x5 FILLER_128_137 ();
 b15zdnd11an1n08x5 FILLER_128_145 ();
 b15zdnd00an1n02x5 FILLER_128_153 ();
 b15zdnd11an1n64x5 FILLER_128_169 ();
 b15zdnd11an1n64x5 FILLER_128_233 ();
 b15zdnd11an1n32x5 FILLER_128_297 ();
 b15zdnd11an1n04x5 FILLER_128_329 ();
 b15zdnd00an1n02x5 FILLER_128_333 ();
 b15zdnd11an1n04x5 FILLER_128_338 ();
 b15zdnd11an1n04x5 FILLER_128_345 ();
 b15zdnd11an1n04x5 FILLER_128_358 ();
 b15zdnd11an1n04x5 FILLER_128_365 ();
 b15zdnd11an1n16x5 FILLER_128_372 ();
 b15zdnd00an1n02x5 FILLER_128_388 ();
 b15zdnd00an1n01x5 FILLER_128_390 ();
 b15zdnd11an1n04x5 FILLER_128_398 ();
 b15zdnd11an1n16x5 FILLER_128_405 ();
 b15zdnd00an1n02x5 FILLER_128_421 ();
 b15zdnd11an1n04x5 FILLER_128_426 ();
 b15zdnd11an1n04x5 FILLER_128_472 ();
 b15zdnd11an1n32x5 FILLER_128_483 ();
 b15zdnd11an1n04x5 FILLER_128_515 ();
 b15zdnd00an1n02x5 FILLER_128_519 ();
 b15zdnd11an1n08x5 FILLER_128_524 ();
 b15zdnd11an1n04x5 FILLER_128_532 ();
 b15zdnd00an1n02x5 FILLER_128_536 ();
 b15zdnd11an1n64x5 FILLER_128_543 ();
 b15zdnd11an1n64x5 FILLER_128_607 ();
 b15zdnd11an1n32x5 FILLER_128_671 ();
 b15zdnd11an1n08x5 FILLER_128_703 ();
 b15zdnd11an1n04x5 FILLER_128_711 ();
 b15zdnd00an1n02x5 FILLER_128_715 ();
 b15zdnd00an1n01x5 FILLER_128_717 ();
 b15zdnd11an1n64x5 FILLER_128_726 ();
 b15zdnd11an1n64x5 FILLER_128_790 ();
 b15zdnd11an1n64x5 FILLER_128_854 ();
 b15zdnd11an1n08x5 FILLER_128_918 ();
 b15zdnd11an1n04x5 FILLER_128_926 ();
 b15zdnd11an1n64x5 FILLER_128_982 ();
 b15zdnd11an1n16x5 FILLER_128_1046 ();
 b15zdnd11an1n08x5 FILLER_128_1062 ();
 b15zdnd11an1n04x5 FILLER_128_1070 ();
 b15zdnd11an1n64x5 FILLER_128_1078 ();
 b15zdnd11an1n64x5 FILLER_128_1142 ();
 b15zdnd11an1n64x5 FILLER_128_1206 ();
 b15zdnd11an1n64x5 FILLER_128_1270 ();
 b15zdnd11an1n64x5 FILLER_128_1334 ();
 b15zdnd11an1n64x5 FILLER_128_1398 ();
 b15zdnd11an1n32x5 FILLER_128_1462 ();
 b15zdnd00an1n02x5 FILLER_128_1494 ();
 b15zdnd11an1n64x5 FILLER_128_1538 ();
 b15zdnd11an1n64x5 FILLER_128_1602 ();
 b15zdnd11an1n64x5 FILLER_128_1666 ();
 b15zdnd11an1n64x5 FILLER_128_1730 ();
 b15zdnd11an1n64x5 FILLER_128_1794 ();
 b15zdnd11an1n64x5 FILLER_128_1858 ();
 b15zdnd11an1n64x5 FILLER_128_1922 ();
 b15zdnd11an1n64x5 FILLER_128_1986 ();
 b15zdnd11an1n64x5 FILLER_128_2050 ();
 b15zdnd11an1n32x5 FILLER_128_2114 ();
 b15zdnd11an1n08x5 FILLER_128_2146 ();
 b15zdnd11an1n16x5 FILLER_128_2162 ();
 b15zdnd11an1n08x5 FILLER_128_2178 ();
 b15zdnd00an1n01x5 FILLER_128_2186 ();
 b15zdnd11an1n32x5 FILLER_128_2220 ();
 b15zdnd11an1n16x5 FILLER_128_2252 ();
 b15zdnd11an1n08x5 FILLER_128_2268 ();
 b15zdnd11an1n08x5 FILLER_129_0 ();
 b15zdnd11an1n04x5 FILLER_129_13 ();
 b15zdnd11an1n04x5 FILLER_129_21 ();
 b15zdnd00an1n02x5 FILLER_129_25 ();
 b15zdnd00an1n01x5 FILLER_129_27 ();
 b15zdnd11an1n04x5 FILLER_129_31 ();
 b15zdnd11an1n04x5 FILLER_129_38 ();
 b15zdnd11an1n32x5 FILLER_129_45 ();
 b15zdnd11an1n08x5 FILLER_129_77 ();
 b15zdnd00an1n02x5 FILLER_129_85 ();
 b15zdnd11an1n64x5 FILLER_129_129 ();
 b15zdnd11an1n64x5 FILLER_129_193 ();
 b15zdnd11an1n64x5 FILLER_129_257 ();
 b15zdnd11an1n32x5 FILLER_129_321 ();
 b15zdnd00an1n01x5 FILLER_129_353 ();
 b15zdnd11an1n64x5 FILLER_129_357 ();
 b15zdnd11an1n08x5 FILLER_129_421 ();
 b15zdnd00an1n02x5 FILLER_129_429 ();
 b15zdnd11an1n04x5 FILLER_129_434 ();
 b15zdnd11an1n04x5 FILLER_129_441 ();
 b15zdnd11an1n08x5 FILLER_129_448 ();
 b15zdnd11an1n04x5 FILLER_129_456 ();
 b15zdnd11an1n32x5 FILLER_129_467 ();
 b15zdnd11an1n08x5 FILLER_129_499 ();
 b15zdnd00an1n02x5 FILLER_129_507 ();
 b15zdnd11an1n04x5 FILLER_129_514 ();
 b15zdnd11an1n64x5 FILLER_129_560 ();
 b15zdnd11an1n64x5 FILLER_129_624 ();
 b15zdnd11an1n64x5 FILLER_129_688 ();
 b15zdnd11an1n64x5 FILLER_129_752 ();
 b15zdnd11an1n32x5 FILLER_129_816 ();
 b15zdnd11an1n16x5 FILLER_129_848 ();
 b15zdnd11an1n08x5 FILLER_129_864 ();
 b15zdnd11an1n04x5 FILLER_129_872 ();
 b15zdnd00an1n02x5 FILLER_129_876 ();
 b15zdnd11an1n32x5 FILLER_129_885 ();
 b15zdnd11an1n16x5 FILLER_129_917 ();
 b15zdnd11an1n08x5 FILLER_129_933 ();
 b15zdnd11an1n04x5 FILLER_129_941 ();
 b15zdnd00an1n02x5 FILLER_129_945 ();
 b15zdnd00an1n01x5 FILLER_129_947 ();
 b15zdnd11an1n04x5 FILLER_129_951 ();
 b15zdnd11an1n64x5 FILLER_129_958 ();
 b15zdnd11an1n16x5 FILLER_129_1022 ();
 b15zdnd11an1n08x5 FILLER_129_1038 ();
 b15zdnd00an1n02x5 FILLER_129_1046 ();
 b15zdnd11an1n04x5 FILLER_129_1070 ();
 b15zdnd11an1n64x5 FILLER_129_1083 ();
 b15zdnd11an1n64x5 FILLER_129_1147 ();
 b15zdnd11an1n64x5 FILLER_129_1211 ();
 b15zdnd11an1n64x5 FILLER_129_1275 ();
 b15zdnd11an1n64x5 FILLER_129_1339 ();
 b15zdnd11an1n32x5 FILLER_129_1403 ();
 b15zdnd00an1n02x5 FILLER_129_1435 ();
 b15zdnd11an1n64x5 FILLER_129_1479 ();
 b15zdnd11an1n16x5 FILLER_129_1543 ();
 b15zdnd11an1n08x5 FILLER_129_1559 ();
 b15zdnd00an1n02x5 FILLER_129_1567 ();
 b15zdnd00an1n01x5 FILLER_129_1569 ();
 b15zdnd11an1n04x5 FILLER_129_1597 ();
 b15zdnd00an1n02x5 FILLER_129_1601 ();
 b15zdnd00an1n01x5 FILLER_129_1603 ();
 b15zdnd11an1n64x5 FILLER_129_1607 ();
 b15zdnd11an1n64x5 FILLER_129_1671 ();
 b15zdnd11an1n64x5 FILLER_129_1735 ();
 b15zdnd11an1n32x5 FILLER_129_1799 ();
 b15zdnd11an1n16x5 FILLER_129_1831 ();
 b15zdnd11an1n04x5 FILLER_129_1847 ();
 b15zdnd00an1n01x5 FILLER_129_1851 ();
 b15zdnd11an1n64x5 FILLER_129_1863 ();
 b15zdnd11an1n64x5 FILLER_129_1927 ();
 b15zdnd11an1n16x5 FILLER_129_1991 ();
 b15zdnd11an1n08x5 FILLER_129_2007 ();
 b15zdnd11an1n04x5 FILLER_129_2015 ();
 b15zdnd00an1n02x5 FILLER_129_2019 ();
 b15zdnd11an1n08x5 FILLER_129_2024 ();
 b15zdnd00an1n01x5 FILLER_129_2032 ();
 b15zdnd11an1n64x5 FILLER_129_2036 ();
 b15zdnd11an1n64x5 FILLER_129_2100 ();
 b15zdnd11an1n64x5 FILLER_129_2164 ();
 b15zdnd11an1n32x5 FILLER_129_2228 ();
 b15zdnd11an1n16x5 FILLER_129_2260 ();
 b15zdnd11an1n08x5 FILLER_129_2276 ();
 b15zdnd11an1n08x5 FILLER_130_8 ();
 b15zdnd00an1n02x5 FILLER_130_16 ();
 b15zdnd00an1n01x5 FILLER_130_18 ();
 b15zdnd11an1n04x5 FILLER_130_22 ();
 b15zdnd11an1n32x5 FILLER_130_29 ();
 b15zdnd11an1n04x5 FILLER_130_61 ();
 b15zdnd00an1n02x5 FILLER_130_65 ();
 b15zdnd00an1n01x5 FILLER_130_67 ();
 b15zdnd11an1n04x5 FILLER_130_74 ();
 b15zdnd11an1n08x5 FILLER_130_83 ();
 b15zdnd11an1n04x5 FILLER_130_91 ();
 b15zdnd11an1n64x5 FILLER_130_137 ();
 b15zdnd11an1n16x5 FILLER_130_201 ();
 b15zdnd11an1n08x5 FILLER_130_217 ();
 b15zdnd00an1n02x5 FILLER_130_225 ();
 b15zdnd00an1n01x5 FILLER_130_227 ();
 b15zdnd11an1n64x5 FILLER_130_242 ();
 b15zdnd11an1n64x5 FILLER_130_306 ();
 b15zdnd11an1n64x5 FILLER_130_370 ();
 b15zdnd00an1n02x5 FILLER_130_434 ();
 b15zdnd00an1n01x5 FILLER_130_436 ();
 b15zdnd11an1n32x5 FILLER_130_448 ();
 b15zdnd11an1n08x5 FILLER_130_480 ();
 b15zdnd11an1n04x5 FILLER_130_488 ();
 b15zdnd00an1n02x5 FILLER_130_492 ();
 b15zdnd11an1n64x5 FILLER_130_546 ();
 b15zdnd11an1n64x5 FILLER_130_610 ();
 b15zdnd11an1n32x5 FILLER_130_674 ();
 b15zdnd11an1n08x5 FILLER_130_706 ();
 b15zdnd11an1n04x5 FILLER_130_714 ();
 b15zdnd11an1n64x5 FILLER_130_726 ();
 b15zdnd11an1n32x5 FILLER_130_790 ();
 b15zdnd11an1n16x5 FILLER_130_822 ();
 b15zdnd11an1n08x5 FILLER_130_838 ();
 b15zdnd11an1n16x5 FILLER_130_888 ();
 b15zdnd11an1n08x5 FILLER_130_904 ();
 b15zdnd00an1n02x5 FILLER_130_912 ();
 b15zdnd00an1n01x5 FILLER_130_914 ();
 b15zdnd11an1n32x5 FILLER_130_919 ();
 b15zdnd11an1n16x5 FILLER_130_951 ();
 b15zdnd11an1n08x5 FILLER_130_967 ();
 b15zdnd11an1n04x5 FILLER_130_975 ();
 b15zdnd11an1n08x5 FILLER_130_994 ();
 b15zdnd11an1n04x5 FILLER_130_1002 ();
 b15zdnd00an1n02x5 FILLER_130_1006 ();
 b15zdnd00an1n01x5 FILLER_130_1008 ();
 b15zdnd11an1n08x5 FILLER_130_1016 ();
 b15zdnd11an1n04x5 FILLER_130_1024 ();
 b15zdnd11an1n16x5 FILLER_130_1032 ();
 b15zdnd11an1n08x5 FILLER_130_1048 ();
 b15zdnd11an1n16x5 FILLER_130_1066 ();
 b15zdnd11an1n08x5 FILLER_130_1082 ();
 b15zdnd00an1n02x5 FILLER_130_1090 ();
 b15zdnd11an1n64x5 FILLER_130_1104 ();
 b15zdnd11an1n32x5 FILLER_130_1168 ();
 b15zdnd11an1n08x5 FILLER_130_1200 ();
 b15zdnd00an1n02x5 FILLER_130_1208 ();
 b15zdnd11an1n64x5 FILLER_130_1219 ();
 b15zdnd11an1n64x5 FILLER_130_1283 ();
 b15zdnd11an1n64x5 FILLER_130_1347 ();
 b15zdnd11an1n64x5 FILLER_130_1411 ();
 b15zdnd11an1n64x5 FILLER_130_1475 ();
 b15zdnd11an1n32x5 FILLER_130_1539 ();
 b15zdnd11an1n08x5 FILLER_130_1571 ();
 b15zdnd11an1n16x5 FILLER_130_1631 ();
 b15zdnd11an1n08x5 FILLER_130_1647 ();
 b15zdnd11an1n16x5 FILLER_130_1664 ();
 b15zdnd00an1n02x5 FILLER_130_1680 ();
 b15zdnd11an1n64x5 FILLER_130_1691 ();
 b15zdnd11an1n64x5 FILLER_130_1755 ();
 b15zdnd11an1n32x5 FILLER_130_1819 ();
 b15zdnd11an1n08x5 FILLER_130_1851 ();
 b15zdnd11an1n04x5 FILLER_130_1859 ();
 b15zdnd00an1n02x5 FILLER_130_1863 ();
 b15zdnd11an1n04x5 FILLER_130_1868 ();
 b15zdnd11an1n64x5 FILLER_130_1875 ();
 b15zdnd11an1n32x5 FILLER_130_1939 ();
 b15zdnd11an1n16x5 FILLER_130_1971 ();
 b15zdnd11an1n08x5 FILLER_130_1987 ();
 b15zdnd11an1n04x5 FILLER_130_1995 ();
 b15zdnd00an1n02x5 FILLER_130_1999 ();
 b15zdnd11an1n64x5 FILLER_130_2053 ();
 b15zdnd11an1n32x5 FILLER_130_2117 ();
 b15zdnd11an1n04x5 FILLER_130_2149 ();
 b15zdnd00an1n01x5 FILLER_130_2153 ();
 b15zdnd11an1n64x5 FILLER_130_2162 ();
 b15zdnd11an1n32x5 FILLER_130_2226 ();
 b15zdnd11an1n16x5 FILLER_130_2258 ();
 b15zdnd00an1n02x5 FILLER_130_2274 ();
 b15zdnd11an1n16x5 FILLER_131_0 ();
 b15zdnd11an1n08x5 FILLER_131_16 ();
 b15zdnd11an1n04x5 FILLER_131_24 ();
 b15zdnd11an1n64x5 FILLER_131_31 ();
 b15zdnd11an1n16x5 FILLER_131_95 ();
 b15zdnd11an1n04x5 FILLER_131_111 ();
 b15zdnd11an1n64x5 FILLER_131_157 ();
 b15zdnd11an1n64x5 FILLER_131_221 ();
 b15zdnd11an1n64x5 FILLER_131_285 ();
 b15zdnd11an1n64x5 FILLER_131_349 ();
 b15zdnd11an1n64x5 FILLER_131_413 ();
 b15zdnd11an1n32x5 FILLER_131_477 ();
 b15zdnd11an1n04x5 FILLER_131_509 ();
 b15zdnd11an1n04x5 FILLER_131_516 ();
 b15zdnd11an1n64x5 FILLER_131_523 ();
 b15zdnd11an1n64x5 FILLER_131_587 ();
 b15zdnd11an1n32x5 FILLER_131_651 ();
 b15zdnd00an1n01x5 FILLER_131_683 ();
 b15zdnd11an1n04x5 FILLER_131_716 ();
 b15zdnd11an1n64x5 FILLER_131_723 ();
 b15zdnd11an1n64x5 FILLER_131_787 ();
 b15zdnd11an1n64x5 FILLER_131_851 ();
 b15zdnd11an1n64x5 FILLER_131_915 ();
 b15zdnd11an1n64x5 FILLER_131_979 ();
 b15zdnd11an1n64x5 FILLER_131_1043 ();
 b15zdnd11an1n64x5 FILLER_131_1107 ();
 b15zdnd11an1n32x5 FILLER_131_1171 ();
 b15zdnd11an1n08x5 FILLER_131_1203 ();
 b15zdnd11an1n04x5 FILLER_131_1211 ();
 b15zdnd11an1n64x5 FILLER_131_1218 ();
 b15zdnd11an1n64x5 FILLER_131_1282 ();
 b15zdnd11an1n64x5 FILLER_131_1346 ();
 b15zdnd11an1n64x5 FILLER_131_1410 ();
 b15zdnd11an1n64x5 FILLER_131_1474 ();
 b15zdnd11an1n32x5 FILLER_131_1538 ();
 b15zdnd11an1n16x5 FILLER_131_1573 ();
 b15zdnd11an1n08x5 FILLER_131_1589 ();
 b15zdnd11an1n04x5 FILLER_131_1597 ();
 b15zdnd11an1n04x5 FILLER_131_1604 ();
 b15zdnd11an1n64x5 FILLER_131_1611 ();
 b15zdnd11an1n64x5 FILLER_131_1675 ();
 b15zdnd11an1n64x5 FILLER_131_1739 ();
 b15zdnd11an1n32x5 FILLER_131_1803 ();
 b15zdnd11an1n04x5 FILLER_131_1835 ();
 b15zdnd00an1n02x5 FILLER_131_1839 ();
 b15zdnd00an1n01x5 FILLER_131_1841 ();
 b15zdnd11an1n64x5 FILLER_131_1894 ();
 b15zdnd11an1n64x5 FILLER_131_1958 ();
 b15zdnd00an1n01x5 FILLER_131_2022 ();
 b15zdnd11an1n64x5 FILLER_131_2026 ();
 b15zdnd11an1n64x5 FILLER_131_2090 ();
 b15zdnd11an1n32x5 FILLER_131_2154 ();
 b15zdnd11an1n16x5 FILLER_131_2186 ();
 b15zdnd11an1n04x5 FILLER_131_2202 ();
 b15zdnd11an1n64x5 FILLER_131_2214 ();
 b15zdnd11an1n04x5 FILLER_131_2278 ();
 b15zdnd00an1n02x5 FILLER_131_2282 ();
 b15zdnd11an1n16x5 FILLER_132_8 ();
 b15zdnd11an1n04x5 FILLER_132_24 ();
 b15zdnd00an1n02x5 FILLER_132_28 ();
 b15zdnd11an1n64x5 FILLER_132_33 ();
 b15zdnd11an1n64x5 FILLER_132_97 ();
 b15zdnd11an1n64x5 FILLER_132_161 ();
 b15zdnd11an1n64x5 FILLER_132_225 ();
 b15zdnd11an1n32x5 FILLER_132_289 ();
 b15zdnd11an1n08x5 FILLER_132_321 ();
 b15zdnd11an1n04x5 FILLER_132_329 ();
 b15zdnd00an1n02x5 FILLER_132_333 ();
 b15zdnd11an1n64x5 FILLER_132_377 ();
 b15zdnd11an1n64x5 FILLER_132_441 ();
 b15zdnd11an1n64x5 FILLER_132_505 ();
 b15zdnd11an1n64x5 FILLER_132_569 ();
 b15zdnd11an1n32x5 FILLER_132_633 ();
 b15zdnd00an1n02x5 FILLER_132_665 ();
 b15zdnd00an1n01x5 FILLER_132_667 ();
 b15zdnd11an1n08x5 FILLER_132_710 ();
 b15zdnd11an1n64x5 FILLER_132_726 ();
 b15zdnd11an1n64x5 FILLER_132_790 ();
 b15zdnd11an1n64x5 FILLER_132_854 ();
 b15zdnd11an1n64x5 FILLER_132_918 ();
 b15zdnd11an1n64x5 FILLER_132_982 ();
 b15zdnd11an1n64x5 FILLER_132_1046 ();
 b15zdnd11an1n64x5 FILLER_132_1110 ();
 b15zdnd11an1n32x5 FILLER_132_1174 ();
 b15zdnd11an1n08x5 FILLER_132_1206 ();
 b15zdnd00an1n01x5 FILLER_132_1214 ();
 b15zdnd11an1n04x5 FILLER_132_1218 ();
 b15zdnd00an1n02x5 FILLER_132_1222 ();
 b15zdnd00an1n01x5 FILLER_132_1224 ();
 b15zdnd11an1n64x5 FILLER_132_1267 ();
 b15zdnd11an1n64x5 FILLER_132_1331 ();
 b15zdnd11an1n64x5 FILLER_132_1395 ();
 b15zdnd11an1n16x5 FILLER_132_1459 ();
 b15zdnd00an1n02x5 FILLER_132_1475 ();
 b15zdnd00an1n01x5 FILLER_132_1477 ();
 b15zdnd11an1n64x5 FILLER_132_1483 ();
 b15zdnd11an1n64x5 FILLER_132_1547 ();
 b15zdnd11an1n64x5 FILLER_132_1611 ();
 b15zdnd11an1n04x5 FILLER_132_1675 ();
 b15zdnd00an1n02x5 FILLER_132_1679 ();
 b15zdnd11an1n64x5 FILLER_132_1690 ();
 b15zdnd11an1n64x5 FILLER_132_1754 ();
 b15zdnd11an1n16x5 FILLER_132_1818 ();
 b15zdnd11an1n08x5 FILLER_132_1834 ();
 b15zdnd11an1n04x5 FILLER_132_1842 ();
 b15zdnd00an1n02x5 FILLER_132_1846 ();
 b15zdnd11an1n04x5 FILLER_132_1859 ();
 b15zdnd00an1n01x5 FILLER_132_1863 ();
 b15zdnd11an1n64x5 FILLER_132_1867 ();
 b15zdnd11an1n64x5 FILLER_132_1931 ();
 b15zdnd11an1n64x5 FILLER_132_1995 ();
 b15zdnd11an1n64x5 FILLER_132_2059 ();
 b15zdnd11an1n16x5 FILLER_132_2123 ();
 b15zdnd11an1n08x5 FILLER_132_2139 ();
 b15zdnd11an1n04x5 FILLER_132_2147 ();
 b15zdnd00an1n02x5 FILLER_132_2151 ();
 b15zdnd00an1n01x5 FILLER_132_2153 ();
 b15zdnd11an1n64x5 FILLER_132_2162 ();
 b15zdnd11an1n32x5 FILLER_132_2226 ();
 b15zdnd11an1n16x5 FILLER_132_2258 ();
 b15zdnd00an1n02x5 FILLER_132_2274 ();
 b15zdnd11an1n32x5 FILLER_133_0 ();
 b15zdnd00an1n02x5 FILLER_133_32 ();
 b15zdnd11an1n64x5 FILLER_133_38 ();
 b15zdnd11an1n16x5 FILLER_133_102 ();
 b15zdnd11an1n08x5 FILLER_133_118 ();
 b15zdnd00an1n01x5 FILLER_133_126 ();
 b15zdnd11an1n08x5 FILLER_133_169 ();
 b15zdnd11an1n04x5 FILLER_133_177 ();
 b15zdnd00an1n01x5 FILLER_133_181 ();
 b15zdnd11an1n64x5 FILLER_133_185 ();
 b15zdnd11an1n64x5 FILLER_133_249 ();
 b15zdnd11an1n64x5 FILLER_133_313 ();
 b15zdnd11an1n64x5 FILLER_133_377 ();
 b15zdnd11an1n64x5 FILLER_133_441 ();
 b15zdnd11an1n64x5 FILLER_133_505 ();
 b15zdnd11an1n32x5 FILLER_133_569 ();
 b15zdnd11an1n16x5 FILLER_133_601 ();
 b15zdnd11an1n04x5 FILLER_133_617 ();
 b15zdnd00an1n01x5 FILLER_133_621 ();
 b15zdnd11an1n16x5 FILLER_133_656 ();
 b15zdnd11an1n04x5 FILLER_133_672 ();
 b15zdnd00an1n01x5 FILLER_133_676 ();
 b15zdnd11an1n64x5 FILLER_133_719 ();
 b15zdnd11an1n64x5 FILLER_133_783 ();
 b15zdnd11an1n32x5 FILLER_133_847 ();
 b15zdnd11an1n64x5 FILLER_133_921 ();
 b15zdnd11an1n64x5 FILLER_133_985 ();
 b15zdnd11an1n08x5 FILLER_133_1049 ();
 b15zdnd11an1n04x5 FILLER_133_1057 ();
 b15zdnd00an1n02x5 FILLER_133_1061 ();
 b15zdnd00an1n01x5 FILLER_133_1063 ();
 b15zdnd11an1n64x5 FILLER_133_1081 ();
 b15zdnd11an1n32x5 FILLER_133_1145 ();
 b15zdnd11an1n08x5 FILLER_133_1177 ();
 b15zdnd11an1n04x5 FILLER_133_1185 ();
 b15zdnd00an1n01x5 FILLER_133_1189 ();
 b15zdnd11an1n04x5 FILLER_133_1242 ();
 b15zdnd11an1n04x5 FILLER_133_1253 ();
 b15zdnd00an1n01x5 FILLER_133_1257 ();
 b15zdnd11an1n04x5 FILLER_133_1261 ();
 b15zdnd00an1n01x5 FILLER_133_1265 ();
 b15zdnd11an1n64x5 FILLER_133_1269 ();
 b15zdnd11an1n64x5 FILLER_133_1333 ();
 b15zdnd11an1n64x5 FILLER_133_1397 ();
 b15zdnd11an1n64x5 FILLER_133_1461 ();
 b15zdnd11an1n64x5 FILLER_133_1525 ();
 b15zdnd11an1n64x5 FILLER_133_1589 ();
 b15zdnd11an1n64x5 FILLER_133_1653 ();
 b15zdnd11an1n64x5 FILLER_133_1717 ();
 b15zdnd11an1n64x5 FILLER_133_1781 ();
 b15zdnd11an1n64x5 FILLER_133_1845 ();
 b15zdnd11an1n64x5 FILLER_133_1909 ();
 b15zdnd11an1n64x5 FILLER_133_1973 ();
 b15zdnd11an1n64x5 FILLER_133_2037 ();
 b15zdnd11an1n64x5 FILLER_133_2101 ();
 b15zdnd11an1n64x5 FILLER_133_2165 ();
 b15zdnd11an1n32x5 FILLER_133_2229 ();
 b15zdnd11an1n16x5 FILLER_133_2261 ();
 b15zdnd11an1n04x5 FILLER_133_2277 ();
 b15zdnd00an1n02x5 FILLER_133_2281 ();
 b15zdnd00an1n01x5 FILLER_133_2283 ();
 b15zdnd11an1n04x5 FILLER_134_8 ();
 b15zdnd00an1n01x5 FILLER_134_12 ();
 b15zdnd11an1n64x5 FILLER_134_55 ();
 b15zdnd11an1n32x5 FILLER_134_119 ();
 b15zdnd11an1n08x5 FILLER_134_151 ();
 b15zdnd00an1n02x5 FILLER_134_159 ();
 b15zdnd11an1n16x5 FILLER_134_203 ();
 b15zdnd11an1n04x5 FILLER_134_219 ();
 b15zdnd00an1n02x5 FILLER_134_223 ();
 b15zdnd11an1n64x5 FILLER_134_267 ();
 b15zdnd11an1n64x5 FILLER_134_331 ();
 b15zdnd11an1n64x5 FILLER_134_395 ();
 b15zdnd11an1n64x5 FILLER_134_459 ();
 b15zdnd11an1n64x5 FILLER_134_523 ();
 b15zdnd11an1n32x5 FILLER_134_587 ();
 b15zdnd11an1n16x5 FILLER_134_619 ();
 b15zdnd11an1n08x5 FILLER_134_635 ();
 b15zdnd11an1n04x5 FILLER_134_643 ();
 b15zdnd00an1n02x5 FILLER_134_647 ();
 b15zdnd00an1n01x5 FILLER_134_649 ();
 b15zdnd11an1n04x5 FILLER_134_653 ();
 b15zdnd11an1n32x5 FILLER_134_660 ();
 b15zdnd11an1n16x5 FILLER_134_692 ();
 b15zdnd11an1n04x5 FILLER_134_708 ();
 b15zdnd00an1n01x5 FILLER_134_712 ();
 b15zdnd00an1n02x5 FILLER_134_716 ();
 b15zdnd11an1n32x5 FILLER_134_726 ();
 b15zdnd11an1n16x5 FILLER_134_758 ();
 b15zdnd11an1n04x5 FILLER_134_774 ();
 b15zdnd11an1n64x5 FILLER_134_820 ();
 b15zdnd11an1n64x5 FILLER_134_884 ();
 b15zdnd11an1n64x5 FILLER_134_948 ();
 b15zdnd11an1n64x5 FILLER_134_1012 ();
 b15zdnd11an1n64x5 FILLER_134_1076 ();
 b15zdnd11an1n32x5 FILLER_134_1140 ();
 b15zdnd11an1n16x5 FILLER_134_1172 ();
 b15zdnd00an1n02x5 FILLER_134_1188 ();
 b15zdnd11an1n04x5 FILLER_134_1242 ();
 b15zdnd00an1n01x5 FILLER_134_1246 ();
 b15zdnd11an1n64x5 FILLER_134_1289 ();
 b15zdnd11an1n64x5 FILLER_134_1353 ();
 b15zdnd11an1n64x5 FILLER_134_1417 ();
 b15zdnd11an1n64x5 FILLER_134_1481 ();
 b15zdnd11an1n32x5 FILLER_134_1545 ();
 b15zdnd11an1n16x5 FILLER_134_1577 ();
 b15zdnd00an1n01x5 FILLER_134_1593 ();
 b15zdnd11an1n64x5 FILLER_134_1597 ();
 b15zdnd11an1n64x5 FILLER_134_1661 ();
 b15zdnd11an1n16x5 FILLER_134_1725 ();
 b15zdnd11an1n08x5 FILLER_134_1741 ();
 b15zdnd11an1n04x5 FILLER_134_1752 ();
 b15zdnd11an1n64x5 FILLER_134_1759 ();
 b15zdnd11an1n64x5 FILLER_134_1823 ();
 b15zdnd11an1n64x5 FILLER_134_1887 ();
 b15zdnd11an1n64x5 FILLER_134_1951 ();
 b15zdnd11an1n64x5 FILLER_134_2015 ();
 b15zdnd11an1n64x5 FILLER_134_2079 ();
 b15zdnd11an1n08x5 FILLER_134_2143 ();
 b15zdnd00an1n02x5 FILLER_134_2151 ();
 b15zdnd00an1n01x5 FILLER_134_2153 ();
 b15zdnd11an1n64x5 FILLER_134_2162 ();
 b15zdnd11an1n32x5 FILLER_134_2226 ();
 b15zdnd11an1n16x5 FILLER_134_2258 ();
 b15zdnd00an1n02x5 FILLER_134_2274 ();
 b15zdnd11an1n16x5 FILLER_135_0 ();
 b15zdnd11an1n08x5 FILLER_135_16 ();
 b15zdnd11an1n04x5 FILLER_135_24 ();
 b15zdnd00an1n02x5 FILLER_135_28 ();
 b15zdnd00an1n01x5 FILLER_135_30 ();
 b15zdnd11an1n64x5 FILLER_135_41 ();
 b15zdnd11an1n32x5 FILLER_135_105 ();
 b15zdnd11an1n16x5 FILLER_135_137 ();
 b15zdnd00an1n02x5 FILLER_135_153 ();
 b15zdnd11an1n64x5 FILLER_135_207 ();
 b15zdnd11an1n64x5 FILLER_135_277 ();
 b15zdnd11an1n64x5 FILLER_135_341 ();
 b15zdnd11an1n64x5 FILLER_135_405 ();
 b15zdnd11an1n64x5 FILLER_135_469 ();
 b15zdnd11an1n64x5 FILLER_135_533 ();
 b15zdnd11an1n64x5 FILLER_135_597 ();
 b15zdnd11an1n32x5 FILLER_135_661 ();
 b15zdnd11an1n08x5 FILLER_135_693 ();
 b15zdnd11an1n64x5 FILLER_135_709 ();
 b15zdnd11an1n16x5 FILLER_135_773 ();
 b15zdnd11an1n64x5 FILLER_135_792 ();
 b15zdnd11an1n08x5 FILLER_135_859 ();
 b15zdnd11an1n04x5 FILLER_135_867 ();
 b15zdnd11an1n64x5 FILLER_135_886 ();
 b15zdnd11an1n64x5 FILLER_135_950 ();
 b15zdnd11an1n64x5 FILLER_135_1014 ();
 b15zdnd11an1n64x5 FILLER_135_1078 ();
 b15zdnd11an1n64x5 FILLER_135_1142 ();
 b15zdnd00an1n02x5 FILLER_135_1206 ();
 b15zdnd11an1n04x5 FILLER_135_1211 ();
 b15zdnd11an1n04x5 FILLER_135_1218 ();
 b15zdnd11an1n08x5 FILLER_135_1225 ();
 b15zdnd00an1n01x5 FILLER_135_1233 ();
 b15zdnd11an1n64x5 FILLER_135_1286 ();
 b15zdnd11an1n64x5 FILLER_135_1350 ();
 b15zdnd11an1n32x5 FILLER_135_1414 ();
 b15zdnd11an1n16x5 FILLER_135_1446 ();
 b15zdnd11an1n04x5 FILLER_135_1462 ();
 b15zdnd11an1n16x5 FILLER_135_1471 ();
 b15zdnd11an1n08x5 FILLER_135_1487 ();
 b15zdnd11an1n04x5 FILLER_135_1495 ();
 b15zdnd11an1n32x5 FILLER_135_1507 ();
 b15zdnd11an1n16x5 FILLER_135_1539 ();
 b15zdnd11an1n08x5 FILLER_135_1555 ();
 b15zdnd11an1n04x5 FILLER_135_1563 ();
 b15zdnd00an1n01x5 FILLER_135_1567 ();
 b15zdnd11an1n64x5 FILLER_135_1620 ();
 b15zdnd11an1n32x5 FILLER_135_1684 ();
 b15zdnd11an1n08x5 FILLER_135_1716 ();
 b15zdnd11an1n04x5 FILLER_135_1724 ();
 b15zdnd00an1n02x5 FILLER_135_1728 ();
 b15zdnd00an1n01x5 FILLER_135_1730 ();
 b15zdnd11an1n64x5 FILLER_135_1783 ();
 b15zdnd11an1n64x5 FILLER_135_1847 ();
 b15zdnd11an1n32x5 FILLER_135_1911 ();
 b15zdnd11an1n16x5 FILLER_135_1943 ();
 b15zdnd00an1n01x5 FILLER_135_1959 ();
 b15zdnd11an1n64x5 FILLER_135_1969 ();
 b15zdnd11an1n64x5 FILLER_135_2033 ();
 b15zdnd11an1n64x5 FILLER_135_2097 ();
 b15zdnd11an1n64x5 FILLER_135_2161 ();
 b15zdnd11an1n32x5 FILLER_135_2225 ();
 b15zdnd11an1n16x5 FILLER_135_2257 ();
 b15zdnd11an1n08x5 FILLER_135_2273 ();
 b15zdnd00an1n02x5 FILLER_135_2281 ();
 b15zdnd00an1n01x5 FILLER_135_2283 ();
 b15zdnd11an1n16x5 FILLER_136_8 ();
 b15zdnd11an1n04x5 FILLER_136_24 ();
 b15zdnd00an1n01x5 FILLER_136_28 ();
 b15zdnd11an1n04x5 FILLER_136_32 ();
 b15zdnd11an1n64x5 FILLER_136_42 ();
 b15zdnd11an1n64x5 FILLER_136_106 ();
 b15zdnd00an1n02x5 FILLER_136_170 ();
 b15zdnd00an1n01x5 FILLER_136_172 ();
 b15zdnd11an1n04x5 FILLER_136_176 ();
 b15zdnd11an1n08x5 FILLER_136_183 ();
 b15zdnd00an1n02x5 FILLER_136_191 ();
 b15zdnd00an1n01x5 FILLER_136_193 ();
 b15zdnd11an1n64x5 FILLER_136_236 ();
 b15zdnd11an1n64x5 FILLER_136_300 ();
 b15zdnd11an1n64x5 FILLER_136_364 ();
 b15zdnd11an1n64x5 FILLER_136_428 ();
 b15zdnd11an1n64x5 FILLER_136_492 ();
 b15zdnd11an1n64x5 FILLER_136_556 ();
 b15zdnd11an1n64x5 FILLER_136_620 ();
 b15zdnd11an1n32x5 FILLER_136_684 ();
 b15zdnd00an1n02x5 FILLER_136_716 ();
 b15zdnd11an1n32x5 FILLER_136_726 ();
 b15zdnd11an1n08x5 FILLER_136_758 ();
 b15zdnd11an1n04x5 FILLER_136_766 ();
 b15zdnd00an1n02x5 FILLER_136_770 ();
 b15zdnd00an1n01x5 FILLER_136_772 ();
 b15zdnd11an1n04x5 FILLER_136_825 ();
 b15zdnd11an1n64x5 FILLER_136_881 ();
 b15zdnd11an1n64x5 FILLER_136_945 ();
 b15zdnd11an1n16x5 FILLER_136_1009 ();
 b15zdnd11an1n08x5 FILLER_136_1025 ();
 b15zdnd00an1n01x5 FILLER_136_1033 ();
 b15zdnd11an1n16x5 FILLER_136_1037 ();
 b15zdnd11an1n04x5 FILLER_136_1053 ();
 b15zdnd11an1n64x5 FILLER_136_1067 ();
 b15zdnd11an1n64x5 FILLER_136_1131 ();
 b15zdnd11an1n16x5 FILLER_136_1195 ();
 b15zdnd11an1n04x5 FILLER_136_1211 ();
 b15zdnd11an1n08x5 FILLER_136_1218 ();
 b15zdnd11an1n04x5 FILLER_136_1226 ();
 b15zdnd00an1n02x5 FILLER_136_1230 ();
 b15zdnd00an1n01x5 FILLER_136_1232 ();
 b15zdnd11an1n04x5 FILLER_136_1242 ();
 b15zdnd11an1n64x5 FILLER_136_1288 ();
 b15zdnd11an1n64x5 FILLER_136_1352 ();
 b15zdnd11an1n64x5 FILLER_136_1416 ();
 b15zdnd11an1n64x5 FILLER_136_1480 ();
 b15zdnd11an1n32x5 FILLER_136_1544 ();
 b15zdnd11an1n16x5 FILLER_136_1576 ();
 b15zdnd00an1n01x5 FILLER_136_1592 ();
 b15zdnd11an1n64x5 FILLER_136_1596 ();
 b15zdnd11an1n64x5 FILLER_136_1660 ();
 b15zdnd11an1n32x5 FILLER_136_1724 ();
 b15zdnd11an1n64x5 FILLER_136_1759 ();
 b15zdnd11an1n64x5 FILLER_136_1823 ();
 b15zdnd11an1n64x5 FILLER_136_1887 ();
 b15zdnd11an1n64x5 FILLER_136_1951 ();
 b15zdnd11an1n64x5 FILLER_136_2015 ();
 b15zdnd11an1n64x5 FILLER_136_2079 ();
 b15zdnd11an1n08x5 FILLER_136_2143 ();
 b15zdnd00an1n02x5 FILLER_136_2151 ();
 b15zdnd00an1n01x5 FILLER_136_2153 ();
 b15zdnd11an1n64x5 FILLER_136_2162 ();
 b15zdnd11an1n32x5 FILLER_136_2226 ();
 b15zdnd11an1n16x5 FILLER_136_2258 ();
 b15zdnd00an1n02x5 FILLER_136_2274 ();
 b15zdnd11an1n04x5 FILLER_137_0 ();
 b15zdnd00an1n01x5 FILLER_137_4 ();
 b15zdnd11an1n16x5 FILLER_137_9 ();
 b15zdnd11an1n04x5 FILLER_137_25 ();
 b15zdnd11an1n04x5 FILLER_137_32 ();
 b15zdnd00an1n02x5 FILLER_137_36 ();
 b15zdnd11an1n64x5 FILLER_137_43 ();
 b15zdnd11an1n64x5 FILLER_137_107 ();
 b15zdnd11an1n64x5 FILLER_137_171 ();
 b15zdnd11an1n08x5 FILLER_137_235 ();
 b15zdnd00an1n01x5 FILLER_137_243 ();
 b15zdnd11an1n64x5 FILLER_137_253 ();
 b15zdnd00an1n02x5 FILLER_137_317 ();
 b15zdnd00an1n01x5 FILLER_137_319 ();
 b15zdnd11an1n64x5 FILLER_137_362 ();
 b15zdnd11an1n64x5 FILLER_137_426 ();
 b15zdnd11an1n08x5 FILLER_137_490 ();
 b15zdnd11an1n04x5 FILLER_137_498 ();
 b15zdnd00an1n01x5 FILLER_137_502 ();
 b15zdnd11an1n32x5 FILLER_137_519 ();
 b15zdnd11an1n08x5 FILLER_137_551 ();
 b15zdnd00an1n02x5 FILLER_137_559 ();
 b15zdnd00an1n01x5 FILLER_137_561 ();
 b15zdnd11an1n32x5 FILLER_137_582 ();
 b15zdnd11an1n08x5 FILLER_137_614 ();
 b15zdnd11an1n04x5 FILLER_137_622 ();
 b15zdnd00an1n02x5 FILLER_137_626 ();
 b15zdnd00an1n01x5 FILLER_137_628 ();
 b15zdnd11an1n64x5 FILLER_137_671 ();
 b15zdnd11an1n64x5 FILLER_137_735 ();
 b15zdnd11an1n64x5 FILLER_137_799 ();
 b15zdnd11an1n64x5 FILLER_137_863 ();
 b15zdnd11an1n64x5 FILLER_137_927 ();
 b15zdnd11an1n16x5 FILLER_137_991 ();
 b15zdnd11an1n08x5 FILLER_137_1007 ();
 b15zdnd11an1n04x5 FILLER_137_1015 ();
 b15zdnd11an1n16x5 FILLER_137_1047 ();
 b15zdnd11an1n04x5 FILLER_137_1063 ();
 b15zdnd00an1n02x5 FILLER_137_1067 ();
 b15zdnd11an1n64x5 FILLER_137_1093 ();
 b15zdnd11an1n64x5 FILLER_137_1157 ();
 b15zdnd11an1n16x5 FILLER_137_1221 ();
 b15zdnd11an1n04x5 FILLER_137_1246 ();
 b15zdnd11an1n64x5 FILLER_137_1292 ();
 b15zdnd11an1n64x5 FILLER_137_1356 ();
 b15zdnd11an1n64x5 FILLER_137_1420 ();
 b15zdnd11an1n64x5 FILLER_137_1484 ();
 b15zdnd11an1n32x5 FILLER_137_1548 ();
 b15zdnd11an1n08x5 FILLER_137_1580 ();
 b15zdnd11an1n04x5 FILLER_137_1588 ();
 b15zdnd00an1n01x5 FILLER_137_1592 ();
 b15zdnd11an1n64x5 FILLER_137_1596 ();
 b15zdnd11an1n32x5 FILLER_137_1660 ();
 b15zdnd11an1n16x5 FILLER_137_1692 ();
 b15zdnd11an1n04x5 FILLER_137_1708 ();
 b15zdnd00an1n02x5 FILLER_137_1712 ();
 b15zdnd00an1n01x5 FILLER_137_1714 ();
 b15zdnd11an1n64x5 FILLER_137_1726 ();
 b15zdnd11an1n64x5 FILLER_137_1790 ();
 b15zdnd11an1n64x5 FILLER_137_1854 ();
 b15zdnd11an1n64x5 FILLER_137_1918 ();
 b15zdnd11an1n64x5 FILLER_137_1982 ();
 b15zdnd11an1n64x5 FILLER_137_2046 ();
 b15zdnd11an1n64x5 FILLER_137_2110 ();
 b15zdnd11an1n64x5 FILLER_137_2174 ();
 b15zdnd11an1n32x5 FILLER_137_2238 ();
 b15zdnd11an1n08x5 FILLER_137_2270 ();
 b15zdnd11an1n04x5 FILLER_137_2278 ();
 b15zdnd00an1n02x5 FILLER_137_2282 ();
 b15zdnd00an1n02x5 FILLER_138_8 ();
 b15zdnd11an1n64x5 FILLER_138_52 ();
 b15zdnd11an1n16x5 FILLER_138_116 ();
 b15zdnd11an1n08x5 FILLER_138_132 ();
 b15zdnd11an1n04x5 FILLER_138_140 ();
 b15zdnd00an1n02x5 FILLER_138_144 ();
 b15zdnd00an1n01x5 FILLER_138_146 ();
 b15zdnd11an1n64x5 FILLER_138_153 ();
 b15zdnd11an1n64x5 FILLER_138_217 ();
 b15zdnd11an1n64x5 FILLER_138_281 ();
 b15zdnd11an1n64x5 FILLER_138_345 ();
 b15zdnd11an1n32x5 FILLER_138_409 ();
 b15zdnd11an1n16x5 FILLER_138_441 ();
 b15zdnd11an1n04x5 FILLER_138_457 ();
 b15zdnd00an1n01x5 FILLER_138_461 ();
 b15zdnd11an1n04x5 FILLER_138_504 ();
 b15zdnd11an1n32x5 FILLER_138_515 ();
 b15zdnd11an1n04x5 FILLER_138_547 ();
 b15zdnd00an1n02x5 FILLER_138_551 ();
 b15zdnd11an1n64x5 FILLER_138_605 ();
 b15zdnd11an1n16x5 FILLER_138_669 ();
 b15zdnd11an1n08x5 FILLER_138_685 ();
 b15zdnd00an1n02x5 FILLER_138_693 ();
 b15zdnd11an1n16x5 FILLER_138_701 ();
 b15zdnd00an1n01x5 FILLER_138_717 ();
 b15zdnd11an1n32x5 FILLER_138_726 ();
 b15zdnd11an1n16x5 FILLER_138_758 ();
 b15zdnd11an1n08x5 FILLER_138_774 ();
 b15zdnd11an1n04x5 FILLER_138_782 ();
 b15zdnd00an1n02x5 FILLER_138_786 ();
 b15zdnd11an1n04x5 FILLER_138_791 ();
 b15zdnd00an1n02x5 FILLER_138_795 ();
 b15zdnd00an1n01x5 FILLER_138_797 ();
 b15zdnd11an1n32x5 FILLER_138_801 ();
 b15zdnd11an1n08x5 FILLER_138_833 ();
 b15zdnd00an1n01x5 FILLER_138_841 ();
 b15zdnd11an1n04x5 FILLER_138_845 ();
 b15zdnd11an1n04x5 FILLER_138_852 ();
 b15zdnd11an1n04x5 FILLER_138_859 ();
 b15zdnd11an1n32x5 FILLER_138_915 ();
 b15zdnd11an1n08x5 FILLER_138_947 ();
 b15zdnd00an1n01x5 FILLER_138_955 ();
 b15zdnd11an1n16x5 FILLER_138_959 ();
 b15zdnd11an1n04x5 FILLER_138_975 ();
 b15zdnd00an1n02x5 FILLER_138_979 ();
 b15zdnd11an1n64x5 FILLER_138_989 ();
 b15zdnd11an1n64x5 FILLER_138_1053 ();
 b15zdnd11an1n64x5 FILLER_138_1117 ();
 b15zdnd11an1n32x5 FILLER_138_1181 ();
 b15zdnd11an1n16x5 FILLER_138_1213 ();
 b15zdnd11an1n08x5 FILLER_138_1229 ();
 b15zdnd00an1n02x5 FILLER_138_1237 ();
 b15zdnd11an1n04x5 FILLER_138_1242 ();
 b15zdnd11an1n64x5 FILLER_138_1288 ();
 b15zdnd11an1n64x5 FILLER_138_1352 ();
 b15zdnd11an1n32x5 FILLER_138_1416 ();
 b15zdnd11an1n08x5 FILLER_138_1448 ();
 b15zdnd11an1n04x5 FILLER_138_1456 ();
 b15zdnd00an1n02x5 FILLER_138_1460 ();
 b15zdnd00an1n01x5 FILLER_138_1462 ();
 b15zdnd11an1n64x5 FILLER_138_1505 ();
 b15zdnd11an1n64x5 FILLER_138_1569 ();
 b15zdnd11an1n64x5 FILLER_138_1633 ();
 b15zdnd11an1n32x5 FILLER_138_1697 ();
 b15zdnd11an1n04x5 FILLER_138_1729 ();
 b15zdnd00an1n01x5 FILLER_138_1733 ();
 b15zdnd11an1n04x5 FILLER_138_1737 ();
 b15zdnd11an1n64x5 FILLER_138_1744 ();
 b15zdnd11an1n64x5 FILLER_138_1808 ();
 b15zdnd11an1n64x5 FILLER_138_1872 ();
 b15zdnd11an1n64x5 FILLER_138_1936 ();
 b15zdnd11an1n64x5 FILLER_138_2000 ();
 b15zdnd11an1n64x5 FILLER_138_2064 ();
 b15zdnd11an1n16x5 FILLER_138_2128 ();
 b15zdnd11an1n08x5 FILLER_138_2144 ();
 b15zdnd00an1n02x5 FILLER_138_2152 ();
 b15zdnd11an1n64x5 FILLER_138_2162 ();
 b15zdnd11an1n32x5 FILLER_138_2226 ();
 b15zdnd11an1n16x5 FILLER_138_2258 ();
 b15zdnd00an1n02x5 FILLER_138_2274 ();
 b15zdnd11an1n64x5 FILLER_139_0 ();
 b15zdnd11an1n64x5 FILLER_139_64 ();
 b15zdnd11an1n08x5 FILLER_139_128 ();
 b15zdnd11an1n04x5 FILLER_139_136 ();
 b15zdnd00an1n02x5 FILLER_139_140 ();
 b15zdnd11an1n64x5 FILLER_139_156 ();
 b15zdnd11an1n64x5 FILLER_139_220 ();
 b15zdnd11an1n64x5 FILLER_139_284 ();
 b15zdnd11an1n64x5 FILLER_139_348 ();
 b15zdnd11an1n64x5 FILLER_139_412 ();
 b15zdnd11an1n64x5 FILLER_139_476 ();
 b15zdnd11an1n32x5 FILLER_139_540 ();
 b15zdnd00an1n01x5 FILLER_139_572 ();
 b15zdnd11an1n04x5 FILLER_139_576 ();
 b15zdnd11an1n64x5 FILLER_139_583 ();
 b15zdnd11an1n64x5 FILLER_139_647 ();
 b15zdnd11an1n64x5 FILLER_139_711 ();
 b15zdnd11an1n08x5 FILLER_139_775 ();
 b15zdnd11an1n04x5 FILLER_139_783 ();
 b15zdnd00an1n01x5 FILLER_139_787 ();
 b15zdnd11an1n64x5 FILLER_139_791 ();
 b15zdnd11an1n04x5 FILLER_139_858 ();
 b15zdnd11an1n64x5 FILLER_139_865 ();
 b15zdnd11an1n64x5 FILLER_139_929 ();
 b15zdnd11an1n64x5 FILLER_139_993 ();
 b15zdnd11an1n08x5 FILLER_139_1057 ();
 b15zdnd11an1n64x5 FILLER_139_1070 ();
 b15zdnd11an1n64x5 FILLER_139_1134 ();
 b15zdnd11an1n16x5 FILLER_139_1198 ();
 b15zdnd11an1n08x5 FILLER_139_1214 ();
 b15zdnd11an1n04x5 FILLER_139_1222 ();
 b15zdnd11an1n04x5 FILLER_139_1258 ();
 b15zdnd11an1n04x5 FILLER_139_1265 ();
 b15zdnd11an1n04x5 FILLER_139_1276 ();
 b15zdnd11an1n64x5 FILLER_139_1283 ();
 b15zdnd11an1n32x5 FILLER_139_1347 ();
 b15zdnd11an1n16x5 FILLER_139_1379 ();
 b15zdnd11an1n08x5 FILLER_139_1395 ();
 b15zdnd11an1n04x5 FILLER_139_1403 ();
 b15zdnd00an1n02x5 FILLER_139_1407 ();
 b15zdnd00an1n01x5 FILLER_139_1409 ();
 b15zdnd11an1n64x5 FILLER_139_1452 ();
 b15zdnd11an1n64x5 FILLER_139_1516 ();
 b15zdnd11an1n64x5 FILLER_139_1580 ();
 b15zdnd11an1n64x5 FILLER_139_1644 ();
 b15zdnd11an1n08x5 FILLER_139_1708 ();
 b15zdnd11an1n64x5 FILLER_139_1768 ();
 b15zdnd11an1n64x5 FILLER_139_1832 ();
 b15zdnd11an1n64x5 FILLER_139_1896 ();
 b15zdnd00an1n01x5 FILLER_139_1960 ();
 b15zdnd11an1n64x5 FILLER_139_1970 ();
 b15zdnd11an1n64x5 FILLER_139_2034 ();
 b15zdnd11an1n64x5 FILLER_139_2098 ();
 b15zdnd11an1n64x5 FILLER_139_2162 ();
 b15zdnd11an1n32x5 FILLER_139_2226 ();
 b15zdnd11an1n16x5 FILLER_139_2258 ();
 b15zdnd11an1n08x5 FILLER_139_2274 ();
 b15zdnd00an1n02x5 FILLER_139_2282 ();
 b15zdnd11an1n64x5 FILLER_140_8 ();
 b15zdnd11an1n64x5 FILLER_140_72 ();
 b15zdnd11an1n08x5 FILLER_140_136 ();
 b15zdnd00an1n02x5 FILLER_140_144 ();
 b15zdnd11an1n64x5 FILLER_140_149 ();
 b15zdnd11an1n16x5 FILLER_140_213 ();
 b15zdnd11an1n08x5 FILLER_140_229 ();
 b15zdnd00an1n01x5 FILLER_140_237 ();
 b15zdnd11an1n04x5 FILLER_140_244 ();
 b15zdnd11an1n16x5 FILLER_140_254 ();
 b15zdnd11an1n32x5 FILLER_140_277 ();
 b15zdnd00an1n02x5 FILLER_140_309 ();
 b15zdnd11an1n64x5 FILLER_140_353 ();
 b15zdnd11an1n64x5 FILLER_140_417 ();
 b15zdnd11an1n64x5 FILLER_140_481 ();
 b15zdnd11an1n32x5 FILLER_140_545 ();
 b15zdnd00an1n01x5 FILLER_140_577 ();
 b15zdnd11an1n64x5 FILLER_140_581 ();
 b15zdnd11an1n32x5 FILLER_140_645 ();
 b15zdnd00an1n01x5 FILLER_140_677 ();
 b15zdnd11an1n16x5 FILLER_140_687 ();
 b15zdnd11an1n08x5 FILLER_140_703 ();
 b15zdnd11an1n04x5 FILLER_140_711 ();
 b15zdnd00an1n02x5 FILLER_140_715 ();
 b15zdnd00an1n01x5 FILLER_140_717 ();
 b15zdnd11an1n32x5 FILLER_140_726 ();
 b15zdnd00an1n02x5 FILLER_140_758 ();
 b15zdnd00an1n01x5 FILLER_140_760 ();
 b15zdnd11an1n64x5 FILLER_140_813 ();
 b15zdnd11an1n64x5 FILLER_140_877 ();
 b15zdnd11an1n64x5 FILLER_140_941 ();
 b15zdnd11an1n64x5 FILLER_140_1005 ();
 b15zdnd11an1n64x5 FILLER_140_1069 ();
 b15zdnd11an1n64x5 FILLER_140_1133 ();
 b15zdnd11an1n32x5 FILLER_140_1197 ();
 b15zdnd11an1n16x5 FILLER_140_1229 ();
 b15zdnd11an1n64x5 FILLER_140_1287 ();
 b15zdnd11an1n64x5 FILLER_140_1351 ();
 b15zdnd11an1n16x5 FILLER_140_1415 ();
 b15zdnd11an1n08x5 FILLER_140_1431 ();
 b15zdnd11an1n04x5 FILLER_140_1439 ();
 b15zdnd11an1n64x5 FILLER_140_1459 ();
 b15zdnd11an1n64x5 FILLER_140_1523 ();
 b15zdnd11an1n64x5 FILLER_140_1587 ();
 b15zdnd11an1n64x5 FILLER_140_1651 ();
 b15zdnd00an1n01x5 FILLER_140_1715 ();
 b15zdnd11an1n04x5 FILLER_140_1719 ();
 b15zdnd00an1n01x5 FILLER_140_1723 ();
 b15zdnd11an1n04x5 FILLER_140_1735 ();
 b15zdnd11an1n04x5 FILLER_140_1742 ();
 b15zdnd11an1n64x5 FILLER_140_1757 ();
 b15zdnd11an1n32x5 FILLER_140_1821 ();
 b15zdnd11an1n08x5 FILLER_140_1853 ();
 b15zdnd11an1n04x5 FILLER_140_1861 ();
 b15zdnd00an1n01x5 FILLER_140_1865 ();
 b15zdnd11an1n32x5 FILLER_140_1893 ();
 b15zdnd11an1n04x5 FILLER_140_1925 ();
 b15zdnd00an1n02x5 FILLER_140_1929 ();
 b15zdnd00an1n01x5 FILLER_140_1931 ();
 b15zdnd11an1n32x5 FILLER_140_1941 ();
 b15zdnd11an1n16x5 FILLER_140_1973 ();
 b15zdnd11an1n08x5 FILLER_140_1989 ();
 b15zdnd11an1n04x5 FILLER_140_1997 ();
 b15zdnd00an1n01x5 FILLER_140_2001 ();
 b15zdnd11an1n64x5 FILLER_140_2013 ();
 b15zdnd11an1n64x5 FILLER_140_2077 ();
 b15zdnd11an1n08x5 FILLER_140_2141 ();
 b15zdnd11an1n04x5 FILLER_140_2149 ();
 b15zdnd00an1n01x5 FILLER_140_2153 ();
 b15zdnd11an1n64x5 FILLER_140_2162 ();
 b15zdnd11an1n32x5 FILLER_140_2226 ();
 b15zdnd11an1n16x5 FILLER_140_2258 ();
 b15zdnd00an1n02x5 FILLER_140_2274 ();
 b15zdnd11an1n64x5 FILLER_141_0 ();
 b15zdnd11an1n64x5 FILLER_141_64 ();
 b15zdnd11an1n64x5 FILLER_141_128 ();
 b15zdnd11an1n16x5 FILLER_141_192 ();
 b15zdnd11an1n08x5 FILLER_141_208 ();
 b15zdnd11an1n04x5 FILLER_141_216 ();
 b15zdnd00an1n02x5 FILLER_141_220 ();
 b15zdnd11an1n08x5 FILLER_141_230 ();
 b15zdnd00an1n02x5 FILLER_141_238 ();
 b15zdnd00an1n01x5 FILLER_141_240 ();
 b15zdnd11an1n64x5 FILLER_141_283 ();
 b15zdnd11an1n64x5 FILLER_141_347 ();
 b15zdnd11an1n64x5 FILLER_141_411 ();
 b15zdnd11an1n64x5 FILLER_141_475 ();
 b15zdnd11an1n64x5 FILLER_141_539 ();
 b15zdnd11an1n64x5 FILLER_141_603 ();
 b15zdnd11an1n64x5 FILLER_141_667 ();
 b15zdnd11an1n32x5 FILLER_141_731 ();
 b15zdnd11an1n16x5 FILLER_141_763 ();
 b15zdnd11an1n04x5 FILLER_141_782 ();
 b15zdnd11an1n64x5 FILLER_141_789 ();
 b15zdnd11an1n64x5 FILLER_141_853 ();
 b15zdnd11an1n32x5 FILLER_141_917 ();
 b15zdnd11an1n16x5 FILLER_141_949 ();
 b15zdnd11an1n08x5 FILLER_141_965 ();
 b15zdnd00an1n01x5 FILLER_141_973 ();
 b15zdnd11an1n64x5 FILLER_141_980 ();
 b15zdnd11an1n64x5 FILLER_141_1044 ();
 b15zdnd11an1n64x5 FILLER_141_1108 ();
 b15zdnd11an1n64x5 FILLER_141_1172 ();
 b15zdnd11an1n04x5 FILLER_141_1268 ();
 b15zdnd11an1n64x5 FILLER_141_1275 ();
 b15zdnd11an1n64x5 FILLER_141_1339 ();
 b15zdnd11an1n64x5 FILLER_141_1403 ();
 b15zdnd11an1n16x5 FILLER_141_1467 ();
 b15zdnd00an1n02x5 FILLER_141_1483 ();
 b15zdnd00an1n01x5 FILLER_141_1485 ();
 b15zdnd11an1n64x5 FILLER_141_1491 ();
 b15zdnd11an1n64x5 FILLER_141_1555 ();
 b15zdnd11an1n64x5 FILLER_141_1619 ();
 b15zdnd11an1n32x5 FILLER_141_1683 ();
 b15zdnd11an1n64x5 FILLER_141_1718 ();
 b15zdnd11an1n64x5 FILLER_141_1782 ();
 b15zdnd11an1n16x5 FILLER_141_1846 ();
 b15zdnd11an1n04x5 FILLER_141_1862 ();
 b15zdnd00an1n02x5 FILLER_141_1866 ();
 b15zdnd00an1n01x5 FILLER_141_1868 ();
 b15zdnd11an1n64x5 FILLER_141_1872 ();
 b15zdnd11an1n64x5 FILLER_141_1936 ();
 b15zdnd11an1n16x5 FILLER_141_2000 ();
 b15zdnd11an1n04x5 FILLER_141_2016 ();
 b15zdnd00an1n02x5 FILLER_141_2020 ();
 b15zdnd11an1n04x5 FILLER_141_2025 ();
 b15zdnd11an1n64x5 FILLER_141_2032 ();
 b15zdnd11an1n64x5 FILLER_141_2096 ();
 b15zdnd11an1n64x5 FILLER_141_2160 ();
 b15zdnd11an1n32x5 FILLER_141_2224 ();
 b15zdnd11an1n16x5 FILLER_141_2256 ();
 b15zdnd11an1n08x5 FILLER_141_2272 ();
 b15zdnd11an1n04x5 FILLER_141_2280 ();
 b15zdnd11an1n64x5 FILLER_142_8 ();
 b15zdnd11an1n64x5 FILLER_142_72 ();
 b15zdnd11an1n64x5 FILLER_142_136 ();
 b15zdnd11an1n16x5 FILLER_142_200 ();
 b15zdnd11an1n08x5 FILLER_142_216 ();
 b15zdnd11an1n04x5 FILLER_142_224 ();
 b15zdnd00an1n01x5 FILLER_142_228 ();
 b15zdnd11an1n04x5 FILLER_142_235 ();
 b15zdnd11an1n64x5 FILLER_142_281 ();
 b15zdnd11an1n64x5 FILLER_142_345 ();
 b15zdnd11an1n64x5 FILLER_142_409 ();
 b15zdnd11an1n64x5 FILLER_142_473 ();
 b15zdnd11an1n64x5 FILLER_142_537 ();
 b15zdnd11an1n64x5 FILLER_142_601 ();
 b15zdnd11an1n32x5 FILLER_142_665 ();
 b15zdnd11an1n16x5 FILLER_142_697 ();
 b15zdnd11an1n04x5 FILLER_142_713 ();
 b15zdnd00an1n01x5 FILLER_142_717 ();
 b15zdnd11an1n64x5 FILLER_142_726 ();
 b15zdnd11an1n64x5 FILLER_142_790 ();
 b15zdnd11an1n64x5 FILLER_142_854 ();
 b15zdnd11an1n16x5 FILLER_142_918 ();
 b15zdnd11an1n08x5 FILLER_142_934 ();
 b15zdnd11an1n04x5 FILLER_142_942 ();
 b15zdnd00an1n01x5 FILLER_142_946 ();
 b15zdnd11an1n64x5 FILLER_142_975 ();
 b15zdnd11an1n64x5 FILLER_142_1039 ();
 b15zdnd11an1n64x5 FILLER_142_1103 ();
 b15zdnd11an1n64x5 FILLER_142_1167 ();
 b15zdnd11an1n16x5 FILLER_142_1231 ();
 b15zdnd11an1n08x5 FILLER_142_1247 ();
 b15zdnd00an1n02x5 FILLER_142_1255 ();
 b15zdnd11an1n64x5 FILLER_142_1260 ();
 b15zdnd11an1n16x5 FILLER_142_1324 ();
 b15zdnd11an1n08x5 FILLER_142_1340 ();
 b15zdnd11an1n04x5 FILLER_142_1348 ();
 b15zdnd11an1n04x5 FILLER_142_1355 ();
 b15zdnd11an1n64x5 FILLER_142_1362 ();
 b15zdnd11an1n64x5 FILLER_142_1426 ();
 b15zdnd11an1n64x5 FILLER_142_1490 ();
 b15zdnd11an1n64x5 FILLER_142_1554 ();
 b15zdnd11an1n64x5 FILLER_142_1618 ();
 b15zdnd11an1n08x5 FILLER_142_1682 ();
 b15zdnd00an1n01x5 FILLER_142_1690 ();
 b15zdnd11an1n64x5 FILLER_142_1743 ();
 b15zdnd11an1n64x5 FILLER_142_1807 ();
 b15zdnd11an1n64x5 FILLER_142_1871 ();
 b15zdnd11an1n64x5 FILLER_142_1935 ();
 b15zdnd11an1n04x5 FILLER_142_1999 ();
 b15zdnd00an1n01x5 FILLER_142_2003 ();
 b15zdnd11an1n64x5 FILLER_142_2056 ();
 b15zdnd11an1n32x5 FILLER_142_2120 ();
 b15zdnd00an1n02x5 FILLER_142_2152 ();
 b15zdnd11an1n64x5 FILLER_142_2162 ();
 b15zdnd11an1n32x5 FILLER_142_2226 ();
 b15zdnd11an1n16x5 FILLER_142_2258 ();
 b15zdnd00an1n02x5 FILLER_142_2274 ();
 b15zdnd11an1n64x5 FILLER_143_0 ();
 b15zdnd11an1n64x5 FILLER_143_64 ();
 b15zdnd11an1n64x5 FILLER_143_128 ();
 b15zdnd11an1n32x5 FILLER_143_192 ();
 b15zdnd11an1n04x5 FILLER_143_224 ();
 b15zdnd00an1n02x5 FILLER_143_228 ();
 b15zdnd11an1n04x5 FILLER_143_236 ();
 b15zdnd00an1n02x5 FILLER_143_240 ();
 b15zdnd11an1n04x5 FILLER_143_251 ();
 b15zdnd11an1n32x5 FILLER_143_297 ();
 b15zdnd11an1n16x5 FILLER_143_329 ();
 b15zdnd11an1n08x5 FILLER_143_345 ();
 b15zdnd11an1n04x5 FILLER_143_353 ();
 b15zdnd00an1n02x5 FILLER_143_357 ();
 b15zdnd11an1n64x5 FILLER_143_365 ();
 b15zdnd11an1n64x5 FILLER_143_429 ();
 b15zdnd11an1n64x5 FILLER_143_493 ();
 b15zdnd11an1n64x5 FILLER_143_557 ();
 b15zdnd11an1n32x5 FILLER_143_621 ();
 b15zdnd11an1n16x5 FILLER_143_653 ();
 b15zdnd11an1n04x5 FILLER_143_669 ();
 b15zdnd00an1n02x5 FILLER_143_673 ();
 b15zdnd11an1n64x5 FILLER_143_697 ();
 b15zdnd11an1n64x5 FILLER_143_761 ();
 b15zdnd11an1n64x5 FILLER_143_825 ();
 b15zdnd11an1n64x5 FILLER_143_889 ();
 b15zdnd11an1n64x5 FILLER_143_953 ();
 b15zdnd11an1n64x5 FILLER_143_1017 ();
 b15zdnd11an1n64x5 FILLER_143_1081 ();
 b15zdnd11an1n64x5 FILLER_143_1145 ();
 b15zdnd11an1n64x5 FILLER_143_1209 ();
 b15zdnd11an1n32x5 FILLER_143_1273 ();
 b15zdnd11an1n16x5 FILLER_143_1305 ();
 b15zdnd11an1n08x5 FILLER_143_1321 ();
 b15zdnd11an1n04x5 FILLER_143_1329 ();
 b15zdnd00an1n02x5 FILLER_143_1333 ();
 b15zdnd00an1n01x5 FILLER_143_1335 ();
 b15zdnd11an1n08x5 FILLER_143_1344 ();
 b15zdnd00an1n01x5 FILLER_143_1352 ();
 b15zdnd11an1n64x5 FILLER_143_1395 ();
 b15zdnd11an1n16x5 FILLER_143_1459 ();
 b15zdnd11an1n04x5 FILLER_143_1475 ();
 b15zdnd11an1n08x5 FILLER_143_1482 ();
 b15zdnd11an1n04x5 FILLER_143_1490 ();
 b15zdnd00an1n01x5 FILLER_143_1494 ();
 b15zdnd11an1n64x5 FILLER_143_1500 ();
 b15zdnd11an1n64x5 FILLER_143_1564 ();
 b15zdnd11an1n64x5 FILLER_143_1628 ();
 b15zdnd11an1n16x5 FILLER_143_1692 ();
 b15zdnd11an1n04x5 FILLER_143_1708 ();
 b15zdnd00an1n02x5 FILLER_143_1712 ();
 b15zdnd11an1n32x5 FILLER_143_1717 ();
 b15zdnd00an1n01x5 FILLER_143_1749 ();
 b15zdnd11an1n64x5 FILLER_143_1761 ();
 b15zdnd11an1n16x5 FILLER_143_1825 ();
 b15zdnd11an1n04x5 FILLER_143_1841 ();
 b15zdnd00an1n02x5 FILLER_143_1845 ();
 b15zdnd00an1n01x5 FILLER_143_1847 ();
 b15zdnd11an1n64x5 FILLER_143_1900 ();
 b15zdnd11an1n32x5 FILLER_143_1964 ();
 b15zdnd11an1n16x5 FILLER_143_1996 ();
 b15zdnd11an1n08x5 FILLER_143_2012 ();
 b15zdnd11an1n04x5 FILLER_143_2020 ();
 b15zdnd00an1n02x5 FILLER_143_2024 ();
 b15zdnd00an1n01x5 FILLER_143_2026 ();
 b15zdnd11an1n04x5 FILLER_143_2030 ();
 b15zdnd11an1n04x5 FILLER_143_2045 ();
 b15zdnd11an1n64x5 FILLER_143_2052 ();
 b15zdnd11an1n64x5 FILLER_143_2116 ();
 b15zdnd11an1n64x5 FILLER_143_2180 ();
 b15zdnd11an1n08x5 FILLER_143_2244 ();
 b15zdnd00an1n02x5 FILLER_143_2252 ();
 b15zdnd11an1n16x5 FILLER_143_2258 ();
 b15zdnd11an1n08x5 FILLER_143_2274 ();
 b15zdnd00an1n02x5 FILLER_143_2282 ();
 b15zdnd11an1n16x5 FILLER_144_8 ();
 b15zdnd00an1n02x5 FILLER_144_24 ();
 b15zdnd11an1n64x5 FILLER_144_46 ();
 b15zdnd11an1n64x5 FILLER_144_110 ();
 b15zdnd11an1n64x5 FILLER_144_174 ();
 b15zdnd11an1n64x5 FILLER_144_238 ();
 b15zdnd11an1n32x5 FILLER_144_302 ();
 b15zdnd11an1n04x5 FILLER_144_334 ();
 b15zdnd00an1n01x5 FILLER_144_338 ();
 b15zdnd11an1n64x5 FILLER_144_351 ();
 b15zdnd11an1n64x5 FILLER_144_415 ();
 b15zdnd11an1n64x5 FILLER_144_479 ();
 b15zdnd11an1n64x5 FILLER_144_543 ();
 b15zdnd11an1n64x5 FILLER_144_607 ();
 b15zdnd11an1n32x5 FILLER_144_671 ();
 b15zdnd11an1n08x5 FILLER_144_703 ();
 b15zdnd11an1n04x5 FILLER_144_711 ();
 b15zdnd00an1n02x5 FILLER_144_715 ();
 b15zdnd00an1n01x5 FILLER_144_717 ();
 b15zdnd11an1n64x5 FILLER_144_726 ();
 b15zdnd11an1n64x5 FILLER_144_790 ();
 b15zdnd11an1n64x5 FILLER_144_854 ();
 b15zdnd11an1n64x5 FILLER_144_918 ();
 b15zdnd11an1n64x5 FILLER_144_982 ();
 b15zdnd11an1n64x5 FILLER_144_1046 ();
 b15zdnd00an1n02x5 FILLER_144_1110 ();
 b15zdnd00an1n01x5 FILLER_144_1112 ();
 b15zdnd11an1n64x5 FILLER_144_1118 ();
 b15zdnd11an1n64x5 FILLER_144_1182 ();
 b15zdnd11an1n64x5 FILLER_144_1246 ();
 b15zdnd11an1n16x5 FILLER_144_1310 ();
 b15zdnd11an1n08x5 FILLER_144_1326 ();
 b15zdnd00an1n02x5 FILLER_144_1334 ();
 b15zdnd00an1n01x5 FILLER_144_1336 ();
 b15zdnd11an1n64x5 FILLER_144_1379 ();
 b15zdnd11an1n16x5 FILLER_144_1443 ();
 b15zdnd11an1n64x5 FILLER_144_1511 ();
 b15zdnd11an1n64x5 FILLER_144_1575 ();
 b15zdnd11an1n64x5 FILLER_144_1639 ();
 b15zdnd11an1n64x5 FILLER_144_1703 ();
 b15zdnd11an1n64x5 FILLER_144_1767 ();
 b15zdnd11an1n32x5 FILLER_144_1831 ();
 b15zdnd11an1n04x5 FILLER_144_1863 ();
 b15zdnd11an1n04x5 FILLER_144_1870 ();
 b15zdnd11an1n04x5 FILLER_144_1877 ();
 b15zdnd11an1n04x5 FILLER_144_1884 ();
 b15zdnd11an1n64x5 FILLER_144_1891 ();
 b15zdnd11an1n16x5 FILLER_144_1955 ();
 b15zdnd00an1n01x5 FILLER_144_1971 ();
 b15zdnd11an1n32x5 FILLER_144_1975 ();
 b15zdnd11an1n08x5 FILLER_144_2007 ();
 b15zdnd11an1n04x5 FILLER_144_2015 ();
 b15zdnd11an1n64x5 FILLER_144_2071 ();
 b15zdnd11an1n16x5 FILLER_144_2135 ();
 b15zdnd00an1n02x5 FILLER_144_2151 ();
 b15zdnd00an1n01x5 FILLER_144_2153 ();
 b15zdnd11an1n64x5 FILLER_144_2162 ();
 b15zdnd11an1n04x5 FILLER_144_2226 ();
 b15zdnd00an1n02x5 FILLER_144_2230 ();
 b15zdnd00an1n02x5 FILLER_144_2274 ();
 b15zdnd11an1n16x5 FILLER_145_0 ();
 b15zdnd11an1n04x5 FILLER_145_16 ();
 b15zdnd11an1n04x5 FILLER_145_23 ();
 b15zdnd11an1n64x5 FILLER_145_30 ();
 b15zdnd11an1n64x5 FILLER_145_94 ();
 b15zdnd11an1n64x5 FILLER_145_158 ();
 b15zdnd11an1n32x5 FILLER_145_222 ();
 b15zdnd00an1n01x5 FILLER_145_254 ();
 b15zdnd11an1n64x5 FILLER_145_297 ();
 b15zdnd11an1n64x5 FILLER_145_361 ();
 b15zdnd11an1n64x5 FILLER_145_425 ();
 b15zdnd11an1n64x5 FILLER_145_489 ();
 b15zdnd11an1n32x5 FILLER_145_553 ();
 b15zdnd11an1n16x5 FILLER_145_585 ();
 b15zdnd00an1n01x5 FILLER_145_601 ();
 b15zdnd11an1n64x5 FILLER_145_608 ();
 b15zdnd11an1n64x5 FILLER_145_672 ();
 b15zdnd11an1n64x5 FILLER_145_736 ();
 b15zdnd11an1n16x5 FILLER_145_800 ();
 b15zdnd11an1n04x5 FILLER_145_816 ();
 b15zdnd00an1n01x5 FILLER_145_820 ();
 b15zdnd11an1n64x5 FILLER_145_830 ();
 b15zdnd11an1n64x5 FILLER_145_894 ();
 b15zdnd11an1n64x5 FILLER_145_958 ();
 b15zdnd11an1n64x5 FILLER_145_1022 ();
 b15zdnd11an1n64x5 FILLER_145_1086 ();
 b15zdnd11an1n64x5 FILLER_145_1150 ();
 b15zdnd11an1n04x5 FILLER_145_1214 ();
 b15zdnd00an1n02x5 FILLER_145_1218 ();
 b15zdnd11an1n64x5 FILLER_145_1247 ();
 b15zdnd11an1n16x5 FILLER_145_1311 ();
 b15zdnd11an1n04x5 FILLER_145_1327 ();
 b15zdnd00an1n02x5 FILLER_145_1331 ();
 b15zdnd00an1n01x5 FILLER_145_1333 ();
 b15zdnd11an1n08x5 FILLER_145_1386 ();
 b15zdnd00an1n01x5 FILLER_145_1394 ();
 b15zdnd11an1n64x5 FILLER_145_1400 ();
 b15zdnd11an1n04x5 FILLER_145_1464 ();
 b15zdnd00an1n01x5 FILLER_145_1468 ();
 b15zdnd11an1n08x5 FILLER_145_1472 ();
 b15zdnd11an1n04x5 FILLER_145_1480 ();
 b15zdnd00an1n01x5 FILLER_145_1484 ();
 b15zdnd11an1n64x5 FILLER_145_1488 ();
 b15zdnd11an1n64x5 FILLER_145_1552 ();
 b15zdnd11an1n32x5 FILLER_145_1616 ();
 b15zdnd11an1n08x5 FILLER_145_1648 ();
 b15zdnd11an1n04x5 FILLER_145_1656 ();
 b15zdnd00an1n01x5 FILLER_145_1660 ();
 b15zdnd11an1n64x5 FILLER_145_1703 ();
 b15zdnd11an1n64x5 FILLER_145_1767 ();
 b15zdnd11an1n16x5 FILLER_145_1831 ();
 b15zdnd11an1n08x5 FILLER_145_1847 ();
 b15zdnd11an1n04x5 FILLER_145_1855 ();
 b15zdnd11an1n64x5 FILLER_145_1901 ();
 b15zdnd11an1n04x5 FILLER_145_1965 ();
 b15zdnd00an1n02x5 FILLER_145_1969 ();
 b15zdnd11an1n04x5 FILLER_145_1974 ();
 b15zdnd11an1n32x5 FILLER_145_1981 ();
 b15zdnd00an1n02x5 FILLER_145_2013 ();
 b15zdnd00an1n01x5 FILLER_145_2015 ();
 b15zdnd11an1n16x5 FILLER_145_2027 ();
 b15zdnd11an1n04x5 FILLER_145_2046 ();
 b15zdnd11an1n16x5 FILLER_145_2053 ();
 b15zdnd11an1n04x5 FILLER_145_2069 ();
 b15zdnd00an1n01x5 FILLER_145_2073 ();
 b15zdnd11an1n64x5 FILLER_145_2116 ();
 b15zdnd11an1n64x5 FILLER_145_2180 ();
 b15zdnd11an1n32x5 FILLER_145_2244 ();
 b15zdnd11an1n08x5 FILLER_145_2276 ();
 b15zdnd11an1n08x5 FILLER_146_8 ();
 b15zdnd11an1n04x5 FILLER_146_16 ();
 b15zdnd11an1n64x5 FILLER_146_23 ();
 b15zdnd11an1n64x5 FILLER_146_87 ();
 b15zdnd11an1n64x5 FILLER_146_151 ();
 b15zdnd11an1n32x5 FILLER_146_215 ();
 b15zdnd11an1n04x5 FILLER_146_247 ();
 b15zdnd00an1n01x5 FILLER_146_251 ();
 b15zdnd11an1n64x5 FILLER_146_294 ();
 b15zdnd11an1n16x5 FILLER_146_358 ();
 b15zdnd00an1n02x5 FILLER_146_374 ();
 b15zdnd00an1n01x5 FILLER_146_376 ();
 b15zdnd11an1n64x5 FILLER_146_383 ();
 b15zdnd11an1n64x5 FILLER_146_447 ();
 b15zdnd11an1n64x5 FILLER_146_511 ();
 b15zdnd11an1n64x5 FILLER_146_575 ();
 b15zdnd11an1n64x5 FILLER_146_639 ();
 b15zdnd11an1n08x5 FILLER_146_703 ();
 b15zdnd11an1n04x5 FILLER_146_711 ();
 b15zdnd00an1n02x5 FILLER_146_715 ();
 b15zdnd00an1n01x5 FILLER_146_717 ();
 b15zdnd11an1n64x5 FILLER_146_726 ();
 b15zdnd11an1n64x5 FILLER_146_790 ();
 b15zdnd11an1n64x5 FILLER_146_854 ();
 b15zdnd11an1n64x5 FILLER_146_918 ();
 b15zdnd11an1n64x5 FILLER_146_982 ();
 b15zdnd11an1n64x5 FILLER_146_1046 ();
 b15zdnd11an1n64x5 FILLER_146_1110 ();
 b15zdnd11an1n32x5 FILLER_146_1174 ();
 b15zdnd11an1n16x5 FILLER_146_1206 ();
 b15zdnd11an1n64x5 FILLER_146_1225 ();
 b15zdnd11an1n32x5 FILLER_146_1289 ();
 b15zdnd11an1n16x5 FILLER_146_1321 ();
 b15zdnd11an1n04x5 FILLER_146_1379 ();
 b15zdnd11an1n04x5 FILLER_146_1386 ();
 b15zdnd11an1n64x5 FILLER_146_1393 ();
 b15zdnd11an1n08x5 FILLER_146_1457 ();
 b15zdnd11an1n04x5 FILLER_146_1465 ();
 b15zdnd00an1n01x5 FILLER_146_1469 ();
 b15zdnd11an1n64x5 FILLER_146_1475 ();
 b15zdnd11an1n64x5 FILLER_146_1539 ();
 b15zdnd11an1n64x5 FILLER_146_1603 ();
 b15zdnd11an1n64x5 FILLER_146_1667 ();
 b15zdnd11an1n64x5 FILLER_146_1731 ();
 b15zdnd11an1n32x5 FILLER_146_1795 ();
 b15zdnd11an1n08x5 FILLER_146_1827 ();
 b15zdnd11an1n04x5 FILLER_146_1835 ();
 b15zdnd00an1n02x5 FILLER_146_1839 ();
 b15zdnd11an1n32x5 FILLER_146_1893 ();
 b15zdnd11an1n16x5 FILLER_146_1925 ();
 b15zdnd11an1n08x5 FILLER_146_1941 ();
 b15zdnd00an1n02x5 FILLER_146_1949 ();
 b15zdnd00an1n01x5 FILLER_146_1951 ();
 b15zdnd11an1n32x5 FILLER_146_2004 ();
 b15zdnd11an1n04x5 FILLER_146_2036 ();
 b15zdnd00an1n01x5 FILLER_146_2040 ();
 b15zdnd11an1n04x5 FILLER_146_2044 ();
 b15zdnd11an1n64x5 FILLER_146_2051 ();
 b15zdnd11an1n32x5 FILLER_146_2115 ();
 b15zdnd11an1n04x5 FILLER_146_2147 ();
 b15zdnd00an1n02x5 FILLER_146_2151 ();
 b15zdnd00an1n01x5 FILLER_146_2153 ();
 b15zdnd11an1n64x5 FILLER_146_2162 ();
 b15zdnd11an1n32x5 FILLER_146_2226 ();
 b15zdnd11an1n16x5 FILLER_146_2258 ();
 b15zdnd00an1n02x5 FILLER_146_2274 ();
 b15zdnd11an1n32x5 FILLER_147_0 ();
 b15zdnd00an1n01x5 FILLER_147_32 ();
 b15zdnd11an1n04x5 FILLER_147_37 ();
 b15zdnd00an1n01x5 FILLER_147_41 ();
 b15zdnd11an1n64x5 FILLER_147_45 ();
 b15zdnd11an1n64x5 FILLER_147_109 ();
 b15zdnd11an1n64x5 FILLER_147_173 ();
 b15zdnd11an1n16x5 FILLER_147_237 ();
 b15zdnd00an1n01x5 FILLER_147_253 ();
 b15zdnd11an1n64x5 FILLER_147_296 ();
 b15zdnd00an1n02x5 FILLER_147_360 ();
 b15zdnd00an1n01x5 FILLER_147_362 ();
 b15zdnd11an1n64x5 FILLER_147_405 ();
 b15zdnd11an1n08x5 FILLER_147_469 ();
 b15zdnd00an1n02x5 FILLER_147_477 ();
 b15zdnd11an1n64x5 FILLER_147_482 ();
 b15zdnd11an1n64x5 FILLER_147_546 ();
 b15zdnd11an1n64x5 FILLER_147_610 ();
 b15zdnd11an1n64x5 FILLER_147_674 ();
 b15zdnd11an1n64x5 FILLER_147_738 ();
 b15zdnd11an1n64x5 FILLER_147_802 ();
 b15zdnd11an1n64x5 FILLER_147_866 ();
 b15zdnd11an1n04x5 FILLER_147_930 ();
 b15zdnd00an1n01x5 FILLER_147_934 ();
 b15zdnd11an1n64x5 FILLER_147_951 ();
 b15zdnd11an1n64x5 FILLER_147_1015 ();
 b15zdnd11an1n64x5 FILLER_147_1079 ();
 b15zdnd11an1n64x5 FILLER_147_1143 ();
 b15zdnd11an1n64x5 FILLER_147_1207 ();
 b15zdnd11an1n64x5 FILLER_147_1271 ();
 b15zdnd11an1n16x5 FILLER_147_1335 ();
 b15zdnd00an1n02x5 FILLER_147_1351 ();
 b15zdnd00an1n01x5 FILLER_147_1353 ();
 b15zdnd11an1n08x5 FILLER_147_1357 ();
 b15zdnd00an1n02x5 FILLER_147_1365 ();
 b15zdnd00an1n01x5 FILLER_147_1367 ();
 b15zdnd11an1n04x5 FILLER_147_1373 ();
 b15zdnd00an1n01x5 FILLER_147_1377 ();
 b15zdnd11an1n64x5 FILLER_147_1430 ();
 b15zdnd11an1n64x5 FILLER_147_1494 ();
 b15zdnd11an1n64x5 FILLER_147_1558 ();
 b15zdnd11an1n64x5 FILLER_147_1622 ();
 b15zdnd11an1n64x5 FILLER_147_1686 ();
 b15zdnd11an1n64x5 FILLER_147_1750 ();
 b15zdnd11an1n32x5 FILLER_147_1814 ();
 b15zdnd11an1n08x5 FILLER_147_1846 ();
 b15zdnd11an1n04x5 FILLER_147_1854 ();
 b15zdnd00an1n01x5 FILLER_147_1858 ();
 b15zdnd11an1n04x5 FILLER_147_1862 ();
 b15zdnd11an1n64x5 FILLER_147_1869 ();
 b15zdnd11an1n32x5 FILLER_147_1933 ();
 b15zdnd11an1n08x5 FILLER_147_1965 ();
 b15zdnd11an1n04x5 FILLER_147_1973 ();
 b15zdnd00an1n01x5 FILLER_147_1977 ();
 b15zdnd11an1n16x5 FILLER_147_1998 ();
 b15zdnd11an1n04x5 FILLER_147_2014 ();
 b15zdnd11an1n64x5 FILLER_147_2070 ();
 b15zdnd11an1n64x5 FILLER_147_2134 ();
 b15zdnd11an1n64x5 FILLER_147_2198 ();
 b15zdnd11an1n16x5 FILLER_147_2262 ();
 b15zdnd11an1n04x5 FILLER_147_2278 ();
 b15zdnd00an1n02x5 FILLER_147_2282 ();
 b15zdnd11an1n08x5 FILLER_148_8 ();
 b15zdnd11an1n04x5 FILLER_148_16 ();
 b15zdnd00an1n02x5 FILLER_148_20 ();
 b15zdnd11an1n64x5 FILLER_148_25 ();
 b15zdnd11an1n64x5 FILLER_148_89 ();
 b15zdnd11an1n64x5 FILLER_148_153 ();
 b15zdnd11an1n32x5 FILLER_148_217 ();
 b15zdnd00an1n02x5 FILLER_148_249 ();
 b15zdnd11an1n64x5 FILLER_148_293 ();
 b15zdnd11an1n16x5 FILLER_148_357 ();
 b15zdnd00an1n02x5 FILLER_148_373 ();
 b15zdnd00an1n01x5 FILLER_148_375 ();
 b15zdnd11an1n32x5 FILLER_148_418 ();
 b15zdnd11an1n04x5 FILLER_148_450 ();
 b15zdnd00an1n02x5 FILLER_148_454 ();
 b15zdnd00an1n01x5 FILLER_148_456 ();
 b15zdnd11an1n04x5 FILLER_148_464 ();
 b15zdnd11an1n08x5 FILLER_148_488 ();
 b15zdnd11an1n04x5 FILLER_148_496 ();
 b15zdnd00an1n02x5 FILLER_148_500 ();
 b15zdnd00an1n01x5 FILLER_148_502 ();
 b15zdnd11an1n64x5 FILLER_148_508 ();
 b15zdnd11an1n64x5 FILLER_148_572 ();
 b15zdnd11an1n64x5 FILLER_148_636 ();
 b15zdnd11an1n16x5 FILLER_148_700 ();
 b15zdnd00an1n02x5 FILLER_148_716 ();
 b15zdnd11an1n64x5 FILLER_148_726 ();
 b15zdnd11an1n08x5 FILLER_148_790 ();
 b15zdnd11an1n04x5 FILLER_148_798 ();
 b15zdnd00an1n02x5 FILLER_148_802 ();
 b15zdnd11an1n64x5 FILLER_148_807 ();
 b15zdnd11an1n16x5 FILLER_148_871 ();
 b15zdnd11an1n08x5 FILLER_148_887 ();
 b15zdnd11an1n04x5 FILLER_148_895 ();
 b15zdnd00an1n01x5 FILLER_148_899 ();
 b15zdnd11an1n32x5 FILLER_148_915 ();
 b15zdnd00an1n01x5 FILLER_148_947 ();
 b15zdnd11an1n16x5 FILLER_148_952 ();
 b15zdnd11an1n04x5 FILLER_148_968 ();
 b15zdnd00an1n02x5 FILLER_148_972 ();
 b15zdnd11an1n64x5 FILLER_148_996 ();
 b15zdnd11an1n64x5 FILLER_148_1060 ();
 b15zdnd11an1n64x5 FILLER_148_1124 ();
 b15zdnd11an1n64x5 FILLER_148_1188 ();
 b15zdnd11an1n64x5 FILLER_148_1252 ();
 b15zdnd11an1n64x5 FILLER_148_1316 ();
 b15zdnd11an1n16x5 FILLER_148_1380 ();
 b15zdnd11an1n04x5 FILLER_148_1396 ();
 b15zdnd11an1n32x5 FILLER_148_1405 ();
 b15zdnd11an1n08x5 FILLER_148_1437 ();
 b15zdnd00an1n02x5 FILLER_148_1445 ();
 b15zdnd11an1n64x5 FILLER_148_1452 ();
 b15zdnd11an1n64x5 FILLER_148_1516 ();
 b15zdnd11an1n64x5 FILLER_148_1580 ();
 b15zdnd11an1n64x5 FILLER_148_1644 ();
 b15zdnd11an1n64x5 FILLER_148_1708 ();
 b15zdnd11an1n64x5 FILLER_148_1772 ();
 b15zdnd11an1n64x5 FILLER_148_1836 ();
 b15zdnd11an1n64x5 FILLER_148_1900 ();
 b15zdnd11an1n64x5 FILLER_148_1964 ();
 b15zdnd11an1n08x5 FILLER_148_2028 ();
 b15zdnd11an1n04x5 FILLER_148_2036 ();
 b15zdnd00an1n01x5 FILLER_148_2040 ();
 b15zdnd11an1n04x5 FILLER_148_2044 ();
 b15zdnd11an1n64x5 FILLER_148_2059 ();
 b15zdnd11an1n16x5 FILLER_148_2123 ();
 b15zdnd11an1n08x5 FILLER_148_2139 ();
 b15zdnd11an1n04x5 FILLER_148_2147 ();
 b15zdnd00an1n02x5 FILLER_148_2151 ();
 b15zdnd00an1n01x5 FILLER_148_2153 ();
 b15zdnd11an1n64x5 FILLER_148_2162 ();
 b15zdnd11an1n32x5 FILLER_148_2226 ();
 b15zdnd11an1n16x5 FILLER_148_2258 ();
 b15zdnd00an1n02x5 FILLER_148_2274 ();
 b15zdnd11an1n64x5 FILLER_149_0 ();
 b15zdnd11an1n64x5 FILLER_149_64 ();
 b15zdnd11an1n64x5 FILLER_149_128 ();
 b15zdnd11an1n64x5 FILLER_149_192 ();
 b15zdnd11an1n64x5 FILLER_149_256 ();
 b15zdnd11an1n32x5 FILLER_149_320 ();
 b15zdnd11an1n16x5 FILLER_149_352 ();
 b15zdnd11an1n04x5 FILLER_149_368 ();
 b15zdnd11an1n04x5 FILLER_149_386 ();
 b15zdnd11an1n16x5 FILLER_149_432 ();
 b15zdnd11an1n04x5 FILLER_149_448 ();
 b15zdnd00an1n02x5 FILLER_149_452 ();
 b15zdnd11an1n04x5 FILLER_149_461 ();
 b15zdnd11an1n64x5 FILLER_149_507 ();
 b15zdnd11an1n64x5 FILLER_149_571 ();
 b15zdnd11an1n64x5 FILLER_149_635 ();
 b15zdnd11an1n64x5 FILLER_149_699 ();
 b15zdnd11an1n64x5 FILLER_149_763 ();
 b15zdnd11an1n64x5 FILLER_149_827 ();
 b15zdnd11an1n64x5 FILLER_149_891 ();
 b15zdnd00an1n02x5 FILLER_149_955 ();
 b15zdnd00an1n01x5 FILLER_149_957 ();
 b15zdnd11an1n04x5 FILLER_149_986 ();
 b15zdnd11an1n04x5 FILLER_149_1021 ();
 b15zdnd11an1n64x5 FILLER_149_1034 ();
 b15zdnd11an1n64x5 FILLER_149_1098 ();
 b15zdnd11an1n64x5 FILLER_149_1162 ();
 b15zdnd11an1n64x5 FILLER_149_1226 ();
 b15zdnd11an1n64x5 FILLER_149_1290 ();
 b15zdnd11an1n32x5 FILLER_149_1354 ();
 b15zdnd11an1n04x5 FILLER_149_1386 ();
 b15zdnd11an1n64x5 FILLER_149_1393 ();
 b15zdnd11an1n64x5 FILLER_149_1457 ();
 b15zdnd11an1n64x5 FILLER_149_1521 ();
 b15zdnd11an1n64x5 FILLER_149_1585 ();
 b15zdnd11an1n64x5 FILLER_149_1649 ();
 b15zdnd11an1n64x5 FILLER_149_1713 ();
 b15zdnd11an1n64x5 FILLER_149_1777 ();
 b15zdnd11an1n64x5 FILLER_149_1841 ();
 b15zdnd11an1n64x5 FILLER_149_1905 ();
 b15zdnd11an1n64x5 FILLER_149_1969 ();
 b15zdnd11an1n64x5 FILLER_149_2033 ();
 b15zdnd11an1n64x5 FILLER_149_2097 ();
 b15zdnd11an1n64x5 FILLER_149_2161 ();
 b15zdnd11an1n32x5 FILLER_149_2225 ();
 b15zdnd11an1n16x5 FILLER_149_2257 ();
 b15zdnd11an1n08x5 FILLER_149_2273 ();
 b15zdnd00an1n02x5 FILLER_149_2281 ();
 b15zdnd00an1n01x5 FILLER_149_2283 ();
 b15zdnd11an1n08x5 FILLER_150_8 ();
 b15zdnd11an1n04x5 FILLER_150_16 ();
 b15zdnd00an1n01x5 FILLER_150_20 ();
 b15zdnd11an1n04x5 FILLER_150_24 ();
 b15zdnd00an1n02x5 FILLER_150_28 ();
 b15zdnd00an1n01x5 FILLER_150_30 ();
 b15zdnd11an1n04x5 FILLER_150_34 ();
 b15zdnd11an1n64x5 FILLER_150_41 ();
 b15zdnd11an1n64x5 FILLER_150_105 ();
 b15zdnd11an1n32x5 FILLER_150_169 ();
 b15zdnd11an1n16x5 FILLER_150_201 ();
 b15zdnd11an1n08x5 FILLER_150_217 ();
 b15zdnd11an1n64x5 FILLER_150_267 ();
 b15zdnd11an1n08x5 FILLER_150_331 ();
 b15zdnd00an1n02x5 FILLER_150_339 ();
 b15zdnd00an1n01x5 FILLER_150_341 ();
 b15zdnd11an1n16x5 FILLER_150_348 ();
 b15zdnd00an1n02x5 FILLER_150_364 ();
 b15zdnd00an1n01x5 FILLER_150_366 ();
 b15zdnd11an1n64x5 FILLER_150_373 ();
 b15zdnd11an1n08x5 FILLER_150_437 ();
 b15zdnd11an1n04x5 FILLER_150_445 ();
 b15zdnd00an1n02x5 FILLER_150_449 ();
 b15zdnd00an1n01x5 FILLER_150_451 ();
 b15zdnd11an1n64x5 FILLER_150_504 ();
 b15zdnd11an1n32x5 FILLER_150_568 ();
 b15zdnd11an1n16x5 FILLER_150_600 ();
 b15zdnd11an1n08x5 FILLER_150_616 ();
 b15zdnd00an1n02x5 FILLER_150_624 ();
 b15zdnd11an1n32x5 FILLER_150_629 ();
 b15zdnd11an1n16x5 FILLER_150_661 ();
 b15zdnd11an1n08x5 FILLER_150_705 ();
 b15zdnd11an1n04x5 FILLER_150_713 ();
 b15zdnd00an1n01x5 FILLER_150_717 ();
 b15zdnd11an1n64x5 FILLER_150_726 ();
 b15zdnd11an1n64x5 FILLER_150_790 ();
 b15zdnd11an1n64x5 FILLER_150_854 ();
 b15zdnd11an1n32x5 FILLER_150_918 ();
 b15zdnd11an1n08x5 FILLER_150_950 ();
 b15zdnd11an1n04x5 FILLER_150_958 ();
 b15zdnd00an1n01x5 FILLER_150_962 ();
 b15zdnd11an1n64x5 FILLER_150_1008 ();
 b15zdnd11an1n64x5 FILLER_150_1072 ();
 b15zdnd11an1n64x5 FILLER_150_1136 ();
 b15zdnd11an1n64x5 FILLER_150_1200 ();
 b15zdnd11an1n64x5 FILLER_150_1264 ();
 b15zdnd11an1n64x5 FILLER_150_1328 ();
 b15zdnd11an1n64x5 FILLER_150_1392 ();
 b15zdnd11an1n64x5 FILLER_150_1456 ();
 b15zdnd11an1n64x5 FILLER_150_1520 ();
 b15zdnd11an1n16x5 FILLER_150_1584 ();
 b15zdnd11an1n08x5 FILLER_150_1600 ();
 b15zdnd11an1n64x5 FILLER_150_1650 ();
 b15zdnd11an1n64x5 FILLER_150_1714 ();
 b15zdnd11an1n64x5 FILLER_150_1778 ();
 b15zdnd11an1n64x5 FILLER_150_1842 ();
 b15zdnd11an1n64x5 FILLER_150_1906 ();
 b15zdnd11an1n64x5 FILLER_150_1970 ();
 b15zdnd11an1n64x5 FILLER_150_2034 ();
 b15zdnd11an1n32x5 FILLER_150_2098 ();
 b15zdnd11an1n16x5 FILLER_150_2130 ();
 b15zdnd11an1n08x5 FILLER_150_2146 ();
 b15zdnd11an1n64x5 FILLER_150_2162 ();
 b15zdnd11an1n32x5 FILLER_150_2226 ();
 b15zdnd11an1n16x5 FILLER_150_2258 ();
 b15zdnd00an1n02x5 FILLER_150_2274 ();
 b15zdnd11an1n16x5 FILLER_151_0 ();
 b15zdnd11an1n08x5 FILLER_151_16 ();
 b15zdnd11an1n04x5 FILLER_151_24 ();
 b15zdnd00an1n02x5 FILLER_151_28 ();
 b15zdnd00an1n01x5 FILLER_151_30 ();
 b15zdnd11an1n64x5 FILLER_151_34 ();
 b15zdnd11an1n64x5 FILLER_151_98 ();
 b15zdnd11an1n64x5 FILLER_151_162 ();
 b15zdnd11an1n32x5 FILLER_151_226 ();
 b15zdnd11an1n08x5 FILLER_151_258 ();
 b15zdnd00an1n02x5 FILLER_151_266 ();
 b15zdnd00an1n01x5 FILLER_151_268 ();
 b15zdnd11an1n08x5 FILLER_151_272 ();
 b15zdnd00an1n02x5 FILLER_151_280 ();
 b15zdnd00an1n01x5 FILLER_151_282 ();
 b15zdnd11an1n64x5 FILLER_151_286 ();
 b15zdnd11an1n08x5 FILLER_151_350 ();
 b15zdnd11an1n04x5 FILLER_151_358 ();
 b15zdnd00an1n02x5 FILLER_151_362 ();
 b15zdnd00an1n01x5 FILLER_151_364 ();
 b15zdnd11an1n04x5 FILLER_151_368 ();
 b15zdnd11an1n32x5 FILLER_151_414 ();
 b15zdnd11an1n16x5 FILLER_151_446 ();
 b15zdnd11an1n08x5 FILLER_151_462 ();
 b15zdnd00an1n01x5 FILLER_151_470 ();
 b15zdnd11an1n04x5 FILLER_151_474 ();
 b15zdnd11an1n64x5 FILLER_151_481 ();
 b15zdnd11an1n16x5 FILLER_151_545 ();
 b15zdnd11an1n08x5 FILLER_151_561 ();
 b15zdnd11an1n04x5 FILLER_151_569 ();
 b15zdnd11an1n16x5 FILLER_151_576 ();
 b15zdnd11an1n04x5 FILLER_151_592 ();
 b15zdnd00an1n02x5 FILLER_151_596 ();
 b15zdnd00an1n01x5 FILLER_151_598 ();
 b15zdnd11an1n32x5 FILLER_151_651 ();
 b15zdnd11an1n08x5 FILLER_151_683 ();
 b15zdnd11an1n04x5 FILLER_151_691 ();
 b15zdnd11an1n04x5 FILLER_151_698 ();
 b15zdnd00an1n01x5 FILLER_151_702 ();
 b15zdnd11an1n64x5 FILLER_151_706 ();
 b15zdnd11an1n64x5 FILLER_151_770 ();
 b15zdnd11an1n64x5 FILLER_151_834 ();
 b15zdnd11an1n32x5 FILLER_151_898 ();
 b15zdnd11an1n16x5 FILLER_151_930 ();
 b15zdnd00an1n02x5 FILLER_151_946 ();
 b15zdnd11an1n32x5 FILLER_151_963 ();
 b15zdnd00an1n01x5 FILLER_151_995 ();
 b15zdnd11an1n16x5 FILLER_151_1010 ();
 b15zdnd00an1n02x5 FILLER_151_1026 ();
 b15zdnd00an1n01x5 FILLER_151_1028 ();
 b15zdnd11an1n64x5 FILLER_151_1040 ();
 b15zdnd11an1n64x5 FILLER_151_1104 ();
 b15zdnd11an1n64x5 FILLER_151_1168 ();
 b15zdnd11an1n64x5 FILLER_151_1232 ();
 b15zdnd11an1n64x5 FILLER_151_1296 ();
 b15zdnd11an1n64x5 FILLER_151_1360 ();
 b15zdnd11an1n64x5 FILLER_151_1424 ();
 b15zdnd11an1n64x5 FILLER_151_1488 ();
 b15zdnd11an1n64x5 FILLER_151_1552 ();
 b15zdnd11an1n64x5 FILLER_151_1616 ();
 b15zdnd11an1n64x5 FILLER_151_1680 ();
 b15zdnd11an1n64x5 FILLER_151_1744 ();
 b15zdnd11an1n64x5 FILLER_151_1808 ();
 b15zdnd11an1n64x5 FILLER_151_1872 ();
 b15zdnd11an1n64x5 FILLER_151_1936 ();
 b15zdnd11an1n64x5 FILLER_151_2000 ();
 b15zdnd11an1n64x5 FILLER_151_2064 ();
 b15zdnd11an1n64x5 FILLER_151_2128 ();
 b15zdnd11an1n64x5 FILLER_151_2192 ();
 b15zdnd11an1n16x5 FILLER_151_2256 ();
 b15zdnd11an1n08x5 FILLER_151_2272 ();
 b15zdnd11an1n04x5 FILLER_151_2280 ();
 b15zdnd11an1n16x5 FILLER_152_8 ();
 b15zdnd11an1n04x5 FILLER_152_24 ();
 b15zdnd00an1n02x5 FILLER_152_28 ();
 b15zdnd11an1n64x5 FILLER_152_33 ();
 b15zdnd11an1n64x5 FILLER_152_97 ();
 b15zdnd11an1n64x5 FILLER_152_161 ();
 b15zdnd00an1n02x5 FILLER_152_225 ();
 b15zdnd00an1n01x5 FILLER_152_227 ();
 b15zdnd11an1n32x5 FILLER_152_280 ();
 b15zdnd11an1n16x5 FILLER_152_312 ();
 b15zdnd11an1n04x5 FILLER_152_328 ();
 b15zdnd00an1n01x5 FILLER_152_332 ();
 b15zdnd11an1n04x5 FILLER_152_339 ();
 b15zdnd11an1n64x5 FILLER_152_395 ();
 b15zdnd11an1n64x5 FILLER_152_459 ();
 b15zdnd11an1n16x5 FILLER_152_523 ();
 b15zdnd11an1n04x5 FILLER_152_539 ();
 b15zdnd00an1n02x5 FILLER_152_543 ();
 b15zdnd00an1n01x5 FILLER_152_545 ();
 b15zdnd11an1n16x5 FILLER_152_598 ();
 b15zdnd11an1n04x5 FILLER_152_614 ();
 b15zdnd11an1n04x5 FILLER_152_621 ();
 b15zdnd11an1n64x5 FILLER_152_628 ();
 b15zdnd11an1n16x5 FILLER_152_692 ();
 b15zdnd11an1n08x5 FILLER_152_708 ();
 b15zdnd00an1n02x5 FILLER_152_716 ();
 b15zdnd11an1n32x5 FILLER_152_726 ();
 b15zdnd00an1n02x5 FILLER_152_758 ();
 b15zdnd11an1n64x5 FILLER_152_764 ();
 b15zdnd00an1n01x5 FILLER_152_828 ();
 b15zdnd11an1n04x5 FILLER_152_838 ();
 b15zdnd00an1n02x5 FILLER_152_842 ();
 b15zdnd00an1n01x5 FILLER_152_844 ();
 b15zdnd11an1n04x5 FILLER_152_879 ();
 b15zdnd11an1n04x5 FILLER_152_916 ();
 b15zdnd11an1n64x5 FILLER_152_934 ();
 b15zdnd11an1n64x5 FILLER_152_998 ();
 b15zdnd11an1n64x5 FILLER_152_1062 ();
 b15zdnd11an1n64x5 FILLER_152_1126 ();
 b15zdnd11an1n64x5 FILLER_152_1190 ();
 b15zdnd11an1n64x5 FILLER_152_1254 ();
 b15zdnd11an1n64x5 FILLER_152_1318 ();
 b15zdnd11an1n64x5 FILLER_152_1382 ();
 b15zdnd11an1n64x5 FILLER_152_1446 ();
 b15zdnd11an1n64x5 FILLER_152_1510 ();
 b15zdnd11an1n64x5 FILLER_152_1574 ();
 b15zdnd11an1n64x5 FILLER_152_1638 ();
 b15zdnd11an1n64x5 FILLER_152_1702 ();
 b15zdnd11an1n32x5 FILLER_152_1766 ();
 b15zdnd11an1n16x5 FILLER_152_1798 ();
 b15zdnd11an1n08x5 FILLER_152_1814 ();
 b15zdnd11an1n04x5 FILLER_152_1822 ();
 b15zdnd00an1n02x5 FILLER_152_1826 ();
 b15zdnd00an1n01x5 FILLER_152_1828 ();
 b15zdnd11an1n64x5 FILLER_152_1871 ();
 b15zdnd11an1n64x5 FILLER_152_1935 ();
 b15zdnd11an1n64x5 FILLER_152_1999 ();
 b15zdnd11an1n64x5 FILLER_152_2063 ();
 b15zdnd11an1n16x5 FILLER_152_2127 ();
 b15zdnd11an1n08x5 FILLER_152_2143 ();
 b15zdnd00an1n02x5 FILLER_152_2151 ();
 b15zdnd00an1n01x5 FILLER_152_2153 ();
 b15zdnd11an1n64x5 FILLER_152_2162 ();
 b15zdnd11an1n32x5 FILLER_152_2226 ();
 b15zdnd11an1n16x5 FILLER_152_2258 ();
 b15zdnd00an1n02x5 FILLER_152_2274 ();
 b15zdnd11an1n64x5 FILLER_153_0 ();
 b15zdnd11an1n64x5 FILLER_153_64 ();
 b15zdnd11an1n64x5 FILLER_153_128 ();
 b15zdnd11an1n32x5 FILLER_153_192 ();
 b15zdnd11an1n08x5 FILLER_153_224 ();
 b15zdnd11an1n32x5 FILLER_153_284 ();
 b15zdnd11an1n16x5 FILLER_153_316 ();
 b15zdnd11an1n04x5 FILLER_153_332 ();
 b15zdnd00an1n01x5 FILLER_153_336 ();
 b15zdnd11an1n08x5 FILLER_153_351 ();
 b15zdnd00an1n02x5 FILLER_153_359 ();
 b15zdnd00an1n01x5 FILLER_153_361 ();
 b15zdnd11an1n04x5 FILLER_153_365 ();
 b15zdnd11an1n32x5 FILLER_153_372 ();
 b15zdnd00an1n02x5 FILLER_153_404 ();
 b15zdnd00an1n01x5 FILLER_153_406 ();
 b15zdnd11an1n64x5 FILLER_153_421 ();
 b15zdnd11an1n64x5 FILLER_153_485 ();
 b15zdnd11an1n08x5 FILLER_153_549 ();
 b15zdnd11an1n04x5 FILLER_153_557 ();
 b15zdnd00an1n02x5 FILLER_153_561 ();
 b15zdnd00an1n01x5 FILLER_153_563 ();
 b15zdnd11an1n04x5 FILLER_153_567 ();
 b15zdnd11an1n08x5 FILLER_153_574 ();
 b15zdnd00an1n02x5 FILLER_153_582 ();
 b15zdnd11an1n64x5 FILLER_153_626 ();
 b15zdnd11an1n64x5 FILLER_153_690 ();
 b15zdnd11an1n04x5 FILLER_153_754 ();
 b15zdnd00an1n02x5 FILLER_153_758 ();
 b15zdnd00an1n01x5 FILLER_153_760 ();
 b15zdnd11an1n32x5 FILLER_153_788 ();
 b15zdnd00an1n01x5 FILLER_153_820 ();
 b15zdnd11an1n64x5 FILLER_153_832 ();
 b15zdnd11an1n64x5 FILLER_153_896 ();
 b15zdnd11an1n64x5 FILLER_153_960 ();
 b15zdnd11an1n16x5 FILLER_153_1024 ();
 b15zdnd11an1n04x5 FILLER_153_1040 ();
 b15zdnd00an1n02x5 FILLER_153_1044 ();
 b15zdnd11an1n04x5 FILLER_153_1049 ();
 b15zdnd11an1n64x5 FILLER_153_1056 ();
 b15zdnd11an1n64x5 FILLER_153_1120 ();
 b15zdnd11an1n64x5 FILLER_153_1184 ();
 b15zdnd11an1n64x5 FILLER_153_1248 ();
 b15zdnd11an1n64x5 FILLER_153_1312 ();
 b15zdnd11an1n64x5 FILLER_153_1376 ();
 b15zdnd11an1n64x5 FILLER_153_1440 ();
 b15zdnd11an1n16x5 FILLER_153_1504 ();
 b15zdnd11an1n08x5 FILLER_153_1520 ();
 b15zdnd11an1n04x5 FILLER_153_1528 ();
 b15zdnd00an1n02x5 FILLER_153_1532 ();
 b15zdnd00an1n01x5 FILLER_153_1534 ();
 b15zdnd11an1n04x5 FILLER_153_1538 ();
 b15zdnd11an1n64x5 FILLER_153_1545 ();
 b15zdnd11an1n64x5 FILLER_153_1609 ();
 b15zdnd11an1n64x5 FILLER_153_1673 ();
 b15zdnd11an1n64x5 FILLER_153_1737 ();
 b15zdnd00an1n02x5 FILLER_153_1801 ();
 b15zdnd00an1n01x5 FILLER_153_1803 ();
 b15zdnd11an1n64x5 FILLER_153_1846 ();
 b15zdnd11an1n64x5 FILLER_153_1910 ();
 b15zdnd11an1n64x5 FILLER_153_1974 ();
 b15zdnd11an1n64x5 FILLER_153_2038 ();
 b15zdnd11an1n64x5 FILLER_153_2102 ();
 b15zdnd11an1n16x5 FILLER_153_2166 ();
 b15zdnd00an1n02x5 FILLER_153_2182 ();
 b15zdnd00an1n01x5 FILLER_153_2184 ();
 b15zdnd11an1n64x5 FILLER_153_2216 ();
 b15zdnd11an1n04x5 FILLER_153_2280 ();
 b15zdnd11an1n08x5 FILLER_154_8 ();
 b15zdnd11an1n04x5 FILLER_154_16 ();
 b15zdnd00an1n02x5 FILLER_154_20 ();
 b15zdnd00an1n01x5 FILLER_154_22 ();
 b15zdnd11an1n64x5 FILLER_154_31 ();
 b15zdnd11an1n32x5 FILLER_154_95 ();
 b15zdnd11an1n64x5 FILLER_154_130 ();
 b15zdnd11an1n32x5 FILLER_154_194 ();
 b15zdnd11an1n16x5 FILLER_154_226 ();
 b15zdnd11an1n08x5 FILLER_154_242 ();
 b15zdnd11an1n04x5 FILLER_154_250 ();
 b15zdnd00an1n01x5 FILLER_154_254 ();
 b15zdnd11an1n04x5 FILLER_154_258 ();
 b15zdnd11an1n16x5 FILLER_154_265 ();
 b15zdnd11an1n64x5 FILLER_154_284 ();
 b15zdnd11an1n64x5 FILLER_154_348 ();
 b15zdnd11an1n64x5 FILLER_154_412 ();
 b15zdnd11an1n04x5 FILLER_154_476 ();
 b15zdnd00an1n01x5 FILLER_154_480 ();
 b15zdnd11an1n64x5 FILLER_154_499 ();
 b15zdnd11an1n64x5 FILLER_154_563 ();
 b15zdnd11an1n64x5 FILLER_154_627 ();
 b15zdnd11an1n16x5 FILLER_154_691 ();
 b15zdnd11an1n08x5 FILLER_154_707 ();
 b15zdnd00an1n02x5 FILLER_154_715 ();
 b15zdnd00an1n01x5 FILLER_154_717 ();
 b15zdnd11an1n32x5 FILLER_154_726 ();
 b15zdnd00an1n02x5 FILLER_154_758 ();
 b15zdnd11an1n32x5 FILLER_154_763 ();
 b15zdnd11an1n08x5 FILLER_154_795 ();
 b15zdnd11an1n04x5 FILLER_154_820 ();
 b15zdnd11an1n08x5 FILLER_154_833 ();
 b15zdnd11an1n16x5 FILLER_154_855 ();
 b15zdnd11an1n08x5 FILLER_154_871 ();
 b15zdnd11an1n04x5 FILLER_154_879 ();
 b15zdnd00an1n02x5 FILLER_154_883 ();
 b15zdnd11an1n64x5 FILLER_154_899 ();
 b15zdnd11an1n32x5 FILLER_154_963 ();
 b15zdnd11an1n16x5 FILLER_154_995 ();
 b15zdnd11an1n08x5 FILLER_154_1011 ();
 b15zdnd00an1n02x5 FILLER_154_1019 ();
 b15zdnd11an1n32x5 FILLER_154_1073 ();
 b15zdnd11an1n16x5 FILLER_154_1105 ();
 b15zdnd11an1n08x5 FILLER_154_1121 ();
 b15zdnd11an1n04x5 FILLER_154_1129 ();
 b15zdnd11an1n64x5 FILLER_154_1136 ();
 b15zdnd11an1n64x5 FILLER_154_1200 ();
 b15zdnd11an1n64x5 FILLER_154_1264 ();
 b15zdnd11an1n64x5 FILLER_154_1328 ();
 b15zdnd11an1n64x5 FILLER_154_1392 ();
 b15zdnd11an1n32x5 FILLER_154_1456 ();
 b15zdnd11an1n16x5 FILLER_154_1488 ();
 b15zdnd11an1n08x5 FILLER_154_1504 ();
 b15zdnd11an1n64x5 FILLER_154_1564 ();
 b15zdnd11an1n32x5 FILLER_154_1628 ();
 b15zdnd00an1n01x5 FILLER_154_1660 ();
 b15zdnd11an1n04x5 FILLER_154_1664 ();
 b15zdnd11an1n64x5 FILLER_154_1671 ();
 b15zdnd11an1n64x5 FILLER_154_1735 ();
 b15zdnd11an1n64x5 FILLER_154_1799 ();
 b15zdnd11an1n64x5 FILLER_154_1863 ();
 b15zdnd11an1n64x5 FILLER_154_1927 ();
 b15zdnd11an1n64x5 FILLER_154_1991 ();
 b15zdnd11an1n64x5 FILLER_154_2055 ();
 b15zdnd11an1n32x5 FILLER_154_2119 ();
 b15zdnd00an1n02x5 FILLER_154_2151 ();
 b15zdnd00an1n01x5 FILLER_154_2153 ();
 b15zdnd11an1n64x5 FILLER_154_2162 ();
 b15zdnd11an1n32x5 FILLER_154_2226 ();
 b15zdnd11an1n16x5 FILLER_154_2258 ();
 b15zdnd00an1n02x5 FILLER_154_2274 ();
 b15zdnd11an1n64x5 FILLER_155_0 ();
 b15zdnd11an1n32x5 FILLER_155_64 ();
 b15zdnd11an1n04x5 FILLER_155_96 ();
 b15zdnd00an1n02x5 FILLER_155_100 ();
 b15zdnd11an1n64x5 FILLER_155_122 ();
 b15zdnd11an1n64x5 FILLER_155_186 ();
 b15zdnd11an1n04x5 FILLER_155_250 ();
 b15zdnd11an1n64x5 FILLER_155_257 ();
 b15zdnd11an1n64x5 FILLER_155_321 ();
 b15zdnd11an1n64x5 FILLER_155_385 ();
 b15zdnd11an1n32x5 FILLER_155_449 ();
 b15zdnd00an1n02x5 FILLER_155_481 ();
 b15zdnd11an1n64x5 FILLER_155_490 ();
 b15zdnd11an1n64x5 FILLER_155_554 ();
 b15zdnd11an1n64x5 FILLER_155_618 ();
 b15zdnd11an1n64x5 FILLER_155_682 ();
 b15zdnd11an1n64x5 FILLER_155_746 ();
 b15zdnd11an1n16x5 FILLER_155_810 ();
 b15zdnd11an1n08x5 FILLER_155_826 ();
 b15zdnd11an1n04x5 FILLER_155_834 ();
 b15zdnd11an1n64x5 FILLER_155_852 ();
 b15zdnd11an1n64x5 FILLER_155_916 ();
 b15zdnd11an1n64x5 FILLER_155_980 ();
 b15zdnd11an1n32x5 FILLER_155_1047 ();
 b15zdnd11an1n16x5 FILLER_155_1079 ();
 b15zdnd11an1n08x5 FILLER_155_1095 ();
 b15zdnd00an1n02x5 FILLER_155_1103 ();
 b15zdnd00an1n01x5 FILLER_155_1105 ();
 b15zdnd11an1n64x5 FILLER_155_1158 ();
 b15zdnd11an1n64x5 FILLER_155_1222 ();
 b15zdnd11an1n64x5 FILLER_155_1286 ();
 b15zdnd11an1n64x5 FILLER_155_1350 ();
 b15zdnd11an1n64x5 FILLER_155_1414 ();
 b15zdnd11an1n64x5 FILLER_155_1478 ();
 b15zdnd00an1n01x5 FILLER_155_1542 ();
 b15zdnd11an1n64x5 FILLER_155_1546 ();
 b15zdnd11an1n32x5 FILLER_155_1610 ();
 b15zdnd00an1n01x5 FILLER_155_1642 ();
 b15zdnd11an1n64x5 FILLER_155_1695 ();
 b15zdnd11an1n64x5 FILLER_155_1759 ();
 b15zdnd11an1n64x5 FILLER_155_1823 ();
 b15zdnd11an1n64x5 FILLER_155_1887 ();
 b15zdnd11an1n64x5 FILLER_155_1951 ();
 b15zdnd11an1n64x5 FILLER_155_2015 ();
 b15zdnd11an1n64x5 FILLER_155_2079 ();
 b15zdnd11an1n64x5 FILLER_155_2143 ();
 b15zdnd11an1n64x5 FILLER_155_2207 ();
 b15zdnd11an1n08x5 FILLER_155_2271 ();
 b15zdnd11an1n04x5 FILLER_155_2279 ();
 b15zdnd00an1n01x5 FILLER_155_2283 ();
 b15zdnd11an1n32x5 FILLER_156_8 ();
 b15zdnd11an1n16x5 FILLER_156_40 ();
 b15zdnd11an1n04x5 FILLER_156_56 ();
 b15zdnd00an1n02x5 FILLER_156_60 ();
 b15zdnd11an1n16x5 FILLER_156_68 ();
 b15zdnd00an1n01x5 FILLER_156_84 ();
 b15zdnd11an1n04x5 FILLER_156_91 ();
 b15zdnd00an1n02x5 FILLER_156_95 ();
 b15zdnd00an1n01x5 FILLER_156_97 ();
 b15zdnd11an1n04x5 FILLER_156_120 ();
 b15zdnd11an1n64x5 FILLER_156_130 ();
 b15zdnd11an1n64x5 FILLER_156_194 ();
 b15zdnd11an1n64x5 FILLER_156_258 ();
 b15zdnd11an1n64x5 FILLER_156_322 ();
 b15zdnd11an1n64x5 FILLER_156_386 ();
 b15zdnd11an1n16x5 FILLER_156_450 ();
 b15zdnd11an1n08x5 FILLER_156_466 ();
 b15zdnd11an1n04x5 FILLER_156_474 ();
 b15zdnd11an1n16x5 FILLER_156_485 ();
 b15zdnd11an1n04x5 FILLER_156_528 ();
 b15zdnd11an1n64x5 FILLER_156_544 ();
 b15zdnd11an1n64x5 FILLER_156_608 ();
 b15zdnd11an1n32x5 FILLER_156_672 ();
 b15zdnd11an1n08x5 FILLER_156_704 ();
 b15zdnd11an1n04x5 FILLER_156_712 ();
 b15zdnd00an1n02x5 FILLER_156_716 ();
 b15zdnd11an1n08x5 FILLER_156_726 ();
 b15zdnd11an1n04x5 FILLER_156_734 ();
 b15zdnd00an1n02x5 FILLER_156_738 ();
 b15zdnd11an1n64x5 FILLER_156_754 ();
 b15zdnd11an1n64x5 FILLER_156_818 ();
 b15zdnd11an1n64x5 FILLER_156_882 ();
 b15zdnd11an1n64x5 FILLER_156_946 ();
 b15zdnd11an1n64x5 FILLER_156_1010 ();
 b15zdnd11an1n32x5 FILLER_156_1074 ();
 b15zdnd11an1n16x5 FILLER_156_1106 ();
 b15zdnd00an1n02x5 FILLER_156_1122 ();
 b15zdnd11an1n04x5 FILLER_156_1127 ();
 b15zdnd11an1n64x5 FILLER_156_1134 ();
 b15zdnd11an1n64x5 FILLER_156_1198 ();
 b15zdnd11an1n64x5 FILLER_156_1262 ();
 b15zdnd11an1n64x5 FILLER_156_1326 ();
 b15zdnd11an1n64x5 FILLER_156_1390 ();
 b15zdnd11an1n64x5 FILLER_156_1454 ();
 b15zdnd11an1n16x5 FILLER_156_1518 ();
 b15zdnd11an1n64x5 FILLER_156_1586 ();
 b15zdnd11an1n16x5 FILLER_156_1650 ();
 b15zdnd00an1n02x5 FILLER_156_1666 ();
 b15zdnd00an1n01x5 FILLER_156_1668 ();
 b15zdnd11an1n64x5 FILLER_156_1672 ();
 b15zdnd11an1n64x5 FILLER_156_1736 ();
 b15zdnd11an1n64x5 FILLER_156_1800 ();
 b15zdnd11an1n64x5 FILLER_156_1864 ();
 b15zdnd11an1n64x5 FILLER_156_1928 ();
 b15zdnd11an1n64x5 FILLER_156_1992 ();
 b15zdnd11an1n64x5 FILLER_156_2056 ();
 b15zdnd11an1n32x5 FILLER_156_2120 ();
 b15zdnd00an1n02x5 FILLER_156_2152 ();
 b15zdnd11an1n64x5 FILLER_156_2162 ();
 b15zdnd11an1n32x5 FILLER_156_2226 ();
 b15zdnd11an1n16x5 FILLER_156_2258 ();
 b15zdnd00an1n02x5 FILLER_156_2274 ();
 b15zdnd11an1n32x5 FILLER_157_0 ();
 b15zdnd11an1n16x5 FILLER_157_32 ();
 b15zdnd11an1n08x5 FILLER_157_48 ();
 b15zdnd11an1n04x5 FILLER_157_56 ();
 b15zdnd11an1n04x5 FILLER_157_66 ();
 b15zdnd00an1n02x5 FILLER_157_70 ();
 b15zdnd00an1n01x5 FILLER_157_72 ();
 b15zdnd11an1n16x5 FILLER_157_94 ();
 b15zdnd11an1n08x5 FILLER_157_110 ();
 b15zdnd00an1n02x5 FILLER_157_118 ();
 b15zdnd00an1n01x5 FILLER_157_120 ();
 b15zdnd11an1n64x5 FILLER_157_139 ();
 b15zdnd11an1n16x5 FILLER_157_203 ();
 b15zdnd11an1n08x5 FILLER_157_219 ();
 b15zdnd00an1n02x5 FILLER_157_227 ();
 b15zdnd11an1n64x5 FILLER_157_232 ();
 b15zdnd11an1n64x5 FILLER_157_296 ();
 b15zdnd11an1n64x5 FILLER_157_360 ();
 b15zdnd11an1n64x5 FILLER_157_424 ();
 b15zdnd11an1n64x5 FILLER_157_488 ();
 b15zdnd11an1n64x5 FILLER_157_552 ();
 b15zdnd11an1n64x5 FILLER_157_616 ();
 b15zdnd11an1n16x5 FILLER_157_680 ();
 b15zdnd00an1n02x5 FILLER_157_696 ();
 b15zdnd00an1n01x5 FILLER_157_698 ();
 b15zdnd11an1n64x5 FILLER_157_730 ();
 b15zdnd11an1n64x5 FILLER_157_794 ();
 b15zdnd11an1n64x5 FILLER_157_858 ();
 b15zdnd11an1n64x5 FILLER_157_922 ();
 b15zdnd11an1n64x5 FILLER_157_986 ();
 b15zdnd11an1n32x5 FILLER_157_1050 ();
 b15zdnd11an1n04x5 FILLER_157_1082 ();
 b15zdnd00an1n01x5 FILLER_157_1086 ();
 b15zdnd11an1n64x5 FILLER_157_1090 ();
 b15zdnd11an1n64x5 FILLER_157_1154 ();
 b15zdnd11an1n16x5 FILLER_157_1218 ();
 b15zdnd11an1n64x5 FILLER_157_1237 ();
 b15zdnd11an1n64x5 FILLER_157_1301 ();
 b15zdnd11an1n64x5 FILLER_157_1365 ();
 b15zdnd11an1n64x5 FILLER_157_1429 ();
 b15zdnd11an1n32x5 FILLER_157_1493 ();
 b15zdnd11an1n16x5 FILLER_157_1525 ();
 b15zdnd11an1n08x5 FILLER_157_1541 ();
 b15zdnd00an1n02x5 FILLER_157_1549 ();
 b15zdnd00an1n01x5 FILLER_157_1551 ();
 b15zdnd11an1n04x5 FILLER_157_1555 ();
 b15zdnd11an1n64x5 FILLER_157_1562 ();
 b15zdnd11an1n64x5 FILLER_157_1626 ();
 b15zdnd11an1n64x5 FILLER_157_1690 ();
 b15zdnd11an1n64x5 FILLER_157_1754 ();
 b15zdnd11an1n64x5 FILLER_157_1818 ();
 b15zdnd11an1n64x5 FILLER_157_1882 ();
 b15zdnd11an1n64x5 FILLER_157_1946 ();
 b15zdnd11an1n64x5 FILLER_157_2010 ();
 b15zdnd11an1n64x5 FILLER_157_2074 ();
 b15zdnd11an1n64x5 FILLER_157_2138 ();
 b15zdnd11an1n64x5 FILLER_157_2202 ();
 b15zdnd11an1n16x5 FILLER_157_2266 ();
 b15zdnd00an1n02x5 FILLER_157_2282 ();
 b15zdnd11an1n64x5 FILLER_158_8 ();
 b15zdnd11an1n08x5 FILLER_158_72 ();
 b15zdnd11an1n04x5 FILLER_158_89 ();
 b15zdnd11an1n64x5 FILLER_158_98 ();
 b15zdnd11an1n32x5 FILLER_158_162 ();
 b15zdnd11an1n08x5 FILLER_158_194 ();
 b15zdnd11an1n64x5 FILLER_158_254 ();
 b15zdnd11an1n64x5 FILLER_158_318 ();
 b15zdnd11an1n16x5 FILLER_158_382 ();
 b15zdnd11an1n08x5 FILLER_158_398 ();
 b15zdnd11an1n04x5 FILLER_158_406 ();
 b15zdnd11an1n64x5 FILLER_158_452 ();
 b15zdnd11an1n64x5 FILLER_158_516 ();
 b15zdnd11an1n64x5 FILLER_158_580 ();
 b15zdnd11an1n64x5 FILLER_158_644 ();
 b15zdnd11an1n08x5 FILLER_158_708 ();
 b15zdnd00an1n02x5 FILLER_158_716 ();
 b15zdnd11an1n64x5 FILLER_158_726 ();
 b15zdnd11an1n64x5 FILLER_158_790 ();
 b15zdnd11an1n64x5 FILLER_158_854 ();
 b15zdnd11an1n64x5 FILLER_158_918 ();
 b15zdnd11an1n64x5 FILLER_158_982 ();
 b15zdnd11an1n32x5 FILLER_158_1046 ();
 b15zdnd11an1n08x5 FILLER_158_1078 ();
 b15zdnd00an1n01x5 FILLER_158_1086 ();
 b15zdnd11an1n64x5 FILLER_158_1114 ();
 b15zdnd11an1n32x5 FILLER_158_1178 ();
 b15zdnd11an1n16x5 FILLER_158_1210 ();
 b15zdnd11an1n08x5 FILLER_158_1226 ();
 b15zdnd00an1n01x5 FILLER_158_1234 ();
 b15zdnd11an1n64x5 FILLER_158_1238 ();
 b15zdnd11an1n64x5 FILLER_158_1302 ();
 b15zdnd11an1n64x5 FILLER_158_1366 ();
 b15zdnd11an1n64x5 FILLER_158_1430 ();
 b15zdnd11an1n64x5 FILLER_158_1494 ();
 b15zdnd00an1n02x5 FILLER_158_1558 ();
 b15zdnd11an1n64x5 FILLER_158_1563 ();
 b15zdnd11an1n64x5 FILLER_158_1627 ();
 b15zdnd11an1n64x5 FILLER_158_1691 ();
 b15zdnd11an1n64x5 FILLER_158_1755 ();
 b15zdnd11an1n64x5 FILLER_158_1819 ();
 b15zdnd11an1n64x5 FILLER_158_1883 ();
 b15zdnd11an1n64x5 FILLER_158_1947 ();
 b15zdnd11an1n32x5 FILLER_158_2011 ();
 b15zdnd11an1n16x5 FILLER_158_2043 ();
 b15zdnd11an1n08x5 FILLER_158_2059 ();
 b15zdnd00an1n01x5 FILLER_158_2067 ();
 b15zdnd11an1n32x5 FILLER_158_2110 ();
 b15zdnd11an1n08x5 FILLER_158_2142 ();
 b15zdnd11an1n04x5 FILLER_158_2150 ();
 b15zdnd11an1n64x5 FILLER_158_2162 ();
 b15zdnd11an1n32x5 FILLER_158_2226 ();
 b15zdnd11an1n16x5 FILLER_158_2258 ();
 b15zdnd00an1n02x5 FILLER_158_2274 ();
 b15zdnd11an1n32x5 FILLER_159_0 ();
 b15zdnd11an1n16x5 FILLER_159_32 ();
 b15zdnd11an1n08x5 FILLER_159_48 ();
 b15zdnd00an1n02x5 FILLER_159_56 ();
 b15zdnd00an1n01x5 FILLER_159_58 ();
 b15zdnd11an1n04x5 FILLER_159_63 ();
 b15zdnd00an1n01x5 FILLER_159_67 ();
 b15zdnd11an1n32x5 FILLER_159_71 ();
 b15zdnd11an1n16x5 FILLER_159_103 ();
 b15zdnd00an1n02x5 FILLER_159_119 ();
 b15zdnd00an1n01x5 FILLER_159_121 ();
 b15zdnd11an1n64x5 FILLER_159_136 ();
 b15zdnd11an1n16x5 FILLER_159_200 ();
 b15zdnd11an1n04x5 FILLER_159_216 ();
 b15zdnd00an1n01x5 FILLER_159_220 ();
 b15zdnd11an1n04x5 FILLER_159_224 ();
 b15zdnd11an1n32x5 FILLER_159_231 ();
 b15zdnd11an1n16x5 FILLER_159_263 ();
 b15zdnd11an1n08x5 FILLER_159_279 ();
 b15zdnd11an1n04x5 FILLER_159_287 ();
 b15zdnd00an1n02x5 FILLER_159_291 ();
 b15zdnd00an1n01x5 FILLER_159_293 ();
 b15zdnd11an1n64x5 FILLER_159_303 ();
 b15zdnd11an1n64x5 FILLER_159_367 ();
 b15zdnd11an1n64x5 FILLER_159_431 ();
 b15zdnd11an1n64x5 FILLER_159_495 ();
 b15zdnd11an1n04x5 FILLER_159_559 ();
 b15zdnd00an1n02x5 FILLER_159_563 ();
 b15zdnd11an1n64x5 FILLER_159_607 ();
 b15zdnd11an1n64x5 FILLER_159_671 ();
 b15zdnd11an1n64x5 FILLER_159_735 ();
 b15zdnd11an1n64x5 FILLER_159_799 ();
 b15zdnd11an1n64x5 FILLER_159_863 ();
 b15zdnd11an1n32x5 FILLER_159_927 ();
 b15zdnd11an1n16x5 FILLER_159_959 ();
 b15zdnd00an1n02x5 FILLER_159_975 ();
 b15zdnd11an1n64x5 FILLER_159_1005 ();
 b15zdnd11an1n64x5 FILLER_159_1069 ();
 b15zdnd11an1n64x5 FILLER_159_1133 ();
 b15zdnd11an1n08x5 FILLER_159_1197 ();
 b15zdnd11an1n04x5 FILLER_159_1205 ();
 b15zdnd00an1n01x5 FILLER_159_1209 ();
 b15zdnd11an1n16x5 FILLER_159_1262 ();
 b15zdnd11an1n04x5 FILLER_159_1278 ();
 b15zdnd00an1n02x5 FILLER_159_1282 ();
 b15zdnd11an1n64x5 FILLER_159_1307 ();
 b15zdnd11an1n64x5 FILLER_159_1371 ();
 b15zdnd11an1n64x5 FILLER_159_1435 ();
 b15zdnd11an1n64x5 FILLER_159_1499 ();
 b15zdnd11an1n08x5 FILLER_159_1563 ();
 b15zdnd11an1n04x5 FILLER_159_1571 ();
 b15zdnd00an1n02x5 FILLER_159_1575 ();
 b15zdnd00an1n01x5 FILLER_159_1577 ();
 b15zdnd11an1n08x5 FILLER_159_1620 ();
 b15zdnd11an1n04x5 FILLER_159_1628 ();
 b15zdnd00an1n02x5 FILLER_159_1632 ();
 b15zdnd11an1n04x5 FILLER_159_1637 ();
 b15zdnd00an1n02x5 FILLER_159_1641 ();
 b15zdnd00an1n01x5 FILLER_159_1643 ();
 b15zdnd11an1n64x5 FILLER_159_1671 ();
 b15zdnd11an1n64x5 FILLER_159_1735 ();
 b15zdnd11an1n64x5 FILLER_159_1799 ();
 b15zdnd11an1n64x5 FILLER_159_1863 ();
 b15zdnd11an1n64x5 FILLER_159_1927 ();
 b15zdnd11an1n64x5 FILLER_159_1991 ();
 b15zdnd11an1n64x5 FILLER_159_2055 ();
 b15zdnd11an1n64x5 FILLER_159_2119 ();
 b15zdnd11an1n64x5 FILLER_159_2183 ();
 b15zdnd11an1n16x5 FILLER_159_2247 ();
 b15zdnd11an1n08x5 FILLER_159_2263 ();
 b15zdnd00an1n01x5 FILLER_159_2271 ();
 b15zdnd11an1n08x5 FILLER_159_2276 ();
 b15zdnd11an1n32x5 FILLER_160_8 ();
 b15zdnd11an1n08x5 FILLER_160_40 ();
 b15zdnd11an1n04x5 FILLER_160_48 ();
 b15zdnd00an1n02x5 FILLER_160_52 ();
 b15zdnd00an1n01x5 FILLER_160_54 ();
 b15zdnd11an1n04x5 FILLER_160_63 ();
 b15zdnd11an1n32x5 FILLER_160_70 ();
 b15zdnd11an1n16x5 FILLER_160_102 ();
 b15zdnd11an1n04x5 FILLER_160_118 ();
 b15zdnd00an1n02x5 FILLER_160_122 ();
 b15zdnd11an1n64x5 FILLER_160_132 ();
 b15zdnd11an1n64x5 FILLER_160_196 ();
 b15zdnd11an1n64x5 FILLER_160_260 ();
 b15zdnd11an1n64x5 FILLER_160_324 ();
 b15zdnd11an1n64x5 FILLER_160_388 ();
 b15zdnd11an1n16x5 FILLER_160_452 ();
 b15zdnd11an1n08x5 FILLER_160_468 ();
 b15zdnd11an1n04x5 FILLER_160_476 ();
 b15zdnd00an1n01x5 FILLER_160_480 ();
 b15zdnd11an1n64x5 FILLER_160_523 ();
 b15zdnd11an1n64x5 FILLER_160_587 ();
 b15zdnd11an1n64x5 FILLER_160_651 ();
 b15zdnd00an1n02x5 FILLER_160_715 ();
 b15zdnd00an1n01x5 FILLER_160_717 ();
 b15zdnd11an1n64x5 FILLER_160_726 ();
 b15zdnd11an1n64x5 FILLER_160_790 ();
 b15zdnd11an1n64x5 FILLER_160_854 ();
 b15zdnd11an1n64x5 FILLER_160_918 ();
 b15zdnd11an1n64x5 FILLER_160_982 ();
 b15zdnd11an1n64x5 FILLER_160_1046 ();
 b15zdnd11an1n64x5 FILLER_160_1110 ();
 b15zdnd11an1n32x5 FILLER_160_1174 ();
 b15zdnd11an1n16x5 FILLER_160_1206 ();
 b15zdnd11an1n08x5 FILLER_160_1222 ();
 b15zdnd11an1n04x5 FILLER_160_1230 ();
 b15zdnd00an1n01x5 FILLER_160_1234 ();
 b15zdnd11an1n64x5 FILLER_160_1238 ();
 b15zdnd11an1n64x5 FILLER_160_1302 ();
 b15zdnd11an1n64x5 FILLER_160_1366 ();
 b15zdnd11an1n64x5 FILLER_160_1430 ();
 b15zdnd11an1n64x5 FILLER_160_1494 ();
 b15zdnd11an1n64x5 FILLER_160_1558 ();
 b15zdnd11an1n64x5 FILLER_160_1622 ();
 b15zdnd11an1n64x5 FILLER_160_1686 ();
 b15zdnd11an1n32x5 FILLER_160_1750 ();
 b15zdnd11an1n08x5 FILLER_160_1782 ();
 b15zdnd11an1n04x5 FILLER_160_1790 ();
 b15zdnd00an1n02x5 FILLER_160_1794 ();
 b15zdnd11an1n64x5 FILLER_160_1799 ();
 b15zdnd11an1n64x5 FILLER_160_1863 ();
 b15zdnd11an1n64x5 FILLER_160_1927 ();
 b15zdnd11an1n64x5 FILLER_160_1991 ();
 b15zdnd11an1n64x5 FILLER_160_2055 ();
 b15zdnd11an1n32x5 FILLER_160_2119 ();
 b15zdnd00an1n02x5 FILLER_160_2151 ();
 b15zdnd00an1n01x5 FILLER_160_2153 ();
 b15zdnd11an1n64x5 FILLER_160_2162 ();
 b15zdnd11an1n32x5 FILLER_160_2226 ();
 b15zdnd11an1n04x5 FILLER_160_2258 ();
 b15zdnd00an1n02x5 FILLER_160_2262 ();
 b15zdnd11an1n08x5 FILLER_160_2268 ();
 b15zdnd11an1n32x5 FILLER_161_0 ();
 b15zdnd11an1n08x5 FILLER_161_32 ();
 b15zdnd11an1n04x5 FILLER_161_40 ();
 b15zdnd00an1n02x5 FILLER_161_44 ();
 b15zdnd00an1n01x5 FILLER_161_46 ();
 b15zdnd11an1n04x5 FILLER_161_65 ();
 b15zdnd11an1n32x5 FILLER_161_73 ();
 b15zdnd11an1n08x5 FILLER_161_105 ();
 b15zdnd11an1n04x5 FILLER_161_113 ();
 b15zdnd11an1n04x5 FILLER_161_121 ();
 b15zdnd11an1n64x5 FILLER_161_131 ();
 b15zdnd11an1n64x5 FILLER_161_195 ();
 b15zdnd11an1n64x5 FILLER_161_259 ();
 b15zdnd11an1n64x5 FILLER_161_323 ();
 b15zdnd11an1n64x5 FILLER_161_387 ();
 b15zdnd11an1n64x5 FILLER_161_451 ();
 b15zdnd11an1n16x5 FILLER_161_515 ();
 b15zdnd11an1n04x5 FILLER_161_531 ();
 b15zdnd00an1n01x5 FILLER_161_535 ();
 b15zdnd11an1n64x5 FILLER_161_578 ();
 b15zdnd11an1n64x5 FILLER_161_642 ();
 b15zdnd11an1n64x5 FILLER_161_706 ();
 b15zdnd11an1n64x5 FILLER_161_770 ();
 b15zdnd11an1n64x5 FILLER_161_834 ();
 b15zdnd11an1n64x5 FILLER_161_898 ();
 b15zdnd11an1n64x5 FILLER_161_962 ();
 b15zdnd11an1n08x5 FILLER_161_1026 ();
 b15zdnd00an1n01x5 FILLER_161_1034 ();
 b15zdnd11an1n64x5 FILLER_161_1046 ();
 b15zdnd11an1n64x5 FILLER_161_1110 ();
 b15zdnd11an1n64x5 FILLER_161_1174 ();
 b15zdnd11an1n64x5 FILLER_161_1238 ();
 b15zdnd11an1n64x5 FILLER_161_1302 ();
 b15zdnd11an1n64x5 FILLER_161_1366 ();
 b15zdnd11an1n64x5 FILLER_161_1430 ();
 b15zdnd11an1n64x5 FILLER_161_1494 ();
 b15zdnd11an1n64x5 FILLER_161_1558 ();
 b15zdnd11an1n64x5 FILLER_161_1622 ();
 b15zdnd11an1n64x5 FILLER_161_1686 ();
 b15zdnd11an1n32x5 FILLER_161_1750 ();
 b15zdnd11an1n08x5 FILLER_161_1782 ();
 b15zdnd11an1n04x5 FILLER_161_1790 ();
 b15zdnd00an1n01x5 FILLER_161_1794 ();
 b15zdnd11an1n04x5 FILLER_161_1798 ();
 b15zdnd11an1n64x5 FILLER_161_1805 ();
 b15zdnd11an1n64x5 FILLER_161_1869 ();
 b15zdnd11an1n64x5 FILLER_161_1933 ();
 b15zdnd11an1n64x5 FILLER_161_1997 ();
 b15zdnd11an1n64x5 FILLER_161_2061 ();
 b15zdnd11an1n64x5 FILLER_161_2125 ();
 b15zdnd11an1n32x5 FILLER_161_2189 ();
 b15zdnd11an1n16x5 FILLER_161_2221 ();
 b15zdnd00an1n02x5 FILLER_161_2237 ();
 b15zdnd00an1n01x5 FILLER_161_2239 ();
 b15zdnd00an1n02x5 FILLER_161_2282 ();
 b15zdnd11an1n32x5 FILLER_162_8 ();
 b15zdnd11an1n08x5 FILLER_162_40 ();
 b15zdnd11an1n04x5 FILLER_162_48 ();
 b15zdnd00an1n02x5 FILLER_162_52 ();
 b15zdnd11an1n64x5 FILLER_162_61 ();
 b15zdnd11an1n64x5 FILLER_162_125 ();
 b15zdnd11an1n64x5 FILLER_162_189 ();
 b15zdnd11an1n64x5 FILLER_162_253 ();
 b15zdnd11an1n64x5 FILLER_162_317 ();
 b15zdnd11an1n64x5 FILLER_162_381 ();
 b15zdnd11an1n32x5 FILLER_162_445 ();
 b15zdnd00an1n01x5 FILLER_162_477 ();
 b15zdnd11an1n64x5 FILLER_162_520 ();
 b15zdnd11an1n64x5 FILLER_162_584 ();
 b15zdnd11an1n64x5 FILLER_162_648 ();
 b15zdnd11an1n04x5 FILLER_162_712 ();
 b15zdnd00an1n02x5 FILLER_162_716 ();
 b15zdnd11an1n64x5 FILLER_162_726 ();
 b15zdnd11an1n64x5 FILLER_162_790 ();
 b15zdnd11an1n64x5 FILLER_162_854 ();
 b15zdnd11an1n64x5 FILLER_162_918 ();
 b15zdnd11an1n16x5 FILLER_162_982 ();
 b15zdnd11an1n04x5 FILLER_162_998 ();
 b15zdnd00an1n02x5 FILLER_162_1002 ();
 b15zdnd00an1n01x5 FILLER_162_1004 ();
 b15zdnd11an1n64x5 FILLER_162_1057 ();
 b15zdnd11an1n64x5 FILLER_162_1121 ();
 b15zdnd11an1n64x5 FILLER_162_1185 ();
 b15zdnd11an1n64x5 FILLER_162_1249 ();
 b15zdnd11an1n64x5 FILLER_162_1313 ();
 b15zdnd11an1n64x5 FILLER_162_1377 ();
 b15zdnd11an1n64x5 FILLER_162_1441 ();
 b15zdnd11an1n64x5 FILLER_162_1505 ();
 b15zdnd11an1n64x5 FILLER_162_1569 ();
 b15zdnd11an1n64x5 FILLER_162_1633 ();
 b15zdnd11an1n64x5 FILLER_162_1697 ();
 b15zdnd11an1n08x5 FILLER_162_1761 ();
 b15zdnd11an1n04x5 FILLER_162_1769 ();
 b15zdnd00an1n02x5 FILLER_162_1773 ();
 b15zdnd00an1n01x5 FILLER_162_1775 ();
 b15zdnd11an1n64x5 FILLER_162_1828 ();
 b15zdnd11an1n32x5 FILLER_162_1892 ();
 b15zdnd11an1n16x5 FILLER_162_1924 ();
 b15zdnd00an1n02x5 FILLER_162_1940 ();
 b15zdnd11an1n64x5 FILLER_162_1945 ();
 b15zdnd11an1n64x5 FILLER_162_2009 ();
 b15zdnd11an1n32x5 FILLER_162_2073 ();
 b15zdnd11an1n08x5 FILLER_162_2105 ();
 b15zdnd11an1n04x5 FILLER_162_2113 ();
 b15zdnd00an1n02x5 FILLER_162_2117 ();
 b15zdnd11an1n08x5 FILLER_162_2146 ();
 b15zdnd11an1n64x5 FILLER_162_2162 ();
 b15zdnd11an1n04x5 FILLER_162_2226 ();
 b15zdnd00an1n02x5 FILLER_162_2230 ();
 b15zdnd00an1n02x5 FILLER_162_2274 ();
 b15zdnd11an1n32x5 FILLER_163_0 ();
 b15zdnd11an1n16x5 FILLER_163_32 ();
 b15zdnd11an1n08x5 FILLER_163_48 ();
 b15zdnd11an1n04x5 FILLER_163_56 ();
 b15zdnd11an1n64x5 FILLER_163_63 ();
 b15zdnd11an1n64x5 FILLER_163_127 ();
 b15zdnd11an1n64x5 FILLER_163_191 ();
 b15zdnd11an1n64x5 FILLER_163_255 ();
 b15zdnd11an1n32x5 FILLER_163_319 ();
 b15zdnd11an1n04x5 FILLER_163_351 ();
 b15zdnd00an1n02x5 FILLER_163_355 ();
 b15zdnd11an1n64x5 FILLER_163_363 ();
 b15zdnd11an1n64x5 FILLER_163_427 ();
 b15zdnd11an1n32x5 FILLER_163_491 ();
 b15zdnd11an1n16x5 FILLER_163_523 ();
 b15zdnd11an1n04x5 FILLER_163_539 ();
 b15zdnd00an1n01x5 FILLER_163_543 ();
 b15zdnd11an1n64x5 FILLER_163_586 ();
 b15zdnd11an1n64x5 FILLER_163_650 ();
 b15zdnd11an1n64x5 FILLER_163_714 ();
 b15zdnd11an1n64x5 FILLER_163_778 ();
 b15zdnd11an1n32x5 FILLER_163_842 ();
 b15zdnd11an1n16x5 FILLER_163_874 ();
 b15zdnd11an1n08x5 FILLER_163_890 ();
 b15zdnd00an1n02x5 FILLER_163_898 ();
 b15zdnd00an1n01x5 FILLER_163_900 ();
 b15zdnd11an1n08x5 FILLER_163_904 ();
 b15zdnd00an1n02x5 FILLER_163_912 ();
 b15zdnd00an1n01x5 FILLER_163_914 ();
 b15zdnd11an1n64x5 FILLER_163_957 ();
 b15zdnd11an1n04x5 FILLER_163_1021 ();
 b15zdnd11an1n04x5 FILLER_163_1028 ();
 b15zdnd11an1n04x5 FILLER_163_1035 ();
 b15zdnd11an1n64x5 FILLER_163_1042 ();
 b15zdnd11an1n64x5 FILLER_163_1106 ();
 b15zdnd11an1n64x5 FILLER_163_1170 ();
 b15zdnd11an1n64x5 FILLER_163_1234 ();
 b15zdnd11an1n64x5 FILLER_163_1298 ();
 b15zdnd11an1n64x5 FILLER_163_1362 ();
 b15zdnd11an1n64x5 FILLER_163_1426 ();
 b15zdnd11an1n64x5 FILLER_163_1490 ();
 b15zdnd11an1n64x5 FILLER_163_1554 ();
 b15zdnd11an1n64x5 FILLER_163_1618 ();
 b15zdnd11an1n64x5 FILLER_163_1682 ();
 b15zdnd11an1n32x5 FILLER_163_1746 ();
 b15zdnd11an1n08x5 FILLER_163_1778 ();
 b15zdnd00an1n02x5 FILLER_163_1786 ();
 b15zdnd11an1n64x5 FILLER_163_1840 ();
 b15zdnd11an1n08x5 FILLER_163_1904 ();
 b15zdnd11an1n04x5 FILLER_163_1912 ();
 b15zdnd11an1n64x5 FILLER_163_1968 ();
 b15zdnd11an1n64x5 FILLER_163_2032 ();
 b15zdnd11an1n08x5 FILLER_163_2096 ();
 b15zdnd11an1n04x5 FILLER_163_2104 ();
 b15zdnd00an1n02x5 FILLER_163_2108 ();
 b15zdnd11an1n64x5 FILLER_163_2137 ();
 b15zdnd11an1n64x5 FILLER_163_2201 ();
 b15zdnd11an1n16x5 FILLER_163_2265 ();
 b15zdnd00an1n02x5 FILLER_163_2281 ();
 b15zdnd00an1n01x5 FILLER_163_2283 ();
 b15zdnd11an1n32x5 FILLER_164_8 ();
 b15zdnd11an1n16x5 FILLER_164_40 ();
 b15zdnd00an1n02x5 FILLER_164_56 ();
 b15zdnd00an1n01x5 FILLER_164_58 ();
 b15zdnd11an1n64x5 FILLER_164_63 ();
 b15zdnd11an1n64x5 FILLER_164_127 ();
 b15zdnd11an1n64x5 FILLER_164_191 ();
 b15zdnd11an1n32x5 FILLER_164_255 ();
 b15zdnd11an1n16x5 FILLER_164_287 ();
 b15zdnd11an1n04x5 FILLER_164_303 ();
 b15zdnd00an1n01x5 FILLER_164_307 ();
 b15zdnd11an1n04x5 FILLER_164_317 ();
 b15zdnd11an1n16x5 FILLER_164_330 ();
 b15zdnd11an1n08x5 FILLER_164_346 ();
 b15zdnd11an1n04x5 FILLER_164_354 ();
 b15zdnd00an1n02x5 FILLER_164_358 ();
 b15zdnd00an1n01x5 FILLER_164_360 ();
 b15zdnd11an1n64x5 FILLER_164_367 ();
 b15zdnd11an1n64x5 FILLER_164_431 ();
 b15zdnd11an1n64x5 FILLER_164_495 ();
 b15zdnd11an1n64x5 FILLER_164_559 ();
 b15zdnd11an1n08x5 FILLER_164_623 ();
 b15zdnd11an1n04x5 FILLER_164_631 ();
 b15zdnd00an1n01x5 FILLER_164_635 ();
 b15zdnd11an1n64x5 FILLER_164_639 ();
 b15zdnd11an1n08x5 FILLER_164_703 ();
 b15zdnd11an1n04x5 FILLER_164_711 ();
 b15zdnd00an1n02x5 FILLER_164_715 ();
 b15zdnd00an1n01x5 FILLER_164_717 ();
 b15zdnd11an1n64x5 FILLER_164_726 ();
 b15zdnd11an1n64x5 FILLER_164_790 ();
 b15zdnd11an1n32x5 FILLER_164_854 ();
 b15zdnd11an1n08x5 FILLER_164_886 ();
 b15zdnd00an1n02x5 FILLER_164_894 ();
 b15zdnd11an1n04x5 FILLER_164_899 ();
 b15zdnd11an1n64x5 FILLER_164_945 ();
 b15zdnd11an1n32x5 FILLER_164_1009 ();
 b15zdnd11an1n16x5 FILLER_164_1041 ();
 b15zdnd11an1n08x5 FILLER_164_1057 ();
 b15zdnd11an1n04x5 FILLER_164_1065 ();
 b15zdnd00an1n02x5 FILLER_164_1069 ();
 b15zdnd11an1n64x5 FILLER_164_1080 ();
 b15zdnd11an1n04x5 FILLER_164_1144 ();
 b15zdnd00an1n01x5 FILLER_164_1148 ();
 b15zdnd11an1n64x5 FILLER_164_1152 ();
 b15zdnd11an1n64x5 FILLER_164_1216 ();
 b15zdnd11an1n64x5 FILLER_164_1280 ();
 b15zdnd11an1n64x5 FILLER_164_1344 ();
 b15zdnd11an1n64x5 FILLER_164_1408 ();
 b15zdnd11an1n64x5 FILLER_164_1472 ();
 b15zdnd11an1n32x5 FILLER_164_1536 ();
 b15zdnd00an1n02x5 FILLER_164_1568 ();
 b15zdnd00an1n01x5 FILLER_164_1570 ();
 b15zdnd11an1n32x5 FILLER_164_1580 ();
 b15zdnd11an1n08x5 FILLER_164_1612 ();
 b15zdnd11an1n04x5 FILLER_164_1620 ();
 b15zdnd00an1n02x5 FILLER_164_1624 ();
 b15zdnd00an1n01x5 FILLER_164_1626 ();
 b15zdnd11an1n64x5 FILLER_164_1636 ();
 b15zdnd11an1n64x5 FILLER_164_1700 ();
 b15zdnd11an1n32x5 FILLER_164_1764 ();
 b15zdnd11an1n08x5 FILLER_164_1796 ();
 b15zdnd00an1n01x5 FILLER_164_1804 ();
 b15zdnd11an1n04x5 FILLER_164_1808 ();
 b15zdnd00an1n01x5 FILLER_164_1812 ();
 b15zdnd11an1n04x5 FILLER_164_1816 ();
 b15zdnd11an1n64x5 FILLER_164_1823 ();
 b15zdnd11an1n32x5 FILLER_164_1887 ();
 b15zdnd11an1n08x5 FILLER_164_1919 ();
 b15zdnd11an1n04x5 FILLER_164_1927 ();
 b15zdnd00an1n02x5 FILLER_164_1931 ();
 b15zdnd11an1n04x5 FILLER_164_1936 ();
 b15zdnd11an1n08x5 FILLER_164_1943 ();
 b15zdnd11an1n64x5 FILLER_164_1993 ();
 b15zdnd11an1n32x5 FILLER_164_2057 ();
 b15zdnd11an1n16x5 FILLER_164_2089 ();
 b15zdnd11an1n04x5 FILLER_164_2105 ();
 b15zdnd00an1n01x5 FILLER_164_2109 ();
 b15zdnd11an1n08x5 FILLER_164_2113 ();
 b15zdnd11an1n16x5 FILLER_164_2124 ();
 b15zdnd11an1n08x5 FILLER_164_2140 ();
 b15zdnd11an1n04x5 FILLER_164_2148 ();
 b15zdnd00an1n02x5 FILLER_164_2152 ();
 b15zdnd11an1n64x5 FILLER_164_2162 ();
 b15zdnd11an1n32x5 FILLER_164_2226 ();
 b15zdnd11an1n16x5 FILLER_164_2258 ();
 b15zdnd00an1n02x5 FILLER_164_2274 ();
 b15zdnd11an1n64x5 FILLER_165_0 ();
 b15zdnd11an1n64x5 FILLER_165_64 ();
 b15zdnd11an1n64x5 FILLER_165_128 ();
 b15zdnd11an1n64x5 FILLER_165_192 ();
 b15zdnd11an1n64x5 FILLER_165_256 ();
 b15zdnd11an1n32x5 FILLER_165_320 ();
 b15zdnd11an1n08x5 FILLER_165_352 ();
 b15zdnd00an1n02x5 FILLER_165_360 ();
 b15zdnd00an1n01x5 FILLER_165_362 ();
 b15zdnd11an1n64x5 FILLER_165_405 ();
 b15zdnd11an1n64x5 FILLER_165_469 ();
 b15zdnd11an1n64x5 FILLER_165_533 ();
 b15zdnd11an1n08x5 FILLER_165_597 ();
 b15zdnd11an1n04x5 FILLER_165_605 ();
 b15zdnd11an1n64x5 FILLER_165_661 ();
 b15zdnd11an1n32x5 FILLER_165_725 ();
 b15zdnd11an1n64x5 FILLER_165_760 ();
 b15zdnd11an1n32x5 FILLER_165_824 ();
 b15zdnd11an1n16x5 FILLER_165_856 ();
 b15zdnd00an1n01x5 FILLER_165_872 ();
 b15zdnd11an1n64x5 FILLER_165_925 ();
 b15zdnd11an1n64x5 FILLER_165_989 ();
 b15zdnd11an1n64x5 FILLER_165_1053 ();
 b15zdnd11an1n04x5 FILLER_165_1117 ();
 b15zdnd00an1n01x5 FILLER_165_1121 ();
 b15zdnd11an1n64x5 FILLER_165_1174 ();
 b15zdnd11an1n64x5 FILLER_165_1238 ();
 b15zdnd11an1n32x5 FILLER_165_1302 ();
 b15zdnd11an1n08x5 FILLER_165_1334 ();
 b15zdnd00an1n02x5 FILLER_165_1342 ();
 b15zdnd00an1n01x5 FILLER_165_1344 ();
 b15zdnd11an1n64x5 FILLER_165_1348 ();
 b15zdnd11an1n64x5 FILLER_165_1412 ();
 b15zdnd11an1n64x5 FILLER_165_1476 ();
 b15zdnd11an1n64x5 FILLER_165_1540 ();
 b15zdnd11an1n08x5 FILLER_165_1604 ();
 b15zdnd11an1n04x5 FILLER_165_1612 ();
 b15zdnd00an1n02x5 FILLER_165_1616 ();
 b15zdnd00an1n01x5 FILLER_165_1618 ();
 b15zdnd11an1n64x5 FILLER_165_1628 ();
 b15zdnd11an1n64x5 FILLER_165_1692 ();
 b15zdnd11an1n16x5 FILLER_165_1756 ();
 b15zdnd11an1n04x5 FILLER_165_1772 ();
 b15zdnd11an1n64x5 FILLER_165_1803 ();
 b15zdnd11an1n32x5 FILLER_165_1867 ();
 b15zdnd11an1n16x5 FILLER_165_1899 ();
 b15zdnd11an1n04x5 FILLER_165_1915 ();
 b15zdnd00an1n02x5 FILLER_165_1919 ();
 b15zdnd00an1n01x5 FILLER_165_1921 ();
 b15zdnd11an1n64x5 FILLER_165_1964 ();
 b15zdnd11an1n32x5 FILLER_165_2028 ();
 b15zdnd11an1n04x5 FILLER_165_2060 ();
 b15zdnd11an1n64x5 FILLER_165_2075 ();
 b15zdnd11an1n64x5 FILLER_165_2139 ();
 b15zdnd11an1n64x5 FILLER_165_2203 ();
 b15zdnd11an1n16x5 FILLER_165_2267 ();
 b15zdnd00an1n01x5 FILLER_165_2283 ();
 b15zdnd11an1n64x5 FILLER_166_8 ();
 b15zdnd11an1n64x5 FILLER_166_72 ();
 b15zdnd11an1n64x5 FILLER_166_136 ();
 b15zdnd11an1n64x5 FILLER_166_200 ();
 b15zdnd11an1n64x5 FILLER_166_264 ();
 b15zdnd11an1n64x5 FILLER_166_328 ();
 b15zdnd11an1n16x5 FILLER_166_392 ();
 b15zdnd11an1n08x5 FILLER_166_408 ();
 b15zdnd11an1n04x5 FILLER_166_416 ();
 b15zdnd00an1n02x5 FILLER_166_420 ();
 b15zdnd00an1n01x5 FILLER_166_422 ();
 b15zdnd11an1n32x5 FILLER_166_431 ();
 b15zdnd11an1n04x5 FILLER_166_463 ();
 b15zdnd00an1n02x5 FILLER_166_467 ();
 b15zdnd11an1n64x5 FILLER_166_481 ();
 b15zdnd11an1n64x5 FILLER_166_545 ();
 b15zdnd11an1n16x5 FILLER_166_609 ();
 b15zdnd00an1n02x5 FILLER_166_625 ();
 b15zdnd00an1n01x5 FILLER_166_627 ();
 b15zdnd11an1n04x5 FILLER_166_631 ();
 b15zdnd11an1n64x5 FILLER_166_638 ();
 b15zdnd11an1n16x5 FILLER_166_702 ();
 b15zdnd11an1n04x5 FILLER_166_726 ();
 b15zdnd11an1n64x5 FILLER_166_782 ();
 b15zdnd11an1n32x5 FILLER_166_846 ();
 b15zdnd11an1n16x5 FILLER_166_878 ();
 b15zdnd00an1n01x5 FILLER_166_894 ();
 b15zdnd11an1n16x5 FILLER_166_898 ();
 b15zdnd11an1n08x5 FILLER_166_914 ();
 b15zdnd00an1n02x5 FILLER_166_922 ();
 b15zdnd11an1n32x5 FILLER_166_952 ();
 b15zdnd00an1n02x5 FILLER_166_984 ();
 b15zdnd00an1n01x5 FILLER_166_986 ();
 b15zdnd11an1n64x5 FILLER_166_998 ();
 b15zdnd11an1n64x5 FILLER_166_1062 ();
 b15zdnd11an1n08x5 FILLER_166_1126 ();
 b15zdnd11an1n04x5 FILLER_166_1134 ();
 b15zdnd00an1n02x5 FILLER_166_1138 ();
 b15zdnd11an1n04x5 FILLER_166_1143 ();
 b15zdnd11an1n64x5 FILLER_166_1150 ();
 b15zdnd11an1n32x5 FILLER_166_1214 ();
 b15zdnd11an1n16x5 FILLER_166_1246 ();
 b15zdnd00an1n01x5 FILLER_166_1262 ();
 b15zdnd11an1n32x5 FILLER_166_1286 ();
 b15zdnd00an1n02x5 FILLER_166_1318 ();
 b15zdnd11an1n32x5 FILLER_166_1372 ();
 b15zdnd11an1n16x5 FILLER_166_1404 ();
 b15zdnd11an1n08x5 FILLER_166_1420 ();
 b15zdnd00an1n01x5 FILLER_166_1428 ();
 b15zdnd11an1n04x5 FILLER_166_1432 ();
 b15zdnd11an1n64x5 FILLER_166_1462 ();
 b15zdnd11an1n64x5 FILLER_166_1526 ();
 b15zdnd11an1n64x5 FILLER_166_1590 ();
 b15zdnd11an1n64x5 FILLER_166_1654 ();
 b15zdnd11an1n32x5 FILLER_166_1718 ();
 b15zdnd11an1n16x5 FILLER_166_1750 ();
 b15zdnd11an1n08x5 FILLER_166_1766 ();
 b15zdnd00an1n02x5 FILLER_166_1774 ();
 b15zdnd00an1n01x5 FILLER_166_1776 ();
 b15zdnd11an1n64x5 FILLER_166_1780 ();
 b15zdnd11an1n64x5 FILLER_166_1844 ();
 b15zdnd11an1n64x5 FILLER_166_1908 ();
 b15zdnd11an1n32x5 FILLER_166_1972 ();
 b15zdnd11an1n16x5 FILLER_166_2004 ();
 b15zdnd11an1n04x5 FILLER_166_2020 ();
 b15zdnd00an1n02x5 FILLER_166_2024 ();
 b15zdnd00an1n01x5 FILLER_166_2026 ();
 b15zdnd11an1n04x5 FILLER_166_2079 ();
 b15zdnd11an1n64x5 FILLER_166_2090 ();
 b15zdnd11an1n32x5 FILLER_166_2162 ();
 b15zdnd11an1n16x5 FILLER_166_2194 ();
 b15zdnd11an1n04x5 FILLER_166_2210 ();
 b15zdnd00an1n01x5 FILLER_166_2214 ();
 b15zdnd11an1n04x5 FILLER_166_2218 ();
 b15zdnd11an1n32x5 FILLER_166_2225 ();
 b15zdnd11an1n16x5 FILLER_166_2257 ();
 b15zdnd00an1n02x5 FILLER_166_2273 ();
 b15zdnd00an1n01x5 FILLER_166_2275 ();
 b15zdnd11an1n64x5 FILLER_167_0 ();
 b15zdnd11an1n64x5 FILLER_167_64 ();
 b15zdnd11an1n08x5 FILLER_167_128 ();
 b15zdnd11an1n64x5 FILLER_167_139 ();
 b15zdnd11an1n64x5 FILLER_167_203 ();
 b15zdnd11an1n64x5 FILLER_167_267 ();
 b15zdnd11an1n64x5 FILLER_167_331 ();
 b15zdnd11an1n32x5 FILLER_167_395 ();
 b15zdnd11an1n16x5 FILLER_167_427 ();
 b15zdnd11an1n08x5 FILLER_167_443 ();
 b15zdnd00an1n02x5 FILLER_167_451 ();
 b15zdnd11an1n04x5 FILLER_167_460 ();
 b15zdnd11an1n04x5 FILLER_167_470 ();
 b15zdnd00an1n01x5 FILLER_167_474 ();
 b15zdnd11an1n64x5 FILLER_167_490 ();
 b15zdnd11an1n04x5 FILLER_167_554 ();
 b15zdnd11an1n08x5 FILLER_167_570 ();
 b15zdnd00an1n02x5 FILLER_167_578 ();
 b15zdnd00an1n01x5 FILLER_167_580 ();
 b15zdnd11an1n64x5 FILLER_167_595 ();
 b15zdnd11an1n64x5 FILLER_167_659 ();
 b15zdnd11an1n16x5 FILLER_167_723 ();
 b15zdnd11an1n08x5 FILLER_167_739 ();
 b15zdnd00an1n02x5 FILLER_167_747 ();
 b15zdnd11an1n04x5 FILLER_167_752 ();
 b15zdnd11an1n64x5 FILLER_167_759 ();
 b15zdnd11an1n16x5 FILLER_167_823 ();
 b15zdnd11an1n04x5 FILLER_167_839 ();
 b15zdnd11an1n04x5 FILLER_167_850 ();
 b15zdnd11an1n32x5 FILLER_167_857 ();
 b15zdnd11an1n16x5 FILLER_167_889 ();
 b15zdnd00an1n01x5 FILLER_167_905 ();
 b15zdnd11an1n64x5 FILLER_167_948 ();
 b15zdnd11an1n64x5 FILLER_167_1012 ();
 b15zdnd11an1n16x5 FILLER_167_1076 ();
 b15zdnd11an1n04x5 FILLER_167_1092 ();
 b15zdnd00an1n01x5 FILLER_167_1096 ();
 b15zdnd11an1n64x5 FILLER_167_1106 ();
 b15zdnd11an1n64x5 FILLER_167_1170 ();
 b15zdnd11an1n64x5 FILLER_167_1234 ();
 b15zdnd11an1n32x5 FILLER_167_1298 ();
 b15zdnd11an1n08x5 FILLER_167_1330 ();
 b15zdnd11an1n04x5 FILLER_167_1341 ();
 b15zdnd11an1n32x5 FILLER_167_1348 ();
 b15zdnd11an1n08x5 FILLER_167_1380 ();
 b15zdnd11an1n08x5 FILLER_167_1412 ();
 b15zdnd11an1n04x5 FILLER_167_1420 ();
 b15zdnd00an1n01x5 FILLER_167_1424 ();
 b15zdnd11an1n04x5 FILLER_167_1428 ();
 b15zdnd11an1n04x5 FILLER_167_1435 ();
 b15zdnd11an1n64x5 FILLER_167_1442 ();
 b15zdnd11an1n64x5 FILLER_167_1506 ();
 b15zdnd11an1n64x5 FILLER_167_1570 ();
 b15zdnd11an1n16x5 FILLER_167_1634 ();
 b15zdnd11an1n04x5 FILLER_167_1650 ();
 b15zdnd00an1n01x5 FILLER_167_1654 ();
 b15zdnd11an1n64x5 FILLER_167_1707 ();
 b15zdnd11an1n64x5 FILLER_167_1771 ();
 b15zdnd11an1n64x5 FILLER_167_1835 ();
 b15zdnd11an1n64x5 FILLER_167_1899 ();
 b15zdnd11an1n64x5 FILLER_167_1963 ();
 b15zdnd11an1n16x5 FILLER_167_2027 ();
 b15zdnd00an1n02x5 FILLER_167_2043 ();
 b15zdnd11an1n64x5 FILLER_167_2097 ();
 b15zdnd11an1n16x5 FILLER_167_2161 ();
 b15zdnd11an1n08x5 FILLER_167_2177 ();
 b15zdnd11an1n04x5 FILLER_167_2185 ();
 b15zdnd00an1n01x5 FILLER_167_2189 ();
 b15zdnd11an1n32x5 FILLER_167_2242 ();
 b15zdnd11an1n08x5 FILLER_167_2274 ();
 b15zdnd00an1n02x5 FILLER_167_2282 ();
 b15zdnd11an1n64x5 FILLER_168_8 ();
 b15zdnd11an1n64x5 FILLER_168_72 ();
 b15zdnd11an1n64x5 FILLER_168_136 ();
 b15zdnd11an1n64x5 FILLER_168_200 ();
 b15zdnd11an1n64x5 FILLER_168_264 ();
 b15zdnd11an1n32x5 FILLER_168_328 ();
 b15zdnd00an1n01x5 FILLER_168_360 ();
 b15zdnd11an1n04x5 FILLER_168_403 ();
 b15zdnd11an1n32x5 FILLER_168_418 ();
 b15zdnd11an1n64x5 FILLER_168_492 ();
 b15zdnd11an1n04x5 FILLER_168_556 ();
 b15zdnd00an1n02x5 FILLER_168_560 ();
 b15zdnd00an1n01x5 FILLER_168_562 ();
 b15zdnd11an1n64x5 FILLER_168_605 ();
 b15zdnd11an1n32x5 FILLER_168_669 ();
 b15zdnd11an1n16x5 FILLER_168_701 ();
 b15zdnd00an1n01x5 FILLER_168_717 ();
 b15zdnd11an1n08x5 FILLER_168_726 ();
 b15zdnd11an1n04x5 FILLER_168_734 ();
 b15zdnd00an1n02x5 FILLER_168_738 ();
 b15zdnd00an1n01x5 FILLER_168_740 ();
 b15zdnd11an1n32x5 FILLER_168_793 ();
 b15zdnd00an1n02x5 FILLER_168_825 ();
 b15zdnd11an1n32x5 FILLER_168_879 ();
 b15zdnd11an1n16x5 FILLER_168_911 ();
 b15zdnd11an1n08x5 FILLER_168_927 ();
 b15zdnd11an1n32x5 FILLER_168_940 ();
 b15zdnd11an1n08x5 FILLER_168_972 ();
 b15zdnd11an1n64x5 FILLER_168_1000 ();
 b15zdnd11an1n32x5 FILLER_168_1064 ();
 b15zdnd00an1n02x5 FILLER_168_1096 ();
 b15zdnd00an1n01x5 FILLER_168_1098 ();
 b15zdnd11an1n64x5 FILLER_168_1108 ();
 b15zdnd11an1n64x5 FILLER_168_1172 ();
 b15zdnd11an1n64x5 FILLER_168_1236 ();
 b15zdnd11an1n32x5 FILLER_168_1300 ();
 b15zdnd11an1n08x5 FILLER_168_1332 ();
 b15zdnd00an1n02x5 FILLER_168_1340 ();
 b15zdnd11an1n08x5 FILLER_168_1345 ();
 b15zdnd11an1n04x5 FILLER_168_1353 ();
 b15zdnd11an1n04x5 FILLER_168_1368 ();
 b15zdnd11an1n16x5 FILLER_168_1383 ();
 b15zdnd11an1n08x5 FILLER_168_1399 ();
 b15zdnd00an1n02x5 FILLER_168_1407 ();
 b15zdnd11an1n64x5 FILLER_168_1461 ();
 b15zdnd11an1n64x5 FILLER_168_1525 ();
 b15zdnd11an1n64x5 FILLER_168_1589 ();
 b15zdnd11an1n16x5 FILLER_168_1653 ();
 b15zdnd11an1n04x5 FILLER_168_1669 ();
 b15zdnd11an1n04x5 FILLER_168_1676 ();
 b15zdnd11an1n64x5 FILLER_168_1683 ();
 b15zdnd11an1n64x5 FILLER_168_1747 ();
 b15zdnd11an1n32x5 FILLER_168_1811 ();
 b15zdnd11an1n04x5 FILLER_168_1843 ();
 b15zdnd00an1n02x5 FILLER_168_1847 ();
 b15zdnd11an1n64x5 FILLER_168_1858 ();
 b15zdnd11an1n64x5 FILLER_168_1922 ();
 b15zdnd11an1n32x5 FILLER_168_1986 ();
 b15zdnd11an1n08x5 FILLER_168_2018 ();
 b15zdnd00an1n02x5 FILLER_168_2026 ();
 b15zdnd11an1n08x5 FILLER_168_2035 ();
 b15zdnd00an1n02x5 FILLER_168_2043 ();
 b15zdnd00an1n01x5 FILLER_168_2045 ();
 b15zdnd11an1n04x5 FILLER_168_2049 ();
 b15zdnd11an1n04x5 FILLER_168_2056 ();
 b15zdnd11an1n04x5 FILLER_168_2063 ();
 b15zdnd11an1n04x5 FILLER_168_2070 ();
 b15zdnd11an1n08x5 FILLER_168_2077 ();
 b15zdnd11an1n16x5 FILLER_168_2127 ();
 b15zdnd11an1n08x5 FILLER_168_2143 ();
 b15zdnd00an1n02x5 FILLER_168_2151 ();
 b15zdnd00an1n01x5 FILLER_168_2153 ();
 b15zdnd11an1n32x5 FILLER_168_2162 ();
 b15zdnd11an1n16x5 FILLER_168_2194 ();
 b15zdnd11an1n04x5 FILLER_168_2210 ();
 b15zdnd00an1n01x5 FILLER_168_2214 ();
 b15zdnd11an1n04x5 FILLER_168_2218 ();
 b15zdnd00an1n01x5 FILLER_168_2222 ();
 b15zdnd11an1n08x5 FILLER_168_2265 ();
 b15zdnd00an1n02x5 FILLER_168_2273 ();
 b15zdnd00an1n01x5 FILLER_168_2275 ();
 b15zdnd11an1n64x5 FILLER_169_0 ();
 b15zdnd11an1n64x5 FILLER_169_64 ();
 b15zdnd11an1n64x5 FILLER_169_128 ();
 b15zdnd11an1n64x5 FILLER_169_192 ();
 b15zdnd11an1n64x5 FILLER_169_256 ();
 b15zdnd11an1n32x5 FILLER_169_320 ();
 b15zdnd00an1n01x5 FILLER_169_352 ();
 b15zdnd11an1n64x5 FILLER_169_356 ();
 b15zdnd00an1n02x5 FILLER_169_420 ();
 b15zdnd00an1n01x5 FILLER_169_422 ();
 b15zdnd11an1n04x5 FILLER_169_465 ();
 b15zdnd11an1n64x5 FILLER_169_481 ();
 b15zdnd11an1n16x5 FILLER_169_545 ();
 b15zdnd11an1n04x5 FILLER_169_561 ();
 b15zdnd00an1n02x5 FILLER_169_565 ();
 b15zdnd00an1n01x5 FILLER_169_567 ();
 b15zdnd11an1n64x5 FILLER_169_610 ();
 b15zdnd11an1n32x5 FILLER_169_674 ();
 b15zdnd11an1n16x5 FILLER_169_706 ();
 b15zdnd11an1n08x5 FILLER_169_722 ();
 b15zdnd00an1n02x5 FILLER_169_730 ();
 b15zdnd11an1n04x5 FILLER_169_774 ();
 b15zdnd11an1n08x5 FILLER_169_781 ();
 b15zdnd00an1n02x5 FILLER_169_789 ();
 b15zdnd11an1n16x5 FILLER_169_833 ();
 b15zdnd11an1n04x5 FILLER_169_849 ();
 b15zdnd11an1n04x5 FILLER_169_856 ();
 b15zdnd11an1n64x5 FILLER_169_863 ();
 b15zdnd11an1n04x5 FILLER_169_927 ();
 b15zdnd00an1n01x5 FILLER_169_931 ();
 b15zdnd11an1n64x5 FILLER_169_949 ();
 b15zdnd11an1n64x5 FILLER_169_1013 ();
 b15zdnd11an1n64x5 FILLER_169_1077 ();
 b15zdnd11an1n64x5 FILLER_169_1141 ();
 b15zdnd11an1n64x5 FILLER_169_1205 ();
 b15zdnd11an1n32x5 FILLER_169_1269 ();
 b15zdnd11an1n08x5 FILLER_169_1301 ();
 b15zdnd11an1n04x5 FILLER_169_1309 ();
 b15zdnd00an1n02x5 FILLER_169_1313 ();
 b15zdnd00an1n01x5 FILLER_169_1315 ();
 b15zdnd11an1n32x5 FILLER_169_1368 ();
 b15zdnd11an1n04x5 FILLER_169_1400 ();
 b15zdnd00an1n02x5 FILLER_169_1404 ();
 b15zdnd00an1n01x5 FILLER_169_1406 ();
 b15zdnd11an1n64x5 FILLER_169_1459 ();
 b15zdnd00an1n01x5 FILLER_169_1523 ();
 b15zdnd11an1n64x5 FILLER_169_1576 ();
 b15zdnd11an1n32x5 FILLER_169_1640 ();
 b15zdnd11an1n08x5 FILLER_169_1672 ();
 b15zdnd11an1n64x5 FILLER_169_1683 ();
 b15zdnd11an1n64x5 FILLER_169_1747 ();
 b15zdnd11an1n64x5 FILLER_169_1811 ();
 b15zdnd11an1n64x5 FILLER_169_1875 ();
 b15zdnd11an1n64x5 FILLER_169_1939 ();
 b15zdnd11an1n32x5 FILLER_169_2003 ();
 b15zdnd11an1n04x5 FILLER_169_2035 ();
 b15zdnd11an1n08x5 FILLER_169_2059 ();
 b15zdnd00an1n02x5 FILLER_169_2067 ();
 b15zdnd00an1n01x5 FILLER_169_2069 ();
 b15zdnd11an1n16x5 FILLER_169_2073 ();
 b15zdnd00an1n01x5 FILLER_169_2089 ();
 b15zdnd11an1n64x5 FILLER_169_2132 ();
 b15zdnd11an1n08x5 FILLER_169_2196 ();
 b15zdnd11an1n04x5 FILLER_169_2204 ();
 b15zdnd11an1n04x5 FILLER_169_2250 ();
 b15zdnd11an1n04x5 FILLER_169_2261 ();
 b15zdnd11an1n08x5 FILLER_169_2272 ();
 b15zdnd11an1n04x5 FILLER_169_2280 ();
 b15zdnd11an1n64x5 FILLER_170_8 ();
 b15zdnd11an1n64x5 FILLER_170_72 ();
 b15zdnd11an1n64x5 FILLER_170_136 ();
 b15zdnd11an1n64x5 FILLER_170_200 ();
 b15zdnd11an1n64x5 FILLER_170_264 ();
 b15zdnd11an1n16x5 FILLER_170_328 ();
 b15zdnd11an1n08x5 FILLER_170_344 ();
 b15zdnd00an1n02x5 FILLER_170_352 ();
 b15zdnd11an1n08x5 FILLER_170_357 ();
 b15zdnd11an1n32x5 FILLER_170_371 ();
 b15zdnd11an1n16x5 FILLER_170_403 ();
 b15zdnd11an1n08x5 FILLER_170_419 ();
 b15zdnd11an1n04x5 FILLER_170_427 ();
 b15zdnd00an1n02x5 FILLER_170_431 ();
 b15zdnd11an1n08x5 FILLER_170_475 ();
 b15zdnd11an1n64x5 FILLER_170_490 ();
 b15zdnd11an1n64x5 FILLER_170_554 ();
 b15zdnd11an1n64x5 FILLER_170_618 ();
 b15zdnd11an1n32x5 FILLER_170_682 ();
 b15zdnd11an1n04x5 FILLER_170_714 ();
 b15zdnd11an1n04x5 FILLER_170_726 ();
 b15zdnd00an1n01x5 FILLER_170_730 ();
 b15zdnd11an1n16x5 FILLER_170_737 ();
 b15zdnd11an1n08x5 FILLER_170_753 ();
 b15zdnd11an1n04x5 FILLER_170_764 ();
 b15zdnd11an1n16x5 FILLER_170_771 ();
 b15zdnd00an1n02x5 FILLER_170_787 ();
 b15zdnd00an1n01x5 FILLER_170_789 ();
 b15zdnd11an1n64x5 FILLER_170_797 ();
 b15zdnd11an1n64x5 FILLER_170_861 ();
 b15zdnd00an1n01x5 FILLER_170_925 ();
 b15zdnd11an1n64x5 FILLER_170_929 ();
 b15zdnd11an1n64x5 FILLER_170_993 ();
 b15zdnd11an1n64x5 FILLER_170_1057 ();
 b15zdnd11an1n64x5 FILLER_170_1121 ();
 b15zdnd11an1n64x5 FILLER_170_1185 ();
 b15zdnd11an1n04x5 FILLER_170_1249 ();
 b15zdnd00an1n01x5 FILLER_170_1253 ();
 b15zdnd11an1n64x5 FILLER_170_1277 ();
 b15zdnd11an1n64x5 FILLER_170_1344 ();
 b15zdnd11an1n16x5 FILLER_170_1408 ();
 b15zdnd11an1n04x5 FILLER_170_1424 ();
 b15zdnd00an1n01x5 FILLER_170_1428 ();
 b15zdnd11an1n04x5 FILLER_170_1432 ();
 b15zdnd11an1n64x5 FILLER_170_1439 ();
 b15zdnd11an1n32x5 FILLER_170_1503 ();
 b15zdnd11an1n08x5 FILLER_170_1535 ();
 b15zdnd11an1n04x5 FILLER_170_1546 ();
 b15zdnd11an1n64x5 FILLER_170_1553 ();
 b15zdnd11an1n64x5 FILLER_170_1617 ();
 b15zdnd11an1n64x5 FILLER_170_1681 ();
 b15zdnd11an1n64x5 FILLER_170_1745 ();
 b15zdnd11an1n64x5 FILLER_170_1809 ();
 b15zdnd11an1n64x5 FILLER_170_1873 ();
 b15zdnd11an1n64x5 FILLER_170_1937 ();
 b15zdnd11an1n64x5 FILLER_170_2001 ();
 b15zdnd11an1n32x5 FILLER_170_2065 ();
 b15zdnd11an1n04x5 FILLER_170_2097 ();
 b15zdnd00an1n01x5 FILLER_170_2101 ();
 b15zdnd11an1n32x5 FILLER_170_2109 ();
 b15zdnd11an1n08x5 FILLER_170_2141 ();
 b15zdnd11an1n04x5 FILLER_170_2149 ();
 b15zdnd00an1n01x5 FILLER_170_2153 ();
 b15zdnd11an1n32x5 FILLER_170_2162 ();
 b15zdnd11an1n16x5 FILLER_170_2194 ();
 b15zdnd11an1n08x5 FILLER_170_2210 ();
 b15zdnd11an1n04x5 FILLER_170_2218 ();
 b15zdnd11an1n04x5 FILLER_170_2228 ();
 b15zdnd00an1n02x5 FILLER_170_2274 ();
 b15zdnd11an1n64x5 FILLER_171_0 ();
 b15zdnd11an1n64x5 FILLER_171_64 ();
 b15zdnd11an1n64x5 FILLER_171_128 ();
 b15zdnd11an1n64x5 FILLER_171_192 ();
 b15zdnd11an1n64x5 FILLER_171_256 ();
 b15zdnd11an1n08x5 FILLER_171_320 ();
 b15zdnd00an1n02x5 FILLER_171_328 ();
 b15zdnd11an1n16x5 FILLER_171_382 ();
 b15zdnd11an1n04x5 FILLER_171_398 ();
 b15zdnd00an1n01x5 FILLER_171_402 ();
 b15zdnd11an1n16x5 FILLER_171_409 ();
 b15zdnd11an1n04x5 FILLER_171_467 ();
 b15zdnd11an1n16x5 FILLER_171_483 ();
 b15zdnd11an1n08x5 FILLER_171_499 ();
 b15zdnd00an1n01x5 FILLER_171_507 ();
 b15zdnd11an1n64x5 FILLER_171_515 ();
 b15zdnd11an1n64x5 FILLER_171_579 ();
 b15zdnd11an1n64x5 FILLER_171_643 ();
 b15zdnd11an1n08x5 FILLER_171_707 ();
 b15zdnd11an1n04x5 FILLER_171_715 ();
 b15zdnd11an1n08x5 FILLER_171_729 ();
 b15zdnd11an1n04x5 FILLER_171_737 ();
 b15zdnd00an1n01x5 FILLER_171_741 ();
 b15zdnd11an1n64x5 FILLER_171_753 ();
 b15zdnd11an1n64x5 FILLER_171_817 ();
 b15zdnd11an1n04x5 FILLER_171_881 ();
 b15zdnd00an1n01x5 FILLER_171_885 ();
 b15zdnd11an1n64x5 FILLER_171_928 ();
 b15zdnd11an1n64x5 FILLER_171_992 ();
 b15zdnd11an1n64x5 FILLER_171_1056 ();
 b15zdnd11an1n64x5 FILLER_171_1120 ();
 b15zdnd11an1n64x5 FILLER_171_1184 ();
 b15zdnd11an1n64x5 FILLER_171_1248 ();
 b15zdnd11an1n16x5 FILLER_171_1312 ();
 b15zdnd11an1n08x5 FILLER_171_1328 ();
 b15zdnd11an1n04x5 FILLER_171_1336 ();
 b15zdnd00an1n02x5 FILLER_171_1340 ();
 b15zdnd11an1n64x5 FILLER_171_1345 ();
 b15zdnd11an1n32x5 FILLER_171_1409 ();
 b15zdnd11an1n08x5 FILLER_171_1441 ();
 b15zdnd11an1n04x5 FILLER_171_1449 ();
 b15zdnd00an1n02x5 FILLER_171_1453 ();
 b15zdnd00an1n01x5 FILLER_171_1455 ();
 b15zdnd11an1n64x5 FILLER_171_1467 ();
 b15zdnd11an1n16x5 FILLER_171_1531 ();
 b15zdnd00an1n02x5 FILLER_171_1547 ();
 b15zdnd11an1n64x5 FILLER_171_1552 ();
 b15zdnd11an1n64x5 FILLER_171_1616 ();
 b15zdnd11an1n64x5 FILLER_171_1680 ();
 b15zdnd11an1n64x5 FILLER_171_1744 ();
 b15zdnd11an1n64x5 FILLER_171_1808 ();
 b15zdnd11an1n64x5 FILLER_171_1872 ();
 b15zdnd11an1n64x5 FILLER_171_1936 ();
 b15zdnd11an1n64x5 FILLER_171_2000 ();
 b15zdnd11an1n64x5 FILLER_171_2064 ();
 b15zdnd11an1n64x5 FILLER_171_2128 ();
 b15zdnd11an1n32x5 FILLER_171_2192 ();
 b15zdnd11an1n04x5 FILLER_171_2224 ();
 b15zdnd00an1n01x5 FILLER_171_2228 ();
 b15zdnd11an1n04x5 FILLER_171_2235 ();
 b15zdnd00an1n01x5 FILLER_171_2239 ();
 b15zdnd00an1n02x5 FILLER_171_2282 ();
 b15zdnd11an1n64x5 FILLER_172_8 ();
 b15zdnd11an1n64x5 FILLER_172_72 ();
 b15zdnd11an1n64x5 FILLER_172_136 ();
 b15zdnd00an1n01x5 FILLER_172_200 ();
 b15zdnd11an1n64x5 FILLER_172_253 ();
 b15zdnd11an1n32x5 FILLER_172_317 ();
 b15zdnd11an1n04x5 FILLER_172_349 ();
 b15zdnd00an1n02x5 FILLER_172_353 ();
 b15zdnd00an1n01x5 FILLER_172_355 ();
 b15zdnd11an1n08x5 FILLER_172_359 ();
 b15zdnd00an1n02x5 FILLER_172_367 ();
 b15zdnd00an1n01x5 FILLER_172_369 ();
 b15zdnd11an1n32x5 FILLER_172_412 ();
 b15zdnd11an1n16x5 FILLER_172_444 ();
 b15zdnd11an1n08x5 FILLER_172_460 ();
 b15zdnd00an1n02x5 FILLER_172_468 ();
 b15zdnd11an1n64x5 FILLER_172_512 ();
 b15zdnd11an1n64x5 FILLER_172_576 ();
 b15zdnd11an1n64x5 FILLER_172_640 ();
 b15zdnd11an1n08x5 FILLER_172_704 ();
 b15zdnd11an1n04x5 FILLER_172_712 ();
 b15zdnd00an1n02x5 FILLER_172_716 ();
 b15zdnd11an1n08x5 FILLER_172_726 ();
 b15zdnd11an1n04x5 FILLER_172_734 ();
 b15zdnd11an1n64x5 FILLER_172_752 ();
 b15zdnd11an1n64x5 FILLER_172_816 ();
 b15zdnd11an1n08x5 FILLER_172_880 ();
 b15zdnd11an1n04x5 FILLER_172_888 ();
 b15zdnd00an1n01x5 FILLER_172_892 ();
 b15zdnd11an1n32x5 FILLER_172_900 ();
 b15zdnd00an1n02x5 FILLER_172_932 ();
 b15zdnd11an1n64x5 FILLER_172_950 ();
 b15zdnd11an1n64x5 FILLER_172_1014 ();
 b15zdnd11an1n64x5 FILLER_172_1078 ();
 b15zdnd11an1n64x5 FILLER_172_1142 ();
 b15zdnd11an1n32x5 FILLER_172_1206 ();
 b15zdnd11an1n16x5 FILLER_172_1238 ();
 b15zdnd11an1n04x5 FILLER_172_1254 ();
 b15zdnd00an1n02x5 FILLER_172_1258 ();
 b15zdnd00an1n01x5 FILLER_172_1260 ();
 b15zdnd11an1n64x5 FILLER_172_1284 ();
 b15zdnd11an1n64x5 FILLER_172_1348 ();
 b15zdnd11an1n64x5 FILLER_172_1412 ();
 b15zdnd11an1n64x5 FILLER_172_1476 ();
 b15zdnd11an1n64x5 FILLER_172_1540 ();
 b15zdnd11an1n64x5 FILLER_172_1604 ();
 b15zdnd11an1n64x5 FILLER_172_1668 ();
 b15zdnd11an1n64x5 FILLER_172_1732 ();
 b15zdnd11an1n64x5 FILLER_172_1796 ();
 b15zdnd11an1n16x5 FILLER_172_1860 ();
 b15zdnd00an1n02x5 FILLER_172_1876 ();
 b15zdnd11an1n64x5 FILLER_172_1887 ();
 b15zdnd11an1n64x5 FILLER_172_1951 ();
 b15zdnd11an1n64x5 FILLER_172_2015 ();
 b15zdnd11an1n64x5 FILLER_172_2079 ();
 b15zdnd11an1n08x5 FILLER_172_2143 ();
 b15zdnd00an1n02x5 FILLER_172_2151 ();
 b15zdnd00an1n01x5 FILLER_172_2153 ();
 b15zdnd11an1n64x5 FILLER_172_2162 ();
 b15zdnd00an1n02x5 FILLER_172_2226 ();
 b15zdnd00an1n01x5 FILLER_172_2228 ();
 b15zdnd00an1n02x5 FILLER_172_2274 ();
 b15zdnd11an1n64x5 FILLER_173_0 ();
 b15zdnd11an1n64x5 FILLER_173_64 ();
 b15zdnd11an1n64x5 FILLER_173_128 ();
 b15zdnd11an1n16x5 FILLER_173_192 ();
 b15zdnd11an1n08x5 FILLER_173_208 ();
 b15zdnd11an1n04x5 FILLER_173_216 ();
 b15zdnd11an1n04x5 FILLER_173_223 ();
 b15zdnd11an1n64x5 FILLER_173_230 ();
 b15zdnd11an1n64x5 FILLER_173_294 ();
 b15zdnd11an1n08x5 FILLER_173_358 ();
 b15zdnd11an1n04x5 FILLER_173_366 ();
 b15zdnd00an1n01x5 FILLER_173_370 ();
 b15zdnd11an1n64x5 FILLER_173_385 ();
 b15zdnd11an1n08x5 FILLER_173_449 ();
 b15zdnd11an1n04x5 FILLER_173_457 ();
 b15zdnd11an1n04x5 FILLER_173_469 ();
 b15zdnd11an1n32x5 FILLER_173_515 ();
 b15zdnd11an1n08x5 FILLER_173_547 ();
 b15zdnd11an1n64x5 FILLER_173_567 ();
 b15zdnd11an1n64x5 FILLER_173_631 ();
 b15zdnd11an1n64x5 FILLER_173_695 ();
 b15zdnd11an1n64x5 FILLER_173_759 ();
 b15zdnd11an1n64x5 FILLER_173_823 ();
 b15zdnd11an1n64x5 FILLER_173_887 ();
 b15zdnd11an1n64x5 FILLER_173_951 ();
 b15zdnd11an1n64x5 FILLER_173_1015 ();
 b15zdnd11an1n64x5 FILLER_173_1079 ();
 b15zdnd11an1n64x5 FILLER_173_1143 ();
 b15zdnd11an1n32x5 FILLER_173_1207 ();
 b15zdnd00an1n02x5 FILLER_173_1239 ();
 b15zdnd00an1n01x5 FILLER_173_1241 ();
 b15zdnd11an1n64x5 FILLER_173_1262 ();
 b15zdnd11an1n32x5 FILLER_173_1326 ();
 b15zdnd11an1n16x5 FILLER_173_1358 ();
 b15zdnd00an1n02x5 FILLER_173_1374 ();
 b15zdnd00an1n01x5 FILLER_173_1376 ();
 b15zdnd11an1n64x5 FILLER_173_1386 ();
 b15zdnd11an1n64x5 FILLER_173_1450 ();
 b15zdnd11an1n32x5 FILLER_173_1514 ();
 b15zdnd11an1n04x5 FILLER_173_1546 ();
 b15zdnd11an1n64x5 FILLER_173_1553 ();
 b15zdnd11an1n16x5 FILLER_173_1617 ();
 b15zdnd11an1n08x5 FILLER_173_1633 ();
 b15zdnd11an1n04x5 FILLER_173_1641 ();
 b15zdnd11an1n32x5 FILLER_173_1653 ();
 b15zdnd11an1n16x5 FILLER_173_1685 ();
 b15zdnd11an1n64x5 FILLER_173_1704 ();
 b15zdnd11an1n64x5 FILLER_173_1768 ();
 b15zdnd11an1n32x5 FILLER_173_1832 ();
 b15zdnd11an1n08x5 FILLER_173_1864 ();
 b15zdnd11an1n04x5 FILLER_173_1872 ();
 b15zdnd00an1n01x5 FILLER_173_1876 ();
 b15zdnd11an1n64x5 FILLER_173_1886 ();
 b15zdnd11an1n32x5 FILLER_173_1950 ();
 b15zdnd11an1n08x5 FILLER_173_1982 ();
 b15zdnd00an1n02x5 FILLER_173_1990 ();
 b15zdnd00an1n01x5 FILLER_173_1992 ();
 b15zdnd11an1n64x5 FILLER_173_2035 ();
 b15zdnd11an1n64x5 FILLER_173_2099 ();
 b15zdnd11an1n64x5 FILLER_173_2163 ();
 b15zdnd11an1n08x5 FILLER_173_2227 ();
 b15zdnd11an1n04x5 FILLER_173_2235 ();
 b15zdnd00an1n01x5 FILLER_173_2239 ();
 b15zdnd00an1n02x5 FILLER_173_2282 ();
 b15zdnd11an1n32x5 FILLER_174_8 ();
 b15zdnd11an1n08x5 FILLER_174_40 ();
 b15zdnd00an1n02x5 FILLER_174_48 ();
 b15zdnd00an1n01x5 FILLER_174_50 ();
 b15zdnd11an1n64x5 FILLER_174_93 ();
 b15zdnd11an1n64x5 FILLER_174_157 ();
 b15zdnd11an1n04x5 FILLER_174_221 ();
 b15zdnd00an1n02x5 FILLER_174_225 ();
 b15zdnd00an1n01x5 FILLER_174_227 ();
 b15zdnd11an1n16x5 FILLER_174_231 ();
 b15zdnd11an1n04x5 FILLER_174_247 ();
 b15zdnd00an1n02x5 FILLER_174_251 ();
 b15zdnd00an1n01x5 FILLER_174_253 ();
 b15zdnd11an1n64x5 FILLER_174_274 ();
 b15zdnd11an1n08x5 FILLER_174_338 ();
 b15zdnd11an1n04x5 FILLER_174_346 ();
 b15zdnd00an1n01x5 FILLER_174_350 ();
 b15zdnd11an1n04x5 FILLER_174_403 ();
 b15zdnd11an1n04x5 FILLER_174_449 ();
 b15zdnd00an1n02x5 FILLER_174_453 ();
 b15zdnd11an1n16x5 FILLER_174_461 ();
 b15zdnd00an1n02x5 FILLER_174_477 ();
 b15zdnd11an1n04x5 FILLER_174_485 ();
 b15zdnd11an1n04x5 FILLER_174_496 ();
 b15zdnd11an1n08x5 FILLER_174_542 ();
 b15zdnd11an1n04x5 FILLER_174_550 ();
 b15zdnd11an1n64x5 FILLER_174_596 ();
 b15zdnd11an1n32x5 FILLER_174_660 ();
 b15zdnd11an1n16x5 FILLER_174_692 ();
 b15zdnd11an1n08x5 FILLER_174_708 ();
 b15zdnd00an1n02x5 FILLER_174_716 ();
 b15zdnd11an1n64x5 FILLER_174_726 ();
 b15zdnd11an1n64x5 FILLER_174_790 ();
 b15zdnd11an1n64x5 FILLER_174_854 ();
 b15zdnd11an1n64x5 FILLER_174_918 ();
 b15zdnd11an1n64x5 FILLER_174_982 ();
 b15zdnd11an1n64x5 FILLER_174_1046 ();
 b15zdnd11an1n64x5 FILLER_174_1110 ();
 b15zdnd11an1n64x5 FILLER_174_1174 ();
 b15zdnd11an1n64x5 FILLER_174_1238 ();
 b15zdnd11an1n64x5 FILLER_174_1302 ();
 b15zdnd11an1n64x5 FILLER_174_1366 ();
 b15zdnd11an1n64x5 FILLER_174_1430 ();
 b15zdnd11an1n32x5 FILLER_174_1494 ();
 b15zdnd11an1n16x5 FILLER_174_1526 ();
 b15zdnd11an1n04x5 FILLER_174_1542 ();
 b15zdnd00an1n02x5 FILLER_174_1546 ();
 b15zdnd00an1n01x5 FILLER_174_1548 ();
 b15zdnd11an1n64x5 FILLER_174_1552 ();
 b15zdnd11an1n32x5 FILLER_174_1616 ();
 b15zdnd11an1n16x5 FILLER_174_1648 ();
 b15zdnd11an1n08x5 FILLER_174_1664 ();
 b15zdnd00an1n02x5 FILLER_174_1672 ();
 b15zdnd11an1n64x5 FILLER_174_1726 ();
 b15zdnd11an1n64x5 FILLER_174_1790 ();
 b15zdnd11an1n64x5 FILLER_174_1854 ();
 b15zdnd11an1n32x5 FILLER_174_1918 ();
 b15zdnd11an1n08x5 FILLER_174_1950 ();
 b15zdnd11an1n04x5 FILLER_174_1958 ();
 b15zdnd00an1n02x5 FILLER_174_1962 ();
 b15zdnd11an1n64x5 FILLER_174_2006 ();
 b15zdnd11an1n08x5 FILLER_174_2070 ();
 b15zdnd11an1n04x5 FILLER_174_2078 ();
 b15zdnd00an1n01x5 FILLER_174_2082 ();
 b15zdnd11an1n16x5 FILLER_174_2125 ();
 b15zdnd11an1n08x5 FILLER_174_2141 ();
 b15zdnd11an1n04x5 FILLER_174_2149 ();
 b15zdnd00an1n01x5 FILLER_174_2153 ();
 b15zdnd11an1n64x5 FILLER_174_2162 ();
 b15zdnd11an1n04x5 FILLER_174_2226 ();
 b15zdnd00an1n02x5 FILLER_174_2230 ();
 b15zdnd00an1n02x5 FILLER_174_2274 ();
 b15zdnd11an1n64x5 FILLER_175_0 ();
 b15zdnd11an1n64x5 FILLER_175_64 ();
 b15zdnd11an1n64x5 FILLER_175_128 ();
 b15zdnd11an1n32x5 FILLER_175_192 ();
 b15zdnd11an1n16x5 FILLER_175_224 ();
 b15zdnd00an1n01x5 FILLER_175_240 ();
 b15zdnd11an1n64x5 FILLER_175_283 ();
 b15zdnd11an1n16x5 FILLER_175_347 ();
 b15zdnd11an1n04x5 FILLER_175_366 ();
 b15zdnd11an1n04x5 FILLER_175_373 ();
 b15zdnd11an1n32x5 FILLER_175_380 ();
 b15zdnd11an1n16x5 FILLER_175_412 ();
 b15zdnd00an1n02x5 FILLER_175_428 ();
 b15zdnd00an1n01x5 FILLER_175_430 ();
 b15zdnd11an1n08x5 FILLER_175_473 ();
 b15zdnd00an1n01x5 FILLER_175_481 ();
 b15zdnd11an1n04x5 FILLER_175_490 ();
 b15zdnd11an1n04x5 FILLER_175_502 ();
 b15zdnd11an1n08x5 FILLER_175_513 ();
 b15zdnd11an1n04x5 FILLER_175_521 ();
 b15zdnd11an1n04x5 FILLER_175_535 ();
 b15zdnd11an1n04x5 FILLER_175_553 ();
 b15zdnd11an1n32x5 FILLER_175_563 ();
 b15zdnd11an1n08x5 FILLER_175_595 ();
 b15zdnd11an1n04x5 FILLER_175_603 ();
 b15zdnd00an1n01x5 FILLER_175_607 ();
 b15zdnd11an1n08x5 FILLER_175_615 ();
 b15zdnd11an1n04x5 FILLER_175_623 ();
 b15zdnd11an1n64x5 FILLER_175_636 ();
 b15zdnd11an1n64x5 FILLER_175_700 ();
 b15zdnd11an1n64x5 FILLER_175_764 ();
 b15zdnd11an1n64x5 FILLER_175_828 ();
 b15zdnd11an1n64x5 FILLER_175_892 ();
 b15zdnd11an1n32x5 FILLER_175_956 ();
 b15zdnd11an1n16x5 FILLER_175_988 ();
 b15zdnd00an1n01x5 FILLER_175_1004 ();
 b15zdnd11an1n64x5 FILLER_175_1050 ();
 b15zdnd11an1n64x5 FILLER_175_1114 ();
 b15zdnd11an1n64x5 FILLER_175_1178 ();
 b15zdnd11an1n64x5 FILLER_175_1242 ();
 b15zdnd11an1n64x5 FILLER_175_1306 ();
 b15zdnd11an1n64x5 FILLER_175_1370 ();
 b15zdnd11an1n64x5 FILLER_175_1434 ();
 b15zdnd11an1n16x5 FILLER_175_1498 ();
 b15zdnd11an1n08x5 FILLER_175_1514 ();
 b15zdnd00an1n02x5 FILLER_175_1522 ();
 b15zdnd11an1n32x5 FILLER_175_1576 ();
 b15zdnd11an1n08x5 FILLER_175_1608 ();
 b15zdnd11an1n04x5 FILLER_175_1616 ();
 b15zdnd11an1n04x5 FILLER_175_1623 ();
 b15zdnd11an1n32x5 FILLER_175_1630 ();
 b15zdnd11an1n08x5 FILLER_175_1662 ();
 b15zdnd11an1n04x5 FILLER_175_1670 ();
 b15zdnd00an1n02x5 FILLER_175_1674 ();
 b15zdnd11an1n04x5 FILLER_175_1696 ();
 b15zdnd11an1n04x5 FILLER_175_1703 ();
 b15zdnd11an1n64x5 FILLER_175_1710 ();
 b15zdnd11an1n64x5 FILLER_175_1774 ();
 b15zdnd11an1n64x5 FILLER_175_1838 ();
 b15zdnd11an1n64x5 FILLER_175_1902 ();
 b15zdnd11an1n64x5 FILLER_175_1966 ();
 b15zdnd11an1n16x5 FILLER_175_2030 ();
 b15zdnd11an1n08x5 FILLER_175_2046 ();
 b15zdnd11an1n64x5 FILLER_175_2096 ();
 b15zdnd11an1n64x5 FILLER_175_2160 ();
 b15zdnd11an1n16x5 FILLER_175_2224 ();
 b15zdnd00an1n02x5 FILLER_175_2282 ();
 b15zdnd11an1n64x5 FILLER_176_8 ();
 b15zdnd11an1n64x5 FILLER_176_72 ();
 b15zdnd11an1n64x5 FILLER_176_136 ();
 b15zdnd11an1n64x5 FILLER_176_200 ();
 b15zdnd11an1n64x5 FILLER_176_264 ();
 b15zdnd11an1n32x5 FILLER_176_328 ();
 b15zdnd11an1n08x5 FILLER_176_360 ();
 b15zdnd11an1n04x5 FILLER_176_368 ();
 b15zdnd00an1n01x5 FILLER_176_372 ();
 b15zdnd11an1n64x5 FILLER_176_425 ();
 b15zdnd11an1n64x5 FILLER_176_489 ();
 b15zdnd11an1n64x5 FILLER_176_553 ();
 b15zdnd11an1n16x5 FILLER_176_617 ();
 b15zdnd11an1n04x5 FILLER_176_633 ();
 b15zdnd00an1n02x5 FILLER_176_637 ();
 b15zdnd00an1n01x5 FILLER_176_639 ();
 b15zdnd11an1n32x5 FILLER_176_660 ();
 b15zdnd11an1n16x5 FILLER_176_692 ();
 b15zdnd11an1n08x5 FILLER_176_708 ();
 b15zdnd00an1n02x5 FILLER_176_716 ();
 b15zdnd11an1n64x5 FILLER_176_726 ();
 b15zdnd11an1n64x5 FILLER_176_790 ();
 b15zdnd11an1n64x5 FILLER_176_854 ();
 b15zdnd00an1n02x5 FILLER_176_918 ();
 b15zdnd11an1n16x5 FILLER_176_936 ();
 b15zdnd11an1n08x5 FILLER_176_952 ();
 b15zdnd11an1n32x5 FILLER_176_971 ();
 b15zdnd11an1n16x5 FILLER_176_1003 ();
 b15zdnd11an1n04x5 FILLER_176_1019 ();
 b15zdnd00an1n01x5 FILLER_176_1023 ();
 b15zdnd11an1n64x5 FILLER_176_1035 ();
 b15zdnd11an1n64x5 FILLER_176_1099 ();
 b15zdnd11an1n64x5 FILLER_176_1163 ();
 b15zdnd11an1n16x5 FILLER_176_1227 ();
 b15zdnd11an1n08x5 FILLER_176_1243 ();
 b15zdnd11an1n04x5 FILLER_176_1251 ();
 b15zdnd00an1n02x5 FILLER_176_1255 ();
 b15zdnd11an1n04x5 FILLER_176_1273 ();
 b15zdnd11an1n64x5 FILLER_176_1293 ();
 b15zdnd11an1n64x5 FILLER_176_1357 ();
 b15zdnd11an1n64x5 FILLER_176_1421 ();
 b15zdnd11an1n64x5 FILLER_176_1485 ();
 b15zdnd11an1n32x5 FILLER_176_1552 ();
 b15zdnd11an1n16x5 FILLER_176_1584 ();
 b15zdnd00an1n02x5 FILLER_176_1600 ();
 b15zdnd11an1n16x5 FILLER_176_1654 ();
 b15zdnd11an1n08x5 FILLER_176_1670 ();
 b15zdnd00an1n01x5 FILLER_176_1678 ();
 b15zdnd11an1n64x5 FILLER_176_1699 ();
 b15zdnd11an1n64x5 FILLER_176_1763 ();
 b15zdnd11an1n64x5 FILLER_176_1827 ();
 b15zdnd11an1n64x5 FILLER_176_1891 ();
 b15zdnd11an1n64x5 FILLER_176_1955 ();
 b15zdnd11an1n64x5 FILLER_176_2019 ();
 b15zdnd11an1n04x5 FILLER_176_2083 ();
 b15zdnd00an1n02x5 FILLER_176_2087 ();
 b15zdnd00an1n01x5 FILLER_176_2089 ();
 b15zdnd11an1n16x5 FILLER_176_2132 ();
 b15zdnd11an1n04x5 FILLER_176_2148 ();
 b15zdnd00an1n02x5 FILLER_176_2152 ();
 b15zdnd11an1n64x5 FILLER_176_2162 ();
 b15zdnd11an1n04x5 FILLER_176_2226 ();
 b15zdnd00an1n02x5 FILLER_176_2230 ();
 b15zdnd00an1n02x5 FILLER_176_2274 ();
 b15zdnd11an1n64x5 FILLER_177_0 ();
 b15zdnd11an1n64x5 FILLER_177_64 ();
 b15zdnd11an1n64x5 FILLER_177_128 ();
 b15zdnd11an1n32x5 FILLER_177_192 ();
 b15zdnd11an1n16x5 FILLER_177_224 ();
 b15zdnd00an1n02x5 FILLER_177_240 ();
 b15zdnd11an1n64x5 FILLER_177_251 ();
 b15zdnd11an1n64x5 FILLER_177_315 ();
 b15zdnd11an1n04x5 FILLER_177_379 ();
 b15zdnd00an1n01x5 FILLER_177_383 ();
 b15zdnd11an1n08x5 FILLER_177_387 ();
 b15zdnd00an1n02x5 FILLER_177_395 ();
 b15zdnd00an1n01x5 FILLER_177_397 ();
 b15zdnd11an1n64x5 FILLER_177_401 ();
 b15zdnd11an1n64x5 FILLER_177_465 ();
 b15zdnd11an1n64x5 FILLER_177_529 ();
 b15zdnd11an1n64x5 FILLER_177_593 ();
 b15zdnd11an1n64x5 FILLER_177_657 ();
 b15zdnd11an1n64x5 FILLER_177_721 ();
 b15zdnd11an1n64x5 FILLER_177_785 ();
 b15zdnd11an1n64x5 FILLER_177_849 ();
 b15zdnd11an1n32x5 FILLER_177_913 ();
 b15zdnd00an1n02x5 FILLER_177_945 ();
 b15zdnd11an1n32x5 FILLER_177_978 ();
 b15zdnd00an1n02x5 FILLER_177_1010 ();
 b15zdnd00an1n01x5 FILLER_177_1012 ();
 b15zdnd11an1n64x5 FILLER_177_1021 ();
 b15zdnd11an1n64x5 FILLER_177_1085 ();
 b15zdnd11an1n64x5 FILLER_177_1149 ();
 b15zdnd11an1n16x5 FILLER_177_1213 ();
 b15zdnd11an1n04x5 FILLER_177_1229 ();
 b15zdnd00an1n02x5 FILLER_177_1233 ();
 b15zdnd11an1n16x5 FILLER_177_1247 ();
 b15zdnd11an1n64x5 FILLER_177_1287 ();
 b15zdnd11an1n64x5 FILLER_177_1351 ();
 b15zdnd11an1n64x5 FILLER_177_1415 ();
 b15zdnd11an1n64x5 FILLER_177_1479 ();
 b15zdnd11an1n64x5 FILLER_177_1543 ();
 b15zdnd11an1n08x5 FILLER_177_1607 ();
 b15zdnd11an1n04x5 FILLER_177_1615 ();
 b15zdnd00an1n01x5 FILLER_177_1619 ();
 b15zdnd11an1n64x5 FILLER_177_1623 ();
 b15zdnd11an1n64x5 FILLER_177_1687 ();
 b15zdnd11an1n64x5 FILLER_177_1751 ();
 b15zdnd11an1n64x5 FILLER_177_1815 ();
 b15zdnd11an1n64x5 FILLER_177_1879 ();
 b15zdnd11an1n64x5 FILLER_177_1943 ();
 b15zdnd11an1n64x5 FILLER_177_2007 ();
 b15zdnd11an1n64x5 FILLER_177_2071 ();
 b15zdnd11an1n64x5 FILLER_177_2135 ();
 b15zdnd11an1n32x5 FILLER_177_2199 ();
 b15zdnd11an1n08x5 FILLER_177_2231 ();
 b15zdnd00an1n01x5 FILLER_177_2239 ();
 b15zdnd00an1n02x5 FILLER_177_2282 ();
 b15zdnd11an1n64x5 FILLER_178_8 ();
 b15zdnd11an1n16x5 FILLER_178_72 ();
 b15zdnd11an1n08x5 FILLER_178_88 ();
 b15zdnd00an1n02x5 FILLER_178_96 ();
 b15zdnd00an1n01x5 FILLER_178_98 ();
 b15zdnd11an1n64x5 FILLER_178_108 ();
 b15zdnd11an1n64x5 FILLER_178_172 ();
 b15zdnd11an1n08x5 FILLER_178_236 ();
 b15zdnd11an1n04x5 FILLER_178_244 ();
 b15zdnd00an1n02x5 FILLER_178_248 ();
 b15zdnd11an1n64x5 FILLER_178_261 ();
 b15zdnd11an1n64x5 FILLER_178_325 ();
 b15zdnd11an1n08x5 FILLER_178_389 ();
 b15zdnd00an1n01x5 FILLER_178_397 ();
 b15zdnd11an1n64x5 FILLER_178_401 ();
 b15zdnd11an1n64x5 FILLER_178_465 ();
 b15zdnd11an1n64x5 FILLER_178_529 ();
 b15zdnd11an1n32x5 FILLER_178_593 ();
 b15zdnd00an1n02x5 FILLER_178_625 ();
 b15zdnd11an1n64x5 FILLER_178_636 ();
 b15zdnd11an1n16x5 FILLER_178_700 ();
 b15zdnd00an1n02x5 FILLER_178_716 ();
 b15zdnd11an1n64x5 FILLER_178_726 ();
 b15zdnd11an1n64x5 FILLER_178_790 ();
 b15zdnd11an1n64x5 FILLER_178_854 ();
 b15zdnd11an1n08x5 FILLER_178_918 ();
 b15zdnd11an1n04x5 FILLER_178_926 ();
 b15zdnd00an1n02x5 FILLER_178_930 ();
 b15zdnd11an1n64x5 FILLER_178_977 ();
 b15zdnd11an1n64x5 FILLER_178_1041 ();
 b15zdnd11an1n64x5 FILLER_178_1105 ();
 b15zdnd11an1n64x5 FILLER_178_1169 ();
 b15zdnd11an1n08x5 FILLER_178_1233 ();
 b15zdnd11an1n04x5 FILLER_178_1241 ();
 b15zdnd00an1n02x5 FILLER_178_1245 ();
 b15zdnd00an1n01x5 FILLER_178_1247 ();
 b15zdnd11an1n64x5 FILLER_178_1272 ();
 b15zdnd11an1n64x5 FILLER_178_1336 ();
 b15zdnd11an1n64x5 FILLER_178_1400 ();
 b15zdnd11an1n64x5 FILLER_178_1464 ();
 b15zdnd11an1n64x5 FILLER_178_1528 ();
 b15zdnd11an1n64x5 FILLER_178_1592 ();
 b15zdnd11an1n64x5 FILLER_178_1656 ();
 b15zdnd11an1n64x5 FILLER_178_1720 ();
 b15zdnd11an1n64x5 FILLER_178_1784 ();
 b15zdnd11an1n64x5 FILLER_178_1848 ();
 b15zdnd11an1n64x5 FILLER_178_1912 ();
 b15zdnd11an1n64x5 FILLER_178_1976 ();
 b15zdnd11an1n64x5 FILLER_178_2040 ();
 b15zdnd11an1n32x5 FILLER_178_2104 ();
 b15zdnd11an1n16x5 FILLER_178_2136 ();
 b15zdnd00an1n02x5 FILLER_178_2152 ();
 b15zdnd11an1n64x5 FILLER_178_2162 ();
 b15zdnd11an1n04x5 FILLER_178_2226 ();
 b15zdnd00an1n02x5 FILLER_178_2230 ();
 b15zdnd00an1n02x5 FILLER_178_2274 ();
 b15zdnd11an1n64x5 FILLER_179_0 ();
 b15zdnd11an1n64x5 FILLER_179_64 ();
 b15zdnd11an1n64x5 FILLER_179_128 ();
 b15zdnd11an1n64x5 FILLER_179_192 ();
 b15zdnd11an1n04x5 FILLER_179_256 ();
 b15zdnd00an1n02x5 FILLER_179_260 ();
 b15zdnd11an1n64x5 FILLER_179_276 ();
 b15zdnd11an1n64x5 FILLER_179_340 ();
 b15zdnd11an1n64x5 FILLER_179_404 ();
 b15zdnd11an1n64x5 FILLER_179_468 ();
 b15zdnd11an1n16x5 FILLER_179_532 ();
 b15zdnd00an1n01x5 FILLER_179_548 ();
 b15zdnd11an1n64x5 FILLER_179_556 ();
 b15zdnd11an1n64x5 FILLER_179_620 ();
 b15zdnd11an1n64x5 FILLER_179_684 ();
 b15zdnd11an1n64x5 FILLER_179_748 ();
 b15zdnd11an1n64x5 FILLER_179_812 ();
 b15zdnd11an1n64x5 FILLER_179_876 ();
 b15zdnd11an1n64x5 FILLER_179_940 ();
 b15zdnd11an1n64x5 FILLER_179_1004 ();
 b15zdnd11an1n64x5 FILLER_179_1068 ();
 b15zdnd11an1n08x5 FILLER_179_1132 ();
 b15zdnd11an1n04x5 FILLER_179_1140 ();
 b15zdnd00an1n01x5 FILLER_179_1144 ();
 b15zdnd11an1n32x5 FILLER_179_1148 ();
 b15zdnd11an1n16x5 FILLER_179_1180 ();
 b15zdnd00an1n01x5 FILLER_179_1196 ();
 b15zdnd11an1n16x5 FILLER_179_1217 ();
 b15zdnd11an1n08x5 FILLER_179_1233 ();
 b15zdnd00an1n01x5 FILLER_179_1241 ();
 b15zdnd11an1n08x5 FILLER_179_1262 ();
 b15zdnd11an1n04x5 FILLER_179_1270 ();
 b15zdnd11an1n64x5 FILLER_179_1284 ();
 b15zdnd11an1n32x5 FILLER_179_1348 ();
 b15zdnd11an1n16x5 FILLER_179_1380 ();
 b15zdnd11an1n08x5 FILLER_179_1396 ();
 b15zdnd11an1n04x5 FILLER_179_1404 ();
 b15zdnd00an1n01x5 FILLER_179_1408 ();
 b15zdnd11an1n64x5 FILLER_179_1418 ();
 b15zdnd11an1n64x5 FILLER_179_1482 ();
 b15zdnd11an1n64x5 FILLER_179_1546 ();
 b15zdnd11an1n64x5 FILLER_179_1610 ();
 b15zdnd11an1n64x5 FILLER_179_1674 ();
 b15zdnd11an1n64x5 FILLER_179_1738 ();
 b15zdnd11an1n64x5 FILLER_179_1802 ();
 b15zdnd11an1n32x5 FILLER_179_1866 ();
 b15zdnd11an1n04x5 FILLER_179_1898 ();
 b15zdnd00an1n02x5 FILLER_179_1902 ();
 b15zdnd00an1n01x5 FILLER_179_1904 ();
 b15zdnd11an1n64x5 FILLER_179_1908 ();
 b15zdnd11an1n64x5 FILLER_179_1972 ();
 b15zdnd11an1n64x5 FILLER_179_2036 ();
 b15zdnd11an1n64x5 FILLER_179_2100 ();
 b15zdnd11an1n32x5 FILLER_179_2164 ();
 b15zdnd11an1n08x5 FILLER_179_2196 ();
 b15zdnd00an1n02x5 FILLER_179_2204 ();
 b15zdnd11an1n16x5 FILLER_179_2209 ();
 b15zdnd11an1n04x5 FILLER_179_2225 ();
 b15zdnd00an1n02x5 FILLER_179_2229 ();
 b15zdnd00an1n01x5 FILLER_179_2231 ();
 b15zdnd11an1n04x5 FILLER_179_2236 ();
 b15zdnd00an1n02x5 FILLER_179_2282 ();
 b15zdnd11an1n64x5 FILLER_180_8 ();
 b15zdnd11an1n64x5 FILLER_180_72 ();
 b15zdnd11an1n08x5 FILLER_180_136 ();
 b15zdnd00an1n02x5 FILLER_180_144 ();
 b15zdnd11an1n64x5 FILLER_180_149 ();
 b15zdnd11an1n32x5 FILLER_180_213 ();
 b15zdnd11an1n04x5 FILLER_180_245 ();
 b15zdnd00an1n02x5 FILLER_180_249 ();
 b15zdnd00an1n01x5 FILLER_180_251 ();
 b15zdnd11an1n64x5 FILLER_180_266 ();
 b15zdnd11an1n64x5 FILLER_180_330 ();
 b15zdnd11an1n64x5 FILLER_180_394 ();
 b15zdnd11an1n32x5 FILLER_180_458 ();
 b15zdnd11an1n16x5 FILLER_180_490 ();
 b15zdnd11an1n08x5 FILLER_180_506 ();
 b15zdnd00an1n01x5 FILLER_180_514 ();
 b15zdnd11an1n08x5 FILLER_180_523 ();
 b15zdnd11an1n04x5 FILLER_180_531 ();
 b15zdnd00an1n02x5 FILLER_180_535 ();
 b15zdnd11an1n64x5 FILLER_180_545 ();
 b15zdnd11an1n64x5 FILLER_180_609 ();
 b15zdnd11an1n32x5 FILLER_180_673 ();
 b15zdnd11an1n08x5 FILLER_180_705 ();
 b15zdnd11an1n04x5 FILLER_180_713 ();
 b15zdnd00an1n01x5 FILLER_180_717 ();
 b15zdnd11an1n64x5 FILLER_180_726 ();
 b15zdnd11an1n64x5 FILLER_180_790 ();
 b15zdnd11an1n04x5 FILLER_180_854 ();
 b15zdnd11an1n64x5 FILLER_180_861 ();
 b15zdnd11an1n64x5 FILLER_180_925 ();
 b15zdnd11an1n16x5 FILLER_180_989 ();
 b15zdnd11an1n08x5 FILLER_180_1005 ();
 b15zdnd00an1n01x5 FILLER_180_1013 ();
 b15zdnd11an1n08x5 FILLER_180_1029 ();
 b15zdnd11an1n04x5 FILLER_180_1037 ();
 b15zdnd11an1n04x5 FILLER_180_1044 ();
 b15zdnd11an1n64x5 FILLER_180_1051 ();
 b15zdnd11an1n16x5 FILLER_180_1115 ();
 b15zdnd11an1n08x5 FILLER_180_1131 ();
 b15zdnd11an1n04x5 FILLER_180_1139 ();
 b15zdnd00an1n02x5 FILLER_180_1143 ();
 b15zdnd11an1n04x5 FILLER_180_1148 ();
 b15zdnd11an1n64x5 FILLER_180_1155 ();
 b15zdnd11an1n32x5 FILLER_180_1219 ();
 b15zdnd11an1n04x5 FILLER_180_1251 ();
 b15zdnd11an1n64x5 FILLER_180_1275 ();
 b15zdnd11an1n64x5 FILLER_180_1339 ();
 b15zdnd11an1n64x5 FILLER_180_1403 ();
 b15zdnd11an1n64x5 FILLER_180_1467 ();
 b15zdnd11an1n64x5 FILLER_180_1531 ();
 b15zdnd11an1n64x5 FILLER_180_1595 ();
 b15zdnd11an1n64x5 FILLER_180_1659 ();
 b15zdnd11an1n64x5 FILLER_180_1723 ();
 b15zdnd11an1n04x5 FILLER_180_1787 ();
 b15zdnd00an1n02x5 FILLER_180_1791 ();
 b15zdnd11an1n04x5 FILLER_180_1796 ();
 b15zdnd11an1n64x5 FILLER_180_1803 ();
 b15zdnd11an1n08x5 FILLER_180_1867 ();
 b15zdnd11an1n04x5 FILLER_180_1875 ();
 b15zdnd11an1n04x5 FILLER_180_1931 ();
 b15zdnd00an1n01x5 FILLER_180_1935 ();
 b15zdnd11an1n04x5 FILLER_180_1939 ();
 b15zdnd11an1n64x5 FILLER_180_1946 ();
 b15zdnd11an1n64x5 FILLER_180_2010 ();
 b15zdnd11an1n64x5 FILLER_180_2074 ();
 b15zdnd11an1n16x5 FILLER_180_2138 ();
 b15zdnd11an1n32x5 FILLER_180_2162 ();
 b15zdnd11an1n08x5 FILLER_180_2194 ();
 b15zdnd11an1n04x5 FILLER_180_2202 ();
 b15zdnd11an1n04x5 FILLER_180_2209 ();
 b15zdnd11an1n04x5 FILLER_180_2216 ();
 b15zdnd00an1n02x5 FILLER_180_2220 ();
 b15zdnd11an1n04x5 FILLER_180_2264 ();
 b15zdnd11an1n04x5 FILLER_180_2272 ();
 b15zdnd11an1n64x5 FILLER_181_0 ();
 b15zdnd11an1n04x5 FILLER_181_64 ();
 b15zdnd00an1n02x5 FILLER_181_68 ();
 b15zdnd00an1n01x5 FILLER_181_70 ();
 b15zdnd11an1n04x5 FILLER_181_74 ();
 b15zdnd11an1n32x5 FILLER_181_81 ();
 b15zdnd11an1n04x5 FILLER_181_113 ();
 b15zdnd00an1n02x5 FILLER_181_117 ();
 b15zdnd11an1n32x5 FILLER_181_171 ();
 b15zdnd11an1n16x5 FILLER_181_203 ();
 b15zdnd11an1n08x5 FILLER_181_219 ();
 b15zdnd00an1n02x5 FILLER_181_227 ();
 b15zdnd00an1n01x5 FILLER_181_229 ();
 b15zdnd11an1n04x5 FILLER_181_233 ();
 b15zdnd11an1n04x5 FILLER_181_264 ();
 b15zdnd11an1n64x5 FILLER_181_310 ();
 b15zdnd11an1n64x5 FILLER_181_374 ();
 b15zdnd11an1n64x5 FILLER_181_438 ();
 b15zdnd11an1n64x5 FILLER_181_502 ();
 b15zdnd11an1n08x5 FILLER_181_566 ();
 b15zdnd00an1n01x5 FILLER_181_574 ();
 b15zdnd11an1n64x5 FILLER_181_617 ();
 b15zdnd11an1n64x5 FILLER_181_681 ();
 b15zdnd11an1n64x5 FILLER_181_745 ();
 b15zdnd11an1n64x5 FILLER_181_809 ();
 b15zdnd11an1n64x5 FILLER_181_873 ();
 b15zdnd11an1n64x5 FILLER_181_937 ();
 b15zdnd11an1n04x5 FILLER_181_1001 ();
 b15zdnd00an1n02x5 FILLER_181_1005 ();
 b15zdnd11an1n04x5 FILLER_181_1018 ();
 b15zdnd11an1n32x5 FILLER_181_1074 ();
 b15zdnd11an1n16x5 FILLER_181_1106 ();
 b15zdnd00an1n02x5 FILLER_181_1122 ();
 b15zdnd00an1n01x5 FILLER_181_1124 ();
 b15zdnd11an1n32x5 FILLER_181_1177 ();
 b15zdnd11an1n16x5 FILLER_181_1209 ();
 b15zdnd11an1n08x5 FILLER_181_1225 ();
 b15zdnd11an1n04x5 FILLER_181_1233 ();
 b15zdnd00an1n01x5 FILLER_181_1237 ();
 b15zdnd11an1n04x5 FILLER_181_1252 ();
 b15zdnd11an1n64x5 FILLER_181_1276 ();
 b15zdnd11an1n64x5 FILLER_181_1340 ();
 b15zdnd11an1n64x5 FILLER_181_1404 ();
 b15zdnd11an1n64x5 FILLER_181_1468 ();
 b15zdnd11an1n64x5 FILLER_181_1532 ();
 b15zdnd11an1n64x5 FILLER_181_1596 ();
 b15zdnd11an1n64x5 FILLER_181_1660 ();
 b15zdnd11an1n32x5 FILLER_181_1724 ();
 b15zdnd11an1n16x5 FILLER_181_1756 ();
 b15zdnd00an1n02x5 FILLER_181_1772 ();
 b15zdnd00an1n01x5 FILLER_181_1774 ();
 b15zdnd11an1n64x5 FILLER_181_1827 ();
 b15zdnd11an1n08x5 FILLER_181_1891 ();
 b15zdnd11an1n04x5 FILLER_181_1899 ();
 b15zdnd00an1n01x5 FILLER_181_1903 ();
 b15zdnd11an1n04x5 FILLER_181_1907 ();
 b15zdnd11an1n04x5 FILLER_181_1914 ();
 b15zdnd11an1n64x5 FILLER_181_1970 ();
 b15zdnd11an1n16x5 FILLER_181_2034 ();
 b15zdnd11an1n08x5 FILLER_181_2050 ();
 b15zdnd00an1n02x5 FILLER_181_2058 ();
 b15zdnd11an1n64x5 FILLER_181_2102 ();
 b15zdnd11an1n08x5 FILLER_181_2166 ();
 b15zdnd11an1n04x5 FILLER_181_2174 ();
 b15zdnd00an1n02x5 FILLER_181_2178 ();
 b15zdnd11an1n04x5 FILLER_181_2232 ();
 b15zdnd00an1n02x5 FILLER_181_2236 ();
 b15zdnd00an1n01x5 FILLER_181_2238 ();
 b15zdnd00an1n02x5 FILLER_181_2281 ();
 b15zdnd00an1n01x5 FILLER_181_2283 ();
 b15zdnd11an1n32x5 FILLER_182_8 ();
 b15zdnd11an1n16x5 FILLER_182_40 ();
 b15zdnd11an1n08x5 FILLER_182_56 ();
 b15zdnd11an1n04x5 FILLER_182_67 ();
 b15zdnd11an1n04x5 FILLER_182_80 ();
 b15zdnd11an1n32x5 FILLER_182_87 ();
 b15zdnd11an1n16x5 FILLER_182_119 ();
 b15zdnd00an1n02x5 FILLER_182_135 ();
 b15zdnd00an1n01x5 FILLER_182_137 ();
 b15zdnd11an1n04x5 FILLER_182_141 ();
 b15zdnd11an1n64x5 FILLER_182_148 ();
 b15zdnd11an1n64x5 FILLER_182_212 ();
 b15zdnd11an1n64x5 FILLER_182_276 ();
 b15zdnd11an1n64x5 FILLER_182_340 ();
 b15zdnd11an1n64x5 FILLER_182_404 ();
 b15zdnd11an1n08x5 FILLER_182_468 ();
 b15zdnd00an1n02x5 FILLER_182_476 ();
 b15zdnd00an1n01x5 FILLER_182_478 ();
 b15zdnd11an1n04x5 FILLER_182_521 ();
 b15zdnd11an1n16x5 FILLER_182_567 ();
 b15zdnd11an1n08x5 FILLER_182_583 ();
 b15zdnd00an1n02x5 FILLER_182_591 ();
 b15zdnd00an1n01x5 FILLER_182_593 ();
 b15zdnd11an1n64x5 FILLER_182_636 ();
 b15zdnd11an1n16x5 FILLER_182_700 ();
 b15zdnd00an1n02x5 FILLER_182_716 ();
 b15zdnd11an1n32x5 FILLER_182_726 ();
 b15zdnd11an1n16x5 FILLER_182_758 ();
 b15zdnd11an1n04x5 FILLER_182_774 ();
 b15zdnd00an1n02x5 FILLER_182_778 ();
 b15zdnd11an1n64x5 FILLER_182_792 ();
 b15zdnd11an1n64x5 FILLER_182_856 ();
 b15zdnd11an1n64x5 FILLER_182_920 ();
 b15zdnd11an1n16x5 FILLER_182_984 ();
 b15zdnd11an1n08x5 FILLER_182_1000 ();
 b15zdnd11an1n08x5 FILLER_182_1019 ();
 b15zdnd11an1n04x5 FILLER_182_1027 ();
 b15zdnd00an1n02x5 FILLER_182_1031 ();
 b15zdnd11an1n16x5 FILLER_182_1085 ();
 b15zdnd11an1n08x5 FILLER_182_1101 ();
 b15zdnd00an1n01x5 FILLER_182_1109 ();
 b15zdnd11an1n64x5 FILLER_182_1162 ();
 b15zdnd11an1n64x5 FILLER_182_1226 ();
 b15zdnd11an1n64x5 FILLER_182_1290 ();
 b15zdnd11an1n64x5 FILLER_182_1354 ();
 b15zdnd11an1n64x5 FILLER_182_1418 ();
 b15zdnd11an1n64x5 FILLER_182_1482 ();
 b15zdnd11an1n64x5 FILLER_182_1546 ();
 b15zdnd11an1n64x5 FILLER_182_1610 ();
 b15zdnd11an1n64x5 FILLER_182_1674 ();
 b15zdnd11an1n32x5 FILLER_182_1738 ();
 b15zdnd11an1n04x5 FILLER_182_1770 ();
 b15zdnd11an1n64x5 FILLER_182_1826 ();
 b15zdnd00an1n01x5 FILLER_182_1890 ();
 b15zdnd11an1n32x5 FILLER_182_1894 ();
 b15zdnd11an1n16x5 FILLER_182_1926 ();
 b15zdnd00an1n01x5 FILLER_182_1942 ();
 b15zdnd11an1n64x5 FILLER_182_1946 ();
 b15zdnd11an1n64x5 FILLER_182_2010 ();
 b15zdnd11an1n08x5 FILLER_182_2074 ();
 b15zdnd11an1n04x5 FILLER_182_2082 ();
 b15zdnd00an1n02x5 FILLER_182_2086 ();
 b15zdnd00an1n01x5 FILLER_182_2088 ();
 b15zdnd11an1n16x5 FILLER_182_2131 ();
 b15zdnd11an1n04x5 FILLER_182_2147 ();
 b15zdnd00an1n02x5 FILLER_182_2151 ();
 b15zdnd00an1n01x5 FILLER_182_2153 ();
 b15zdnd11an1n16x5 FILLER_182_2162 ();
 b15zdnd11an1n04x5 FILLER_182_2178 ();
 b15zdnd00an1n02x5 FILLER_182_2182 ();
 b15zdnd00an1n01x5 FILLER_182_2184 ();
 b15zdnd11an1n04x5 FILLER_182_2227 ();
 b15zdnd00an1n02x5 FILLER_182_2273 ();
 b15zdnd00an1n01x5 FILLER_182_2275 ();
 b15zdnd11an1n32x5 FILLER_183_0 ();
 b15zdnd11an1n16x5 FILLER_183_32 ();
 b15zdnd11an1n64x5 FILLER_183_100 ();
 b15zdnd11an1n32x5 FILLER_183_164 ();
 b15zdnd11an1n08x5 FILLER_183_196 ();
 b15zdnd11an1n04x5 FILLER_183_204 ();
 b15zdnd00an1n02x5 FILLER_183_208 ();
 b15zdnd11an1n64x5 FILLER_183_219 ();
 b15zdnd11an1n16x5 FILLER_183_283 ();
 b15zdnd11an1n08x5 FILLER_183_299 ();
 b15zdnd11an1n64x5 FILLER_183_349 ();
 b15zdnd11an1n64x5 FILLER_183_413 ();
 b15zdnd11an1n32x5 FILLER_183_477 ();
 b15zdnd11an1n16x5 FILLER_183_509 ();
 b15zdnd00an1n01x5 FILLER_183_525 ();
 b15zdnd11an1n64x5 FILLER_183_533 ();
 b15zdnd11an1n08x5 FILLER_183_597 ();
 b15zdnd00an1n01x5 FILLER_183_605 ();
 b15zdnd11an1n64x5 FILLER_183_658 ();
 b15zdnd11an1n32x5 FILLER_183_722 ();
 b15zdnd00an1n01x5 FILLER_183_754 ();
 b15zdnd11an1n64x5 FILLER_183_758 ();
 b15zdnd11an1n64x5 FILLER_183_822 ();
 b15zdnd11an1n04x5 FILLER_183_886 ();
 b15zdnd00an1n02x5 FILLER_183_890 ();
 b15zdnd00an1n01x5 FILLER_183_892 ();
 b15zdnd11an1n64x5 FILLER_183_909 ();
 b15zdnd11an1n64x5 FILLER_183_973 ();
 b15zdnd11an1n08x5 FILLER_183_1037 ();
 b15zdnd00an1n01x5 FILLER_183_1045 ();
 b15zdnd11an1n04x5 FILLER_183_1049 ();
 b15zdnd11an1n04x5 FILLER_183_1056 ();
 b15zdnd11an1n64x5 FILLER_183_1063 ();
 b15zdnd00an1n02x5 FILLER_183_1127 ();
 b15zdnd00an1n01x5 FILLER_183_1129 ();
 b15zdnd11an1n04x5 FILLER_183_1133 ();
 b15zdnd11an1n64x5 FILLER_183_1140 ();
 b15zdnd11an1n64x5 FILLER_183_1204 ();
 b15zdnd11an1n64x5 FILLER_183_1268 ();
 b15zdnd11an1n64x5 FILLER_183_1332 ();
 b15zdnd11an1n08x5 FILLER_183_1396 ();
 b15zdnd00an1n01x5 FILLER_183_1404 ();
 b15zdnd11an1n64x5 FILLER_183_1414 ();
 b15zdnd11an1n64x5 FILLER_183_1478 ();
 b15zdnd11an1n64x5 FILLER_183_1542 ();
 b15zdnd11an1n64x5 FILLER_183_1606 ();
 b15zdnd11an1n64x5 FILLER_183_1670 ();
 b15zdnd11an1n32x5 FILLER_183_1734 ();
 b15zdnd11an1n16x5 FILLER_183_1766 ();
 b15zdnd11an1n08x5 FILLER_183_1782 ();
 b15zdnd00an1n02x5 FILLER_183_1790 ();
 b15zdnd00an1n01x5 FILLER_183_1792 ();
 b15zdnd11an1n04x5 FILLER_183_1796 ();
 b15zdnd11an1n32x5 FILLER_183_1803 ();
 b15zdnd11an1n16x5 FILLER_183_1835 ();
 b15zdnd11an1n08x5 FILLER_183_1851 ();
 b15zdnd11an1n04x5 FILLER_183_1859 ();
 b15zdnd00an1n02x5 FILLER_183_1863 ();
 b15zdnd11an1n64x5 FILLER_183_1917 ();
 b15zdnd11an1n32x5 FILLER_183_1981 ();
 b15zdnd11an1n16x5 FILLER_183_2013 ();
 b15zdnd11an1n04x5 FILLER_183_2029 ();
 b15zdnd00an1n01x5 FILLER_183_2033 ();
 b15zdnd11an1n04x5 FILLER_183_2037 ();
 b15zdnd11an1n64x5 FILLER_183_2044 ();
 b15zdnd11an1n16x5 FILLER_183_2108 ();
 b15zdnd00an1n02x5 FILLER_183_2124 ();
 b15zdnd00an1n01x5 FILLER_183_2126 ();
 b15zdnd11an1n08x5 FILLER_183_2136 ();
 b15zdnd11an1n04x5 FILLER_183_2144 ();
 b15zdnd00an1n02x5 FILLER_183_2148 ();
 b15zdnd11an1n04x5 FILLER_183_2192 ();
 b15zdnd00an1n01x5 FILLER_183_2196 ();
 b15zdnd11an1n04x5 FILLER_183_2201 ();
 b15zdnd11an1n04x5 FILLER_183_2209 ();
 b15zdnd11an1n04x5 FILLER_183_2258 ();
 b15zdnd11an1n04x5 FILLER_183_2269 ();
 b15zdnd11an1n04x5 FILLER_183_2277 ();
 b15zdnd00an1n02x5 FILLER_183_2281 ();
 b15zdnd00an1n01x5 FILLER_183_2283 ();
 b15zdnd11an1n32x5 FILLER_184_8 ();
 b15zdnd11an1n04x5 FILLER_184_40 ();
 b15zdnd11an1n04x5 FILLER_184_47 ();
 b15zdnd11an1n08x5 FILLER_184_103 ();
 b15zdnd11an1n32x5 FILLER_184_120 ();
 b15zdnd11an1n08x5 FILLER_184_152 ();
 b15zdnd00an1n02x5 FILLER_184_160 ();
 b15zdnd00an1n01x5 FILLER_184_162 ();
 b15zdnd11an1n64x5 FILLER_184_190 ();
 b15zdnd11an1n64x5 FILLER_184_254 ();
 b15zdnd11an1n08x5 FILLER_184_318 ();
 b15zdnd11an1n04x5 FILLER_184_326 ();
 b15zdnd00an1n02x5 FILLER_184_330 ();
 b15zdnd00an1n01x5 FILLER_184_332 ();
 b15zdnd11an1n64x5 FILLER_184_375 ();
 b15zdnd11an1n32x5 FILLER_184_439 ();
 b15zdnd11an1n08x5 FILLER_184_471 ();
 b15zdnd00an1n02x5 FILLER_184_479 ();
 b15zdnd11an1n64x5 FILLER_184_489 ();
 b15zdnd11an1n64x5 FILLER_184_553 ();
 b15zdnd11an1n08x5 FILLER_184_617 ();
 b15zdnd00an1n01x5 FILLER_184_625 ();
 b15zdnd11an1n04x5 FILLER_184_629 ();
 b15zdnd11an1n64x5 FILLER_184_636 ();
 b15zdnd11an1n16x5 FILLER_184_700 ();
 b15zdnd00an1n02x5 FILLER_184_716 ();
 b15zdnd11an1n64x5 FILLER_184_726 ();
 b15zdnd11an1n32x5 FILLER_184_790 ();
 b15zdnd11an1n16x5 FILLER_184_822 ();
 b15zdnd11an1n08x5 FILLER_184_838 ();
 b15zdnd11an1n04x5 FILLER_184_846 ();
 b15zdnd11an1n64x5 FILLER_184_862 ();
 b15zdnd11an1n64x5 FILLER_184_926 ();
 b15zdnd11an1n64x5 FILLER_184_990 ();
 b15zdnd11an1n04x5 FILLER_184_1054 ();
 b15zdnd00an1n01x5 FILLER_184_1058 ();
 b15zdnd11an1n64x5 FILLER_184_1062 ();
 b15zdnd11an1n08x5 FILLER_184_1126 ();
 b15zdnd00an1n02x5 FILLER_184_1134 ();
 b15zdnd11an1n64x5 FILLER_184_1139 ();
 b15zdnd11an1n64x5 FILLER_184_1203 ();
 b15zdnd11an1n64x5 FILLER_184_1267 ();
 b15zdnd11an1n08x5 FILLER_184_1331 ();
 b15zdnd00an1n02x5 FILLER_184_1339 ();
 b15zdnd11an1n64x5 FILLER_184_1344 ();
 b15zdnd11an1n64x5 FILLER_184_1408 ();
 b15zdnd11an1n64x5 FILLER_184_1472 ();
 b15zdnd11an1n64x5 FILLER_184_1536 ();
 b15zdnd11an1n64x5 FILLER_184_1600 ();
 b15zdnd11an1n64x5 FILLER_184_1664 ();
 b15zdnd11an1n64x5 FILLER_184_1728 ();
 b15zdnd00an1n01x5 FILLER_184_1792 ();
 b15zdnd11an1n04x5 FILLER_184_1796 ();
 b15zdnd11an1n64x5 FILLER_184_1803 ();
 b15zdnd11an1n16x5 FILLER_184_1867 ();
 b15zdnd11an1n04x5 FILLER_184_1883 ();
 b15zdnd00an1n02x5 FILLER_184_1887 ();
 b15zdnd00an1n01x5 FILLER_184_1889 ();
 b15zdnd11an1n64x5 FILLER_184_1893 ();
 b15zdnd11an1n32x5 FILLER_184_1957 ();
 b15zdnd11an1n16x5 FILLER_184_1989 ();
 b15zdnd11an1n08x5 FILLER_184_2005 ();
 b15zdnd00an1n02x5 FILLER_184_2013 ();
 b15zdnd11an1n64x5 FILLER_184_2067 ();
 b15zdnd11an1n16x5 FILLER_184_2131 ();
 b15zdnd11an1n04x5 FILLER_184_2147 ();
 b15zdnd00an1n02x5 FILLER_184_2151 ();
 b15zdnd00an1n01x5 FILLER_184_2153 ();
 b15zdnd00an1n02x5 FILLER_184_2162 ();
 b15zdnd11an1n04x5 FILLER_184_2206 ();
 b15zdnd11an1n04x5 FILLER_184_2215 ();
 b15zdnd00an1n01x5 FILLER_184_2219 ();
 b15zdnd11an1n04x5 FILLER_184_2227 ();
 b15zdnd00an1n02x5 FILLER_184_2273 ();
 b15zdnd00an1n01x5 FILLER_184_2275 ();
 b15zdnd11an1n16x5 FILLER_185_0 ();
 b15zdnd11an1n04x5 FILLER_185_16 ();
 b15zdnd11an1n04x5 FILLER_185_23 ();
 b15zdnd00an1n02x5 FILLER_185_27 ();
 b15zdnd11an1n04x5 FILLER_185_33 ();
 b15zdnd00an1n02x5 FILLER_185_37 ();
 b15zdnd11an1n64x5 FILLER_185_91 ();
 b15zdnd11an1n08x5 FILLER_185_155 ();
 b15zdnd11an1n64x5 FILLER_185_166 ();
 b15zdnd11an1n64x5 FILLER_185_230 ();
 b15zdnd11an1n08x5 FILLER_185_294 ();
 b15zdnd11an1n64x5 FILLER_185_344 ();
 b15zdnd11an1n32x5 FILLER_185_408 ();
 b15zdnd11an1n04x5 FILLER_185_440 ();
 b15zdnd00an1n01x5 FILLER_185_444 ();
 b15zdnd11an1n64x5 FILLER_185_487 ();
 b15zdnd11an1n64x5 FILLER_185_551 ();
 b15zdnd11an1n16x5 FILLER_185_615 ();
 b15zdnd00an1n02x5 FILLER_185_631 ();
 b15zdnd11an1n64x5 FILLER_185_636 ();
 b15zdnd11an1n32x5 FILLER_185_700 ();
 b15zdnd11an1n16x5 FILLER_185_732 ();
 b15zdnd11an1n04x5 FILLER_185_748 ();
 b15zdnd00an1n02x5 FILLER_185_752 ();
 b15zdnd11an1n08x5 FILLER_185_771 ();
 b15zdnd00an1n01x5 FILLER_185_779 ();
 b15zdnd11an1n16x5 FILLER_185_808 ();
 b15zdnd11an1n08x5 FILLER_185_824 ();
 b15zdnd11an1n32x5 FILLER_185_846 ();
 b15zdnd11an1n16x5 FILLER_185_878 ();
 b15zdnd11an1n04x5 FILLER_185_894 ();
 b15zdnd11an1n32x5 FILLER_185_924 ();
 b15zdnd11an1n08x5 FILLER_185_956 ();
 b15zdnd11an1n04x5 FILLER_185_964 ();
 b15zdnd00an1n02x5 FILLER_185_968 ();
 b15zdnd00an1n01x5 FILLER_185_970 ();
 b15zdnd11an1n64x5 FILLER_185_999 ();
 b15zdnd11an1n64x5 FILLER_185_1063 ();
 b15zdnd11an1n64x5 FILLER_185_1127 ();
 b15zdnd11an1n32x5 FILLER_185_1191 ();
 b15zdnd11an1n16x5 FILLER_185_1223 ();
 b15zdnd11an1n08x5 FILLER_185_1239 ();
 b15zdnd11an1n08x5 FILLER_185_1251 ();
 b15zdnd11an1n04x5 FILLER_185_1259 ();
 b15zdnd00an1n02x5 FILLER_185_1263 ();
 b15zdnd00an1n01x5 FILLER_185_1265 ();
 b15zdnd11an1n32x5 FILLER_185_1274 ();
 b15zdnd11an1n16x5 FILLER_185_1306 ();
 b15zdnd11an1n04x5 FILLER_185_1322 ();
 b15zdnd00an1n02x5 FILLER_185_1326 ();
 b15zdnd00an1n01x5 FILLER_185_1328 ();
 b15zdnd11an1n64x5 FILLER_185_1356 ();
 b15zdnd11an1n64x5 FILLER_185_1420 ();
 b15zdnd11an1n64x5 FILLER_185_1484 ();
 b15zdnd11an1n64x5 FILLER_185_1548 ();
 b15zdnd11an1n64x5 FILLER_185_1612 ();
 b15zdnd11an1n64x5 FILLER_185_1676 ();
 b15zdnd11an1n64x5 FILLER_185_1740 ();
 b15zdnd11an1n64x5 FILLER_185_1804 ();
 b15zdnd11an1n16x5 FILLER_185_1868 ();
 b15zdnd11an1n04x5 FILLER_185_1884 ();
 b15zdnd00an1n01x5 FILLER_185_1888 ();
 b15zdnd11an1n64x5 FILLER_185_1892 ();
 b15zdnd11an1n32x5 FILLER_185_1956 ();
 b15zdnd11an1n16x5 FILLER_185_1988 ();
 b15zdnd00an1n02x5 FILLER_185_2004 ();
 b15zdnd00an1n01x5 FILLER_185_2006 ();
 b15zdnd11an1n04x5 FILLER_185_2014 ();
 b15zdnd11an1n32x5 FILLER_185_2060 ();
 b15zdnd11an1n16x5 FILLER_185_2092 ();
 b15zdnd11an1n04x5 FILLER_185_2108 ();
 b15zdnd00an1n01x5 FILLER_185_2112 ();
 b15zdnd11an1n04x5 FILLER_185_2155 ();
 b15zdnd11an1n04x5 FILLER_185_2201 ();
 b15zdnd00an1n02x5 FILLER_185_2205 ();
 b15zdnd00an1n01x5 FILLER_185_2207 ();
 b15zdnd11an1n04x5 FILLER_185_2250 ();
 b15zdnd11an1n04x5 FILLER_185_2278 ();
 b15zdnd00an1n02x5 FILLER_185_2282 ();
 b15zdnd00an1n02x5 FILLER_186_8 ();
 b15zdnd11an1n08x5 FILLER_186_52 ();
 b15zdnd00an1n02x5 FILLER_186_60 ();
 b15zdnd11an1n04x5 FILLER_186_65 ();
 b15zdnd11an1n04x5 FILLER_186_72 ();
 b15zdnd11an1n64x5 FILLER_186_79 ();
 b15zdnd11an1n64x5 FILLER_186_143 ();
 b15zdnd11an1n64x5 FILLER_186_207 ();
 b15zdnd11an1n64x5 FILLER_186_271 ();
 b15zdnd11an1n64x5 FILLER_186_335 ();
 b15zdnd11an1n32x5 FILLER_186_399 ();
 b15zdnd11an1n16x5 FILLER_186_431 ();
 b15zdnd00an1n02x5 FILLER_186_447 ();
 b15zdnd00an1n01x5 FILLER_186_449 ();
 b15zdnd11an1n16x5 FILLER_186_492 ();
 b15zdnd11an1n08x5 FILLER_186_508 ();
 b15zdnd11an1n04x5 FILLER_186_516 ();
 b15zdnd11an1n16x5 FILLER_186_562 ();
 b15zdnd11an1n04x5 FILLER_186_578 ();
 b15zdnd00an1n01x5 FILLER_186_582 ();
 b15zdnd11an1n64x5 FILLER_186_625 ();
 b15zdnd11an1n16x5 FILLER_186_689 ();
 b15zdnd11an1n08x5 FILLER_186_705 ();
 b15zdnd11an1n04x5 FILLER_186_713 ();
 b15zdnd00an1n01x5 FILLER_186_717 ();
 b15zdnd11an1n08x5 FILLER_186_726 ();
 b15zdnd11an1n04x5 FILLER_186_734 ();
 b15zdnd00an1n02x5 FILLER_186_738 ();
 b15zdnd11an1n64x5 FILLER_186_772 ();
 b15zdnd11an1n16x5 FILLER_186_836 ();
 b15zdnd11an1n64x5 FILLER_186_888 ();
 b15zdnd11an1n64x5 FILLER_186_952 ();
 b15zdnd11an1n64x5 FILLER_186_1016 ();
 b15zdnd11an1n64x5 FILLER_186_1080 ();
 b15zdnd11an1n64x5 FILLER_186_1144 ();
 b15zdnd11an1n64x5 FILLER_186_1208 ();
 b15zdnd11an1n32x5 FILLER_186_1272 ();
 b15zdnd11an1n08x5 FILLER_186_1304 ();
 b15zdnd11an1n04x5 FILLER_186_1312 ();
 b15zdnd11an1n64x5 FILLER_186_1368 ();
 b15zdnd11an1n64x5 FILLER_186_1432 ();
 b15zdnd11an1n64x5 FILLER_186_1496 ();
 b15zdnd11an1n64x5 FILLER_186_1560 ();
 b15zdnd11an1n64x5 FILLER_186_1624 ();
 b15zdnd11an1n64x5 FILLER_186_1688 ();
 b15zdnd11an1n64x5 FILLER_186_1752 ();
 b15zdnd11an1n64x5 FILLER_186_1816 ();
 b15zdnd11an1n64x5 FILLER_186_1880 ();
 b15zdnd11an1n64x5 FILLER_186_1944 ();
 b15zdnd11an1n08x5 FILLER_186_2008 ();
 b15zdnd00an1n02x5 FILLER_186_2016 ();
 b15zdnd11an1n64x5 FILLER_186_2060 ();
 b15zdnd11an1n16x5 FILLER_186_2124 ();
 b15zdnd11an1n08x5 FILLER_186_2140 ();
 b15zdnd11an1n04x5 FILLER_186_2148 ();
 b15zdnd00an1n02x5 FILLER_186_2152 ();
 b15zdnd11an1n04x5 FILLER_186_2162 ();
 b15zdnd00an1n02x5 FILLER_186_2166 ();
 b15zdnd00an1n01x5 FILLER_186_2168 ();
 b15zdnd11an1n04x5 FILLER_186_2221 ();
 b15zdnd11an1n04x5 FILLER_186_2228 ();
 b15zdnd00an1n02x5 FILLER_186_2274 ();
 b15zdnd11an1n16x5 FILLER_187_0 ();
 b15zdnd11an1n08x5 FILLER_187_16 ();
 b15zdnd11an1n04x5 FILLER_187_24 ();
 b15zdnd11an1n32x5 FILLER_187_31 ();
 b15zdnd11an1n08x5 FILLER_187_63 ();
 b15zdnd11an1n04x5 FILLER_187_71 ();
 b15zdnd00an1n02x5 FILLER_187_75 ();
 b15zdnd11an1n64x5 FILLER_187_80 ();
 b15zdnd11an1n64x5 FILLER_187_144 ();
 b15zdnd11an1n64x5 FILLER_187_208 ();
 b15zdnd11an1n64x5 FILLER_187_272 ();
 b15zdnd11an1n64x5 FILLER_187_336 ();
 b15zdnd11an1n64x5 FILLER_187_400 ();
 b15zdnd00an1n02x5 FILLER_187_464 ();
 b15zdnd11an1n32x5 FILLER_187_472 ();
 b15zdnd11an1n16x5 FILLER_187_504 ();
 b15zdnd00an1n02x5 FILLER_187_520 ();
 b15zdnd00an1n01x5 FILLER_187_522 ();
 b15zdnd11an1n08x5 FILLER_187_527 ();
 b15zdnd11an1n04x5 FILLER_187_535 ();
 b15zdnd00an1n02x5 FILLER_187_539 ();
 b15zdnd11an1n64x5 FILLER_187_583 ();
 b15zdnd11an1n16x5 FILLER_187_647 ();
 b15zdnd11an1n08x5 FILLER_187_663 ();
 b15zdnd11an1n04x5 FILLER_187_671 ();
 b15zdnd00an1n02x5 FILLER_187_675 ();
 b15zdnd00an1n01x5 FILLER_187_677 ();
 b15zdnd11an1n64x5 FILLER_187_681 ();
 b15zdnd11an1n08x5 FILLER_187_745 ();
 b15zdnd11an1n64x5 FILLER_187_764 ();
 b15zdnd11an1n64x5 FILLER_187_828 ();
 b15zdnd11an1n64x5 FILLER_187_892 ();
 b15zdnd11an1n64x5 FILLER_187_956 ();
 b15zdnd11an1n64x5 FILLER_187_1020 ();
 b15zdnd11an1n64x5 FILLER_187_1084 ();
 b15zdnd11an1n64x5 FILLER_187_1148 ();
 b15zdnd11an1n64x5 FILLER_187_1212 ();
 b15zdnd11an1n32x5 FILLER_187_1276 ();
 b15zdnd11an1n16x5 FILLER_187_1308 ();
 b15zdnd11an1n04x5 FILLER_187_1324 ();
 b15zdnd00an1n01x5 FILLER_187_1328 ();
 b15zdnd11an1n04x5 FILLER_187_1332 ();
 b15zdnd00an1n02x5 FILLER_187_1336 ();
 b15zdnd00an1n01x5 FILLER_187_1338 ();
 b15zdnd11an1n04x5 FILLER_187_1342 ();
 b15zdnd11an1n04x5 FILLER_187_1349 ();
 b15zdnd00an1n02x5 FILLER_187_1353 ();
 b15zdnd11an1n64x5 FILLER_187_1363 ();
 b15zdnd11an1n64x5 FILLER_187_1427 ();
 b15zdnd11an1n64x5 FILLER_187_1491 ();
 b15zdnd11an1n64x5 FILLER_187_1555 ();
 b15zdnd11an1n64x5 FILLER_187_1619 ();
 b15zdnd11an1n64x5 FILLER_187_1683 ();
 b15zdnd11an1n64x5 FILLER_187_1747 ();
 b15zdnd11an1n64x5 FILLER_187_1811 ();
 b15zdnd11an1n64x5 FILLER_187_1875 ();
 b15zdnd11an1n64x5 FILLER_187_1939 ();
 b15zdnd11an1n32x5 FILLER_187_2003 ();
 b15zdnd11an1n04x5 FILLER_187_2035 ();
 b15zdnd11an1n32x5 FILLER_187_2042 ();
 b15zdnd11an1n16x5 FILLER_187_2074 ();
 b15zdnd11an1n08x5 FILLER_187_2090 ();
 b15zdnd00an1n01x5 FILLER_187_2098 ();
 b15zdnd11an1n32x5 FILLER_187_2108 ();
 b15zdnd11an1n16x5 FILLER_187_2140 ();
 b15zdnd11an1n08x5 FILLER_187_2156 ();
 b15zdnd11an1n04x5 FILLER_187_2164 ();
 b15zdnd00an1n02x5 FILLER_187_2168 ();
 b15zdnd00an1n01x5 FILLER_187_2170 ();
 b15zdnd11an1n04x5 FILLER_187_2174 ();
 b15zdnd11an1n04x5 FILLER_187_2181 ();
 b15zdnd11an1n04x5 FILLER_187_2227 ();
 b15zdnd00an1n01x5 FILLER_187_2231 ();
 b15zdnd11an1n04x5 FILLER_187_2236 ();
 b15zdnd00an1n02x5 FILLER_187_2282 ();
 b15zdnd11an1n64x5 FILLER_188_8 ();
 b15zdnd11an1n64x5 FILLER_188_72 ();
 b15zdnd11an1n64x5 FILLER_188_136 ();
 b15zdnd11an1n64x5 FILLER_188_200 ();
 b15zdnd11an1n64x5 FILLER_188_264 ();
 b15zdnd11an1n64x5 FILLER_188_328 ();
 b15zdnd11an1n64x5 FILLER_188_392 ();
 b15zdnd11an1n32x5 FILLER_188_456 ();
 b15zdnd11an1n08x5 FILLER_188_488 ();
 b15zdnd00an1n01x5 FILLER_188_496 ();
 b15zdnd11an1n04x5 FILLER_188_539 ();
 b15zdnd00an1n02x5 FILLER_188_543 ();
 b15zdnd00an1n01x5 FILLER_188_545 ();
 b15zdnd11an1n64x5 FILLER_188_560 ();
 b15zdnd11an1n16x5 FILLER_188_624 ();
 b15zdnd11an1n08x5 FILLER_188_640 ();
 b15zdnd00an1n02x5 FILLER_188_648 ();
 b15zdnd00an1n01x5 FILLER_188_650 ();
 b15zdnd11an1n08x5 FILLER_188_703 ();
 b15zdnd11an1n04x5 FILLER_188_711 ();
 b15zdnd00an1n02x5 FILLER_188_715 ();
 b15zdnd00an1n01x5 FILLER_188_717 ();
 b15zdnd11an1n16x5 FILLER_188_726 ();
 b15zdnd11an1n04x5 FILLER_188_742 ();
 b15zdnd11an1n08x5 FILLER_188_753 ();
 b15zdnd11an1n32x5 FILLER_188_764 ();
 b15zdnd11an1n16x5 FILLER_188_796 ();
 b15zdnd11an1n08x5 FILLER_188_812 ();
 b15zdnd11an1n04x5 FILLER_188_820 ();
 b15zdnd00an1n02x5 FILLER_188_824 ();
 b15zdnd00an1n01x5 FILLER_188_826 ();
 b15zdnd11an1n64x5 FILLER_188_858 ();
 b15zdnd11an1n64x5 FILLER_188_922 ();
 b15zdnd11an1n64x5 FILLER_188_986 ();
 b15zdnd11an1n64x5 FILLER_188_1050 ();
 b15zdnd11an1n64x5 FILLER_188_1114 ();
 b15zdnd11an1n64x5 FILLER_188_1178 ();
 b15zdnd11an1n64x5 FILLER_188_1242 ();
 b15zdnd11an1n64x5 FILLER_188_1306 ();
 b15zdnd11an1n64x5 FILLER_188_1370 ();
 b15zdnd11an1n04x5 FILLER_188_1434 ();
 b15zdnd11an1n64x5 FILLER_188_1490 ();
 b15zdnd11an1n64x5 FILLER_188_1554 ();
 b15zdnd11an1n64x5 FILLER_188_1618 ();
 b15zdnd11an1n64x5 FILLER_188_1682 ();
 b15zdnd11an1n64x5 FILLER_188_1746 ();
 b15zdnd11an1n64x5 FILLER_188_1810 ();
 b15zdnd11an1n64x5 FILLER_188_1874 ();
 b15zdnd11an1n64x5 FILLER_188_1938 ();
 b15zdnd11an1n64x5 FILLER_188_2002 ();
 b15zdnd11an1n64x5 FILLER_188_2066 ();
 b15zdnd11an1n16x5 FILLER_188_2130 ();
 b15zdnd11an1n08x5 FILLER_188_2146 ();
 b15zdnd11an1n16x5 FILLER_188_2162 ();
 b15zdnd11an1n04x5 FILLER_188_2178 ();
 b15zdnd00an1n01x5 FILLER_188_2182 ();
 b15zdnd11an1n04x5 FILLER_188_2187 ();
 b15zdnd11an1n04x5 FILLER_188_2233 ();
 b15zdnd11an1n04x5 FILLER_188_2270 ();
 b15zdnd00an1n02x5 FILLER_188_2274 ();
 b15zdnd11an1n64x5 FILLER_189_0 ();
 b15zdnd11an1n64x5 FILLER_189_64 ();
 b15zdnd11an1n64x5 FILLER_189_128 ();
 b15zdnd11an1n64x5 FILLER_189_192 ();
 b15zdnd11an1n64x5 FILLER_189_256 ();
 b15zdnd11an1n64x5 FILLER_189_320 ();
 b15zdnd11an1n64x5 FILLER_189_384 ();
 b15zdnd11an1n32x5 FILLER_189_448 ();
 b15zdnd11an1n16x5 FILLER_189_480 ();
 b15zdnd11an1n04x5 FILLER_189_496 ();
 b15zdnd00an1n02x5 FILLER_189_500 ();
 b15zdnd11an1n32x5 FILLER_189_544 ();
 b15zdnd11an1n16x5 FILLER_189_576 ();
 b15zdnd00an1n02x5 FILLER_189_592 ();
 b15zdnd00an1n01x5 FILLER_189_594 ();
 b15zdnd11an1n32x5 FILLER_189_637 ();
 b15zdnd11an1n04x5 FILLER_189_672 ();
 b15zdnd11an1n64x5 FILLER_189_679 ();
 b15zdnd11an1n16x5 FILLER_189_743 ();
 b15zdnd11an1n04x5 FILLER_189_759 ();
 b15zdnd00an1n02x5 FILLER_189_763 ();
 b15zdnd00an1n01x5 FILLER_189_765 ();
 b15zdnd11an1n04x5 FILLER_189_772 ();
 b15zdnd11an1n32x5 FILLER_189_787 ();
 b15zdnd00an1n01x5 FILLER_189_819 ();
 b15zdnd11an1n16x5 FILLER_189_844 ();
 b15zdnd00an1n02x5 FILLER_189_860 ();
 b15zdnd11an1n64x5 FILLER_189_869 ();
 b15zdnd11an1n32x5 FILLER_189_933 ();
 b15zdnd11an1n08x5 FILLER_189_965 ();
 b15zdnd11an1n04x5 FILLER_189_973 ();
 b15zdnd00an1n02x5 FILLER_189_977 ();
 b15zdnd00an1n01x5 FILLER_189_979 ();
 b15zdnd11an1n16x5 FILLER_189_1004 ();
 b15zdnd11an1n04x5 FILLER_189_1020 ();
 b15zdnd11an1n32x5 FILLER_189_1066 ();
 b15zdnd11an1n16x5 FILLER_189_1098 ();
 b15zdnd11an1n08x5 FILLER_189_1114 ();
 b15zdnd11an1n04x5 FILLER_189_1122 ();
 b15zdnd00an1n02x5 FILLER_189_1126 ();
 b15zdnd11an1n64x5 FILLER_189_1170 ();
 b15zdnd11an1n64x5 FILLER_189_1234 ();
 b15zdnd11an1n64x5 FILLER_189_1298 ();
 b15zdnd11an1n32x5 FILLER_189_1362 ();
 b15zdnd11an1n16x5 FILLER_189_1394 ();
 b15zdnd11an1n08x5 FILLER_189_1410 ();
 b15zdnd11an1n04x5 FILLER_189_1418 ();
 b15zdnd11an1n04x5 FILLER_189_1474 ();
 b15zdnd11an1n64x5 FILLER_189_1481 ();
 b15zdnd11an1n64x5 FILLER_189_1545 ();
 b15zdnd11an1n64x5 FILLER_189_1609 ();
 b15zdnd11an1n64x5 FILLER_189_1673 ();
 b15zdnd11an1n64x5 FILLER_189_1737 ();
 b15zdnd11an1n64x5 FILLER_189_1801 ();
 b15zdnd11an1n64x5 FILLER_189_1865 ();
 b15zdnd11an1n64x5 FILLER_189_1929 ();
 b15zdnd11an1n64x5 FILLER_189_1993 ();
 b15zdnd11an1n64x5 FILLER_189_2057 ();
 b15zdnd11an1n32x5 FILLER_189_2121 ();
 b15zdnd11an1n16x5 FILLER_189_2153 ();
 b15zdnd11an1n04x5 FILLER_189_2169 ();
 b15zdnd00an1n02x5 FILLER_189_2173 ();
 b15zdnd11an1n04x5 FILLER_189_2206 ();
 b15zdnd11an1n04x5 FILLER_189_2252 ();
 b15zdnd11an1n04x5 FILLER_189_2280 ();
 b15zdnd11an1n64x5 FILLER_190_8 ();
 b15zdnd11an1n64x5 FILLER_190_72 ();
 b15zdnd11an1n64x5 FILLER_190_136 ();
 b15zdnd11an1n64x5 FILLER_190_200 ();
 b15zdnd11an1n64x5 FILLER_190_264 ();
 b15zdnd11an1n64x5 FILLER_190_328 ();
 b15zdnd11an1n64x5 FILLER_190_392 ();
 b15zdnd11an1n64x5 FILLER_190_456 ();
 b15zdnd11an1n04x5 FILLER_190_520 ();
 b15zdnd00an1n01x5 FILLER_190_524 ();
 b15zdnd11an1n64x5 FILLER_190_539 ();
 b15zdnd11an1n64x5 FILLER_190_603 ();
 b15zdnd11an1n32x5 FILLER_190_667 ();
 b15zdnd11an1n16x5 FILLER_190_699 ();
 b15zdnd00an1n02x5 FILLER_190_715 ();
 b15zdnd00an1n01x5 FILLER_190_717 ();
 b15zdnd11an1n64x5 FILLER_190_726 ();
 b15zdnd11an1n32x5 FILLER_190_790 ();
 b15zdnd00an1n02x5 FILLER_190_822 ();
 b15zdnd11an1n64x5 FILLER_190_876 ();
 b15zdnd11an1n32x5 FILLER_190_940 ();
 b15zdnd11an1n08x5 FILLER_190_972 ();
 b15zdnd00an1n02x5 FILLER_190_980 ();
 b15zdnd11an1n04x5 FILLER_190_988 ();
 b15zdnd11an1n64x5 FILLER_190_995 ();
 b15zdnd11an1n64x5 FILLER_190_1059 ();
 b15zdnd11an1n16x5 FILLER_190_1123 ();
 b15zdnd11an1n08x5 FILLER_190_1139 ();
 b15zdnd11an1n64x5 FILLER_190_1150 ();
 b15zdnd11an1n16x5 FILLER_190_1214 ();
 b15zdnd11an1n04x5 FILLER_190_1230 ();
 b15zdnd00an1n02x5 FILLER_190_1234 ();
 b15zdnd00an1n01x5 FILLER_190_1236 ();
 b15zdnd11an1n64x5 FILLER_190_1260 ();
 b15zdnd11an1n64x5 FILLER_190_1324 ();
 b15zdnd11an1n32x5 FILLER_190_1388 ();
 b15zdnd11an1n16x5 FILLER_190_1420 ();
 b15zdnd11an1n04x5 FILLER_190_1436 ();
 b15zdnd11an1n04x5 FILLER_190_1443 ();
 b15zdnd11an1n08x5 FILLER_190_1450 ();
 b15zdnd11an1n04x5 FILLER_190_1458 ();
 b15zdnd00an1n01x5 FILLER_190_1462 ();
 b15zdnd11an1n04x5 FILLER_190_1466 ();
 b15zdnd11an1n64x5 FILLER_190_1473 ();
 b15zdnd11an1n64x5 FILLER_190_1537 ();
 b15zdnd11an1n64x5 FILLER_190_1601 ();
 b15zdnd11an1n16x5 FILLER_190_1665 ();
 b15zdnd11an1n08x5 FILLER_190_1681 ();
 b15zdnd00an1n02x5 FILLER_190_1689 ();
 b15zdnd00an1n01x5 FILLER_190_1691 ();
 b15zdnd11an1n32x5 FILLER_190_1712 ();
 b15zdnd11an1n08x5 FILLER_190_1744 ();
 b15zdnd11an1n04x5 FILLER_190_1752 ();
 b15zdnd00an1n01x5 FILLER_190_1756 ();
 b15zdnd11an1n64x5 FILLER_190_1788 ();
 b15zdnd11an1n64x5 FILLER_190_1852 ();
 b15zdnd11an1n64x5 FILLER_190_1916 ();
 b15zdnd11an1n64x5 FILLER_190_1980 ();
 b15zdnd11an1n64x5 FILLER_190_2044 ();
 b15zdnd11an1n32x5 FILLER_190_2108 ();
 b15zdnd11an1n08x5 FILLER_190_2140 ();
 b15zdnd11an1n04x5 FILLER_190_2148 ();
 b15zdnd00an1n02x5 FILLER_190_2152 ();
 b15zdnd11an1n04x5 FILLER_190_2162 ();
 b15zdnd00an1n01x5 FILLER_190_2166 ();
 b15zdnd11an1n04x5 FILLER_190_2185 ();
 b15zdnd11an1n04x5 FILLER_190_2222 ();
 b15zdnd11an1n08x5 FILLER_190_2268 ();
 b15zdnd11an1n64x5 FILLER_191_0 ();
 b15zdnd11an1n64x5 FILLER_191_64 ();
 b15zdnd11an1n64x5 FILLER_191_128 ();
 b15zdnd11an1n32x5 FILLER_191_192 ();
 b15zdnd11an1n64x5 FILLER_191_233 ();
 b15zdnd11an1n64x5 FILLER_191_297 ();
 b15zdnd11an1n64x5 FILLER_191_361 ();
 b15zdnd11an1n32x5 FILLER_191_425 ();
 b15zdnd11an1n16x5 FILLER_191_457 ();
 b15zdnd00an1n02x5 FILLER_191_473 ();
 b15zdnd11an1n64x5 FILLER_191_517 ();
 b15zdnd11an1n64x5 FILLER_191_581 ();
 b15zdnd11an1n64x5 FILLER_191_645 ();
 b15zdnd11an1n64x5 FILLER_191_709 ();
 b15zdnd11an1n64x5 FILLER_191_773 ();
 b15zdnd11an1n32x5 FILLER_191_837 ();
 b15zdnd11an1n16x5 FILLER_191_869 ();
 b15zdnd11an1n04x5 FILLER_191_885 ();
 b15zdnd00an1n02x5 FILLER_191_889 ();
 b15zdnd00an1n01x5 FILLER_191_891 ();
 b15zdnd11an1n64x5 FILLER_191_902 ();
 b15zdnd11an1n64x5 FILLER_191_966 ();
 b15zdnd11an1n64x5 FILLER_191_1030 ();
 b15zdnd11an1n64x5 FILLER_191_1094 ();
 b15zdnd11an1n64x5 FILLER_191_1158 ();
 b15zdnd11an1n64x5 FILLER_191_1222 ();
 b15zdnd11an1n64x5 FILLER_191_1286 ();
 b15zdnd11an1n64x5 FILLER_191_1350 ();
 b15zdnd11an1n32x5 FILLER_191_1414 ();
 b15zdnd11an1n64x5 FILLER_191_1449 ();
 b15zdnd11an1n64x5 FILLER_191_1513 ();
 b15zdnd11an1n64x5 FILLER_191_1577 ();
 b15zdnd11an1n64x5 FILLER_191_1641 ();
 b15zdnd11an1n64x5 FILLER_191_1705 ();
 b15zdnd11an1n64x5 FILLER_191_1769 ();
 b15zdnd11an1n64x5 FILLER_191_1833 ();
 b15zdnd11an1n64x5 FILLER_191_1897 ();
 b15zdnd11an1n64x5 FILLER_191_1961 ();
 b15zdnd11an1n64x5 FILLER_191_2025 ();
 b15zdnd11an1n32x5 FILLER_191_2089 ();
 b15zdnd11an1n16x5 FILLER_191_2121 ();
 b15zdnd11an1n04x5 FILLER_191_2137 ();
 b15zdnd00an1n02x5 FILLER_191_2141 ();
 b15zdnd00an1n01x5 FILLER_191_2143 ();
 b15zdnd11an1n08x5 FILLER_191_2186 ();
 b15zdnd11an1n04x5 FILLER_191_2236 ();
 b15zdnd00an1n02x5 FILLER_191_2282 ();
 b15zdnd11an1n64x5 FILLER_192_8 ();
 b15zdnd11an1n64x5 FILLER_192_72 ();
 b15zdnd11an1n64x5 FILLER_192_136 ();
 b15zdnd11an1n08x5 FILLER_192_200 ();
 b15zdnd00an1n02x5 FILLER_192_208 ();
 b15zdnd11an1n16x5 FILLER_192_219 ();
 b15zdnd11an1n08x5 FILLER_192_235 ();
 b15zdnd11an1n04x5 FILLER_192_243 ();
 b15zdnd00an1n01x5 FILLER_192_247 ();
 b15zdnd11an1n64x5 FILLER_192_260 ();
 b15zdnd11an1n64x5 FILLER_192_324 ();
 b15zdnd11an1n64x5 FILLER_192_388 ();
 b15zdnd11an1n64x5 FILLER_192_452 ();
 b15zdnd11an1n32x5 FILLER_192_516 ();
 b15zdnd11an1n16x5 FILLER_192_548 ();
 b15zdnd11an1n08x5 FILLER_192_564 ();
 b15zdnd00an1n02x5 FILLER_192_572 ();
 b15zdnd11an1n08x5 FILLER_192_582 ();
 b15zdnd11an1n04x5 FILLER_192_590 ();
 b15zdnd11an1n64x5 FILLER_192_608 ();
 b15zdnd11an1n32x5 FILLER_192_672 ();
 b15zdnd11an1n08x5 FILLER_192_704 ();
 b15zdnd11an1n04x5 FILLER_192_712 ();
 b15zdnd00an1n02x5 FILLER_192_716 ();
 b15zdnd11an1n64x5 FILLER_192_726 ();
 b15zdnd11an1n64x5 FILLER_192_790 ();
 b15zdnd11an1n16x5 FILLER_192_854 ();
 b15zdnd11an1n08x5 FILLER_192_870 ();
 b15zdnd11an1n04x5 FILLER_192_878 ();
 b15zdnd00an1n02x5 FILLER_192_882 ();
 b15zdnd11an1n64x5 FILLER_192_918 ();
 b15zdnd11an1n64x5 FILLER_192_982 ();
 b15zdnd11an1n64x5 FILLER_192_1046 ();
 b15zdnd11an1n64x5 FILLER_192_1110 ();
 b15zdnd11an1n64x5 FILLER_192_1174 ();
 b15zdnd11an1n64x5 FILLER_192_1238 ();
 b15zdnd11an1n64x5 FILLER_192_1302 ();
 b15zdnd11an1n32x5 FILLER_192_1366 ();
 b15zdnd11an1n16x5 FILLER_192_1398 ();
 b15zdnd11an1n08x5 FILLER_192_1414 ();
 b15zdnd11an1n04x5 FILLER_192_1422 ();
 b15zdnd00an1n02x5 FILLER_192_1426 ();
 b15zdnd11an1n64x5 FILLER_192_1480 ();
 b15zdnd11an1n64x5 FILLER_192_1544 ();
 b15zdnd11an1n64x5 FILLER_192_1608 ();
 b15zdnd11an1n64x5 FILLER_192_1672 ();
 b15zdnd11an1n64x5 FILLER_192_1736 ();
 b15zdnd11an1n64x5 FILLER_192_1800 ();
 b15zdnd11an1n64x5 FILLER_192_1864 ();
 b15zdnd11an1n64x5 FILLER_192_1928 ();
 b15zdnd11an1n64x5 FILLER_192_1992 ();
 b15zdnd11an1n32x5 FILLER_192_2056 ();
 b15zdnd11an1n16x5 FILLER_192_2088 ();
 b15zdnd11an1n08x5 FILLER_192_2104 ();
 b15zdnd11an1n04x5 FILLER_192_2112 ();
 b15zdnd00an1n02x5 FILLER_192_2116 ();
 b15zdnd00an1n01x5 FILLER_192_2118 ();
 b15zdnd11an1n32x5 FILLER_192_2122 ();
 b15zdnd00an1n02x5 FILLER_192_2162 ();
 b15zdnd11an1n08x5 FILLER_192_2206 ();
 b15zdnd00an1n02x5 FILLER_192_2214 ();
 b15zdnd11an1n04x5 FILLER_192_2220 ();
 b15zdnd11an1n04x5 FILLER_192_2228 ();
 b15zdnd00an1n02x5 FILLER_192_2274 ();
 b15zdnd11an1n64x5 FILLER_193_0 ();
 b15zdnd11an1n64x5 FILLER_193_64 ();
 b15zdnd11an1n32x5 FILLER_193_128 ();
 b15zdnd11an1n08x5 FILLER_193_160 ();
 b15zdnd11an1n04x5 FILLER_193_168 ();
 b15zdnd11an1n04x5 FILLER_193_212 ();
 b15zdnd11an1n04x5 FILLER_193_219 ();
 b15zdnd11an1n16x5 FILLER_193_226 ();
 b15zdnd11an1n04x5 FILLER_193_242 ();
 b15zdnd00an1n02x5 FILLER_193_246 ();
 b15zdnd00an1n01x5 FILLER_193_248 ();
 b15zdnd11an1n64x5 FILLER_193_252 ();
 b15zdnd11an1n64x5 FILLER_193_316 ();
 b15zdnd11an1n32x5 FILLER_193_380 ();
 b15zdnd11an1n16x5 FILLER_193_412 ();
 b15zdnd11an1n08x5 FILLER_193_428 ();
 b15zdnd00an1n01x5 FILLER_193_436 ();
 b15zdnd11an1n32x5 FILLER_193_442 ();
 b15zdnd00an1n02x5 FILLER_193_474 ();
 b15zdnd00an1n01x5 FILLER_193_476 ();
 b15zdnd11an1n64x5 FILLER_193_489 ();
 b15zdnd11an1n64x5 FILLER_193_553 ();
 b15zdnd11an1n64x5 FILLER_193_617 ();
 b15zdnd11an1n64x5 FILLER_193_681 ();
 b15zdnd11an1n32x5 FILLER_193_745 ();
 b15zdnd11an1n16x5 FILLER_193_777 ();
 b15zdnd11an1n08x5 FILLER_193_793 ();
 b15zdnd11an1n04x5 FILLER_193_801 ();
 b15zdnd00an1n02x5 FILLER_193_805 ();
 b15zdnd00an1n01x5 FILLER_193_807 ();
 b15zdnd11an1n64x5 FILLER_193_822 ();
 b15zdnd11an1n64x5 FILLER_193_886 ();
 b15zdnd11an1n64x5 FILLER_193_950 ();
 b15zdnd11an1n64x5 FILLER_193_1014 ();
 b15zdnd11an1n32x5 FILLER_193_1078 ();
 b15zdnd11an1n16x5 FILLER_193_1110 ();
 b15zdnd11an1n08x5 FILLER_193_1126 ();
 b15zdnd11an1n04x5 FILLER_193_1134 ();
 b15zdnd00an1n02x5 FILLER_193_1138 ();
 b15zdnd00an1n01x5 FILLER_193_1140 ();
 b15zdnd11an1n32x5 FILLER_193_1169 ();
 b15zdnd00an1n01x5 FILLER_193_1201 ();
 b15zdnd11an1n64x5 FILLER_193_1210 ();
 b15zdnd11an1n64x5 FILLER_193_1274 ();
 b15zdnd11an1n64x5 FILLER_193_1338 ();
 b15zdnd11an1n32x5 FILLER_193_1402 ();
 b15zdnd11an1n08x5 FILLER_193_1434 ();
 b15zdnd11an1n04x5 FILLER_193_1442 ();
 b15zdnd00an1n01x5 FILLER_193_1446 ();
 b15zdnd11an1n04x5 FILLER_193_1450 ();
 b15zdnd11an1n64x5 FILLER_193_1457 ();
 b15zdnd11an1n64x5 FILLER_193_1521 ();
 b15zdnd11an1n64x5 FILLER_193_1585 ();
 b15zdnd11an1n64x5 FILLER_193_1649 ();
 b15zdnd11an1n64x5 FILLER_193_1713 ();
 b15zdnd11an1n64x5 FILLER_193_1777 ();
 b15zdnd11an1n64x5 FILLER_193_1841 ();
 b15zdnd11an1n64x5 FILLER_193_1905 ();
 b15zdnd11an1n32x5 FILLER_193_1969 ();
 b15zdnd11an1n08x5 FILLER_193_2001 ();
 b15zdnd11an1n08x5 FILLER_193_2016 ();
 b15zdnd11an1n32x5 FILLER_193_2036 ();
 b15zdnd11an1n16x5 FILLER_193_2068 ();
 b15zdnd11an1n08x5 FILLER_193_2084 ();
 b15zdnd00an1n01x5 FILLER_193_2092 ();
 b15zdnd11an1n04x5 FILLER_193_2145 ();
 b15zdnd11an1n08x5 FILLER_193_2191 ();
 b15zdnd11an1n04x5 FILLER_193_2199 ();
 b15zdnd00an1n02x5 FILLER_193_2203 ();
 b15zdnd11an1n04x5 FILLER_193_2236 ();
 b15zdnd00an1n02x5 FILLER_193_2282 ();
 b15zdnd11an1n64x5 FILLER_194_8 ();
 b15zdnd11an1n64x5 FILLER_194_72 ();
 b15zdnd11an1n64x5 FILLER_194_136 ();
 b15zdnd11an1n64x5 FILLER_194_200 ();
 b15zdnd11an1n64x5 FILLER_194_264 ();
 b15zdnd11an1n64x5 FILLER_194_328 ();
 b15zdnd11an1n16x5 FILLER_194_392 ();
 b15zdnd00an1n01x5 FILLER_194_408 ();
 b15zdnd11an1n64x5 FILLER_194_412 ();
 b15zdnd11an1n04x5 FILLER_194_476 ();
 b15zdnd11an1n64x5 FILLER_194_486 ();
 b15zdnd11an1n04x5 FILLER_194_550 ();
 b15zdnd00an1n02x5 FILLER_194_554 ();
 b15zdnd11an1n64x5 FILLER_194_564 ();
 b15zdnd11an1n64x5 FILLER_194_628 ();
 b15zdnd11an1n16x5 FILLER_194_692 ();
 b15zdnd11an1n08x5 FILLER_194_708 ();
 b15zdnd00an1n02x5 FILLER_194_716 ();
 b15zdnd11an1n32x5 FILLER_194_726 ();
 b15zdnd11an1n08x5 FILLER_194_758 ();
 b15zdnd11an1n04x5 FILLER_194_766 ();
 b15zdnd00an1n01x5 FILLER_194_770 ();
 b15zdnd11an1n64x5 FILLER_194_816 ();
 b15zdnd11an1n08x5 FILLER_194_880 ();
 b15zdnd11an1n04x5 FILLER_194_888 ();
 b15zdnd00an1n02x5 FILLER_194_892 ();
 b15zdnd11an1n04x5 FILLER_194_905 ();
 b15zdnd11an1n32x5 FILLER_194_931 ();
 b15zdnd11an1n04x5 FILLER_194_963 ();
 b15zdnd00an1n01x5 FILLER_194_967 ();
 b15zdnd11an1n64x5 FILLER_194_985 ();
 b15zdnd11an1n64x5 FILLER_194_1049 ();
 b15zdnd11an1n08x5 FILLER_194_1113 ();
 b15zdnd11an1n04x5 FILLER_194_1121 ();
 b15zdnd00an1n02x5 FILLER_194_1125 ();
 b15zdnd00an1n01x5 FILLER_194_1127 ();
 b15zdnd11an1n64x5 FILLER_194_1170 ();
 b15zdnd11an1n64x5 FILLER_194_1234 ();
 b15zdnd11an1n64x5 FILLER_194_1298 ();
 b15zdnd11an1n64x5 FILLER_194_1362 ();
 b15zdnd11an1n16x5 FILLER_194_1426 ();
 b15zdnd11an1n08x5 FILLER_194_1442 ();
 b15zdnd00an1n02x5 FILLER_194_1450 ();
 b15zdnd00an1n01x5 FILLER_194_1452 ();
 b15zdnd11an1n64x5 FILLER_194_1456 ();
 b15zdnd11an1n64x5 FILLER_194_1520 ();
 b15zdnd00an1n01x5 FILLER_194_1584 ();
 b15zdnd11an1n64x5 FILLER_194_1588 ();
 b15zdnd11an1n32x5 FILLER_194_1652 ();
 b15zdnd11an1n08x5 FILLER_194_1684 ();
 b15zdnd11an1n04x5 FILLER_194_1692 ();
 b15zdnd00an1n01x5 FILLER_194_1696 ();
 b15zdnd11an1n04x5 FILLER_194_1700 ();
 b15zdnd11an1n64x5 FILLER_194_1707 ();
 b15zdnd11an1n64x5 FILLER_194_1771 ();
 b15zdnd11an1n64x5 FILLER_194_1835 ();
 b15zdnd11an1n64x5 FILLER_194_1899 ();
 b15zdnd11an1n32x5 FILLER_194_1963 ();
 b15zdnd11an1n64x5 FILLER_194_2037 ();
 b15zdnd00an1n02x5 FILLER_194_2101 ();
 b15zdnd00an1n01x5 FILLER_194_2103 ();
 b15zdnd11an1n04x5 FILLER_194_2107 ();
 b15zdnd11an1n04x5 FILLER_194_2117 ();
 b15zdnd11an1n16x5 FILLER_194_2124 ();
 b15zdnd11an1n04x5 FILLER_194_2140 ();
 b15zdnd00an1n01x5 FILLER_194_2144 ();
 b15zdnd00an1n02x5 FILLER_194_2152 ();
 b15zdnd11an1n64x5 FILLER_194_2162 ();
 b15zdnd11an1n08x5 FILLER_194_2268 ();
 b15zdnd11an1n64x5 FILLER_195_0 ();
 b15zdnd11an1n64x5 FILLER_195_64 ();
 b15zdnd11an1n64x5 FILLER_195_128 ();
 b15zdnd11an1n64x5 FILLER_195_192 ();
 b15zdnd11an1n64x5 FILLER_195_256 ();
 b15zdnd11an1n64x5 FILLER_195_320 ();
 b15zdnd11an1n08x5 FILLER_195_384 ();
 b15zdnd11an1n16x5 FILLER_195_444 ();
 b15zdnd11an1n08x5 FILLER_195_460 ();
 b15zdnd00an1n01x5 FILLER_195_468 ();
 b15zdnd11an1n08x5 FILLER_195_472 ();
 b15zdnd11an1n64x5 FILLER_195_483 ();
 b15zdnd11an1n64x5 FILLER_195_547 ();
 b15zdnd11an1n64x5 FILLER_195_611 ();
 b15zdnd11an1n32x5 FILLER_195_675 ();
 b15zdnd11an1n04x5 FILLER_195_707 ();
 b15zdnd00an1n01x5 FILLER_195_711 ();
 b15zdnd11an1n32x5 FILLER_195_754 ();
 b15zdnd11an1n16x5 FILLER_195_786 ();
 b15zdnd11an1n04x5 FILLER_195_805 ();
 b15zdnd11an1n64x5 FILLER_195_821 ();
 b15zdnd11an1n64x5 FILLER_195_885 ();
 b15zdnd11an1n16x5 FILLER_195_949 ();
 b15zdnd11an1n08x5 FILLER_195_965 ();
 b15zdnd00an1n01x5 FILLER_195_973 ();
 b15zdnd11an1n04x5 FILLER_195_980 ();
 b15zdnd11an1n04x5 FILLER_195_987 ();
 b15zdnd11an1n64x5 FILLER_195_1019 ();
 b15zdnd11an1n04x5 FILLER_195_1083 ();
 b15zdnd00an1n02x5 FILLER_195_1087 ();
 b15zdnd00an1n01x5 FILLER_195_1089 ();
 b15zdnd11an1n64x5 FILLER_195_1101 ();
 b15zdnd11an1n64x5 FILLER_195_1165 ();
 b15zdnd11an1n64x5 FILLER_195_1229 ();
 b15zdnd11an1n64x5 FILLER_195_1293 ();
 b15zdnd11an1n64x5 FILLER_195_1357 ();
 b15zdnd11an1n64x5 FILLER_195_1421 ();
 b15zdnd11an1n64x5 FILLER_195_1485 ();
 b15zdnd11an1n32x5 FILLER_195_1549 ();
 b15zdnd00an1n02x5 FILLER_195_1581 ();
 b15zdnd00an1n01x5 FILLER_195_1583 ();
 b15zdnd11an1n04x5 FILLER_195_1587 ();
 b15zdnd11an1n32x5 FILLER_195_1594 ();
 b15zdnd11an1n16x5 FILLER_195_1626 ();
 b15zdnd11an1n04x5 FILLER_195_1645 ();
 b15zdnd11an1n16x5 FILLER_195_1652 ();
 b15zdnd11an1n08x5 FILLER_195_1668 ();
 b15zdnd00an1n02x5 FILLER_195_1676 ();
 b15zdnd00an1n01x5 FILLER_195_1678 ();
 b15zdnd11an1n64x5 FILLER_195_1731 ();
 b15zdnd11an1n64x5 FILLER_195_1795 ();
 b15zdnd11an1n64x5 FILLER_195_1859 ();
 b15zdnd11an1n32x5 FILLER_195_1923 ();
 b15zdnd11an1n08x5 FILLER_195_1955 ();
 b15zdnd00an1n02x5 FILLER_195_1963 ();
 b15zdnd00an1n01x5 FILLER_195_1965 ();
 b15zdnd11an1n32x5 FILLER_195_2008 ();
 b15zdnd00an1n01x5 FILLER_195_2040 ();
 b15zdnd11an1n32x5 FILLER_195_2044 ();
 b15zdnd11an1n16x5 FILLER_195_2076 ();
 b15zdnd00an1n02x5 FILLER_195_2092 ();
 b15zdnd11an1n08x5 FILLER_195_2100 ();
 b15zdnd11an1n04x5 FILLER_195_2108 ();
 b15zdnd00an1n02x5 FILLER_195_2112 ();
 b15zdnd11an1n32x5 FILLER_195_2156 ();
 b15zdnd11an1n16x5 FILLER_195_2188 ();
 b15zdnd00an1n02x5 FILLER_195_2204 ();
 b15zdnd11an1n16x5 FILLER_195_2211 ();
 b15zdnd11an1n08x5 FILLER_195_2227 ();
 b15zdnd11an1n04x5 FILLER_195_2235 ();
 b15zdnd00an1n01x5 FILLER_195_2239 ();
 b15zdnd00an1n02x5 FILLER_195_2282 ();
 b15zdnd11an1n64x5 FILLER_196_8 ();
 b15zdnd11an1n64x5 FILLER_196_72 ();
 b15zdnd11an1n64x5 FILLER_196_136 ();
 b15zdnd11an1n64x5 FILLER_196_200 ();
 b15zdnd11an1n32x5 FILLER_196_264 ();
 b15zdnd11an1n08x5 FILLER_196_296 ();
 b15zdnd11an1n04x5 FILLER_196_304 ();
 b15zdnd00an1n01x5 FILLER_196_308 ();
 b15zdnd11an1n32x5 FILLER_196_361 ();
 b15zdnd11an1n16x5 FILLER_196_393 ();
 b15zdnd11an1n04x5 FILLER_196_409 ();
 b15zdnd00an1n02x5 FILLER_196_413 ();
 b15zdnd11an1n32x5 FILLER_196_418 ();
 b15zdnd11an1n04x5 FILLER_196_450 ();
 b15zdnd00an1n02x5 FILLER_196_454 ();
 b15zdnd00an1n01x5 FILLER_196_456 ();
 b15zdnd11an1n04x5 FILLER_196_460 ();
 b15zdnd00an1n02x5 FILLER_196_464 ();
 b15zdnd00an1n01x5 FILLER_196_466 ();
 b15zdnd11an1n64x5 FILLER_196_509 ();
 b15zdnd11an1n16x5 FILLER_196_573 ();
 b15zdnd00an1n01x5 FILLER_196_589 ();
 b15zdnd11an1n04x5 FILLER_196_598 ();
 b15zdnd11an1n64x5 FILLER_196_608 ();
 b15zdnd11an1n32x5 FILLER_196_672 ();
 b15zdnd11an1n08x5 FILLER_196_704 ();
 b15zdnd11an1n04x5 FILLER_196_712 ();
 b15zdnd00an1n02x5 FILLER_196_716 ();
 b15zdnd11an1n32x5 FILLER_196_726 ();
 b15zdnd11an1n16x5 FILLER_196_758 ();
 b15zdnd00an1n01x5 FILLER_196_774 ();
 b15zdnd11an1n64x5 FILLER_196_827 ();
 b15zdnd11an1n64x5 FILLER_196_891 ();
 b15zdnd11an1n08x5 FILLER_196_955 ();
 b15zdnd11an1n04x5 FILLER_196_963 ();
 b15zdnd11an1n64x5 FILLER_196_1012 ();
 b15zdnd11an1n32x5 FILLER_196_1076 ();
 b15zdnd11an1n16x5 FILLER_196_1108 ();
 b15zdnd11an1n04x5 FILLER_196_1124 ();
 b15zdnd11an1n64x5 FILLER_196_1143 ();
 b15zdnd11an1n08x5 FILLER_196_1207 ();
 b15zdnd11an1n04x5 FILLER_196_1215 ();
 b15zdnd11an1n64x5 FILLER_196_1224 ();
 b15zdnd11an1n64x5 FILLER_196_1288 ();
 b15zdnd11an1n64x5 FILLER_196_1352 ();
 b15zdnd11an1n64x5 FILLER_196_1416 ();
 b15zdnd11an1n64x5 FILLER_196_1480 ();
 b15zdnd11an1n16x5 FILLER_196_1544 ();
 b15zdnd11an1n04x5 FILLER_196_1560 ();
 b15zdnd00an1n01x5 FILLER_196_1564 ();
 b15zdnd11an1n04x5 FILLER_196_1617 ();
 b15zdnd11an1n16x5 FILLER_196_1673 ();
 b15zdnd11an1n08x5 FILLER_196_1689 ();
 b15zdnd11an1n04x5 FILLER_196_1697 ();
 b15zdnd00an1n02x5 FILLER_196_1701 ();
 b15zdnd00an1n01x5 FILLER_196_1703 ();
 b15zdnd11an1n64x5 FILLER_196_1707 ();
 b15zdnd11an1n64x5 FILLER_196_1771 ();
 b15zdnd11an1n64x5 FILLER_196_1835 ();
 b15zdnd11an1n64x5 FILLER_196_1899 ();
 b15zdnd11an1n32x5 FILLER_196_1963 ();
 b15zdnd11an1n16x5 FILLER_196_1995 ();
 b15zdnd11an1n04x5 FILLER_196_2011 ();
 b15zdnd00an1n02x5 FILLER_196_2015 ();
 b15zdnd00an1n01x5 FILLER_196_2017 ();
 b15zdnd11an1n64x5 FILLER_196_2060 ();
 b15zdnd11an1n08x5 FILLER_196_2124 ();
 b15zdnd00an1n02x5 FILLER_196_2132 ();
 b15zdnd11an1n08x5 FILLER_196_2143 ();
 b15zdnd00an1n02x5 FILLER_196_2151 ();
 b15zdnd00an1n01x5 FILLER_196_2153 ();
 b15zdnd11an1n16x5 FILLER_196_2162 ();
 b15zdnd11an1n04x5 FILLER_196_2178 ();
 b15zdnd00an1n01x5 FILLER_196_2182 ();
 b15zdnd11an1n16x5 FILLER_196_2225 ();
 b15zdnd00an1n02x5 FILLER_196_2241 ();
 b15zdnd00an1n01x5 FILLER_196_2243 ();
 b15zdnd11an1n04x5 FILLER_196_2248 ();
 b15zdnd11an1n04x5 FILLER_196_2256 ();
 b15zdnd11an1n04x5 FILLER_196_2264 ();
 b15zdnd11an1n04x5 FILLER_196_2272 ();
 b15zdnd11an1n64x5 FILLER_197_0 ();
 b15zdnd11an1n64x5 FILLER_197_64 ();
 b15zdnd11an1n64x5 FILLER_197_128 ();
 b15zdnd11an1n64x5 FILLER_197_192 ();
 b15zdnd00an1n02x5 FILLER_197_256 ();
 b15zdnd11an1n32x5 FILLER_197_285 ();
 b15zdnd00an1n02x5 FILLER_197_317 ();
 b15zdnd00an1n01x5 FILLER_197_319 ();
 b15zdnd11an1n04x5 FILLER_197_323 ();
 b15zdnd11an1n04x5 FILLER_197_330 ();
 b15zdnd11an1n64x5 FILLER_197_337 ();
 b15zdnd11an1n04x5 FILLER_197_401 ();
 b15zdnd00an1n02x5 FILLER_197_405 ();
 b15zdnd11an1n08x5 FILLER_197_410 ();
 b15zdnd11an1n04x5 FILLER_197_460 ();
 b15zdnd11an1n64x5 FILLER_197_516 ();
 b15zdnd11an1n16x5 FILLER_197_580 ();
 b15zdnd11an1n64x5 FILLER_197_638 ();
 b15zdnd11an1n64x5 FILLER_197_702 ();
 b15zdnd11an1n16x5 FILLER_197_766 ();
 b15zdnd11an1n08x5 FILLER_197_782 ();
 b15zdnd11an1n04x5 FILLER_197_790 ();
 b15zdnd11an1n04x5 FILLER_197_797 ();
 b15zdnd11an1n64x5 FILLER_197_804 ();
 b15zdnd11an1n64x5 FILLER_197_868 ();
 b15zdnd11an1n08x5 FILLER_197_932 ();
 b15zdnd11an1n16x5 FILLER_197_951 ();
 b15zdnd11an1n04x5 FILLER_197_967 ();
 b15zdnd00an1n01x5 FILLER_197_971 ();
 b15zdnd11an1n08x5 FILLER_197_984 ();
 b15zdnd11an1n04x5 FILLER_197_992 ();
 b15zdnd00an1n02x5 FILLER_197_996 ();
 b15zdnd00an1n01x5 FILLER_197_998 ();
 b15zdnd11an1n08x5 FILLER_197_1010 ();
 b15zdnd11an1n04x5 FILLER_197_1018 ();
 b15zdnd00an1n01x5 FILLER_197_1022 ();
 b15zdnd11an1n64x5 FILLER_197_1027 ();
 b15zdnd11an1n32x5 FILLER_197_1091 ();
 b15zdnd11an1n08x5 FILLER_197_1123 ();
 b15zdnd11an1n04x5 FILLER_197_1131 ();
 b15zdnd00an1n01x5 FILLER_197_1135 ();
 b15zdnd11an1n08x5 FILLER_197_1156 ();
 b15zdnd11an1n04x5 FILLER_197_1164 ();
 b15zdnd00an1n02x5 FILLER_197_1168 ();
 b15zdnd11an1n64x5 FILLER_197_1176 ();
 b15zdnd11an1n16x5 FILLER_197_1240 ();
 b15zdnd00an1n02x5 FILLER_197_1256 ();
 b15zdnd11an1n04x5 FILLER_197_1261 ();
 b15zdnd11an1n64x5 FILLER_197_1268 ();
 b15zdnd11an1n64x5 FILLER_197_1332 ();
 b15zdnd11an1n32x5 FILLER_197_1396 ();
 b15zdnd11an1n04x5 FILLER_197_1428 ();
 b15zdnd11an1n64x5 FILLER_197_1441 ();
 b15zdnd11an1n64x5 FILLER_197_1505 ();
 b15zdnd11an1n16x5 FILLER_197_1621 ();
 b15zdnd11an1n04x5 FILLER_197_1637 ();
 b15zdnd00an1n01x5 FILLER_197_1641 ();
 b15zdnd11an1n64x5 FILLER_197_1645 ();
 b15zdnd11an1n64x5 FILLER_197_1709 ();
 b15zdnd11an1n64x5 FILLER_197_1773 ();
 b15zdnd11an1n64x5 FILLER_197_1837 ();
 b15zdnd11an1n64x5 FILLER_197_1901 ();
 b15zdnd11an1n32x5 FILLER_197_1965 ();
 b15zdnd11an1n16x5 FILLER_197_1997 ();
 b15zdnd00an1n01x5 FILLER_197_2013 ();
 b15zdnd11an1n64x5 FILLER_197_2066 ();
 b15zdnd11an1n08x5 FILLER_197_2130 ();
 b15zdnd00an1n02x5 FILLER_197_2138 ();
 b15zdnd11an1n04x5 FILLER_197_2182 ();
 b15zdnd11an1n08x5 FILLER_197_2228 ();
 b15zdnd11an1n04x5 FILLER_197_2236 ();
 b15zdnd00an1n02x5 FILLER_197_2282 ();
 b15zdnd11an1n64x5 FILLER_198_8 ();
 b15zdnd11an1n64x5 FILLER_198_72 ();
 b15zdnd11an1n64x5 FILLER_198_136 ();
 b15zdnd11an1n32x5 FILLER_198_200 ();
 b15zdnd11an1n16x5 FILLER_198_232 ();
 b15zdnd11an1n08x5 FILLER_198_248 ();
 b15zdnd00an1n02x5 FILLER_198_256 ();
 b15zdnd11an1n64x5 FILLER_198_261 ();
 b15zdnd11an1n64x5 FILLER_198_325 ();
 b15zdnd11an1n32x5 FILLER_198_389 ();
 b15zdnd11an1n16x5 FILLER_198_421 ();
 b15zdnd11an1n04x5 FILLER_198_437 ();
 b15zdnd00an1n02x5 FILLER_198_441 ();
 b15zdnd11an1n04x5 FILLER_198_495 ();
 b15zdnd11an1n16x5 FILLER_198_502 ();
 b15zdnd00an1n02x5 FILLER_198_518 ();
 b15zdnd00an1n01x5 FILLER_198_520 ();
 b15zdnd11an1n64x5 FILLER_198_529 ();
 b15zdnd11an1n32x5 FILLER_198_593 ();
 b15zdnd11an1n16x5 FILLER_198_625 ();
 b15zdnd11an1n04x5 FILLER_198_641 ();
 b15zdnd00an1n01x5 FILLER_198_645 ();
 b15zdnd11an1n16x5 FILLER_198_688 ();
 b15zdnd11an1n08x5 FILLER_198_704 ();
 b15zdnd11an1n04x5 FILLER_198_712 ();
 b15zdnd00an1n02x5 FILLER_198_716 ();
 b15zdnd11an1n64x5 FILLER_198_726 ();
 b15zdnd11an1n64x5 FILLER_198_790 ();
 b15zdnd11an1n64x5 FILLER_198_854 ();
 b15zdnd11an1n32x5 FILLER_198_918 ();
 b15zdnd11an1n16x5 FILLER_198_950 ();
 b15zdnd00an1n02x5 FILLER_198_966 ();
 b15zdnd00an1n01x5 FILLER_198_968 ();
 b15zdnd11an1n16x5 FILLER_198_1003 ();
 b15zdnd11an1n04x5 FILLER_198_1019 ();
 b15zdnd11an1n64x5 FILLER_198_1034 ();
 b15zdnd11an1n16x5 FILLER_198_1098 ();
 b15zdnd11an1n08x5 FILLER_198_1114 ();
 b15zdnd00an1n02x5 FILLER_198_1122 ();
 b15zdnd00an1n01x5 FILLER_198_1124 ();
 b15zdnd11an1n64x5 FILLER_198_1170 ();
 b15zdnd11an1n04x5 FILLER_198_1234 ();
 b15zdnd00an1n02x5 FILLER_198_1238 ();
 b15zdnd11an1n64x5 FILLER_198_1292 ();
 b15zdnd11an1n64x5 FILLER_198_1356 ();
 b15zdnd11an1n64x5 FILLER_198_1420 ();
 b15zdnd11an1n64x5 FILLER_198_1484 ();
 b15zdnd11an1n32x5 FILLER_198_1548 ();
 b15zdnd11an1n04x5 FILLER_198_1580 ();
 b15zdnd00an1n02x5 FILLER_198_1584 ();
 b15zdnd00an1n01x5 FILLER_198_1586 ();
 b15zdnd11an1n04x5 FILLER_198_1590 ();
 b15zdnd11an1n64x5 FILLER_198_1597 ();
 b15zdnd11an1n64x5 FILLER_198_1661 ();
 b15zdnd11an1n64x5 FILLER_198_1725 ();
 b15zdnd11an1n64x5 FILLER_198_1789 ();
 b15zdnd11an1n64x5 FILLER_198_1853 ();
 b15zdnd11an1n64x5 FILLER_198_1917 ();
 b15zdnd11an1n32x5 FILLER_198_1981 ();
 b15zdnd11an1n04x5 FILLER_198_2013 ();
 b15zdnd11an1n04x5 FILLER_198_2024 ();
 b15zdnd11an1n64x5 FILLER_198_2073 ();
 b15zdnd11an1n16x5 FILLER_198_2137 ();
 b15zdnd00an1n01x5 FILLER_198_2153 ();
 b15zdnd11an1n32x5 FILLER_198_2162 ();
 b15zdnd11an1n16x5 FILLER_198_2194 ();
 b15zdnd11an1n08x5 FILLER_198_2210 ();
 b15zdnd00an1n02x5 FILLER_198_2218 ();
 b15zdnd11an1n04x5 FILLER_198_2227 ();
 b15zdnd00an1n01x5 FILLER_198_2231 ();
 b15zdnd00an1n02x5 FILLER_198_2274 ();
 b15zdnd11an1n64x5 FILLER_199_0 ();
 b15zdnd11an1n64x5 FILLER_199_64 ();
 b15zdnd11an1n64x5 FILLER_199_128 ();
 b15zdnd11an1n64x5 FILLER_199_192 ();
 b15zdnd11an1n64x5 FILLER_199_256 ();
 b15zdnd11an1n64x5 FILLER_199_320 ();
 b15zdnd11an1n64x5 FILLER_199_384 ();
 b15zdnd11an1n08x5 FILLER_199_448 ();
 b15zdnd11an1n04x5 FILLER_199_456 ();
 b15zdnd00an1n02x5 FILLER_199_460 ();
 b15zdnd11an1n04x5 FILLER_199_465 ();
 b15zdnd11an1n32x5 FILLER_199_511 ();
 b15zdnd11an1n16x5 FILLER_199_543 ();
 b15zdnd11an1n04x5 FILLER_199_559 ();
 b15zdnd00an1n01x5 FILLER_199_563 ();
 b15zdnd11an1n04x5 FILLER_199_606 ();
 b15zdnd11an1n64x5 FILLER_199_627 ();
 b15zdnd11an1n64x5 FILLER_199_733 ();
 b15zdnd11an1n64x5 FILLER_199_797 ();
 b15zdnd11an1n64x5 FILLER_199_861 ();
 b15zdnd11an1n04x5 FILLER_199_925 ();
 b15zdnd00an1n02x5 FILLER_199_929 ();
 b15zdnd00an1n01x5 FILLER_199_931 ();
 b15zdnd11an1n04x5 FILLER_199_974 ();
 b15zdnd00an1n02x5 FILLER_199_978 ();
 b15zdnd00an1n01x5 FILLER_199_980 ();
 b15zdnd11an1n64x5 FILLER_199_992 ();
 b15zdnd11an1n64x5 FILLER_199_1056 ();
 b15zdnd11an1n32x5 FILLER_199_1120 ();
 b15zdnd11an1n16x5 FILLER_199_1152 ();
 b15zdnd11an1n04x5 FILLER_199_1168 ();
 b15zdnd00an1n01x5 FILLER_199_1172 ();
 b15zdnd11an1n64x5 FILLER_199_1184 ();
 b15zdnd11an1n16x5 FILLER_199_1248 ();
 b15zdnd11an1n04x5 FILLER_199_1267 ();
 b15zdnd11an1n64x5 FILLER_199_1297 ();
 b15zdnd11an1n64x5 FILLER_199_1361 ();
 b15zdnd11an1n64x5 FILLER_199_1425 ();
 b15zdnd11an1n64x5 FILLER_199_1489 ();
 b15zdnd11an1n32x5 FILLER_199_1553 ();
 b15zdnd11an1n04x5 FILLER_199_1585 ();
 b15zdnd00an1n02x5 FILLER_199_1589 ();
 b15zdnd00an1n01x5 FILLER_199_1591 ();
 b15zdnd11an1n64x5 FILLER_199_1595 ();
 b15zdnd11an1n64x5 FILLER_199_1659 ();
 b15zdnd11an1n64x5 FILLER_199_1723 ();
 b15zdnd11an1n64x5 FILLER_199_1787 ();
 b15zdnd11an1n64x5 FILLER_199_1851 ();
 b15zdnd11an1n32x5 FILLER_199_1915 ();
 b15zdnd11an1n16x5 FILLER_199_1947 ();
 b15zdnd11an1n04x5 FILLER_199_1963 ();
 b15zdnd00an1n02x5 FILLER_199_1967 ();
 b15zdnd11an1n04x5 FILLER_199_2011 ();
 b15zdnd00an1n02x5 FILLER_199_2015 ();
 b15zdnd11an1n16x5 FILLER_199_2059 ();
 b15zdnd11an1n08x5 FILLER_199_2075 ();
 b15zdnd11an1n04x5 FILLER_199_2083 ();
 b15zdnd00an1n02x5 FILLER_199_2087 ();
 b15zdnd00an1n01x5 FILLER_199_2089 ();
 b15zdnd11an1n64x5 FILLER_199_2097 ();
 b15zdnd11an1n16x5 FILLER_199_2161 ();
 b15zdnd11an1n08x5 FILLER_199_2177 ();
 b15zdnd00an1n02x5 FILLER_199_2185 ();
 b15zdnd00an1n01x5 FILLER_199_2187 ();
 b15zdnd11an1n16x5 FILLER_199_2219 ();
 b15zdnd11an1n04x5 FILLER_199_2235 ();
 b15zdnd00an1n01x5 FILLER_199_2239 ();
 b15zdnd00an1n02x5 FILLER_199_2282 ();
 b15zdnd11an1n64x5 FILLER_200_8 ();
 b15zdnd11an1n64x5 FILLER_200_72 ();
 b15zdnd11an1n32x5 FILLER_200_136 ();
 b15zdnd11an1n08x5 FILLER_200_168 ();
 b15zdnd00an1n02x5 FILLER_200_176 ();
 b15zdnd00an1n01x5 FILLER_200_178 ();
 b15zdnd11an1n64x5 FILLER_200_206 ();
 b15zdnd11an1n64x5 FILLER_200_270 ();
 b15zdnd11an1n64x5 FILLER_200_334 ();
 b15zdnd11an1n64x5 FILLER_200_398 ();
 b15zdnd11an1n08x5 FILLER_200_462 ();
 b15zdnd11an1n04x5 FILLER_200_477 ();
 b15zdnd00an1n02x5 FILLER_200_481 ();
 b15zdnd00an1n01x5 FILLER_200_483 ();
 b15zdnd11an1n64x5 FILLER_200_487 ();
 b15zdnd11an1n32x5 FILLER_200_551 ();
 b15zdnd11an1n08x5 FILLER_200_583 ();
 b15zdnd11an1n04x5 FILLER_200_591 ();
 b15zdnd00an1n02x5 FILLER_200_595 ();
 b15zdnd00an1n01x5 FILLER_200_597 ();
 b15zdnd11an1n64x5 FILLER_200_605 ();
 b15zdnd11an1n32x5 FILLER_200_669 ();
 b15zdnd11an1n16x5 FILLER_200_701 ();
 b15zdnd00an1n01x5 FILLER_200_717 ();
 b15zdnd11an1n64x5 FILLER_200_726 ();
 b15zdnd11an1n64x5 FILLER_200_790 ();
 b15zdnd11an1n64x5 FILLER_200_854 ();
 b15zdnd11an1n08x5 FILLER_200_918 ();
 b15zdnd11an1n04x5 FILLER_200_926 ();
 b15zdnd00an1n02x5 FILLER_200_930 ();
 b15zdnd00an1n01x5 FILLER_200_932 ();
 b15zdnd11an1n32x5 FILLER_200_940 ();
 b15zdnd11an1n16x5 FILLER_200_972 ();
 b15zdnd11an1n16x5 FILLER_200_997 ();
 b15zdnd00an1n02x5 FILLER_200_1013 ();
 b15zdnd11an1n08x5 FILLER_200_1029 ();
 b15zdnd00an1n02x5 FILLER_200_1037 ();
 b15zdnd00an1n01x5 FILLER_200_1039 ();
 b15zdnd11an1n04x5 FILLER_200_1050 ();
 b15zdnd11an1n32x5 FILLER_200_1085 ();
 b15zdnd11an1n16x5 FILLER_200_1117 ();
 b15zdnd00an1n02x5 FILLER_200_1133 ();
 b15zdnd11an1n64x5 FILLER_200_1140 ();
 b15zdnd11an1n16x5 FILLER_200_1204 ();
 b15zdnd11an1n08x5 FILLER_200_1220 ();
 b15zdnd00an1n01x5 FILLER_200_1228 ();
 b15zdnd11an1n04x5 FILLER_200_1241 ();
 b15zdnd11an1n64x5 FILLER_200_1262 ();
 b15zdnd11an1n64x5 FILLER_200_1326 ();
 b15zdnd11an1n64x5 FILLER_200_1390 ();
 b15zdnd11an1n32x5 FILLER_200_1454 ();
 b15zdnd11an1n08x5 FILLER_200_1486 ();
 b15zdnd11an1n04x5 FILLER_200_1494 ();
 b15zdnd11an1n64x5 FILLER_200_1515 ();
 b15zdnd11an1n64x5 FILLER_200_1579 ();
 b15zdnd11an1n64x5 FILLER_200_1643 ();
 b15zdnd11an1n64x5 FILLER_200_1707 ();
 b15zdnd11an1n64x5 FILLER_200_1771 ();
 b15zdnd11an1n64x5 FILLER_200_1835 ();
 b15zdnd11an1n64x5 FILLER_200_1899 ();
 b15zdnd11an1n32x5 FILLER_200_1963 ();
 b15zdnd00an1n02x5 FILLER_200_1995 ();
 b15zdnd00an1n01x5 FILLER_200_1997 ();
 b15zdnd11an1n04x5 FILLER_200_2040 ();
 b15zdnd00an1n02x5 FILLER_200_2044 ();
 b15zdnd11an1n64x5 FILLER_200_2049 ();
 b15zdnd11an1n32x5 FILLER_200_2113 ();
 b15zdnd11an1n08x5 FILLER_200_2145 ();
 b15zdnd00an1n01x5 FILLER_200_2153 ();
 b15zdnd11an1n64x5 FILLER_200_2162 ();
 b15zdnd11an1n04x5 FILLER_200_2226 ();
 b15zdnd00an1n02x5 FILLER_200_2230 ();
 b15zdnd00an1n02x5 FILLER_200_2274 ();
 b15zdnd11an1n64x5 FILLER_201_0 ();
 b15zdnd11an1n64x5 FILLER_201_64 ();
 b15zdnd11an1n32x5 FILLER_201_128 ();
 b15zdnd11an1n16x5 FILLER_201_160 ();
 b15zdnd00an1n02x5 FILLER_201_176 ();
 b15zdnd11an1n64x5 FILLER_201_181 ();
 b15zdnd11an1n64x5 FILLER_201_245 ();
 b15zdnd11an1n64x5 FILLER_201_309 ();
 b15zdnd11an1n64x5 FILLER_201_373 ();
 b15zdnd11an1n64x5 FILLER_201_437 ();
 b15zdnd11an1n64x5 FILLER_201_501 ();
 b15zdnd11an1n32x5 FILLER_201_565 ();
 b15zdnd11an1n16x5 FILLER_201_597 ();
 b15zdnd11an1n08x5 FILLER_201_613 ();
 b15zdnd00an1n02x5 FILLER_201_621 ();
 b15zdnd00an1n01x5 FILLER_201_623 ();
 b15zdnd11an1n64x5 FILLER_201_666 ();
 b15zdnd11an1n64x5 FILLER_201_730 ();
 b15zdnd11an1n64x5 FILLER_201_794 ();
 b15zdnd11an1n64x5 FILLER_201_858 ();
 b15zdnd11an1n32x5 FILLER_201_922 ();
 b15zdnd11an1n04x5 FILLER_201_954 ();
 b15zdnd00an1n02x5 FILLER_201_958 ();
 b15zdnd00an1n01x5 FILLER_201_960 ();
 b15zdnd11an1n16x5 FILLER_201_993 ();
 b15zdnd11an1n08x5 FILLER_201_1009 ();
 b15zdnd00an1n02x5 FILLER_201_1017 ();
 b15zdnd11an1n04x5 FILLER_201_1030 ();
 b15zdnd11an1n04x5 FILLER_201_1062 ();
 b15zdnd11an1n64x5 FILLER_201_1077 ();
 b15zdnd11an1n64x5 FILLER_201_1141 ();
 b15zdnd11an1n16x5 FILLER_201_1205 ();
 b15zdnd11an1n04x5 FILLER_201_1221 ();
 b15zdnd11an1n64x5 FILLER_201_1245 ();
 b15zdnd11an1n08x5 FILLER_201_1309 ();
 b15zdnd11an1n04x5 FILLER_201_1317 ();
 b15zdnd11an1n32x5 FILLER_201_1331 ();
 b15zdnd11an1n64x5 FILLER_201_1377 ();
 b15zdnd11an1n64x5 FILLER_201_1441 ();
 b15zdnd11an1n64x5 FILLER_201_1505 ();
 b15zdnd00an1n01x5 FILLER_201_1569 ();
 b15zdnd11an1n64x5 FILLER_201_1587 ();
 b15zdnd11an1n64x5 FILLER_201_1651 ();
 b15zdnd11an1n64x5 FILLER_201_1715 ();
 b15zdnd11an1n64x5 FILLER_201_1779 ();
 b15zdnd11an1n64x5 FILLER_201_1843 ();
 b15zdnd11an1n32x5 FILLER_201_1907 ();
 b15zdnd11an1n16x5 FILLER_201_1939 ();
 b15zdnd11an1n08x5 FILLER_201_1955 ();
 b15zdnd11an1n04x5 FILLER_201_1963 ();
 b15zdnd00an1n01x5 FILLER_201_1967 ();
 b15zdnd11an1n08x5 FILLER_201_2010 ();
 b15zdnd11an1n04x5 FILLER_201_2018 ();
 b15zdnd00an1n02x5 FILLER_201_2022 ();
 b15zdnd11an1n04x5 FILLER_201_2030 ();
 b15zdnd11an1n64x5 FILLER_201_2037 ();
 b15zdnd11an1n64x5 FILLER_201_2101 ();
 b15zdnd11an1n64x5 FILLER_201_2165 ();
 b15zdnd11an1n16x5 FILLER_201_2229 ();
 b15zdnd11an1n08x5 FILLER_201_2245 ();
 b15zdnd11an1n04x5 FILLER_201_2253 ();
 b15zdnd00an1n02x5 FILLER_201_2257 ();
 b15zdnd00an1n01x5 FILLER_201_2259 ();
 b15zdnd11an1n04x5 FILLER_201_2264 ();
 b15zdnd11an1n08x5 FILLER_201_2272 ();
 b15zdnd11an1n04x5 FILLER_201_2280 ();
 b15zdnd11an1n64x5 FILLER_202_8 ();
 b15zdnd11an1n64x5 FILLER_202_72 ();
 b15zdnd11an1n64x5 FILLER_202_136 ();
 b15zdnd11an1n64x5 FILLER_202_200 ();
 b15zdnd11an1n64x5 FILLER_202_264 ();
 b15zdnd11an1n32x5 FILLER_202_328 ();
 b15zdnd11an1n16x5 FILLER_202_360 ();
 b15zdnd00an1n01x5 FILLER_202_376 ();
 b15zdnd11an1n64x5 FILLER_202_386 ();
 b15zdnd11an1n16x5 FILLER_202_450 ();
 b15zdnd11an1n04x5 FILLER_202_466 ();
 b15zdnd00an1n02x5 FILLER_202_470 ();
 b15zdnd00an1n01x5 FILLER_202_472 ();
 b15zdnd11an1n08x5 FILLER_202_515 ();
 b15zdnd00an1n01x5 FILLER_202_523 ();
 b15zdnd11an1n64x5 FILLER_202_532 ();
 b15zdnd11an1n64x5 FILLER_202_596 ();
 b15zdnd11an1n32x5 FILLER_202_660 ();
 b15zdnd11an1n16x5 FILLER_202_692 ();
 b15zdnd11an1n08x5 FILLER_202_708 ();
 b15zdnd00an1n02x5 FILLER_202_716 ();
 b15zdnd11an1n64x5 FILLER_202_726 ();
 b15zdnd11an1n64x5 FILLER_202_790 ();
 b15zdnd11an1n64x5 FILLER_202_854 ();
 b15zdnd11an1n08x5 FILLER_202_918 ();
 b15zdnd00an1n02x5 FILLER_202_926 ();
 b15zdnd11an1n32x5 FILLER_202_939 ();
 b15zdnd11an1n16x5 FILLER_202_971 ();
 b15zdnd11an1n08x5 FILLER_202_987 ();
 b15zdnd11an1n04x5 FILLER_202_995 ();
 b15zdnd11an1n32x5 FILLER_202_1027 ();
 b15zdnd11an1n08x5 FILLER_202_1059 ();
 b15zdnd11an1n04x5 FILLER_202_1067 ();
 b15zdnd11an1n64x5 FILLER_202_1080 ();
 b15zdnd11an1n64x5 FILLER_202_1144 ();
 b15zdnd11an1n64x5 FILLER_202_1208 ();
 b15zdnd11an1n04x5 FILLER_202_1272 ();
 b15zdnd11an1n16x5 FILLER_202_1308 ();
 b15zdnd11an1n64x5 FILLER_202_1331 ();
 b15zdnd11an1n64x5 FILLER_202_1395 ();
 b15zdnd11an1n64x5 FILLER_202_1459 ();
 b15zdnd11an1n64x5 FILLER_202_1523 ();
 b15zdnd11an1n32x5 FILLER_202_1587 ();
 b15zdnd11an1n08x5 FILLER_202_1619 ();
 b15zdnd11an1n64x5 FILLER_202_1636 ();
 b15zdnd11an1n16x5 FILLER_202_1700 ();
 b15zdnd11an1n08x5 FILLER_202_1716 ();
 b15zdnd11an1n04x5 FILLER_202_1724 ();
 b15zdnd00an1n02x5 FILLER_202_1728 ();
 b15zdnd11an1n64x5 FILLER_202_1750 ();
 b15zdnd11an1n64x5 FILLER_202_1814 ();
 b15zdnd11an1n64x5 FILLER_202_1878 ();
 b15zdnd11an1n32x5 FILLER_202_1942 ();
 b15zdnd11an1n16x5 FILLER_202_1974 ();
 b15zdnd11an1n04x5 FILLER_202_1990 ();
 b15zdnd00an1n02x5 FILLER_202_1994 ();
 b15zdnd00an1n01x5 FILLER_202_1996 ();
 b15zdnd11an1n16x5 FILLER_202_2039 ();
 b15zdnd11an1n04x5 FILLER_202_2055 ();
 b15zdnd11an1n04x5 FILLER_202_2062 ();
 b15zdnd11an1n32x5 FILLER_202_2069 ();
 b15zdnd11an1n16x5 FILLER_202_2101 ();
 b15zdnd11an1n08x5 FILLER_202_2117 ();
 b15zdnd00an1n02x5 FILLER_202_2125 ();
 b15zdnd11an1n04x5 FILLER_202_2136 ();
 b15zdnd11an1n04x5 FILLER_202_2149 ();
 b15zdnd00an1n01x5 FILLER_202_2153 ();
 b15zdnd11an1n64x5 FILLER_202_2162 ();
 b15zdnd11an1n04x5 FILLER_202_2226 ();
 b15zdnd00an1n02x5 FILLER_202_2230 ();
 b15zdnd00an1n02x5 FILLER_202_2274 ();
 b15zdnd11an1n64x5 FILLER_203_0 ();
 b15zdnd11an1n08x5 FILLER_203_64 ();
 b15zdnd11an1n04x5 FILLER_203_72 ();
 b15zdnd00an1n02x5 FILLER_203_76 ();
 b15zdnd00an1n01x5 FILLER_203_78 ();
 b15zdnd11an1n64x5 FILLER_203_89 ();
 b15zdnd11an1n64x5 FILLER_203_153 ();
 b15zdnd11an1n64x5 FILLER_203_217 ();
 b15zdnd11an1n64x5 FILLER_203_281 ();
 b15zdnd11an1n64x5 FILLER_203_345 ();
 b15zdnd11an1n64x5 FILLER_203_409 ();
 b15zdnd11an1n64x5 FILLER_203_473 ();
 b15zdnd11an1n64x5 FILLER_203_537 ();
 b15zdnd11an1n64x5 FILLER_203_601 ();
 b15zdnd11an1n64x5 FILLER_203_665 ();
 b15zdnd11an1n64x5 FILLER_203_729 ();
 b15zdnd11an1n64x5 FILLER_203_793 ();
 b15zdnd11an1n64x5 FILLER_203_857 ();
 b15zdnd11an1n64x5 FILLER_203_921 ();
 b15zdnd11an1n64x5 FILLER_203_985 ();
 b15zdnd11an1n64x5 FILLER_203_1049 ();
 b15zdnd11an1n64x5 FILLER_203_1113 ();
 b15zdnd11an1n64x5 FILLER_203_1177 ();
 b15zdnd11an1n32x5 FILLER_203_1241 ();
 b15zdnd11an1n16x5 FILLER_203_1273 ();
 b15zdnd00an1n02x5 FILLER_203_1289 ();
 b15zdnd11an1n16x5 FILLER_203_1311 ();
 b15zdnd11an1n08x5 FILLER_203_1327 ();
 b15zdnd11an1n04x5 FILLER_203_1335 ();
 b15zdnd11an1n16x5 FILLER_203_1359 ();
 b15zdnd11an1n08x5 FILLER_203_1375 ();
 b15zdnd11an1n04x5 FILLER_203_1383 ();
 b15zdnd00an1n01x5 FILLER_203_1387 ();
 b15zdnd11an1n64x5 FILLER_203_1402 ();
 b15zdnd11an1n64x5 FILLER_203_1466 ();
 b15zdnd11an1n64x5 FILLER_203_1530 ();
 b15zdnd11an1n64x5 FILLER_203_1594 ();
 b15zdnd11an1n32x5 FILLER_203_1658 ();
 b15zdnd11an1n16x5 FILLER_203_1690 ();
 b15zdnd11an1n04x5 FILLER_203_1706 ();
 b15zdnd11an1n64x5 FILLER_203_1713 ();
 b15zdnd11an1n64x5 FILLER_203_1777 ();
 b15zdnd11an1n64x5 FILLER_203_1841 ();
 b15zdnd11an1n16x5 FILLER_203_1905 ();
 b15zdnd11an1n04x5 FILLER_203_1924 ();
 b15zdnd11an1n64x5 FILLER_203_1931 ();
 b15zdnd11an1n32x5 FILLER_203_1995 ();
 b15zdnd11an1n08x5 FILLER_203_2027 ();
 b15zdnd11an1n04x5 FILLER_203_2035 ();
 b15zdnd00an1n02x5 FILLER_203_2039 ();
 b15zdnd11an1n64x5 FILLER_203_2093 ();
 b15zdnd11an1n64x5 FILLER_203_2157 ();
 b15zdnd11an1n16x5 FILLER_203_2221 ();
 b15zdnd00an1n02x5 FILLER_203_2237 ();
 b15zdnd00an1n01x5 FILLER_203_2239 ();
 b15zdnd00an1n02x5 FILLER_203_2282 ();
 b15zdnd11an1n32x5 FILLER_204_8 ();
 b15zdnd11an1n16x5 FILLER_204_40 ();
 b15zdnd11an1n08x5 FILLER_204_56 ();
 b15zdnd00an1n01x5 FILLER_204_64 ();
 b15zdnd11an1n64x5 FILLER_204_69 ();
 b15zdnd11an1n16x5 FILLER_204_133 ();
 b15zdnd11an1n08x5 FILLER_204_149 ();
 b15zdnd00an1n01x5 FILLER_204_157 ();
 b15zdnd11an1n64x5 FILLER_204_161 ();
 b15zdnd11an1n64x5 FILLER_204_225 ();
 b15zdnd11an1n64x5 FILLER_204_289 ();
 b15zdnd11an1n64x5 FILLER_204_353 ();
 b15zdnd11an1n64x5 FILLER_204_417 ();
 b15zdnd11an1n32x5 FILLER_204_481 ();
 b15zdnd11an1n16x5 FILLER_204_513 ();
 b15zdnd11an1n04x5 FILLER_204_529 ();
 b15zdnd00an1n02x5 FILLER_204_533 ();
 b15zdnd00an1n01x5 FILLER_204_535 ();
 b15zdnd11an1n64x5 FILLER_204_578 ();
 b15zdnd11an1n32x5 FILLER_204_642 ();
 b15zdnd11an1n16x5 FILLER_204_674 ();
 b15zdnd11an1n04x5 FILLER_204_690 ();
 b15zdnd00an1n02x5 FILLER_204_716 ();
 b15zdnd11an1n64x5 FILLER_204_726 ();
 b15zdnd11an1n64x5 FILLER_204_790 ();
 b15zdnd11an1n16x5 FILLER_204_854 ();
 b15zdnd11an1n04x5 FILLER_204_870 ();
 b15zdnd00an1n01x5 FILLER_204_874 ();
 b15zdnd11an1n64x5 FILLER_204_893 ();
 b15zdnd11an1n64x5 FILLER_204_957 ();
 b15zdnd11an1n64x5 FILLER_204_1021 ();
 b15zdnd11an1n64x5 FILLER_204_1085 ();
 b15zdnd11an1n64x5 FILLER_204_1149 ();
 b15zdnd11an1n64x5 FILLER_204_1213 ();
 b15zdnd11an1n64x5 FILLER_204_1277 ();
 b15zdnd11an1n32x5 FILLER_204_1341 ();
 b15zdnd11an1n16x5 FILLER_204_1373 ();
 b15zdnd11an1n08x5 FILLER_204_1389 ();
 b15zdnd11an1n04x5 FILLER_204_1397 ();
 b15zdnd00an1n02x5 FILLER_204_1401 ();
 b15zdnd11an1n64x5 FILLER_204_1423 ();
 b15zdnd11an1n64x5 FILLER_204_1487 ();
 b15zdnd11an1n64x5 FILLER_204_1551 ();
 b15zdnd11an1n64x5 FILLER_204_1615 ();
 b15zdnd11an1n32x5 FILLER_204_1679 ();
 b15zdnd11an1n64x5 FILLER_204_1714 ();
 b15zdnd11an1n32x5 FILLER_204_1778 ();
 b15zdnd11an1n04x5 FILLER_204_1810 ();
 b15zdnd00an1n01x5 FILLER_204_1814 ();
 b15zdnd11an1n04x5 FILLER_204_1818 ();
 b15zdnd11an1n16x5 FILLER_204_1874 ();
 b15zdnd11an1n08x5 FILLER_204_1890 ();
 b15zdnd00an1n02x5 FILLER_204_1898 ();
 b15zdnd11an1n64x5 FILLER_204_1952 ();
 b15zdnd11an1n32x5 FILLER_204_2016 ();
 b15zdnd11an1n16x5 FILLER_204_2048 ();
 b15zdnd00an1n02x5 FILLER_204_2064 ();
 b15zdnd00an1n01x5 FILLER_204_2066 ();
 b15zdnd11an1n64x5 FILLER_204_2070 ();
 b15zdnd11an1n16x5 FILLER_204_2134 ();
 b15zdnd11an1n04x5 FILLER_204_2150 ();
 b15zdnd11an1n32x5 FILLER_204_2162 ();
 b15zdnd11an1n08x5 FILLER_204_2194 ();
 b15zdnd00an1n01x5 FILLER_204_2202 ();
 b15zdnd11an1n16x5 FILLER_204_2208 ();
 b15zdnd11an1n08x5 FILLER_204_2224 ();
 b15zdnd00an1n02x5 FILLER_204_2274 ();
 b15zdnd11an1n64x5 FILLER_205_0 ();
 b15zdnd11an1n32x5 FILLER_205_73 ();
 b15zdnd11an1n16x5 FILLER_205_105 ();
 b15zdnd11an1n08x5 FILLER_205_121 ();
 b15zdnd00an1n02x5 FILLER_205_129 ();
 b15zdnd11an1n04x5 FILLER_205_163 ();
 b15zdnd11an1n16x5 FILLER_205_170 ();
 b15zdnd11an1n04x5 FILLER_205_186 ();
 b15zdnd00an1n02x5 FILLER_205_190 ();
 b15zdnd11an1n64x5 FILLER_205_195 ();
 b15zdnd11an1n64x5 FILLER_205_259 ();
 b15zdnd11an1n64x5 FILLER_205_323 ();
 b15zdnd11an1n64x5 FILLER_205_387 ();
 b15zdnd11an1n64x5 FILLER_205_451 ();
 b15zdnd11an1n16x5 FILLER_205_515 ();
 b15zdnd11an1n08x5 FILLER_205_531 ();
 b15zdnd11an1n64x5 FILLER_205_546 ();
 b15zdnd11an1n64x5 FILLER_205_610 ();
 b15zdnd11an1n32x5 FILLER_205_674 ();
 b15zdnd11an1n16x5 FILLER_205_706 ();
 b15zdnd11an1n08x5 FILLER_205_722 ();
 b15zdnd00an1n02x5 FILLER_205_730 ();
 b15zdnd00an1n01x5 FILLER_205_732 ();
 b15zdnd11an1n04x5 FILLER_205_741 ();
 b15zdnd11an1n64x5 FILLER_205_759 ();
 b15zdnd11an1n64x5 FILLER_205_823 ();
 b15zdnd11an1n64x5 FILLER_205_887 ();
 b15zdnd11an1n64x5 FILLER_205_951 ();
 b15zdnd11an1n64x5 FILLER_205_1015 ();
 b15zdnd11an1n16x5 FILLER_205_1079 ();
 b15zdnd11an1n04x5 FILLER_205_1095 ();
 b15zdnd11an1n04x5 FILLER_205_1119 ();
 b15zdnd11an1n08x5 FILLER_205_1140 ();
 b15zdnd11an1n04x5 FILLER_205_1148 ();
 b15zdnd00an1n02x5 FILLER_205_1152 ();
 b15zdnd11an1n64x5 FILLER_205_1158 ();
 b15zdnd11an1n64x5 FILLER_205_1222 ();
 b15zdnd11an1n16x5 FILLER_205_1286 ();
 b15zdnd11an1n04x5 FILLER_205_1302 ();
 b15zdnd11an1n64x5 FILLER_205_1324 ();
 b15zdnd11an1n64x5 FILLER_205_1388 ();
 b15zdnd11an1n64x5 FILLER_205_1452 ();
 b15zdnd11an1n64x5 FILLER_205_1516 ();
 b15zdnd11an1n64x5 FILLER_205_1580 ();
 b15zdnd11an1n32x5 FILLER_205_1644 ();
 b15zdnd11an1n08x5 FILLER_205_1676 ();
 b15zdnd00an1n02x5 FILLER_205_1684 ();
 b15zdnd11an1n32x5 FILLER_205_1738 ();
 b15zdnd11an1n16x5 FILLER_205_1770 ();
 b15zdnd11an1n04x5 FILLER_205_1786 ();
 b15zdnd11an1n04x5 FILLER_205_1842 ();
 b15zdnd11an1n32x5 FILLER_205_1849 ();
 b15zdnd11an1n08x5 FILLER_205_1881 ();
 b15zdnd11an1n04x5 FILLER_205_1889 ();
 b15zdnd00an1n01x5 FILLER_205_1893 ();
 b15zdnd11an1n64x5 FILLER_205_1946 ();
 b15zdnd11an1n64x5 FILLER_205_2010 ();
 b15zdnd11an1n32x5 FILLER_205_2074 ();
 b15zdnd11an1n16x5 FILLER_205_2106 ();
 b15zdnd11an1n08x5 FILLER_205_2122 ();
 b15zdnd11an1n04x5 FILLER_205_2130 ();
 b15zdnd00an1n01x5 FILLER_205_2134 ();
 b15zdnd11an1n32x5 FILLER_205_2177 ();
 b15zdnd11an1n16x5 FILLER_205_2209 ();
 b15zdnd11an1n04x5 FILLER_205_2225 ();
 b15zdnd00an1n02x5 FILLER_205_2229 ();
 b15zdnd00an1n01x5 FILLER_205_2231 ();
 b15zdnd11an1n04x5 FILLER_205_2236 ();
 b15zdnd00an1n02x5 FILLER_205_2282 ();
 b15zdnd11an1n32x5 FILLER_206_8 ();
 b15zdnd11an1n16x5 FILLER_206_40 ();
 b15zdnd11an1n04x5 FILLER_206_65 ();
 b15zdnd11an1n64x5 FILLER_206_79 ();
 b15zdnd11an1n16x5 FILLER_206_143 ();
 b15zdnd11an1n04x5 FILLER_206_159 ();
 b15zdnd00an1n01x5 FILLER_206_163 ();
 b15zdnd11an1n04x5 FILLER_206_196 ();
 b15zdnd00an1n02x5 FILLER_206_200 ();
 b15zdnd11an1n64x5 FILLER_206_244 ();
 b15zdnd11an1n64x5 FILLER_206_308 ();
 b15zdnd11an1n64x5 FILLER_206_372 ();
 b15zdnd11an1n08x5 FILLER_206_436 ();
 b15zdnd11an1n04x5 FILLER_206_444 ();
 b15zdnd11an1n64x5 FILLER_206_490 ();
 b15zdnd00an1n02x5 FILLER_206_554 ();
 b15zdnd00an1n01x5 FILLER_206_556 ();
 b15zdnd11an1n16x5 FILLER_206_565 ();
 b15zdnd11an1n04x5 FILLER_206_581 ();
 b15zdnd11an1n64x5 FILLER_206_592 ();
 b15zdnd11an1n32x5 FILLER_206_656 ();
 b15zdnd11an1n16x5 FILLER_206_688 ();
 b15zdnd11an1n08x5 FILLER_206_704 ();
 b15zdnd11an1n04x5 FILLER_206_712 ();
 b15zdnd00an1n02x5 FILLER_206_716 ();
 b15zdnd11an1n64x5 FILLER_206_726 ();
 b15zdnd11an1n64x5 FILLER_206_790 ();
 b15zdnd11an1n64x5 FILLER_206_854 ();
 b15zdnd11an1n64x5 FILLER_206_918 ();
 b15zdnd11an1n32x5 FILLER_206_982 ();
 b15zdnd11an1n08x5 FILLER_206_1014 ();
 b15zdnd11an1n04x5 FILLER_206_1022 ();
 b15zdnd11an1n16x5 FILLER_206_1054 ();
 b15zdnd11an1n04x5 FILLER_206_1070 ();
 b15zdnd00an1n02x5 FILLER_206_1074 ();
 b15zdnd00an1n01x5 FILLER_206_1076 ();
 b15zdnd11an1n04x5 FILLER_206_1122 ();
 b15zdnd11an1n64x5 FILLER_206_1137 ();
 b15zdnd11an1n32x5 FILLER_206_1201 ();
 b15zdnd00an1n01x5 FILLER_206_1233 ();
 b15zdnd11an1n64x5 FILLER_206_1242 ();
 b15zdnd11an1n64x5 FILLER_206_1306 ();
 b15zdnd11an1n32x5 FILLER_206_1370 ();
 b15zdnd11an1n16x5 FILLER_206_1402 ();
 b15zdnd00an1n01x5 FILLER_206_1418 ();
 b15zdnd11an1n64x5 FILLER_206_1433 ();
 b15zdnd11an1n32x5 FILLER_206_1497 ();
 b15zdnd11an1n16x5 FILLER_206_1529 ();
 b15zdnd11an1n04x5 FILLER_206_1545 ();
 b15zdnd00an1n02x5 FILLER_206_1549 ();
 b15zdnd11an1n64x5 FILLER_206_1582 ();
 b15zdnd11an1n64x5 FILLER_206_1646 ();
 b15zdnd00an1n01x5 FILLER_206_1710 ();
 b15zdnd11an1n64x5 FILLER_206_1714 ();
 b15zdnd11an1n32x5 FILLER_206_1778 ();
 b15zdnd00an1n02x5 FILLER_206_1810 ();
 b15zdnd00an1n01x5 FILLER_206_1812 ();
 b15zdnd11an1n16x5 FILLER_206_1816 ();
 b15zdnd11an1n08x5 FILLER_206_1832 ();
 b15zdnd11an1n04x5 FILLER_206_1840 ();
 b15zdnd11an1n64x5 FILLER_206_1847 ();
 b15zdnd00an1n01x5 FILLER_206_1911 ();
 b15zdnd11an1n04x5 FILLER_206_1915 ();
 b15zdnd11an1n04x5 FILLER_206_1922 ();
 b15zdnd11an1n04x5 FILLER_206_1929 ();
 b15zdnd11an1n64x5 FILLER_206_1936 ();
 b15zdnd11an1n64x5 FILLER_206_2000 ();
 b15zdnd11an1n32x5 FILLER_206_2064 ();
 b15zdnd11an1n04x5 FILLER_206_2096 ();
 b15zdnd00an1n01x5 FILLER_206_2100 ();
 b15zdnd11an1n08x5 FILLER_206_2143 ();
 b15zdnd00an1n02x5 FILLER_206_2151 ();
 b15zdnd00an1n01x5 FILLER_206_2153 ();
 b15zdnd11an1n16x5 FILLER_206_2162 ();
 b15zdnd11an1n08x5 FILLER_206_2220 ();
 b15zdnd11an1n04x5 FILLER_206_2228 ();
 b15zdnd00an1n02x5 FILLER_206_2274 ();
 b15zdnd11an1n32x5 FILLER_207_0 ();
 b15zdnd11an1n16x5 FILLER_207_32 ();
 b15zdnd11an1n08x5 FILLER_207_48 ();
 b15zdnd00an1n01x5 FILLER_207_56 ();
 b15zdnd11an1n64x5 FILLER_207_73 ();
 b15zdnd11an1n16x5 FILLER_207_137 ();
 b15zdnd00an1n02x5 FILLER_207_153 ();
 b15zdnd11an1n16x5 FILLER_207_164 ();
 b15zdnd11an1n08x5 FILLER_207_180 ();
 b15zdnd11an1n04x5 FILLER_207_188 ();
 b15zdnd00an1n01x5 FILLER_207_192 ();
 b15zdnd11an1n64x5 FILLER_207_196 ();
 b15zdnd11an1n64x5 FILLER_207_260 ();
 b15zdnd11an1n64x5 FILLER_207_324 ();
 b15zdnd11an1n16x5 FILLER_207_388 ();
 b15zdnd11an1n08x5 FILLER_207_404 ();
 b15zdnd11an1n04x5 FILLER_207_412 ();
 b15zdnd00an1n02x5 FILLER_207_416 ();
 b15zdnd00an1n01x5 FILLER_207_418 ();
 b15zdnd11an1n04x5 FILLER_207_428 ();
 b15zdnd11an1n64x5 FILLER_207_441 ();
 b15zdnd11an1n64x5 FILLER_207_505 ();
 b15zdnd11an1n04x5 FILLER_207_569 ();
 b15zdnd00an1n02x5 FILLER_207_573 ();
 b15zdnd00an1n01x5 FILLER_207_575 ();
 b15zdnd11an1n64x5 FILLER_207_618 ();
 b15zdnd11an1n04x5 FILLER_207_682 ();
 b15zdnd00an1n02x5 FILLER_207_686 ();
 b15zdnd11an1n64x5 FILLER_207_730 ();
 b15zdnd11an1n64x5 FILLER_207_794 ();
 b15zdnd11an1n64x5 FILLER_207_858 ();
 b15zdnd11an1n64x5 FILLER_207_922 ();
 b15zdnd11an1n64x5 FILLER_207_986 ();
 b15zdnd11an1n08x5 FILLER_207_1050 ();
 b15zdnd11an1n04x5 FILLER_207_1058 ();
 b15zdnd00an1n01x5 FILLER_207_1062 ();
 b15zdnd11an1n16x5 FILLER_207_1074 ();
 b15zdnd11an1n08x5 FILLER_207_1090 ();
 b15zdnd11an1n04x5 FILLER_207_1098 ();
 b15zdnd11an1n16x5 FILLER_207_1106 ();
 b15zdnd11an1n04x5 FILLER_207_1122 ();
 b15zdnd11an1n64x5 FILLER_207_1147 ();
 b15zdnd11an1n64x5 FILLER_207_1211 ();
 b15zdnd11an1n64x5 FILLER_207_1275 ();
 b15zdnd11an1n64x5 FILLER_207_1339 ();
 b15zdnd11an1n64x5 FILLER_207_1403 ();
 b15zdnd11an1n64x5 FILLER_207_1467 ();
 b15zdnd11an1n64x5 FILLER_207_1531 ();
 b15zdnd11an1n64x5 FILLER_207_1595 ();
 b15zdnd11an1n64x5 FILLER_207_1659 ();
 b15zdnd11an1n64x5 FILLER_207_1723 ();
 b15zdnd11an1n16x5 FILLER_207_1787 ();
 b15zdnd11an1n08x5 FILLER_207_1803 ();
 b15zdnd00an1n02x5 FILLER_207_1811 ();
 b15zdnd11an1n16x5 FILLER_207_1816 ();
 b15zdnd11an1n08x5 FILLER_207_1832 ();
 b15zdnd00an1n02x5 FILLER_207_1840 ();
 b15zdnd11an1n04x5 FILLER_207_1845 ();
 b15zdnd11an1n64x5 FILLER_207_1858 ();
 b15zdnd11an1n64x5 FILLER_207_1922 ();
 b15zdnd11an1n64x5 FILLER_207_1986 ();
 b15zdnd11an1n64x5 FILLER_207_2050 ();
 b15zdnd11an1n32x5 FILLER_207_2114 ();
 b15zdnd11an1n08x5 FILLER_207_2146 ();
 b15zdnd11an1n04x5 FILLER_207_2154 ();
 b15zdnd11an1n04x5 FILLER_207_2200 ();
 b15zdnd11an1n04x5 FILLER_207_2221 ();
 b15zdnd00an1n01x5 FILLER_207_2225 ();
 b15zdnd11an1n04x5 FILLER_207_2233 ();
 b15zdnd11an1n04x5 FILLER_207_2279 ();
 b15zdnd00an1n01x5 FILLER_207_2283 ();
 b15zdnd11an1n64x5 FILLER_208_8 ();
 b15zdnd11an1n64x5 FILLER_208_72 ();
 b15zdnd11an1n64x5 FILLER_208_136 ();
 b15zdnd11an1n64x5 FILLER_208_200 ();
 b15zdnd11an1n64x5 FILLER_208_264 ();
 b15zdnd11an1n64x5 FILLER_208_328 ();
 b15zdnd11an1n64x5 FILLER_208_392 ();
 b15zdnd11an1n64x5 FILLER_208_456 ();
 b15zdnd11an1n64x5 FILLER_208_520 ();
 b15zdnd11an1n16x5 FILLER_208_584 ();
 b15zdnd00an1n02x5 FILLER_208_600 ();
 b15zdnd00an1n01x5 FILLER_208_602 ();
 b15zdnd11an1n64x5 FILLER_208_645 ();
 b15zdnd11an1n08x5 FILLER_208_709 ();
 b15zdnd00an1n01x5 FILLER_208_717 ();
 b15zdnd11an1n32x5 FILLER_208_726 ();
 b15zdnd11an1n16x5 FILLER_208_758 ();
 b15zdnd11an1n04x5 FILLER_208_774 ();
 b15zdnd00an1n02x5 FILLER_208_778 ();
 b15zdnd11an1n64x5 FILLER_208_832 ();
 b15zdnd11an1n64x5 FILLER_208_896 ();
 b15zdnd11an1n64x5 FILLER_208_960 ();
 b15zdnd11an1n64x5 FILLER_208_1024 ();
 b15zdnd11an1n16x5 FILLER_208_1088 ();
 b15zdnd11an1n04x5 FILLER_208_1104 ();
 b15zdnd11an1n64x5 FILLER_208_1129 ();
 b15zdnd11an1n32x5 FILLER_208_1193 ();
 b15zdnd11an1n16x5 FILLER_208_1225 ();
 b15zdnd11an1n04x5 FILLER_208_1241 ();
 b15zdnd00an1n02x5 FILLER_208_1245 ();
 b15zdnd00an1n01x5 FILLER_208_1247 ();
 b15zdnd11an1n64x5 FILLER_208_1258 ();
 b15zdnd11an1n64x5 FILLER_208_1322 ();
 b15zdnd11an1n04x5 FILLER_208_1386 ();
 b15zdnd11an1n64x5 FILLER_208_1410 ();
 b15zdnd11an1n16x5 FILLER_208_1474 ();
 b15zdnd00an1n01x5 FILLER_208_1490 ();
 b15zdnd11an1n64x5 FILLER_208_1511 ();
 b15zdnd11an1n64x5 FILLER_208_1575 ();
 b15zdnd11an1n16x5 FILLER_208_1639 ();
 b15zdnd00an1n02x5 FILLER_208_1655 ();
 b15zdnd00an1n01x5 FILLER_208_1657 ();
 b15zdnd11an1n64x5 FILLER_208_1667 ();
 b15zdnd11an1n64x5 FILLER_208_1731 ();
 b15zdnd11an1n64x5 FILLER_208_1795 ();
 b15zdnd11an1n64x5 FILLER_208_1859 ();
 b15zdnd11an1n64x5 FILLER_208_1923 ();
 b15zdnd11an1n64x5 FILLER_208_1987 ();
 b15zdnd11an1n64x5 FILLER_208_2051 ();
 b15zdnd11an1n32x5 FILLER_208_2115 ();
 b15zdnd11an1n04x5 FILLER_208_2147 ();
 b15zdnd00an1n02x5 FILLER_208_2151 ();
 b15zdnd00an1n01x5 FILLER_208_2153 ();
 b15zdnd11an1n32x5 FILLER_208_2162 ();
 b15zdnd11an1n04x5 FILLER_208_2197 ();
 b15zdnd11an1n08x5 FILLER_208_2204 ();
 b15zdnd00an1n01x5 FILLER_208_2212 ();
 b15zdnd11an1n04x5 FILLER_208_2217 ();
 b15zdnd11an1n04x5 FILLER_208_2263 ();
 b15zdnd11an1n04x5 FILLER_208_2271 ();
 b15zdnd00an1n01x5 FILLER_208_2275 ();
 b15zdnd11an1n64x5 FILLER_209_0 ();
 b15zdnd11an1n64x5 FILLER_209_64 ();
 b15zdnd11an1n64x5 FILLER_209_128 ();
 b15zdnd11an1n64x5 FILLER_209_192 ();
 b15zdnd11an1n64x5 FILLER_209_256 ();
 b15zdnd11an1n32x5 FILLER_209_320 ();
 b15zdnd11an1n08x5 FILLER_209_352 ();
 b15zdnd00an1n01x5 FILLER_209_360 ();
 b15zdnd11an1n64x5 FILLER_209_364 ();
 b15zdnd11an1n64x5 FILLER_209_428 ();
 b15zdnd11an1n64x5 FILLER_209_492 ();
 b15zdnd11an1n64x5 FILLER_209_556 ();
 b15zdnd11an1n64x5 FILLER_209_620 ();
 b15zdnd00an1n02x5 FILLER_209_684 ();
 b15zdnd00an1n01x5 FILLER_209_686 ();
 b15zdnd11an1n16x5 FILLER_209_690 ();
 b15zdnd11an1n08x5 FILLER_209_706 ();
 b15zdnd00an1n02x5 FILLER_209_714 ();
 b15zdnd00an1n01x5 FILLER_209_716 ();
 b15zdnd11an1n32x5 FILLER_209_759 ();
 b15zdnd11an1n08x5 FILLER_209_791 ();
 b15zdnd00an1n01x5 FILLER_209_799 ();
 b15zdnd11an1n04x5 FILLER_209_803 ();
 b15zdnd11an1n64x5 FILLER_209_810 ();
 b15zdnd11an1n64x5 FILLER_209_874 ();
 b15zdnd11an1n64x5 FILLER_209_938 ();
 b15zdnd11an1n64x5 FILLER_209_1002 ();
 b15zdnd11an1n64x5 FILLER_209_1066 ();
 b15zdnd00an1n01x5 FILLER_209_1130 ();
 b15zdnd11an1n64x5 FILLER_209_1135 ();
 b15zdnd11an1n32x5 FILLER_209_1199 ();
 b15zdnd11an1n04x5 FILLER_209_1231 ();
 b15zdnd00an1n02x5 FILLER_209_1235 ();
 b15zdnd11an1n64x5 FILLER_209_1249 ();
 b15zdnd11an1n64x5 FILLER_209_1313 ();
 b15zdnd11an1n32x5 FILLER_209_1377 ();
 b15zdnd11an1n16x5 FILLER_209_1409 ();
 b15zdnd11an1n04x5 FILLER_209_1425 ();
 b15zdnd00an1n01x5 FILLER_209_1429 ();
 b15zdnd11an1n64x5 FILLER_209_1447 ();
 b15zdnd11an1n64x5 FILLER_209_1511 ();
 b15zdnd11an1n64x5 FILLER_209_1575 ();
 b15zdnd11an1n64x5 FILLER_209_1639 ();
 b15zdnd11an1n64x5 FILLER_209_1703 ();
 b15zdnd11an1n64x5 FILLER_209_1767 ();
 b15zdnd11an1n32x5 FILLER_209_1831 ();
 b15zdnd11an1n16x5 FILLER_209_1863 ();
 b15zdnd11an1n08x5 FILLER_209_1879 ();
 b15zdnd00an1n02x5 FILLER_209_1887 ();
 b15zdnd00an1n01x5 FILLER_209_1889 ();
 b15zdnd11an1n64x5 FILLER_209_1932 ();
 b15zdnd11an1n64x5 FILLER_209_1996 ();
 b15zdnd11an1n64x5 FILLER_209_2060 ();
 b15zdnd11an1n32x5 FILLER_209_2124 ();
 b15zdnd11an1n16x5 FILLER_209_2156 ();
 b15zdnd11an1n08x5 FILLER_209_2172 ();
 b15zdnd00an1n02x5 FILLER_209_2180 ();
 b15zdnd00an1n01x5 FILLER_209_2182 ();
 b15zdnd11an1n04x5 FILLER_209_2235 ();
 b15zdnd00an1n02x5 FILLER_209_2281 ();
 b15zdnd00an1n01x5 FILLER_209_2283 ();
 b15zdnd11an1n64x5 FILLER_210_8 ();
 b15zdnd11an1n64x5 FILLER_210_72 ();
 b15zdnd11an1n64x5 FILLER_210_136 ();
 b15zdnd11an1n64x5 FILLER_210_200 ();
 b15zdnd11an1n64x5 FILLER_210_264 ();
 b15zdnd11an1n08x5 FILLER_210_328 ();
 b15zdnd11an1n64x5 FILLER_210_388 ();
 b15zdnd11an1n64x5 FILLER_210_452 ();
 b15zdnd11an1n08x5 FILLER_210_516 ();
 b15zdnd11an1n04x5 FILLER_210_524 ();
 b15zdnd00an1n01x5 FILLER_210_528 ();
 b15zdnd11an1n64x5 FILLER_210_537 ();
 b15zdnd11an1n32x5 FILLER_210_601 ();
 b15zdnd11an1n16x5 FILLER_210_633 ();
 b15zdnd11an1n08x5 FILLER_210_649 ();
 b15zdnd11an1n04x5 FILLER_210_657 ();
 b15zdnd00an1n02x5 FILLER_210_661 ();
 b15zdnd00an1n01x5 FILLER_210_663 ();
 b15zdnd00an1n02x5 FILLER_210_716 ();
 b15zdnd11an1n64x5 FILLER_210_726 ();
 b15zdnd11an1n08x5 FILLER_210_790 ();
 b15zdnd00an1n02x5 FILLER_210_798 ();
 b15zdnd00an1n01x5 FILLER_210_800 ();
 b15zdnd11an1n64x5 FILLER_210_804 ();
 b15zdnd11an1n08x5 FILLER_210_868 ();
 b15zdnd11an1n04x5 FILLER_210_876 ();
 b15zdnd00an1n02x5 FILLER_210_880 ();
 b15zdnd11an1n64x5 FILLER_210_914 ();
 b15zdnd11an1n64x5 FILLER_210_978 ();
 b15zdnd11an1n64x5 FILLER_210_1042 ();
 b15zdnd11an1n04x5 FILLER_210_1106 ();
 b15zdnd00an1n01x5 FILLER_210_1110 ();
 b15zdnd11an1n16x5 FILLER_210_1119 ();
 b15zdnd11an1n08x5 FILLER_210_1135 ();
 b15zdnd00an1n02x5 FILLER_210_1143 ();
 b15zdnd11an1n64x5 FILLER_210_1156 ();
 b15zdnd11an1n64x5 FILLER_210_1220 ();
 b15zdnd11an1n64x5 FILLER_210_1284 ();
 b15zdnd11an1n32x5 FILLER_210_1348 ();
 b15zdnd11an1n08x5 FILLER_210_1380 ();
 b15zdnd11an1n04x5 FILLER_210_1388 ();
 b15zdnd00an1n02x5 FILLER_210_1392 ();
 b15zdnd11an1n64x5 FILLER_210_1408 ();
 b15zdnd11an1n64x5 FILLER_210_1472 ();
 b15zdnd11an1n64x5 FILLER_210_1536 ();
 b15zdnd11an1n64x5 FILLER_210_1600 ();
 b15zdnd11an1n64x5 FILLER_210_1664 ();
 b15zdnd11an1n64x5 FILLER_210_1728 ();
 b15zdnd11an1n64x5 FILLER_210_1792 ();
 b15zdnd11an1n64x5 FILLER_210_1856 ();
 b15zdnd11an1n64x5 FILLER_210_1920 ();
 b15zdnd11an1n64x5 FILLER_210_1984 ();
 b15zdnd11an1n64x5 FILLER_210_2048 ();
 b15zdnd11an1n32x5 FILLER_210_2112 ();
 b15zdnd11an1n08x5 FILLER_210_2144 ();
 b15zdnd00an1n02x5 FILLER_210_2152 ();
 b15zdnd11an1n32x5 FILLER_210_2162 ();
 b15zdnd00an1n02x5 FILLER_210_2194 ();
 b15zdnd00an1n01x5 FILLER_210_2196 ();
 b15zdnd11an1n04x5 FILLER_210_2200 ();
 b15zdnd11an1n04x5 FILLER_210_2246 ();
 b15zdnd11an1n04x5 FILLER_210_2254 ();
 b15zdnd11an1n08x5 FILLER_210_2262 ();
 b15zdnd00an1n02x5 FILLER_210_2274 ();
 b15zdnd11an1n64x5 FILLER_211_0 ();
 b15zdnd11an1n64x5 FILLER_211_64 ();
 b15zdnd11an1n64x5 FILLER_211_128 ();
 b15zdnd11an1n64x5 FILLER_211_192 ();
 b15zdnd11an1n64x5 FILLER_211_256 ();
 b15zdnd11an1n32x5 FILLER_211_320 ();
 b15zdnd00an1n01x5 FILLER_211_352 ();
 b15zdnd11an1n04x5 FILLER_211_356 ();
 b15zdnd11an1n64x5 FILLER_211_363 ();
 b15zdnd11an1n64x5 FILLER_211_427 ();
 b15zdnd11an1n32x5 FILLER_211_491 ();
 b15zdnd00an1n01x5 FILLER_211_523 ();
 b15zdnd11an1n64x5 FILLER_211_566 ();
 b15zdnd11an1n32x5 FILLER_211_630 ();
 b15zdnd11an1n16x5 FILLER_211_662 ();
 b15zdnd11an1n04x5 FILLER_211_678 ();
 b15zdnd00an1n02x5 FILLER_211_682 ();
 b15zdnd00an1n01x5 FILLER_211_684 ();
 b15zdnd11an1n04x5 FILLER_211_688 ();
 b15zdnd11an1n08x5 FILLER_211_695 ();
 b15zdnd00an1n02x5 FILLER_211_703 ();
 b15zdnd00an1n01x5 FILLER_211_705 ();
 b15zdnd11an1n64x5 FILLER_211_758 ();
 b15zdnd11an1n64x5 FILLER_211_822 ();
 b15zdnd11an1n64x5 FILLER_211_886 ();
 b15zdnd11an1n64x5 FILLER_211_950 ();
 b15zdnd11an1n64x5 FILLER_211_1014 ();
 b15zdnd11an1n16x5 FILLER_211_1078 ();
 b15zdnd11an1n08x5 FILLER_211_1094 ();
 b15zdnd11an1n04x5 FILLER_211_1102 ();
 b15zdnd00an1n02x5 FILLER_211_1106 ();
 b15zdnd11an1n64x5 FILLER_211_1144 ();
 b15zdnd11an1n16x5 FILLER_211_1208 ();
 b15zdnd11an1n08x5 FILLER_211_1224 ();
 b15zdnd11an1n04x5 FILLER_211_1232 ();
 b15zdnd11an1n04x5 FILLER_211_1248 ();
 b15zdnd00an1n02x5 FILLER_211_1252 ();
 b15zdnd11an1n64x5 FILLER_211_1270 ();
 b15zdnd11an1n64x5 FILLER_211_1334 ();
 b15zdnd11an1n64x5 FILLER_211_1398 ();
 b15zdnd11an1n64x5 FILLER_211_1462 ();
 b15zdnd11an1n64x5 FILLER_211_1526 ();
 b15zdnd11an1n64x5 FILLER_211_1590 ();
 b15zdnd00an1n01x5 FILLER_211_1654 ();
 b15zdnd11an1n64x5 FILLER_211_1664 ();
 b15zdnd11an1n64x5 FILLER_211_1728 ();
 b15zdnd11an1n64x5 FILLER_211_1792 ();
 b15zdnd11an1n64x5 FILLER_211_1856 ();
 b15zdnd11an1n64x5 FILLER_211_1920 ();
 b15zdnd11an1n64x5 FILLER_211_1984 ();
 b15zdnd11an1n64x5 FILLER_211_2048 ();
 b15zdnd11an1n64x5 FILLER_211_2112 ();
 b15zdnd11an1n16x5 FILLER_211_2176 ();
 b15zdnd00an1n02x5 FILLER_211_2192 ();
 b15zdnd11an1n04x5 FILLER_211_2236 ();
 b15zdnd00an1n02x5 FILLER_211_2282 ();
 b15zdnd11an1n04x5 FILLER_212_8 ();
 b15zdnd00an1n02x5 FILLER_212_12 ();
 b15zdnd11an1n32x5 FILLER_212_18 ();
 b15zdnd11an1n04x5 FILLER_212_50 ();
 b15zdnd00an1n02x5 FILLER_212_54 ();
 b15zdnd11an1n64x5 FILLER_212_59 ();
 b15zdnd11an1n64x5 FILLER_212_123 ();
 b15zdnd11an1n64x5 FILLER_212_187 ();
 b15zdnd11an1n64x5 FILLER_212_251 ();
 b15zdnd11an1n64x5 FILLER_212_315 ();
 b15zdnd11an1n64x5 FILLER_212_379 ();
 b15zdnd11an1n64x5 FILLER_212_443 ();
 b15zdnd11an1n32x5 FILLER_212_507 ();
 b15zdnd11an1n08x5 FILLER_212_539 ();
 b15zdnd00an1n02x5 FILLER_212_547 ();
 b15zdnd00an1n01x5 FILLER_212_549 ();
 b15zdnd11an1n16x5 FILLER_212_592 ();
 b15zdnd00an1n01x5 FILLER_212_608 ();
 b15zdnd11an1n16x5 FILLER_212_651 ();
 b15zdnd11an1n04x5 FILLER_212_667 ();
 b15zdnd00an1n02x5 FILLER_212_671 ();
 b15zdnd00an1n01x5 FILLER_212_673 ();
 b15zdnd00an1n02x5 FILLER_212_716 ();
 b15zdnd00an1n02x5 FILLER_212_726 ();
 b15zdnd00an1n01x5 FILLER_212_728 ();
 b15zdnd11an1n04x5 FILLER_212_732 ();
 b15zdnd11an1n04x5 FILLER_212_739 ();
 b15zdnd00an1n02x5 FILLER_212_743 ();
 b15zdnd00an1n01x5 FILLER_212_745 ();
 b15zdnd11an1n64x5 FILLER_212_788 ();
 b15zdnd11an1n64x5 FILLER_212_852 ();
 b15zdnd11an1n64x5 FILLER_212_916 ();
 b15zdnd11an1n64x5 FILLER_212_980 ();
 b15zdnd11an1n64x5 FILLER_212_1044 ();
 b15zdnd11an1n32x5 FILLER_212_1108 ();
 b15zdnd00an1n02x5 FILLER_212_1140 ();
 b15zdnd00an1n01x5 FILLER_212_1142 ();
 b15zdnd11an1n64x5 FILLER_212_1154 ();
 b15zdnd11an1n64x5 FILLER_212_1218 ();
 b15zdnd11an1n32x5 FILLER_212_1282 ();
 b15zdnd00an1n01x5 FILLER_212_1314 ();
 b15zdnd11an1n32x5 FILLER_212_1335 ();
 b15zdnd00an1n02x5 FILLER_212_1367 ();
 b15zdnd00an1n01x5 FILLER_212_1369 ();
 b15zdnd11an1n64x5 FILLER_212_1384 ();
 b15zdnd11an1n64x5 FILLER_212_1448 ();
 b15zdnd11an1n32x5 FILLER_212_1512 ();
 b15zdnd11an1n04x5 FILLER_212_1544 ();
 b15zdnd00an1n02x5 FILLER_212_1548 ();
 b15zdnd00an1n01x5 FILLER_212_1550 ();
 b15zdnd11an1n64x5 FILLER_212_1571 ();
 b15zdnd11an1n64x5 FILLER_212_1635 ();
 b15zdnd11an1n64x5 FILLER_212_1699 ();
 b15zdnd11an1n64x5 FILLER_212_1763 ();
 b15zdnd11an1n64x5 FILLER_212_1827 ();
 b15zdnd11an1n16x5 FILLER_212_1891 ();
 b15zdnd11an1n08x5 FILLER_212_1907 ();
 b15zdnd11an1n04x5 FILLER_212_1915 ();
 b15zdnd00an1n02x5 FILLER_212_1919 ();
 b15zdnd11an1n64x5 FILLER_212_1963 ();
 b15zdnd11an1n64x5 FILLER_212_2027 ();
 b15zdnd11an1n32x5 FILLER_212_2091 ();
 b15zdnd11an1n16x5 FILLER_212_2123 ();
 b15zdnd11an1n08x5 FILLER_212_2139 ();
 b15zdnd11an1n04x5 FILLER_212_2147 ();
 b15zdnd00an1n02x5 FILLER_212_2151 ();
 b15zdnd00an1n01x5 FILLER_212_2153 ();
 b15zdnd11an1n16x5 FILLER_212_2162 ();
 b15zdnd11an1n08x5 FILLER_212_2178 ();
 b15zdnd11an1n04x5 FILLER_212_2228 ();
 b15zdnd00an1n02x5 FILLER_212_2274 ();
 b15zdnd00an1n02x5 FILLER_213_0 ();
 b15zdnd00an1n01x5 FILLER_213_2 ();
 b15zdnd11an1n64x5 FILLER_213_45 ();
 b15zdnd11an1n32x5 FILLER_213_109 ();
 b15zdnd11an1n16x5 FILLER_213_141 ();
 b15zdnd00an1n02x5 FILLER_213_157 ();
 b15zdnd11an1n64x5 FILLER_213_168 ();
 b15zdnd11an1n32x5 FILLER_213_232 ();
 b15zdnd11an1n16x5 FILLER_213_264 ();
 b15zdnd11an1n08x5 FILLER_213_280 ();
 b15zdnd00an1n02x5 FILLER_213_288 ();
 b15zdnd11an1n64x5 FILLER_213_332 ();
 b15zdnd11an1n04x5 FILLER_213_396 ();
 b15zdnd00an1n02x5 FILLER_213_400 ();
 b15zdnd00an1n01x5 FILLER_213_402 ();
 b15zdnd11an1n64x5 FILLER_213_406 ();
 b15zdnd11an1n64x5 FILLER_213_470 ();
 b15zdnd11an1n16x5 FILLER_213_534 ();
 b15zdnd11an1n08x5 FILLER_213_550 ();
 b15zdnd00an1n02x5 FILLER_213_558 ();
 b15zdnd00an1n01x5 FILLER_213_560 ();
 b15zdnd11an1n64x5 FILLER_213_568 ();
 b15zdnd11an1n64x5 FILLER_213_632 ();
 b15zdnd11an1n32x5 FILLER_213_696 ();
 b15zdnd11an1n04x5 FILLER_213_728 ();
 b15zdnd11an1n64x5 FILLER_213_735 ();
 b15zdnd11an1n64x5 FILLER_213_799 ();
 b15zdnd11an1n64x5 FILLER_213_863 ();
 b15zdnd11an1n64x5 FILLER_213_927 ();
 b15zdnd11an1n64x5 FILLER_213_991 ();
 b15zdnd11an1n64x5 FILLER_213_1055 ();
 b15zdnd11an1n64x5 FILLER_213_1119 ();
 b15zdnd11an1n64x5 FILLER_213_1183 ();
 b15zdnd11an1n64x5 FILLER_213_1247 ();
 b15zdnd11an1n64x5 FILLER_213_1311 ();
 b15zdnd11an1n64x5 FILLER_213_1375 ();
 b15zdnd11an1n64x5 FILLER_213_1439 ();
 b15zdnd11an1n16x5 FILLER_213_1503 ();
 b15zdnd11an1n04x5 FILLER_213_1519 ();
 b15zdnd00an1n02x5 FILLER_213_1523 ();
 b15zdnd00an1n01x5 FILLER_213_1525 ();
 b15zdnd11an1n64x5 FILLER_213_1535 ();
 b15zdnd11an1n64x5 FILLER_213_1599 ();
 b15zdnd11an1n64x5 FILLER_213_1663 ();
 b15zdnd11an1n64x5 FILLER_213_1727 ();
 b15zdnd11an1n64x5 FILLER_213_1791 ();
 b15zdnd11an1n64x5 FILLER_213_1855 ();
 b15zdnd11an1n16x5 FILLER_213_1919 ();
 b15zdnd11an1n08x5 FILLER_213_1935 ();
 b15zdnd11an1n04x5 FILLER_213_1943 ();
 b15zdnd00an1n02x5 FILLER_213_1947 ();
 b15zdnd00an1n01x5 FILLER_213_1949 ();
 b15zdnd11an1n64x5 FILLER_213_1992 ();
 b15zdnd11an1n64x5 FILLER_213_2056 ();
 b15zdnd11an1n32x5 FILLER_213_2120 ();
 b15zdnd11an1n16x5 FILLER_213_2152 ();
 b15zdnd11an1n08x5 FILLER_213_2168 ();
 b15zdnd11an1n04x5 FILLER_213_2176 ();
 b15zdnd00an1n02x5 FILLER_213_2180 ();
 b15zdnd00an1n01x5 FILLER_213_2182 ();
 b15zdnd11an1n04x5 FILLER_213_2225 ();
 b15zdnd11an1n04x5 FILLER_213_2233 ();
 b15zdnd00an1n02x5 FILLER_213_2237 ();
 b15zdnd00an1n02x5 FILLER_213_2281 ();
 b15zdnd00an1n01x5 FILLER_213_2283 ();
 b15zdnd11an1n32x5 FILLER_214_8 ();
 b15zdnd11an1n16x5 FILLER_214_40 ();
 b15zdnd11an1n04x5 FILLER_214_56 ();
 b15zdnd00an1n02x5 FILLER_214_60 ();
 b15zdnd11an1n04x5 FILLER_214_67 ();
 b15zdnd11an1n64x5 FILLER_214_78 ();
 b15zdnd11an1n64x5 FILLER_214_142 ();
 b15zdnd11an1n32x5 FILLER_214_206 ();
 b15zdnd11an1n16x5 FILLER_214_238 ();
 b15zdnd11an1n04x5 FILLER_214_254 ();
 b15zdnd00an1n01x5 FILLER_214_258 ();
 b15zdnd11an1n64x5 FILLER_214_275 ();
 b15zdnd11an1n32x5 FILLER_214_339 ();
 b15zdnd11an1n08x5 FILLER_214_371 ();
 b15zdnd00an1n02x5 FILLER_214_379 ();
 b15zdnd11an1n04x5 FILLER_214_433 ();
 b15zdnd11an1n32x5 FILLER_214_444 ();
 b15zdnd11an1n16x5 FILLER_214_476 ();
 b15zdnd11an1n04x5 FILLER_214_492 ();
 b15zdnd11an1n04x5 FILLER_214_538 ();
 b15zdnd00an1n02x5 FILLER_214_542 ();
 b15zdnd11an1n04x5 FILLER_214_550 ();
 b15zdnd11an1n64x5 FILLER_214_562 ();
 b15zdnd11an1n16x5 FILLER_214_626 ();
 b15zdnd11an1n04x5 FILLER_214_642 ();
 b15zdnd00an1n02x5 FILLER_214_646 ();
 b15zdnd00an1n01x5 FILLER_214_648 ();
 b15zdnd11an1n16x5 FILLER_214_691 ();
 b15zdnd11an1n08x5 FILLER_214_707 ();
 b15zdnd00an1n02x5 FILLER_214_715 ();
 b15zdnd00an1n01x5 FILLER_214_717 ();
 b15zdnd11an1n64x5 FILLER_214_726 ();
 b15zdnd11an1n64x5 FILLER_214_790 ();
 b15zdnd11an1n64x5 FILLER_214_854 ();
 b15zdnd11an1n64x5 FILLER_214_918 ();
 b15zdnd11an1n64x5 FILLER_214_982 ();
 b15zdnd11an1n32x5 FILLER_214_1046 ();
 b15zdnd11an1n16x5 FILLER_214_1078 ();
 b15zdnd11an1n08x5 FILLER_214_1094 ();
 b15zdnd00an1n02x5 FILLER_214_1102 ();
 b15zdnd11an1n64x5 FILLER_214_1146 ();
 b15zdnd11an1n64x5 FILLER_214_1210 ();
 b15zdnd11an1n32x5 FILLER_214_1274 ();
 b15zdnd11an1n16x5 FILLER_214_1306 ();
 b15zdnd11an1n08x5 FILLER_214_1322 ();
 b15zdnd11an1n04x5 FILLER_214_1330 ();
 b15zdnd11an1n16x5 FILLER_214_1348 ();
 b15zdnd11an1n16x5 FILLER_214_1381 ();
 b15zdnd11an1n08x5 FILLER_214_1397 ();
 b15zdnd11an1n04x5 FILLER_214_1405 ();
 b15zdnd11an1n32x5 FILLER_214_1429 ();
 b15zdnd11an1n16x5 FILLER_214_1461 ();
 b15zdnd11an1n08x5 FILLER_214_1477 ();
 b15zdnd00an1n02x5 FILLER_214_1485 ();
 b15zdnd00an1n01x5 FILLER_214_1487 ();
 b15zdnd11an1n64x5 FILLER_214_1508 ();
 b15zdnd11an1n64x5 FILLER_214_1572 ();
 b15zdnd11an1n64x5 FILLER_214_1636 ();
 b15zdnd11an1n64x5 FILLER_214_1700 ();
 b15zdnd11an1n64x5 FILLER_214_1764 ();
 b15zdnd11an1n64x5 FILLER_214_1828 ();
 b15zdnd11an1n64x5 FILLER_214_1892 ();
 b15zdnd11an1n64x5 FILLER_214_1956 ();
 b15zdnd11an1n64x5 FILLER_214_2020 ();
 b15zdnd11an1n64x5 FILLER_214_2084 ();
 b15zdnd11an1n04x5 FILLER_214_2148 ();
 b15zdnd00an1n02x5 FILLER_214_2152 ();
 b15zdnd11an1n16x5 FILLER_214_2162 ();
 b15zdnd00an1n01x5 FILLER_214_2178 ();
 b15zdnd11an1n04x5 FILLER_214_2221 ();
 b15zdnd11an1n08x5 FILLER_214_2267 ();
 b15zdnd00an1n01x5 FILLER_214_2275 ();
 b15zdnd11an1n64x5 FILLER_215_0 ();
 b15zdnd11an1n64x5 FILLER_215_64 ();
 b15zdnd11an1n64x5 FILLER_215_128 ();
 b15zdnd11an1n64x5 FILLER_215_192 ();
 b15zdnd11an1n32x5 FILLER_215_256 ();
 b15zdnd11an1n08x5 FILLER_215_288 ();
 b15zdnd00an1n02x5 FILLER_215_296 ();
 b15zdnd00an1n01x5 FILLER_215_298 ();
 b15zdnd11an1n64x5 FILLER_215_325 ();
 b15zdnd11an1n08x5 FILLER_215_389 ();
 b15zdnd11an1n04x5 FILLER_215_400 ();
 b15zdnd11an1n32x5 FILLER_215_407 ();
 b15zdnd11an1n16x5 FILLER_215_439 ();
 b15zdnd00an1n01x5 FILLER_215_455 ();
 b15zdnd11an1n08x5 FILLER_215_508 ();
 b15zdnd00an1n02x5 FILLER_215_516 ();
 b15zdnd00an1n01x5 FILLER_215_518 ();
 b15zdnd11an1n08x5 FILLER_215_525 ();
 b15zdnd11an1n04x5 FILLER_215_533 ();
 b15zdnd11an1n64x5 FILLER_215_579 ();
 b15zdnd11an1n64x5 FILLER_215_643 ();
 b15zdnd11an1n64x5 FILLER_215_707 ();
 b15zdnd11an1n64x5 FILLER_215_771 ();
 b15zdnd11an1n64x5 FILLER_215_835 ();
 b15zdnd11an1n64x5 FILLER_215_899 ();
 b15zdnd11an1n64x5 FILLER_215_963 ();
 b15zdnd11an1n32x5 FILLER_215_1027 ();
 b15zdnd11an1n16x5 FILLER_215_1059 ();
 b15zdnd00an1n02x5 FILLER_215_1075 ();
 b15zdnd11an1n64x5 FILLER_215_1101 ();
 b15zdnd11an1n64x5 FILLER_215_1165 ();
 b15zdnd11an1n64x5 FILLER_215_1229 ();
 b15zdnd11an1n64x5 FILLER_215_1293 ();
 b15zdnd11an1n16x5 FILLER_215_1357 ();
 b15zdnd11an1n04x5 FILLER_215_1373 ();
 b15zdnd00an1n02x5 FILLER_215_1377 ();
 b15zdnd00an1n01x5 FILLER_215_1379 ();
 b15zdnd11an1n04x5 FILLER_215_1400 ();
 b15zdnd11an1n64x5 FILLER_215_1416 ();
 b15zdnd11an1n64x5 FILLER_215_1480 ();
 b15zdnd11an1n64x5 FILLER_215_1544 ();
 b15zdnd11an1n64x5 FILLER_215_1608 ();
 b15zdnd11an1n64x5 FILLER_215_1672 ();
 b15zdnd11an1n64x5 FILLER_215_1736 ();
 b15zdnd11an1n64x5 FILLER_215_1800 ();
 b15zdnd11an1n04x5 FILLER_215_1864 ();
 b15zdnd00an1n02x5 FILLER_215_1868 ();
 b15zdnd00an1n01x5 FILLER_215_1870 ();
 b15zdnd11an1n64x5 FILLER_215_1880 ();
 b15zdnd11an1n64x5 FILLER_215_1944 ();
 b15zdnd11an1n32x5 FILLER_215_2008 ();
 b15zdnd11an1n04x5 FILLER_215_2040 ();
 b15zdnd00an1n02x5 FILLER_215_2044 ();
 b15zdnd00an1n01x5 FILLER_215_2046 ();
 b15zdnd11an1n08x5 FILLER_215_2089 ();
 b15zdnd00an1n02x5 FILLER_215_2097 ();
 b15zdnd11an1n16x5 FILLER_215_2108 ();
 b15zdnd11an1n08x5 FILLER_215_2124 ();
 b15zdnd11an1n04x5 FILLER_215_2132 ();
 b15zdnd00an1n01x5 FILLER_215_2136 ();
 b15zdnd11an1n04x5 FILLER_215_2179 ();
 b15zdnd00an1n01x5 FILLER_215_2183 ();
 b15zdnd11an1n04x5 FILLER_215_2204 ();
 b15zdnd11an1n04x5 FILLER_215_2250 ();
 b15zdnd11an1n04x5 FILLER_215_2274 ();
 b15zdnd00an1n02x5 FILLER_215_2282 ();
 b15zdnd11an1n32x5 FILLER_216_8 ();
 b15zdnd11an1n16x5 FILLER_216_40 ();
 b15zdnd11an1n08x5 FILLER_216_56 ();
 b15zdnd11an1n04x5 FILLER_216_64 ();
 b15zdnd00an1n01x5 FILLER_216_68 ();
 b15zdnd11an1n64x5 FILLER_216_87 ();
 b15zdnd11an1n04x5 FILLER_216_151 ();
 b15zdnd11an1n04x5 FILLER_216_164 ();
 b15zdnd00an1n02x5 FILLER_216_168 ();
 b15zdnd11an1n64x5 FILLER_216_212 ();
 b15zdnd11an1n64x5 FILLER_216_276 ();
 b15zdnd11an1n64x5 FILLER_216_340 ();
 b15zdnd11an1n16x5 FILLER_216_404 ();
 b15zdnd11an1n08x5 FILLER_216_420 ();
 b15zdnd11an1n04x5 FILLER_216_428 ();
 b15zdnd00an1n02x5 FILLER_216_432 ();
 b15zdnd00an1n01x5 FILLER_216_434 ();
 b15zdnd11an1n08x5 FILLER_216_477 ();
 b15zdnd11an1n32x5 FILLER_216_527 ();
 b15zdnd00an1n02x5 FILLER_216_559 ();
 b15zdnd11an1n08x5 FILLER_216_568 ();
 b15zdnd11an1n04x5 FILLER_216_582 ();
 b15zdnd11an1n64x5 FILLER_216_594 ();
 b15zdnd11an1n32x5 FILLER_216_658 ();
 b15zdnd11an1n16x5 FILLER_216_690 ();
 b15zdnd11an1n08x5 FILLER_216_706 ();
 b15zdnd11an1n04x5 FILLER_216_714 ();
 b15zdnd11an1n64x5 FILLER_216_726 ();
 b15zdnd11an1n64x5 FILLER_216_790 ();
 b15zdnd11an1n64x5 FILLER_216_854 ();
 b15zdnd11an1n64x5 FILLER_216_918 ();
 b15zdnd11an1n64x5 FILLER_216_982 ();
 b15zdnd11an1n64x5 FILLER_216_1046 ();
 b15zdnd11an1n64x5 FILLER_216_1110 ();
 b15zdnd11an1n64x5 FILLER_216_1174 ();
 b15zdnd11an1n64x5 FILLER_216_1238 ();
 b15zdnd11an1n32x5 FILLER_216_1302 ();
 b15zdnd00an1n02x5 FILLER_216_1334 ();
 b15zdnd11an1n08x5 FILLER_216_1356 ();
 b15zdnd00an1n02x5 FILLER_216_1364 ();
 b15zdnd11an1n64x5 FILLER_216_1386 ();
 b15zdnd11an1n32x5 FILLER_216_1450 ();
 b15zdnd11an1n64x5 FILLER_216_1499 ();
 b15zdnd11an1n64x5 FILLER_216_1563 ();
 b15zdnd11an1n64x5 FILLER_216_1627 ();
 b15zdnd11an1n64x5 FILLER_216_1691 ();
 b15zdnd11an1n64x5 FILLER_216_1755 ();
 b15zdnd11an1n32x5 FILLER_216_1819 ();
 b15zdnd11an1n16x5 FILLER_216_1851 ();
 b15zdnd11an1n08x5 FILLER_216_1867 ();
 b15zdnd00an1n02x5 FILLER_216_1875 ();
 b15zdnd11an1n64x5 FILLER_216_1886 ();
 b15zdnd11an1n64x5 FILLER_216_1950 ();
 b15zdnd11an1n32x5 FILLER_216_2014 ();
 b15zdnd11an1n16x5 FILLER_216_2046 ();
 b15zdnd11an1n08x5 FILLER_216_2062 ();
 b15zdnd11an1n04x5 FILLER_216_2070 ();
 b15zdnd00an1n02x5 FILLER_216_2074 ();
 b15zdnd11an1n32x5 FILLER_216_2118 ();
 b15zdnd11an1n04x5 FILLER_216_2150 ();
 b15zdnd11an1n16x5 FILLER_216_2162 ();
 b15zdnd11an1n08x5 FILLER_216_2178 ();
 b15zdnd11an1n04x5 FILLER_216_2228 ();
 b15zdnd00an1n02x5 FILLER_216_2274 ();
 b15zdnd11an1n64x5 FILLER_217_0 ();
 b15zdnd11an1n08x5 FILLER_217_64 ();
 b15zdnd00an1n02x5 FILLER_217_72 ();
 b15zdnd00an1n01x5 FILLER_217_74 ();
 b15zdnd11an1n64x5 FILLER_217_84 ();
 b15zdnd11an1n64x5 FILLER_217_148 ();
 b15zdnd11an1n32x5 FILLER_217_212 ();
 b15zdnd11an1n16x5 FILLER_217_244 ();
 b15zdnd11an1n64x5 FILLER_217_288 ();
 b15zdnd11an1n64x5 FILLER_217_352 ();
 b15zdnd11an1n32x5 FILLER_217_416 ();
 b15zdnd11an1n08x5 FILLER_217_448 ();
 b15zdnd00an1n02x5 FILLER_217_456 ();
 b15zdnd00an1n01x5 FILLER_217_458 ();
 b15zdnd11an1n04x5 FILLER_217_462 ();
 b15zdnd11an1n04x5 FILLER_217_469 ();
 b15zdnd11an1n04x5 FILLER_217_476 ();
 b15zdnd11an1n04x5 FILLER_217_483 ();
 b15zdnd00an1n02x5 FILLER_217_487 ();
 b15zdnd00an1n01x5 FILLER_217_489 ();
 b15zdnd11an1n08x5 FILLER_217_493 ();
 b15zdnd00an1n02x5 FILLER_217_501 ();
 b15zdnd00an1n01x5 FILLER_217_503 ();
 b15zdnd11an1n04x5 FILLER_217_546 ();
 b15zdnd11an1n04x5 FILLER_217_556 ();
 b15zdnd00an1n02x5 FILLER_217_560 ();
 b15zdnd11an1n64x5 FILLER_217_604 ();
 b15zdnd11an1n64x5 FILLER_217_668 ();
 b15zdnd11an1n64x5 FILLER_217_732 ();
 b15zdnd11an1n64x5 FILLER_217_796 ();
 b15zdnd11an1n32x5 FILLER_217_860 ();
 b15zdnd11an1n16x5 FILLER_217_892 ();
 b15zdnd11an1n08x5 FILLER_217_908 ();
 b15zdnd00an1n02x5 FILLER_217_916 ();
 b15zdnd00an1n01x5 FILLER_217_918 ();
 b15zdnd11an1n64x5 FILLER_217_922 ();
 b15zdnd11an1n64x5 FILLER_217_986 ();
 b15zdnd11an1n64x5 FILLER_217_1050 ();
 b15zdnd11an1n64x5 FILLER_217_1114 ();
 b15zdnd11an1n64x5 FILLER_217_1178 ();
 b15zdnd11an1n64x5 FILLER_217_1242 ();
 b15zdnd11an1n08x5 FILLER_217_1306 ();
 b15zdnd11an1n04x5 FILLER_217_1321 ();
 b15zdnd11an1n64x5 FILLER_217_1339 ();
 b15zdnd11an1n64x5 FILLER_217_1403 ();
 b15zdnd11an1n08x5 FILLER_217_1467 ();
 b15zdnd11an1n04x5 FILLER_217_1475 ();
 b15zdnd00an1n01x5 FILLER_217_1479 ();
 b15zdnd11an1n64x5 FILLER_217_1494 ();
 b15zdnd11an1n32x5 FILLER_217_1558 ();
 b15zdnd11an1n16x5 FILLER_217_1590 ();
 b15zdnd11an1n04x5 FILLER_217_1606 ();
 b15zdnd00an1n02x5 FILLER_217_1610 ();
 b15zdnd00an1n01x5 FILLER_217_1612 ();
 b15zdnd11an1n64x5 FILLER_217_1640 ();
 b15zdnd11an1n64x5 FILLER_217_1704 ();
 b15zdnd11an1n64x5 FILLER_217_1768 ();
 b15zdnd11an1n64x5 FILLER_217_1832 ();
 b15zdnd11an1n64x5 FILLER_217_1896 ();
 b15zdnd11an1n64x5 FILLER_217_1960 ();
 b15zdnd11an1n16x5 FILLER_217_2024 ();
 b15zdnd11an1n08x5 FILLER_217_2040 ();
 b15zdnd00an1n02x5 FILLER_217_2048 ();
 b15zdnd11an1n08x5 FILLER_217_2053 ();
 b15zdnd11an1n04x5 FILLER_217_2061 ();
 b15zdnd00an1n02x5 FILLER_217_2065 ();
 b15zdnd00an1n01x5 FILLER_217_2067 ();
 b15zdnd11an1n08x5 FILLER_217_2071 ();
 b15zdnd11an1n04x5 FILLER_217_2079 ();
 b15zdnd11an1n08x5 FILLER_217_2125 ();
 b15zdnd11an1n04x5 FILLER_217_2133 ();
 b15zdnd00an1n01x5 FILLER_217_2137 ();
 b15zdnd11an1n08x5 FILLER_217_2180 ();
 b15zdnd11an1n04x5 FILLER_217_2188 ();
 b15zdnd00an1n02x5 FILLER_217_2192 ();
 b15zdnd11an1n04x5 FILLER_217_2236 ();
 b15zdnd00an1n02x5 FILLER_217_2282 ();
 b15zdnd11an1n64x5 FILLER_218_8 ();
 b15zdnd11an1n04x5 FILLER_218_72 ();
 b15zdnd11an1n64x5 FILLER_218_81 ();
 b15zdnd11an1n16x5 FILLER_218_145 ();
 b15zdnd11an1n08x5 FILLER_218_161 ();
 b15zdnd00an1n01x5 FILLER_218_169 ();
 b15zdnd11an1n16x5 FILLER_218_198 ();
 b15zdnd11an1n08x5 FILLER_218_214 ();
 b15zdnd11an1n04x5 FILLER_218_222 ();
 b15zdnd00an1n01x5 FILLER_218_226 ();
 b15zdnd11an1n08x5 FILLER_218_269 ();
 b15zdnd11an1n04x5 FILLER_218_277 ();
 b15zdnd11an1n08x5 FILLER_218_284 ();
 b15zdnd11an1n64x5 FILLER_218_295 ();
 b15zdnd11an1n64x5 FILLER_218_359 ();
 b15zdnd11an1n32x5 FILLER_218_423 ();
 b15zdnd11an1n08x5 FILLER_218_455 ();
 b15zdnd00an1n01x5 FILLER_218_463 ();
 b15zdnd11an1n04x5 FILLER_218_516 ();
 b15zdnd00an1n01x5 FILLER_218_520 ();
 b15zdnd11an1n04x5 FILLER_218_563 ();
 b15zdnd11an1n16x5 FILLER_218_609 ();
 b15zdnd11an1n08x5 FILLER_218_625 ();
 b15zdnd11an1n04x5 FILLER_218_633 ();
 b15zdnd00an1n02x5 FILLER_218_637 ();
 b15zdnd11an1n64x5 FILLER_218_642 ();
 b15zdnd11an1n08x5 FILLER_218_706 ();
 b15zdnd11an1n04x5 FILLER_218_714 ();
 b15zdnd11an1n64x5 FILLER_218_726 ();
 b15zdnd11an1n64x5 FILLER_218_790 ();
 b15zdnd11an1n32x5 FILLER_218_854 ();
 b15zdnd11an1n08x5 FILLER_218_886 ();
 b15zdnd11an1n04x5 FILLER_218_894 ();
 b15zdnd00an1n01x5 FILLER_218_898 ();
 b15zdnd11an1n04x5 FILLER_218_913 ();
 b15zdnd11an1n16x5 FILLER_218_920 ();
 b15zdnd11an1n08x5 FILLER_218_936 ();
 b15zdnd00an1n01x5 FILLER_218_944 ();
 b15zdnd11an1n64x5 FILLER_218_948 ();
 b15zdnd11an1n64x5 FILLER_218_1012 ();
 b15zdnd11an1n64x5 FILLER_218_1076 ();
 b15zdnd11an1n64x5 FILLER_218_1140 ();
 b15zdnd11an1n64x5 FILLER_218_1204 ();
 b15zdnd00an1n02x5 FILLER_218_1268 ();
 b15zdnd00an1n01x5 FILLER_218_1270 ();
 b15zdnd11an1n32x5 FILLER_218_1285 ();
 b15zdnd11an1n08x5 FILLER_218_1317 ();
 b15zdnd11an1n64x5 FILLER_218_1345 ();
 b15zdnd11an1n64x5 FILLER_218_1409 ();
 b15zdnd11an1n64x5 FILLER_218_1473 ();
 b15zdnd11an1n32x5 FILLER_218_1537 ();
 b15zdnd00an1n01x5 FILLER_218_1569 ();
 b15zdnd11an1n32x5 FILLER_218_1622 ();
 b15zdnd11an1n16x5 FILLER_218_1654 ();
 b15zdnd11an1n08x5 FILLER_218_1670 ();
 b15zdnd00an1n02x5 FILLER_218_1678 ();
 b15zdnd11an1n04x5 FILLER_218_1683 ();
 b15zdnd11an1n64x5 FILLER_218_1690 ();
 b15zdnd11an1n64x5 FILLER_218_1754 ();
 b15zdnd11an1n64x5 FILLER_218_1818 ();
 b15zdnd11an1n64x5 FILLER_218_1882 ();
 b15zdnd11an1n64x5 FILLER_218_1946 ();
 b15zdnd11an1n16x5 FILLER_218_2010 ();
 b15zdnd00an1n01x5 FILLER_218_2026 ();
 b15zdnd11an1n04x5 FILLER_218_2034 ();
 b15zdnd00an1n02x5 FILLER_218_2038 ();
 b15zdnd00an1n01x5 FILLER_218_2040 ();
 b15zdnd11an1n04x5 FILLER_218_2093 ();
 b15zdnd11an1n04x5 FILLER_218_2104 ();
 b15zdnd11an1n04x5 FILLER_218_2115 ();
 b15zdnd11an1n16x5 FILLER_218_2126 ();
 b15zdnd11an1n08x5 FILLER_218_2142 ();
 b15zdnd11an1n04x5 FILLER_218_2150 ();
 b15zdnd11an1n16x5 FILLER_218_2162 ();
 b15zdnd11an1n04x5 FILLER_218_2202 ();
 b15zdnd11an1n04x5 FILLER_218_2248 ();
 b15zdnd11an1n04x5 FILLER_218_2256 ();
 b15zdnd11an1n04x5 FILLER_218_2264 ();
 b15zdnd00an1n02x5 FILLER_218_2268 ();
 b15zdnd00an1n02x5 FILLER_218_2274 ();
 b15zdnd11an1n64x5 FILLER_219_0 ();
 b15zdnd11an1n08x5 FILLER_219_64 ();
 b15zdnd11an1n04x5 FILLER_219_72 ();
 b15zdnd11an1n32x5 FILLER_219_80 ();
 b15zdnd11an1n04x5 FILLER_219_112 ();
 b15zdnd11an1n04x5 FILLER_219_119 ();
 b15zdnd11an1n04x5 FILLER_219_126 ();
 b15zdnd11an1n16x5 FILLER_219_133 ();
 b15zdnd11an1n08x5 FILLER_219_149 ();
 b15zdnd00an1n02x5 FILLER_219_157 ();
 b15zdnd11an1n04x5 FILLER_219_191 ();
 b15zdnd11an1n04x5 FILLER_219_198 ();
 b15zdnd00an1n02x5 FILLER_219_202 ();
 b15zdnd00an1n01x5 FILLER_219_204 ();
 b15zdnd11an1n32x5 FILLER_219_208 ();
 b15zdnd11an1n04x5 FILLER_219_240 ();
 b15zdnd00an1n02x5 FILLER_219_244 ();
 b15zdnd11an1n64x5 FILLER_219_288 ();
 b15zdnd11an1n64x5 FILLER_219_352 ();
 b15zdnd11an1n32x5 FILLER_219_416 ();
 b15zdnd11an1n16x5 FILLER_219_448 ();
 b15zdnd11an1n08x5 FILLER_219_467 ();
 b15zdnd11an1n32x5 FILLER_219_517 ();
 b15zdnd11an1n16x5 FILLER_219_549 ();
 b15zdnd00an1n01x5 FILLER_219_565 ();
 b15zdnd11an1n32x5 FILLER_219_573 ();
 b15zdnd11an1n04x5 FILLER_219_605 ();
 b15zdnd00an1n02x5 FILLER_219_609 ();
 b15zdnd00an1n01x5 FILLER_219_611 ();
 b15zdnd11an1n64x5 FILLER_219_664 ();
 b15zdnd11an1n64x5 FILLER_219_728 ();
 b15zdnd11an1n32x5 FILLER_219_792 ();
 b15zdnd11an1n08x5 FILLER_219_824 ();
 b15zdnd00an1n01x5 FILLER_219_832 ();
 b15zdnd11an1n16x5 FILLER_219_875 ();
 b15zdnd11an1n04x5 FILLER_219_891 ();
 b15zdnd11an1n04x5 FILLER_219_947 ();
 b15zdnd11an1n64x5 FILLER_219_954 ();
 b15zdnd11an1n64x5 FILLER_219_1018 ();
 b15zdnd11an1n64x5 FILLER_219_1082 ();
 b15zdnd11an1n32x5 FILLER_219_1146 ();
 b15zdnd11an1n04x5 FILLER_219_1178 ();
 b15zdnd00an1n02x5 FILLER_219_1182 ();
 b15zdnd11an1n64x5 FILLER_219_1204 ();
 b15zdnd11an1n64x5 FILLER_219_1268 ();
 b15zdnd11an1n64x5 FILLER_219_1332 ();
 b15zdnd11an1n64x5 FILLER_219_1396 ();
 b15zdnd11an1n64x5 FILLER_219_1460 ();
 b15zdnd11an1n32x5 FILLER_219_1524 ();
 b15zdnd11an1n04x5 FILLER_219_1556 ();
 b15zdnd11an1n08x5 FILLER_219_1577 ();
 b15zdnd00an1n02x5 FILLER_219_1585 ();
 b15zdnd00an1n01x5 FILLER_219_1587 ();
 b15zdnd11an1n04x5 FILLER_219_1591 ();
 b15zdnd11an1n16x5 FILLER_219_1598 ();
 b15zdnd00an1n01x5 FILLER_219_1614 ();
 b15zdnd11an1n32x5 FILLER_219_1618 ();
 b15zdnd00an1n02x5 FILLER_219_1650 ();
 b15zdnd00an1n01x5 FILLER_219_1652 ();
 b15zdnd11an1n64x5 FILLER_219_1705 ();
 b15zdnd11an1n64x5 FILLER_219_1769 ();
 b15zdnd11an1n64x5 FILLER_219_1833 ();
 b15zdnd11an1n64x5 FILLER_219_1897 ();
 b15zdnd11an1n64x5 FILLER_219_1961 ();
 b15zdnd11an1n04x5 FILLER_219_2077 ();
 b15zdnd11an1n04x5 FILLER_219_2085 ();
 b15zdnd11an1n08x5 FILLER_219_2131 ();
 b15zdnd00an1n02x5 FILLER_219_2139 ();
 b15zdnd11an1n04x5 FILLER_219_2183 ();
 b15zdnd11an1n04x5 FILLER_219_2239 ();
 b15zdnd11an1n04x5 FILLER_219_2250 ();
 b15zdnd11an1n04x5 FILLER_219_2258 ();
 b15zdnd11an1n04x5 FILLER_219_2266 ();
 b15zdnd11an1n04x5 FILLER_219_2274 ();
 b15zdnd00an1n02x5 FILLER_219_2282 ();
 b15zdnd00an1n02x5 FILLER_220_8 ();
 b15zdnd11an1n08x5 FILLER_220_36 ();
 b15zdnd11an1n04x5 FILLER_220_44 ();
 b15zdnd00an1n01x5 FILLER_220_48 ();
 b15zdnd11an1n04x5 FILLER_220_75 ();
 b15zdnd11an1n08x5 FILLER_220_88 ();
 b15zdnd00an1n01x5 FILLER_220_96 ();
 b15zdnd11an1n32x5 FILLER_220_149 ();
 b15zdnd11an1n04x5 FILLER_220_184 ();
 b15zdnd11an1n32x5 FILLER_220_191 ();
 b15zdnd00an1n02x5 FILLER_220_223 ();
 b15zdnd00an1n01x5 FILLER_220_225 ();
 b15zdnd11an1n16x5 FILLER_220_268 ();
 b15zdnd11an1n04x5 FILLER_220_284 ();
 b15zdnd00an1n02x5 FILLER_220_288 ();
 b15zdnd11an1n64x5 FILLER_220_293 ();
 b15zdnd11an1n64x5 FILLER_220_357 ();
 b15zdnd11an1n64x5 FILLER_220_421 ();
 b15zdnd11an1n64x5 FILLER_220_485 ();
 b15zdnd11an1n64x5 FILLER_220_549 ();
 b15zdnd11an1n16x5 FILLER_220_613 ();
 b15zdnd11an1n08x5 FILLER_220_629 ();
 b15zdnd11an1n04x5 FILLER_220_640 ();
 b15zdnd11an1n64x5 FILLER_220_647 ();
 b15zdnd11an1n04x5 FILLER_220_711 ();
 b15zdnd00an1n02x5 FILLER_220_715 ();
 b15zdnd00an1n01x5 FILLER_220_717 ();
 b15zdnd11an1n64x5 FILLER_220_726 ();
 b15zdnd00an1n02x5 FILLER_220_790 ();
 b15zdnd00an1n01x5 FILLER_220_792 ();
 b15zdnd11an1n64x5 FILLER_220_845 ();
 b15zdnd11an1n08x5 FILLER_220_909 ();
 b15zdnd00an1n02x5 FILLER_220_917 ();
 b15zdnd11an1n64x5 FILLER_220_971 ();
 b15zdnd11an1n64x5 FILLER_220_1035 ();
 b15zdnd11an1n64x5 FILLER_220_1099 ();
 b15zdnd11an1n64x5 FILLER_220_1163 ();
 b15zdnd11an1n32x5 FILLER_220_1227 ();
 b15zdnd00an1n02x5 FILLER_220_1259 ();
 b15zdnd11an1n64x5 FILLER_220_1281 ();
 b15zdnd11an1n64x5 FILLER_220_1345 ();
 b15zdnd11an1n64x5 FILLER_220_1409 ();
 b15zdnd11an1n64x5 FILLER_220_1473 ();
 b15zdnd11an1n04x5 FILLER_220_1537 ();
 b15zdnd00an1n02x5 FILLER_220_1541 ();
 b15zdnd00an1n01x5 FILLER_220_1543 ();
 b15zdnd11an1n16x5 FILLER_220_1564 ();
 b15zdnd11an1n08x5 FILLER_220_1580 ();
 b15zdnd11an1n04x5 FILLER_220_1588 ();
 b15zdnd00an1n02x5 FILLER_220_1592 ();
 b15zdnd11an1n32x5 FILLER_220_1597 ();
 b15zdnd11an1n16x5 FILLER_220_1629 ();
 b15zdnd11an1n08x5 FILLER_220_1645 ();
 b15zdnd11an1n04x5 FILLER_220_1653 ();
 b15zdnd00an1n02x5 FILLER_220_1657 ();
 b15zdnd11an1n64x5 FILLER_220_1711 ();
 b15zdnd11an1n16x5 FILLER_220_1775 ();
 b15zdnd11an1n04x5 FILLER_220_1791 ();
 b15zdnd00an1n01x5 FILLER_220_1795 ();
 b15zdnd11an1n04x5 FILLER_220_1799 ();
 b15zdnd11an1n64x5 FILLER_220_1806 ();
 b15zdnd11an1n64x5 FILLER_220_1870 ();
 b15zdnd11an1n64x5 FILLER_220_1934 ();
 b15zdnd11an1n32x5 FILLER_220_1998 ();
 b15zdnd11an1n08x5 FILLER_220_2030 ();
 b15zdnd11an1n04x5 FILLER_220_2038 ();
 b15zdnd00an1n02x5 FILLER_220_2042 ();
 b15zdnd00an1n01x5 FILLER_220_2044 ();
 b15zdnd11an1n04x5 FILLER_220_2048 ();
 b15zdnd11an1n04x5 FILLER_220_2055 ();
 b15zdnd11an1n04x5 FILLER_220_2062 ();
 b15zdnd00an1n01x5 FILLER_220_2066 ();
 b15zdnd11an1n08x5 FILLER_220_2070 ();
 b15zdnd11an1n04x5 FILLER_220_2078 ();
 b15zdnd00an1n01x5 FILLER_220_2082 ();
 b15zdnd11an1n16x5 FILLER_220_2125 ();
 b15zdnd11an1n08x5 FILLER_220_2141 ();
 b15zdnd11an1n04x5 FILLER_220_2149 ();
 b15zdnd00an1n01x5 FILLER_220_2153 ();
 b15zdnd00an1n02x5 FILLER_220_2162 ();
 b15zdnd00an1n01x5 FILLER_220_2164 ();
 b15zdnd11an1n04x5 FILLER_220_2168 ();
 b15zdnd11an1n04x5 FILLER_220_2175 ();
 b15zdnd11an1n04x5 FILLER_220_2182 ();
 b15zdnd11an1n04x5 FILLER_220_2228 ();
 b15zdnd00an1n02x5 FILLER_220_2274 ();
 b15zdnd11an1n64x5 FILLER_221_0 ();
 b15zdnd11an1n08x5 FILLER_221_64 ();
 b15zdnd00an1n02x5 FILLER_221_72 ();
 b15zdnd00an1n01x5 FILLER_221_74 ();
 b15zdnd11an1n32x5 FILLER_221_82 ();
 b15zdnd11an1n08x5 FILLER_221_114 ();
 b15zdnd00an1n01x5 FILLER_221_122 ();
 b15zdnd11an1n64x5 FILLER_221_175 ();
 b15zdnd11an1n64x5 FILLER_221_239 ();
 b15zdnd11an1n64x5 FILLER_221_303 ();
 b15zdnd11an1n64x5 FILLER_221_367 ();
 b15zdnd11an1n64x5 FILLER_221_431 ();
 b15zdnd11an1n64x5 FILLER_221_495 ();
 b15zdnd11an1n64x5 FILLER_221_559 ();
 b15zdnd11an1n64x5 FILLER_221_623 ();
 b15zdnd11an1n64x5 FILLER_221_687 ();
 b15zdnd11an1n32x5 FILLER_221_751 ();
 b15zdnd11an1n16x5 FILLER_221_783 ();
 b15zdnd11an1n04x5 FILLER_221_799 ();
 b15zdnd00an1n01x5 FILLER_221_803 ();
 b15zdnd11an1n32x5 FILLER_221_846 ();
 b15zdnd11an1n04x5 FILLER_221_890 ();
 b15zdnd11an1n04x5 FILLER_221_946 ();
 b15zdnd11an1n64x5 FILLER_221_953 ();
 b15zdnd11an1n64x5 FILLER_221_1017 ();
 b15zdnd11an1n64x5 FILLER_221_1081 ();
 b15zdnd11an1n32x5 FILLER_221_1145 ();
 b15zdnd11an1n08x5 FILLER_221_1177 ();
 b15zdnd11an1n04x5 FILLER_221_1185 ();
 b15zdnd11an1n64x5 FILLER_221_1192 ();
 b15zdnd00an1n02x5 FILLER_221_1256 ();
 b15zdnd00an1n01x5 FILLER_221_1258 ();
 b15zdnd11an1n64x5 FILLER_221_1273 ();
 b15zdnd11an1n64x5 FILLER_221_1337 ();
 b15zdnd11an1n32x5 FILLER_221_1401 ();
 b15zdnd00an1n02x5 FILLER_221_1433 ();
 b15zdnd00an1n01x5 FILLER_221_1435 ();
 b15zdnd11an1n16x5 FILLER_221_1457 ();
 b15zdnd11an1n08x5 FILLER_221_1473 ();
 b15zdnd00an1n02x5 FILLER_221_1481 ();
 b15zdnd00an1n01x5 FILLER_221_1483 ();
 b15zdnd11an1n64x5 FILLER_221_1504 ();
 b15zdnd11an1n64x5 FILLER_221_1568 ();
 b15zdnd11an1n32x5 FILLER_221_1632 ();
 b15zdnd11an1n04x5 FILLER_221_1664 ();
 b15zdnd00an1n02x5 FILLER_221_1668 ();
 b15zdnd00an1n01x5 FILLER_221_1670 ();
 b15zdnd11an1n04x5 FILLER_221_1674 ();
 b15zdnd11an1n04x5 FILLER_221_1681 ();
 b15zdnd11an1n64x5 FILLER_221_1688 ();
 b15zdnd11an1n16x5 FILLER_221_1752 ();
 b15zdnd11an1n08x5 FILLER_221_1768 ();
 b15zdnd00an1n02x5 FILLER_221_1776 ();
 b15zdnd11an1n32x5 FILLER_221_1830 ();
 b15zdnd11an1n16x5 FILLER_221_1862 ();
 b15zdnd11an1n08x5 FILLER_221_1878 ();
 b15zdnd00an1n02x5 FILLER_221_1886 ();
 b15zdnd11an1n64x5 FILLER_221_1940 ();
 b15zdnd11an1n64x5 FILLER_221_2004 ();
 b15zdnd11an1n64x5 FILLER_221_2068 ();
 b15zdnd11an1n16x5 FILLER_221_2132 ();
 b15zdnd11an1n04x5 FILLER_221_2148 ();
 b15zdnd11an1n08x5 FILLER_221_2194 ();
 b15zdnd00an1n01x5 FILLER_221_2202 ();
 b15zdnd11an1n04x5 FILLER_221_2236 ();
 b15zdnd00an1n02x5 FILLER_221_2282 ();
 b15zdnd11an1n64x5 FILLER_222_8 ();
 b15zdnd11an1n04x5 FILLER_222_72 ();
 b15zdnd11an1n64x5 FILLER_222_79 ();
 b15zdnd11an1n04x5 FILLER_222_146 ();
 b15zdnd11an1n04x5 FILLER_222_153 ();
 b15zdnd11an1n64x5 FILLER_222_160 ();
 b15zdnd11an1n64x5 FILLER_222_224 ();
 b15zdnd11an1n64x5 FILLER_222_288 ();
 b15zdnd11an1n64x5 FILLER_222_352 ();
 b15zdnd11an1n64x5 FILLER_222_416 ();
 b15zdnd11an1n64x5 FILLER_222_480 ();
 b15zdnd11an1n64x5 FILLER_222_544 ();
 b15zdnd11an1n64x5 FILLER_222_608 ();
 b15zdnd11an1n32x5 FILLER_222_672 ();
 b15zdnd11an1n08x5 FILLER_222_704 ();
 b15zdnd11an1n04x5 FILLER_222_712 ();
 b15zdnd00an1n02x5 FILLER_222_716 ();
 b15zdnd11an1n64x5 FILLER_222_726 ();
 b15zdnd11an1n16x5 FILLER_222_790 ();
 b15zdnd11an1n04x5 FILLER_222_806 ();
 b15zdnd00an1n02x5 FILLER_222_810 ();
 b15zdnd00an1n01x5 FILLER_222_812 ();
 b15zdnd11an1n04x5 FILLER_222_816 ();
 b15zdnd11an1n04x5 FILLER_222_823 ();
 b15zdnd11an1n64x5 FILLER_222_830 ();
 b15zdnd11an1n16x5 FILLER_222_894 ();
 b15zdnd11an1n04x5 FILLER_222_910 ();
 b15zdnd00an1n01x5 FILLER_222_914 ();
 b15zdnd11an1n04x5 FILLER_222_918 ();
 b15zdnd11an1n04x5 FILLER_222_925 ();
 b15zdnd11an1n64x5 FILLER_222_932 ();
 b15zdnd11an1n64x5 FILLER_222_996 ();
 b15zdnd11an1n04x5 FILLER_222_1060 ();
 b15zdnd00an1n01x5 FILLER_222_1064 ();
 b15zdnd11an1n64x5 FILLER_222_1085 ();
 b15zdnd11an1n32x5 FILLER_222_1149 ();
 b15zdnd00an1n02x5 FILLER_222_1181 ();
 b15zdnd11an1n04x5 FILLER_222_1186 ();
 b15zdnd11an1n64x5 FILLER_222_1193 ();
 b15zdnd11an1n64x5 FILLER_222_1257 ();
 b15zdnd11an1n64x5 FILLER_222_1321 ();
 b15zdnd11an1n32x5 FILLER_222_1385 ();
 b15zdnd11an1n16x5 FILLER_222_1417 ();
 b15zdnd11an1n08x5 FILLER_222_1433 ();
 b15zdnd00an1n02x5 FILLER_222_1441 ();
 b15zdnd11an1n08x5 FILLER_222_1457 ();
 b15zdnd11an1n04x5 FILLER_222_1465 ();
 b15zdnd11an1n64x5 FILLER_222_1476 ();
 b15zdnd11an1n64x5 FILLER_222_1540 ();
 b15zdnd11an1n64x5 FILLER_222_1604 ();
 b15zdnd11an1n16x5 FILLER_222_1668 ();
 b15zdnd00an1n01x5 FILLER_222_1684 ();
 b15zdnd11an1n64x5 FILLER_222_1688 ();
 b15zdnd11an1n16x5 FILLER_222_1752 ();
 b15zdnd11an1n04x5 FILLER_222_1768 ();
 b15zdnd00an1n02x5 FILLER_222_1772 ();
 b15zdnd11an1n16x5 FILLER_222_1777 ();
 b15zdnd11an1n08x5 FILLER_222_1793 ();
 b15zdnd00an1n02x5 FILLER_222_1801 ();
 b15zdnd11an1n64x5 FILLER_222_1806 ();
 b15zdnd11an1n32x5 FILLER_222_1870 ();
 b15zdnd11an1n04x5 FILLER_222_1902 ();
 b15zdnd11an1n04x5 FILLER_222_1909 ();
 b15zdnd11an1n64x5 FILLER_222_1916 ();
 b15zdnd11an1n64x5 FILLER_222_1980 ();
 b15zdnd11an1n08x5 FILLER_222_2044 ();
 b15zdnd11an1n04x5 FILLER_222_2052 ();
 b15zdnd00an1n02x5 FILLER_222_2056 ();
 b15zdnd11an1n32x5 FILLER_222_2100 ();
 b15zdnd11an1n16x5 FILLER_222_2132 ();
 b15zdnd11an1n04x5 FILLER_222_2148 ();
 b15zdnd00an1n02x5 FILLER_222_2152 ();
 b15zdnd11an1n04x5 FILLER_222_2162 ();
 b15zdnd00an1n01x5 FILLER_222_2166 ();
 b15zdnd11an1n04x5 FILLER_222_2209 ();
 b15zdnd11an1n04x5 FILLER_222_2228 ();
 b15zdnd00an1n02x5 FILLER_222_2274 ();
 b15zdnd11an1n64x5 FILLER_223_0 ();
 b15zdnd11an1n64x5 FILLER_223_64 ();
 b15zdnd11an1n64x5 FILLER_223_128 ();
 b15zdnd11an1n64x5 FILLER_223_192 ();
 b15zdnd11an1n64x5 FILLER_223_256 ();
 b15zdnd11an1n64x5 FILLER_223_320 ();
 b15zdnd11an1n64x5 FILLER_223_384 ();
 b15zdnd11an1n64x5 FILLER_223_448 ();
 b15zdnd11an1n64x5 FILLER_223_512 ();
 b15zdnd11an1n64x5 FILLER_223_576 ();
 b15zdnd11an1n64x5 FILLER_223_640 ();
 b15zdnd11an1n64x5 FILLER_223_704 ();
 b15zdnd11an1n64x5 FILLER_223_768 ();
 b15zdnd11an1n64x5 FILLER_223_832 ();
 b15zdnd11an1n16x5 FILLER_223_896 ();
 b15zdnd11an1n04x5 FILLER_223_912 ();
 b15zdnd00an1n02x5 FILLER_223_916 ();
 b15zdnd00an1n01x5 FILLER_223_918 ();
 b15zdnd11an1n64x5 FILLER_223_922 ();
 b15zdnd11an1n64x5 FILLER_223_986 ();
 b15zdnd11an1n08x5 FILLER_223_1050 ();
 b15zdnd11an1n04x5 FILLER_223_1058 ();
 b15zdnd00an1n02x5 FILLER_223_1062 ();
 b15zdnd11an1n32x5 FILLER_223_1116 ();
 b15zdnd11an1n16x5 FILLER_223_1148 ();
 b15zdnd00an1n01x5 FILLER_223_1164 ();
 b15zdnd11an1n04x5 FILLER_223_1217 ();
 b15zdnd11an1n08x5 FILLER_223_1229 ();
 b15zdnd11an1n64x5 FILLER_223_1249 ();
 b15zdnd11an1n32x5 FILLER_223_1313 ();
 b15zdnd11an1n16x5 FILLER_223_1345 ();
 b15zdnd00an1n01x5 FILLER_223_1361 ();
 b15zdnd11an1n64x5 FILLER_223_1379 ();
 b15zdnd11an1n32x5 FILLER_223_1443 ();
 b15zdnd00an1n01x5 FILLER_223_1475 ();
 b15zdnd11an1n64x5 FILLER_223_1493 ();
 b15zdnd11an1n64x5 FILLER_223_1557 ();
 b15zdnd11an1n64x5 FILLER_223_1621 ();
 b15zdnd11an1n64x5 FILLER_223_1685 ();
 b15zdnd11an1n16x5 FILLER_223_1749 ();
 b15zdnd11an1n08x5 FILLER_223_1765 ();
 b15zdnd11an1n64x5 FILLER_223_1800 ();
 b15zdnd11an1n32x5 FILLER_223_1864 ();
 b15zdnd11an1n16x5 FILLER_223_1896 ();
 b15zdnd11an1n16x5 FILLER_223_1915 ();
 b15zdnd00an1n02x5 FILLER_223_1931 ();
 b15zdnd00an1n01x5 FILLER_223_1933 ();
 b15zdnd11an1n04x5 FILLER_223_1937 ();
 b15zdnd11an1n64x5 FILLER_223_1944 ();
 b15zdnd11an1n32x5 FILLER_223_2008 ();
 b15zdnd11an1n08x5 FILLER_223_2040 ();
 b15zdnd00an1n01x5 FILLER_223_2048 ();
 b15zdnd11an1n32x5 FILLER_223_2091 ();
 b15zdnd11an1n08x5 FILLER_223_2123 ();
 b15zdnd00an1n02x5 FILLER_223_2131 ();
 b15zdnd00an1n01x5 FILLER_223_2133 ();
 b15zdnd11an1n08x5 FILLER_223_2186 ();
 b15zdnd11an1n04x5 FILLER_223_2236 ();
 b15zdnd00an1n02x5 FILLER_223_2282 ();
 b15zdnd11an1n64x5 FILLER_224_8 ();
 b15zdnd00an1n02x5 FILLER_224_72 ();
 b15zdnd11an1n64x5 FILLER_224_82 ();
 b15zdnd11an1n64x5 FILLER_224_146 ();
 b15zdnd11an1n64x5 FILLER_224_210 ();
 b15zdnd11an1n64x5 FILLER_224_274 ();
 b15zdnd11an1n32x5 FILLER_224_338 ();
 b15zdnd11an1n16x5 FILLER_224_370 ();
 b15zdnd00an1n02x5 FILLER_224_386 ();
 b15zdnd00an1n01x5 FILLER_224_388 ();
 b15zdnd11an1n64x5 FILLER_224_392 ();
 b15zdnd11an1n64x5 FILLER_224_456 ();
 b15zdnd11an1n64x5 FILLER_224_520 ();
 b15zdnd11an1n64x5 FILLER_224_584 ();
 b15zdnd11an1n64x5 FILLER_224_648 ();
 b15zdnd11an1n04x5 FILLER_224_712 ();
 b15zdnd00an1n02x5 FILLER_224_716 ();
 b15zdnd11an1n64x5 FILLER_224_726 ();
 b15zdnd11an1n64x5 FILLER_224_790 ();
 b15zdnd11an1n64x5 FILLER_224_854 ();
 b15zdnd11an1n64x5 FILLER_224_918 ();
 b15zdnd11an1n64x5 FILLER_224_982 ();
 b15zdnd00an1n02x5 FILLER_224_1046 ();
 b15zdnd11an1n04x5 FILLER_224_1100 ();
 b15zdnd11an1n64x5 FILLER_224_1107 ();
 b15zdnd11an1n32x5 FILLER_224_1171 ();
 b15zdnd11an1n04x5 FILLER_224_1203 ();
 b15zdnd11an1n16x5 FILLER_224_1215 ();
 b15zdnd11an1n08x5 FILLER_224_1231 ();
 b15zdnd11an1n04x5 FILLER_224_1239 ();
 b15zdnd11an1n64x5 FILLER_224_1251 ();
 b15zdnd11an1n64x5 FILLER_224_1315 ();
 b15zdnd11an1n32x5 FILLER_224_1379 ();
 b15zdnd11an1n16x5 FILLER_224_1411 ();
 b15zdnd00an1n02x5 FILLER_224_1427 ();
 b15zdnd11an1n64x5 FILLER_224_1441 ();
 b15zdnd11an1n64x5 FILLER_224_1505 ();
 b15zdnd11an1n64x5 FILLER_224_1569 ();
 b15zdnd11an1n64x5 FILLER_224_1633 ();
 b15zdnd11an1n64x5 FILLER_224_1697 ();
 b15zdnd11an1n64x5 FILLER_224_1761 ();
 b15zdnd11an1n64x5 FILLER_224_1825 ();
 b15zdnd11an1n16x5 FILLER_224_1889 ();
 b15zdnd11an1n04x5 FILLER_224_1905 ();
 b15zdnd00an1n02x5 FILLER_224_1909 ();
 b15zdnd11an1n64x5 FILLER_224_1963 ();
 b15zdnd11an1n04x5 FILLER_224_2027 ();
 b15zdnd00an1n02x5 FILLER_224_2031 ();
 b15zdnd00an1n01x5 FILLER_224_2033 ();
 b15zdnd11an1n08x5 FILLER_224_2076 ();
 b15zdnd00an1n02x5 FILLER_224_2084 ();
 b15zdnd00an1n01x5 FILLER_224_2086 ();
 b15zdnd11an1n16x5 FILLER_224_2129 ();
 b15zdnd11an1n04x5 FILLER_224_2145 ();
 b15zdnd00an1n02x5 FILLER_224_2152 ();
 b15zdnd00an1n02x5 FILLER_224_2162 ();
 b15zdnd00an1n01x5 FILLER_224_2164 ();
 b15zdnd11an1n04x5 FILLER_224_2172 ();
 b15zdnd11an1n04x5 FILLER_224_2218 ();
 b15zdnd11an1n04x5 FILLER_224_2228 ();
 b15zdnd00an1n02x5 FILLER_224_2274 ();
 b15zdnd11an1n64x5 FILLER_225_0 ();
 b15zdnd11an1n64x5 FILLER_225_64 ();
 b15zdnd00an1n02x5 FILLER_225_128 ();
 b15zdnd00an1n01x5 FILLER_225_130 ();
 b15zdnd11an1n64x5 FILLER_225_173 ();
 b15zdnd11an1n32x5 FILLER_225_237 ();
 b15zdnd11an1n16x5 FILLER_225_269 ();
 b15zdnd00an1n02x5 FILLER_225_285 ();
 b15zdnd00an1n01x5 FILLER_225_287 ();
 b15zdnd11an1n16x5 FILLER_225_340 ();
 b15zdnd11an1n04x5 FILLER_225_356 ();
 b15zdnd00an1n02x5 FILLER_225_360 ();
 b15zdnd11an1n64x5 FILLER_225_414 ();
 b15zdnd11an1n08x5 FILLER_225_478 ();
 b15zdnd11an1n04x5 FILLER_225_486 ();
 b15zdnd00an1n02x5 FILLER_225_490 ();
 b15zdnd11an1n16x5 FILLER_225_498 ();
 b15zdnd11an1n08x5 FILLER_225_514 ();
 b15zdnd11an1n04x5 FILLER_225_522 ();
 b15zdnd11an1n08x5 FILLER_225_532 ();
 b15zdnd11an1n04x5 FILLER_225_540 ();
 b15zdnd00an1n02x5 FILLER_225_544 ();
 b15zdnd00an1n01x5 FILLER_225_546 ();
 b15zdnd11an1n64x5 FILLER_225_561 ();
 b15zdnd11an1n64x5 FILLER_225_625 ();
 b15zdnd11an1n64x5 FILLER_225_689 ();
 b15zdnd11an1n64x5 FILLER_225_753 ();
 b15zdnd11an1n64x5 FILLER_225_817 ();
 b15zdnd11an1n64x5 FILLER_225_881 ();
 b15zdnd11an1n64x5 FILLER_225_945 ();
 b15zdnd11an1n32x5 FILLER_225_1009 ();
 b15zdnd11an1n16x5 FILLER_225_1041 ();
 b15zdnd11an1n08x5 FILLER_225_1057 ();
 b15zdnd11an1n08x5 FILLER_225_1068 ();
 b15zdnd00an1n02x5 FILLER_225_1076 ();
 b15zdnd11an1n04x5 FILLER_225_1081 ();
 b15zdnd11an1n04x5 FILLER_225_1088 ();
 b15zdnd11an1n64x5 FILLER_225_1095 ();
 b15zdnd11an1n16x5 FILLER_225_1159 ();
 b15zdnd11an1n04x5 FILLER_225_1175 ();
 b15zdnd00an1n02x5 FILLER_225_1179 ();
 b15zdnd00an1n01x5 FILLER_225_1181 ();
 b15zdnd11an1n04x5 FILLER_225_1185 ();
 b15zdnd11an1n64x5 FILLER_225_1192 ();
 b15zdnd11an1n64x5 FILLER_225_1256 ();
 b15zdnd11an1n64x5 FILLER_225_1320 ();
 b15zdnd00an1n02x5 FILLER_225_1384 ();
 b15zdnd00an1n01x5 FILLER_225_1386 ();
 b15zdnd11an1n64x5 FILLER_225_1407 ();
 b15zdnd11an1n64x5 FILLER_225_1471 ();
 b15zdnd11an1n64x5 FILLER_225_1535 ();
 b15zdnd11an1n64x5 FILLER_225_1599 ();
 b15zdnd11an1n64x5 FILLER_225_1663 ();
 b15zdnd11an1n64x5 FILLER_225_1727 ();
 b15zdnd11an1n64x5 FILLER_225_1791 ();
 b15zdnd11an1n32x5 FILLER_225_1855 ();
 b15zdnd11an1n16x5 FILLER_225_1887 ();
 b15zdnd11an1n04x5 FILLER_225_1903 ();
 b15zdnd11an1n64x5 FILLER_225_1959 ();
 b15zdnd11an1n32x5 FILLER_225_2023 ();
 b15zdnd11an1n08x5 FILLER_225_2055 ();
 b15zdnd11an1n32x5 FILLER_225_2105 ();
 b15zdnd11an1n16x5 FILLER_225_2137 ();
 b15zdnd00an1n01x5 FILLER_225_2153 ();
 b15zdnd11an1n04x5 FILLER_225_2157 ();
 b15zdnd11an1n04x5 FILLER_225_2203 ();
 b15zdnd11an1n08x5 FILLER_225_2249 ();
 b15zdnd00an1n02x5 FILLER_225_2257 ();
 b15zdnd00an1n01x5 FILLER_225_2259 ();
 b15zdnd11an1n04x5 FILLER_225_2264 ();
 b15zdnd11an1n04x5 FILLER_225_2272 ();
 b15zdnd11an1n04x5 FILLER_225_2280 ();
 b15zdnd11an1n64x5 FILLER_226_8 ();
 b15zdnd11an1n64x5 FILLER_226_72 ();
 b15zdnd11an1n08x5 FILLER_226_136 ();
 b15zdnd11an1n04x5 FILLER_226_144 ();
 b15zdnd00an1n02x5 FILLER_226_148 ();
 b15zdnd00an1n01x5 FILLER_226_150 ();
 b15zdnd11an1n64x5 FILLER_226_193 ();
 b15zdnd11an1n32x5 FILLER_226_257 ();
 b15zdnd11an1n16x5 FILLER_226_289 ();
 b15zdnd00an1n02x5 FILLER_226_305 ();
 b15zdnd00an1n01x5 FILLER_226_307 ();
 b15zdnd11an1n04x5 FILLER_226_311 ();
 b15zdnd11an1n04x5 FILLER_226_318 ();
 b15zdnd11an1n32x5 FILLER_226_325 ();
 b15zdnd11an1n16x5 FILLER_226_357 ();
 b15zdnd11an1n04x5 FILLER_226_373 ();
 b15zdnd00an1n02x5 FILLER_226_377 ();
 b15zdnd00an1n01x5 FILLER_226_379 ();
 b15zdnd11an1n04x5 FILLER_226_383 ();
 b15zdnd11an1n32x5 FILLER_226_390 ();
 b15zdnd11an1n08x5 FILLER_226_422 ();
 b15zdnd00an1n02x5 FILLER_226_430 ();
 b15zdnd11an1n04x5 FILLER_226_441 ();
 b15zdnd00an1n02x5 FILLER_226_445 ();
 b15zdnd00an1n01x5 FILLER_226_447 ();
 b15zdnd11an1n64x5 FILLER_226_456 ();
 b15zdnd11an1n64x5 FILLER_226_520 ();
 b15zdnd11an1n04x5 FILLER_226_584 ();
 b15zdnd00an1n01x5 FILLER_226_588 ();
 b15zdnd11an1n64x5 FILLER_226_597 ();
 b15zdnd11an1n32x5 FILLER_226_661 ();
 b15zdnd11an1n16x5 FILLER_226_693 ();
 b15zdnd11an1n08x5 FILLER_226_709 ();
 b15zdnd00an1n01x5 FILLER_226_717 ();
 b15zdnd11an1n64x5 FILLER_226_726 ();
 b15zdnd11an1n64x5 FILLER_226_790 ();
 b15zdnd11an1n64x5 FILLER_226_854 ();
 b15zdnd11an1n64x5 FILLER_226_918 ();
 b15zdnd11an1n64x5 FILLER_226_982 ();
 b15zdnd11an1n16x5 FILLER_226_1046 ();
 b15zdnd11an1n04x5 FILLER_226_1062 ();
 b15zdnd00an1n02x5 FILLER_226_1066 ();
 b15zdnd11an1n32x5 FILLER_226_1071 ();
 b15zdnd11an1n16x5 FILLER_226_1103 ();
 b15zdnd11an1n08x5 FILLER_226_1119 ();
 b15zdnd11an1n16x5 FILLER_226_1136 ();
 b15zdnd11an1n08x5 FILLER_226_1152 ();
 b15zdnd11an1n04x5 FILLER_226_1160 ();
 b15zdnd11an1n64x5 FILLER_226_1216 ();
 b15zdnd11an1n64x5 FILLER_226_1280 ();
 b15zdnd11an1n16x5 FILLER_226_1344 ();
 b15zdnd11an1n08x5 FILLER_226_1360 ();
 b15zdnd00an1n02x5 FILLER_226_1368 ();
 b15zdnd00an1n01x5 FILLER_226_1370 ();
 b15zdnd11an1n64x5 FILLER_226_1383 ();
 b15zdnd11an1n64x5 FILLER_226_1447 ();
 b15zdnd00an1n02x5 FILLER_226_1511 ();
 b15zdnd11an1n64x5 FILLER_226_1530 ();
 b15zdnd11an1n64x5 FILLER_226_1594 ();
 b15zdnd11an1n64x5 FILLER_226_1658 ();
 b15zdnd11an1n64x5 FILLER_226_1722 ();
 b15zdnd11an1n64x5 FILLER_226_1786 ();
 b15zdnd11an1n64x5 FILLER_226_1850 ();
 b15zdnd11an1n08x5 FILLER_226_1914 ();
 b15zdnd00an1n02x5 FILLER_226_1922 ();
 b15zdnd00an1n01x5 FILLER_226_1924 ();
 b15zdnd11an1n04x5 FILLER_226_1928 ();
 b15zdnd11an1n04x5 FILLER_226_1935 ();
 b15zdnd11an1n64x5 FILLER_226_1942 ();
 b15zdnd11an1n64x5 FILLER_226_2006 ();
 b15zdnd11an1n64x5 FILLER_226_2070 ();
 b15zdnd11an1n16x5 FILLER_226_2134 ();
 b15zdnd11an1n04x5 FILLER_226_2150 ();
 b15zdnd11an1n04x5 FILLER_226_2162 ();
 b15zdnd00an1n02x5 FILLER_226_2166 ();
 b15zdnd11an1n04x5 FILLER_226_2210 ();
 b15zdnd11an1n04x5 FILLER_226_2259 ();
 b15zdnd11an1n08x5 FILLER_226_2267 ();
 b15zdnd00an1n01x5 FILLER_226_2275 ();
 b15zdnd11an1n64x5 FILLER_227_0 ();
 b15zdnd11an1n32x5 FILLER_227_64 ();
 b15zdnd11an1n16x5 FILLER_227_96 ();
 b15zdnd11an1n64x5 FILLER_227_154 ();
 b15zdnd11an1n64x5 FILLER_227_218 ();
 b15zdnd11an1n64x5 FILLER_227_282 ();
 b15zdnd11an1n64x5 FILLER_227_346 ();
 b15zdnd11an1n64x5 FILLER_227_410 ();
 b15zdnd11an1n64x5 FILLER_227_474 ();
 b15zdnd11an1n64x5 FILLER_227_538 ();
 b15zdnd11an1n64x5 FILLER_227_602 ();
 b15zdnd11an1n64x5 FILLER_227_666 ();
 b15zdnd11an1n64x5 FILLER_227_730 ();
 b15zdnd11an1n64x5 FILLER_227_794 ();
 b15zdnd11an1n64x5 FILLER_227_858 ();
 b15zdnd11an1n64x5 FILLER_227_922 ();
 b15zdnd11an1n32x5 FILLER_227_986 ();
 b15zdnd11an1n04x5 FILLER_227_1018 ();
 b15zdnd11an1n64x5 FILLER_227_1033 ();
 b15zdnd11an1n64x5 FILLER_227_1097 ();
 b15zdnd11an1n16x5 FILLER_227_1161 ();
 b15zdnd11an1n08x5 FILLER_227_1177 ();
 b15zdnd11an1n04x5 FILLER_227_1185 ();
 b15zdnd00an1n01x5 FILLER_227_1189 ();
 b15zdnd11an1n64x5 FILLER_227_1193 ();
 b15zdnd11an1n64x5 FILLER_227_1257 ();
 b15zdnd11an1n64x5 FILLER_227_1321 ();
 b15zdnd11an1n32x5 FILLER_227_1385 ();
 b15zdnd11an1n04x5 FILLER_227_1417 ();
 b15zdnd00an1n01x5 FILLER_227_1421 ();
 b15zdnd11an1n64x5 FILLER_227_1442 ();
 b15zdnd11an1n64x5 FILLER_227_1506 ();
 b15zdnd11an1n64x5 FILLER_227_1570 ();
 b15zdnd11an1n64x5 FILLER_227_1634 ();
 b15zdnd11an1n64x5 FILLER_227_1698 ();
 b15zdnd11an1n64x5 FILLER_227_1762 ();
 b15zdnd11an1n64x5 FILLER_227_1826 ();
 b15zdnd11an1n32x5 FILLER_227_1890 ();
 b15zdnd11an1n08x5 FILLER_227_1922 ();
 b15zdnd11an1n04x5 FILLER_227_1930 ();
 b15zdnd00an1n02x5 FILLER_227_1934 ();
 b15zdnd00an1n01x5 FILLER_227_1936 ();
 b15zdnd11an1n64x5 FILLER_227_1940 ();
 b15zdnd11an1n64x5 FILLER_227_2004 ();
 b15zdnd11an1n64x5 FILLER_227_2068 ();
 b15zdnd11an1n32x5 FILLER_227_2132 ();
 b15zdnd11an1n08x5 FILLER_227_2167 ();
 b15zdnd11an1n04x5 FILLER_227_2175 ();
 b15zdnd00an1n01x5 FILLER_227_2179 ();
 b15zdnd11an1n04x5 FILLER_227_2222 ();
 b15zdnd11an1n04x5 FILLER_227_2268 ();
 b15zdnd11an1n08x5 FILLER_227_2276 ();
 b15zdnd11an1n64x5 FILLER_228_8 ();
 b15zdnd11an1n64x5 FILLER_228_72 ();
 b15zdnd11an1n64x5 FILLER_228_136 ();
 b15zdnd11an1n08x5 FILLER_228_200 ();
 b15zdnd11an1n04x5 FILLER_228_208 ();
 b15zdnd11an1n64x5 FILLER_228_254 ();
 b15zdnd11an1n32x5 FILLER_228_318 ();
 b15zdnd11an1n16x5 FILLER_228_350 ();
 b15zdnd11an1n08x5 FILLER_228_366 ();
 b15zdnd00an1n02x5 FILLER_228_374 ();
 b15zdnd00an1n01x5 FILLER_228_376 ();
 b15zdnd11an1n64x5 FILLER_228_419 ();
 b15zdnd11an1n64x5 FILLER_228_483 ();
 b15zdnd11an1n64x5 FILLER_228_547 ();
 b15zdnd11an1n04x5 FILLER_228_611 ();
 b15zdnd00an1n02x5 FILLER_228_615 ();
 b15zdnd11an1n64x5 FILLER_228_623 ();
 b15zdnd11an1n16x5 FILLER_228_687 ();
 b15zdnd11an1n08x5 FILLER_228_703 ();
 b15zdnd11an1n04x5 FILLER_228_711 ();
 b15zdnd00an1n02x5 FILLER_228_715 ();
 b15zdnd00an1n01x5 FILLER_228_717 ();
 b15zdnd11an1n64x5 FILLER_228_726 ();
 b15zdnd11an1n64x5 FILLER_228_790 ();
 b15zdnd11an1n64x5 FILLER_228_854 ();
 b15zdnd11an1n64x5 FILLER_228_918 ();
 b15zdnd11an1n64x5 FILLER_228_982 ();
 b15zdnd11an1n64x5 FILLER_228_1046 ();
 b15zdnd11an1n64x5 FILLER_228_1110 ();
 b15zdnd11an1n64x5 FILLER_228_1174 ();
 b15zdnd11an1n64x5 FILLER_228_1238 ();
 b15zdnd11an1n32x5 FILLER_228_1302 ();
 b15zdnd11an1n16x5 FILLER_228_1334 ();
 b15zdnd00an1n02x5 FILLER_228_1350 ();
 b15zdnd11an1n64x5 FILLER_228_1372 ();
 b15zdnd11an1n64x5 FILLER_228_1436 ();
 b15zdnd11an1n64x5 FILLER_228_1500 ();
 b15zdnd11an1n64x5 FILLER_228_1564 ();
 b15zdnd11an1n64x5 FILLER_228_1628 ();
 b15zdnd11an1n64x5 FILLER_228_1692 ();
 b15zdnd11an1n64x5 FILLER_228_1756 ();
 b15zdnd11an1n32x5 FILLER_228_1820 ();
 b15zdnd11an1n04x5 FILLER_228_1852 ();
 b15zdnd00an1n02x5 FILLER_228_1856 ();
 b15zdnd00an1n01x5 FILLER_228_1858 ();
 b15zdnd11an1n64x5 FILLER_228_1901 ();
 b15zdnd11an1n64x5 FILLER_228_1965 ();
 b15zdnd11an1n64x5 FILLER_228_2029 ();
 b15zdnd11an1n32x5 FILLER_228_2093 ();
 b15zdnd11an1n16x5 FILLER_228_2125 ();
 b15zdnd11an1n08x5 FILLER_228_2141 ();
 b15zdnd11an1n04x5 FILLER_228_2149 ();
 b15zdnd00an1n01x5 FILLER_228_2153 ();
 b15zdnd11an1n16x5 FILLER_228_2162 ();
 b15zdnd11an1n08x5 FILLER_228_2178 ();
 b15zdnd11an1n04x5 FILLER_228_2228 ();
 b15zdnd00an1n02x5 FILLER_228_2274 ();
 b15zdnd11an1n64x5 FILLER_229_0 ();
 b15zdnd00an1n01x5 FILLER_229_64 ();
 b15zdnd11an1n08x5 FILLER_229_75 ();
 b15zdnd11an1n04x5 FILLER_229_83 ();
 b15zdnd11an1n64x5 FILLER_229_101 ();
 b15zdnd11an1n64x5 FILLER_229_165 ();
 b15zdnd11an1n64x5 FILLER_229_229 ();
 b15zdnd11an1n64x5 FILLER_229_293 ();
 b15zdnd11an1n64x5 FILLER_229_357 ();
 b15zdnd11an1n64x5 FILLER_229_421 ();
 b15zdnd11an1n64x5 FILLER_229_485 ();
 b15zdnd11an1n64x5 FILLER_229_549 ();
 b15zdnd11an1n64x5 FILLER_229_613 ();
 b15zdnd11an1n64x5 FILLER_229_677 ();
 b15zdnd11an1n16x5 FILLER_229_741 ();
 b15zdnd11an1n08x5 FILLER_229_757 ();
 b15zdnd00an1n02x5 FILLER_229_765 ();
 b15zdnd00an1n01x5 FILLER_229_767 ();
 b15zdnd11an1n64x5 FILLER_229_820 ();
 b15zdnd11an1n64x5 FILLER_229_884 ();
 b15zdnd11an1n64x5 FILLER_229_948 ();
 b15zdnd11an1n64x5 FILLER_229_1012 ();
 b15zdnd11an1n64x5 FILLER_229_1076 ();
 b15zdnd11an1n64x5 FILLER_229_1140 ();
 b15zdnd11an1n64x5 FILLER_229_1204 ();
 b15zdnd11an1n64x5 FILLER_229_1268 ();
 b15zdnd11an1n64x5 FILLER_229_1332 ();
 b15zdnd11an1n64x5 FILLER_229_1396 ();
 b15zdnd11an1n64x5 FILLER_229_1460 ();
 b15zdnd11an1n64x5 FILLER_229_1524 ();
 b15zdnd11an1n64x5 FILLER_229_1588 ();
 b15zdnd11an1n64x5 FILLER_229_1652 ();
 b15zdnd11an1n64x5 FILLER_229_1716 ();
 b15zdnd11an1n64x5 FILLER_229_1780 ();
 b15zdnd11an1n64x5 FILLER_229_1844 ();
 b15zdnd11an1n64x5 FILLER_229_1908 ();
 b15zdnd11an1n64x5 FILLER_229_1972 ();
 b15zdnd11an1n16x5 FILLER_229_2036 ();
 b15zdnd00an1n01x5 FILLER_229_2052 ();
 b15zdnd11an1n64x5 FILLER_229_2095 ();
 b15zdnd11an1n08x5 FILLER_229_2159 ();
 b15zdnd11an1n04x5 FILLER_229_2167 ();
 b15zdnd00an1n02x5 FILLER_229_2171 ();
 b15zdnd11an1n04x5 FILLER_229_2190 ();
 b15zdnd11an1n04x5 FILLER_229_2236 ();
 b15zdnd00an1n02x5 FILLER_229_2282 ();
 b15zdnd11an1n64x5 FILLER_230_8 ();
 b15zdnd00an1n01x5 FILLER_230_72 ();
 b15zdnd11an1n64x5 FILLER_230_115 ();
 b15zdnd11an1n64x5 FILLER_230_179 ();
 b15zdnd11an1n16x5 FILLER_230_243 ();
 b15zdnd11an1n04x5 FILLER_230_259 ();
 b15zdnd00an1n02x5 FILLER_230_263 ();
 b15zdnd11an1n64x5 FILLER_230_307 ();
 b15zdnd11an1n64x5 FILLER_230_371 ();
 b15zdnd11an1n64x5 FILLER_230_435 ();
 b15zdnd11an1n64x5 FILLER_230_499 ();
 b15zdnd11an1n64x5 FILLER_230_563 ();
 b15zdnd11an1n64x5 FILLER_230_627 ();
 b15zdnd11an1n16x5 FILLER_230_691 ();
 b15zdnd11an1n08x5 FILLER_230_707 ();
 b15zdnd00an1n02x5 FILLER_230_715 ();
 b15zdnd00an1n01x5 FILLER_230_717 ();
 b15zdnd11an1n32x5 FILLER_230_726 ();
 b15zdnd11an1n16x5 FILLER_230_758 ();
 b15zdnd11an1n08x5 FILLER_230_774 ();
 b15zdnd00an1n02x5 FILLER_230_782 ();
 b15zdnd11an1n64x5 FILLER_230_826 ();
 b15zdnd11an1n64x5 FILLER_230_890 ();
 b15zdnd11an1n64x5 FILLER_230_954 ();
 b15zdnd11an1n64x5 FILLER_230_1018 ();
 b15zdnd11an1n64x5 FILLER_230_1082 ();
 b15zdnd11an1n64x5 FILLER_230_1146 ();
 b15zdnd11an1n64x5 FILLER_230_1210 ();
 b15zdnd11an1n64x5 FILLER_230_1274 ();
 b15zdnd11an1n16x5 FILLER_230_1338 ();
 b15zdnd11an1n08x5 FILLER_230_1354 ();
 b15zdnd00an1n02x5 FILLER_230_1362 ();
 b15zdnd00an1n01x5 FILLER_230_1364 ();
 b15zdnd11an1n64x5 FILLER_230_1385 ();
 b15zdnd11an1n64x5 FILLER_230_1449 ();
 b15zdnd11an1n64x5 FILLER_230_1513 ();
 b15zdnd11an1n32x5 FILLER_230_1577 ();
 b15zdnd11an1n08x5 FILLER_230_1609 ();
 b15zdnd11an1n04x5 FILLER_230_1617 ();
 b15zdnd00an1n01x5 FILLER_230_1621 ();
 b15zdnd11an1n32x5 FILLER_230_1646 ();
 b15zdnd11an1n16x5 FILLER_230_1678 ();
 b15zdnd11an1n08x5 FILLER_230_1694 ();
 b15zdnd00an1n02x5 FILLER_230_1702 ();
 b15zdnd11an1n64x5 FILLER_230_1724 ();
 b15zdnd11an1n64x5 FILLER_230_1788 ();
 b15zdnd11an1n64x5 FILLER_230_1852 ();
 b15zdnd11an1n64x5 FILLER_230_1916 ();
 b15zdnd11an1n64x5 FILLER_230_1980 ();
 b15zdnd11an1n64x5 FILLER_230_2044 ();
 b15zdnd11an1n32x5 FILLER_230_2108 ();
 b15zdnd11an1n08x5 FILLER_230_2140 ();
 b15zdnd11an1n04x5 FILLER_230_2148 ();
 b15zdnd00an1n02x5 FILLER_230_2152 ();
 b15zdnd11an1n16x5 FILLER_230_2162 ();
 b15zdnd00an1n02x5 FILLER_230_2178 ();
 b15zdnd00an1n01x5 FILLER_230_2180 ();
 b15zdnd11an1n04x5 FILLER_230_2223 ();
 b15zdnd11an1n04x5 FILLER_230_2269 ();
 b15zdnd00an1n02x5 FILLER_230_2273 ();
 b15zdnd00an1n01x5 FILLER_230_2275 ();
 b15zdnd11an1n64x5 FILLER_231_0 ();
 b15zdnd11an1n08x5 FILLER_231_64 ();
 b15zdnd11an1n04x5 FILLER_231_72 ();
 b15zdnd00an1n02x5 FILLER_231_76 ();
 b15zdnd00an1n01x5 FILLER_231_78 ();
 b15zdnd11an1n08x5 FILLER_231_94 ();
 b15zdnd11an1n64x5 FILLER_231_144 ();
 b15zdnd11an1n64x5 FILLER_231_208 ();
 b15zdnd11an1n64x5 FILLER_231_272 ();
 b15zdnd11an1n64x5 FILLER_231_336 ();
 b15zdnd11an1n64x5 FILLER_231_400 ();
 b15zdnd11an1n16x5 FILLER_231_464 ();
 b15zdnd11an1n04x5 FILLER_231_480 ();
 b15zdnd00an1n01x5 FILLER_231_484 ();
 b15zdnd11an1n64x5 FILLER_231_491 ();
 b15zdnd11an1n64x5 FILLER_231_555 ();
 b15zdnd11an1n64x5 FILLER_231_619 ();
 b15zdnd11an1n64x5 FILLER_231_683 ();
 b15zdnd11an1n32x5 FILLER_231_747 ();
 b15zdnd11an1n08x5 FILLER_231_779 ();
 b15zdnd00an1n01x5 FILLER_231_787 ();
 b15zdnd11an1n04x5 FILLER_231_791 ();
 b15zdnd11an1n64x5 FILLER_231_798 ();
 b15zdnd11an1n64x5 FILLER_231_862 ();
 b15zdnd11an1n64x5 FILLER_231_926 ();
 b15zdnd11an1n64x5 FILLER_231_990 ();
 b15zdnd11an1n64x5 FILLER_231_1054 ();
 b15zdnd11an1n64x5 FILLER_231_1118 ();
 b15zdnd11an1n64x5 FILLER_231_1182 ();
 b15zdnd11an1n64x5 FILLER_231_1246 ();
 b15zdnd11an1n16x5 FILLER_231_1310 ();
 b15zdnd11an1n08x5 FILLER_231_1326 ();
 b15zdnd11an1n04x5 FILLER_231_1334 ();
 b15zdnd00an1n01x5 FILLER_231_1338 ();
 b15zdnd11an1n64x5 FILLER_231_1359 ();
 b15zdnd11an1n64x5 FILLER_231_1423 ();
 b15zdnd11an1n64x5 FILLER_231_1487 ();
 b15zdnd11an1n64x5 FILLER_231_1551 ();
 b15zdnd11an1n64x5 FILLER_231_1615 ();
 b15zdnd11an1n08x5 FILLER_231_1679 ();
 b15zdnd11an1n04x5 FILLER_231_1687 ();
 b15zdnd00an1n01x5 FILLER_231_1691 ();
 b15zdnd11an1n64x5 FILLER_231_1716 ();
 b15zdnd11an1n64x5 FILLER_231_1780 ();
 b15zdnd11an1n64x5 FILLER_231_1844 ();
 b15zdnd11an1n64x5 FILLER_231_1908 ();
 b15zdnd11an1n64x5 FILLER_231_1972 ();
 b15zdnd11an1n64x5 FILLER_231_2036 ();
 b15zdnd11an1n64x5 FILLER_231_2100 ();
 b15zdnd11an1n08x5 FILLER_231_2164 ();
 b15zdnd11an1n04x5 FILLER_231_2172 ();
 b15zdnd00an1n02x5 FILLER_231_2176 ();
 b15zdnd11an1n04x5 FILLER_231_2190 ();
 b15zdnd11an1n04x5 FILLER_231_2236 ();
 b15zdnd00an1n02x5 FILLER_231_2282 ();
 b15zdnd11an1n64x5 FILLER_232_8 ();
 b15zdnd11an1n64x5 FILLER_232_72 ();
 b15zdnd11an1n64x5 FILLER_232_136 ();
 b15zdnd11an1n64x5 FILLER_232_200 ();
 b15zdnd11an1n64x5 FILLER_232_264 ();
 b15zdnd11an1n64x5 FILLER_232_328 ();
 b15zdnd11an1n04x5 FILLER_232_392 ();
 b15zdnd00an1n02x5 FILLER_232_396 ();
 b15zdnd11an1n64x5 FILLER_232_414 ();
 b15zdnd11an1n64x5 FILLER_232_478 ();
 b15zdnd11an1n64x5 FILLER_232_542 ();
 b15zdnd11an1n64x5 FILLER_232_606 ();
 b15zdnd11an1n32x5 FILLER_232_670 ();
 b15zdnd11an1n16x5 FILLER_232_702 ();
 b15zdnd11an1n32x5 FILLER_232_726 ();
 b15zdnd11an1n16x5 FILLER_232_758 ();
 b15zdnd11an1n08x5 FILLER_232_774 ();
 b15zdnd11an1n04x5 FILLER_232_782 ();
 b15zdnd00an1n02x5 FILLER_232_786 ();
 b15zdnd00an1n01x5 FILLER_232_788 ();
 b15zdnd11an1n64x5 FILLER_232_792 ();
 b15zdnd11an1n64x5 FILLER_232_856 ();
 b15zdnd11an1n64x5 FILLER_232_920 ();
 b15zdnd11an1n64x5 FILLER_232_984 ();
 b15zdnd11an1n64x5 FILLER_232_1048 ();
 b15zdnd11an1n64x5 FILLER_232_1112 ();
 b15zdnd11an1n64x5 FILLER_232_1176 ();
 b15zdnd11an1n64x5 FILLER_232_1240 ();
 b15zdnd11an1n64x5 FILLER_232_1304 ();
 b15zdnd11an1n64x5 FILLER_232_1368 ();
 b15zdnd11an1n64x5 FILLER_232_1432 ();
 b15zdnd11an1n64x5 FILLER_232_1496 ();
 b15zdnd11an1n64x5 FILLER_232_1560 ();
 b15zdnd11an1n64x5 FILLER_232_1624 ();
 b15zdnd11an1n64x5 FILLER_232_1688 ();
 b15zdnd11an1n64x5 FILLER_232_1752 ();
 b15zdnd11an1n64x5 FILLER_232_1816 ();
 b15zdnd11an1n64x5 FILLER_232_1880 ();
 b15zdnd11an1n64x5 FILLER_232_1944 ();
 b15zdnd11an1n64x5 FILLER_232_2008 ();
 b15zdnd11an1n64x5 FILLER_232_2072 ();
 b15zdnd11an1n16x5 FILLER_232_2136 ();
 b15zdnd00an1n02x5 FILLER_232_2152 ();
 b15zdnd11an1n16x5 FILLER_232_2162 ();
 b15zdnd11an1n08x5 FILLER_232_2178 ();
 b15zdnd11an1n04x5 FILLER_232_2228 ();
 b15zdnd00an1n02x5 FILLER_232_2274 ();
 b15zdnd11an1n64x5 FILLER_233_0 ();
 b15zdnd11an1n64x5 FILLER_233_64 ();
 b15zdnd11an1n32x5 FILLER_233_128 ();
 b15zdnd11an1n08x5 FILLER_233_160 ();
 b15zdnd11an1n64x5 FILLER_233_186 ();
 b15zdnd11an1n64x5 FILLER_233_250 ();
 b15zdnd11an1n64x5 FILLER_233_314 ();
 b15zdnd11an1n64x5 FILLER_233_378 ();
 b15zdnd11an1n64x5 FILLER_233_442 ();
 b15zdnd11an1n64x5 FILLER_233_506 ();
 b15zdnd11an1n64x5 FILLER_233_570 ();
 b15zdnd11an1n32x5 FILLER_233_634 ();
 b15zdnd11an1n16x5 FILLER_233_666 ();
 b15zdnd11an1n08x5 FILLER_233_685 ();
 b15zdnd00an1n02x5 FILLER_233_693 ();
 b15zdnd11an1n64x5 FILLER_233_737 ();
 b15zdnd11an1n64x5 FILLER_233_801 ();
 b15zdnd11an1n64x5 FILLER_233_865 ();
 b15zdnd11an1n64x5 FILLER_233_929 ();
 b15zdnd11an1n64x5 FILLER_233_993 ();
 b15zdnd11an1n64x5 FILLER_233_1057 ();
 b15zdnd11an1n64x5 FILLER_233_1121 ();
 b15zdnd11an1n64x5 FILLER_233_1185 ();
 b15zdnd11an1n64x5 FILLER_233_1249 ();
 b15zdnd11an1n64x5 FILLER_233_1313 ();
 b15zdnd11an1n32x5 FILLER_233_1377 ();
 b15zdnd11an1n16x5 FILLER_233_1409 ();
 b15zdnd11an1n04x5 FILLER_233_1425 ();
 b15zdnd00an1n02x5 FILLER_233_1429 ();
 b15zdnd11an1n64x5 FILLER_233_1445 ();
 b15zdnd11an1n64x5 FILLER_233_1509 ();
 b15zdnd11an1n64x5 FILLER_233_1573 ();
 b15zdnd11an1n64x5 FILLER_233_1637 ();
 b15zdnd11an1n64x5 FILLER_233_1701 ();
 b15zdnd11an1n64x5 FILLER_233_1765 ();
 b15zdnd11an1n64x5 FILLER_233_1829 ();
 b15zdnd11an1n64x5 FILLER_233_1893 ();
 b15zdnd11an1n64x5 FILLER_233_1957 ();
 b15zdnd11an1n16x5 FILLER_233_2021 ();
 b15zdnd11an1n64x5 FILLER_233_2061 ();
 b15zdnd11an1n08x5 FILLER_233_2125 ();
 b15zdnd11an1n04x5 FILLER_233_2133 ();
 b15zdnd00an1n02x5 FILLER_233_2137 ();
 b15zdnd00an1n01x5 FILLER_233_2139 ();
 b15zdnd11an1n08x5 FILLER_233_2182 ();
 b15zdnd00an1n01x5 FILLER_233_2190 ();
 b15zdnd11an1n04x5 FILLER_233_2233 ();
 b15zdnd11an1n04x5 FILLER_233_2279 ();
 b15zdnd00an1n01x5 FILLER_233_2283 ();
 b15zdnd11an1n64x5 FILLER_234_8 ();
 b15zdnd00an1n02x5 FILLER_234_72 ();
 b15zdnd00an1n01x5 FILLER_234_74 ();
 b15zdnd11an1n64x5 FILLER_234_89 ();
 b15zdnd11an1n16x5 FILLER_234_153 ();
 b15zdnd00an1n01x5 FILLER_234_169 ();
 b15zdnd11an1n64x5 FILLER_234_190 ();
 b15zdnd11an1n64x5 FILLER_234_254 ();
 b15zdnd11an1n64x5 FILLER_234_318 ();
 b15zdnd11an1n64x5 FILLER_234_382 ();
 b15zdnd11an1n64x5 FILLER_234_446 ();
 b15zdnd11an1n64x5 FILLER_234_510 ();
 b15zdnd11an1n64x5 FILLER_234_574 ();
 b15zdnd11an1n16x5 FILLER_234_638 ();
 b15zdnd00an1n01x5 FILLER_234_654 ();
 b15zdnd11an1n08x5 FILLER_234_707 ();
 b15zdnd00an1n02x5 FILLER_234_715 ();
 b15zdnd00an1n01x5 FILLER_234_717 ();
 b15zdnd00an1n02x5 FILLER_234_726 ();
 b15zdnd11an1n64x5 FILLER_234_770 ();
 b15zdnd11an1n64x5 FILLER_234_834 ();
 b15zdnd11an1n32x5 FILLER_234_898 ();
 b15zdnd00an1n02x5 FILLER_234_930 ();
 b15zdnd11an1n64x5 FILLER_234_941 ();
 b15zdnd11an1n64x5 FILLER_234_1005 ();
 b15zdnd11an1n64x5 FILLER_234_1069 ();
 b15zdnd11an1n04x5 FILLER_234_1133 ();
 b15zdnd00an1n02x5 FILLER_234_1137 ();
 b15zdnd11an1n64x5 FILLER_234_1148 ();
 b15zdnd11an1n64x5 FILLER_234_1212 ();
 b15zdnd11an1n32x5 FILLER_234_1276 ();
 b15zdnd11an1n08x5 FILLER_234_1308 ();
 b15zdnd11an1n04x5 FILLER_234_1316 ();
 b15zdnd00an1n01x5 FILLER_234_1320 ();
 b15zdnd11an1n16x5 FILLER_234_1338 ();
 b15zdnd11an1n04x5 FILLER_234_1354 ();
 b15zdnd00an1n02x5 FILLER_234_1358 ();
 b15zdnd11an1n16x5 FILLER_234_1377 ();
 b15zdnd11an1n04x5 FILLER_234_1393 ();
 b15zdnd00an1n01x5 FILLER_234_1397 ();
 b15zdnd11an1n08x5 FILLER_234_1415 ();
 b15zdnd00an1n02x5 FILLER_234_1423 ();
 b15zdnd11an1n64x5 FILLER_234_1445 ();
 b15zdnd11an1n64x5 FILLER_234_1509 ();
 b15zdnd11an1n64x5 FILLER_234_1573 ();
 b15zdnd11an1n64x5 FILLER_234_1637 ();
 b15zdnd11an1n64x5 FILLER_234_1701 ();
 b15zdnd11an1n64x5 FILLER_234_1765 ();
 b15zdnd11an1n64x5 FILLER_234_1829 ();
 b15zdnd11an1n64x5 FILLER_234_1893 ();
 b15zdnd11an1n64x5 FILLER_234_1957 ();
 b15zdnd11an1n32x5 FILLER_234_2021 ();
 b15zdnd11an1n08x5 FILLER_234_2053 ();
 b15zdnd00an1n02x5 FILLER_234_2061 ();
 b15zdnd00an1n01x5 FILLER_234_2063 ();
 b15zdnd11an1n64x5 FILLER_234_2067 ();
 b15zdnd11an1n16x5 FILLER_234_2131 ();
 b15zdnd11an1n04x5 FILLER_234_2147 ();
 b15zdnd00an1n02x5 FILLER_234_2151 ();
 b15zdnd00an1n01x5 FILLER_234_2153 ();
 b15zdnd11an1n16x5 FILLER_234_2162 ();
 b15zdnd11an1n08x5 FILLER_234_2178 ();
 b15zdnd11an1n04x5 FILLER_234_2228 ();
 b15zdnd00an1n02x5 FILLER_234_2274 ();
 b15zdnd11an1n32x5 FILLER_235_0 ();
 b15zdnd11an1n16x5 FILLER_235_32 ();
 b15zdnd00an1n02x5 FILLER_235_48 ();
 b15zdnd00an1n01x5 FILLER_235_50 ();
 b15zdnd11an1n64x5 FILLER_235_93 ();
 b15zdnd11an1n64x5 FILLER_235_157 ();
 b15zdnd11an1n64x5 FILLER_235_221 ();
 b15zdnd11an1n64x5 FILLER_235_285 ();
 b15zdnd11an1n32x5 FILLER_235_349 ();
 b15zdnd11an1n16x5 FILLER_235_381 ();
 b15zdnd11an1n08x5 FILLER_235_397 ();
 b15zdnd11an1n04x5 FILLER_235_405 ();
 b15zdnd00an1n02x5 FILLER_235_409 ();
 b15zdnd11an1n64x5 FILLER_235_426 ();
 b15zdnd11an1n64x5 FILLER_235_490 ();
 b15zdnd11an1n64x5 FILLER_235_554 ();
 b15zdnd11an1n32x5 FILLER_235_618 ();
 b15zdnd11an1n08x5 FILLER_235_650 ();
 b15zdnd11an1n04x5 FILLER_235_658 ();
 b15zdnd00an1n02x5 FILLER_235_662 ();
 b15zdnd11an1n04x5 FILLER_235_706 ();
 b15zdnd11an1n64x5 FILLER_235_762 ();
 b15zdnd11an1n64x5 FILLER_235_826 ();
 b15zdnd11an1n32x5 FILLER_235_890 ();
 b15zdnd11an1n08x5 FILLER_235_922 ();
 b15zdnd11an1n04x5 FILLER_235_944 ();
 b15zdnd11an1n64x5 FILLER_235_951 ();
 b15zdnd11an1n64x5 FILLER_235_1015 ();
 b15zdnd11an1n32x5 FILLER_235_1079 ();
 b15zdnd11an1n16x5 FILLER_235_1111 ();
 b15zdnd11an1n64x5 FILLER_235_1136 ();
 b15zdnd11an1n64x5 FILLER_235_1200 ();
 b15zdnd11an1n16x5 FILLER_235_1264 ();
 b15zdnd11an1n08x5 FILLER_235_1280 ();
 b15zdnd00an1n02x5 FILLER_235_1288 ();
 b15zdnd00an1n01x5 FILLER_235_1290 ();
 b15zdnd11an1n64x5 FILLER_235_1308 ();
 b15zdnd11an1n32x5 FILLER_235_1372 ();
 b15zdnd11an1n16x5 FILLER_235_1404 ();
 b15zdnd11an1n64x5 FILLER_235_1432 ();
 b15zdnd11an1n64x5 FILLER_235_1496 ();
 b15zdnd11an1n64x5 FILLER_235_1560 ();
 b15zdnd11an1n64x5 FILLER_235_1624 ();
 b15zdnd11an1n64x5 FILLER_235_1688 ();
 b15zdnd11an1n64x5 FILLER_235_1752 ();
 b15zdnd11an1n64x5 FILLER_235_1816 ();
 b15zdnd11an1n64x5 FILLER_235_1880 ();
 b15zdnd11an1n64x5 FILLER_235_1944 ();
 b15zdnd11an1n32x5 FILLER_235_2008 ();
 b15zdnd00an1n02x5 FILLER_235_2040 ();
 b15zdnd00an1n01x5 FILLER_235_2042 ();
 b15zdnd11an1n64x5 FILLER_235_2085 ();
 b15zdnd11an1n32x5 FILLER_235_2149 ();
 b15zdnd11an1n08x5 FILLER_235_2181 ();
 b15zdnd11an1n04x5 FILLER_235_2189 ();
 b15zdnd00an1n01x5 FILLER_235_2193 ();
 b15zdnd11an1n04x5 FILLER_235_2236 ();
 b15zdnd00an1n02x5 FILLER_235_2282 ();
 b15zdnd11an1n64x5 FILLER_236_8 ();
 b15zdnd11an1n16x5 FILLER_236_72 ();
 b15zdnd00an1n02x5 FILLER_236_88 ();
 b15zdnd11an1n16x5 FILLER_236_132 ();
 b15zdnd11an1n64x5 FILLER_236_190 ();
 b15zdnd11an1n64x5 FILLER_236_254 ();
 b15zdnd11an1n64x5 FILLER_236_318 ();
 b15zdnd11an1n64x5 FILLER_236_382 ();
 b15zdnd11an1n08x5 FILLER_236_446 ();
 b15zdnd11an1n04x5 FILLER_236_454 ();
 b15zdnd00an1n02x5 FILLER_236_458 ();
 b15zdnd00an1n01x5 FILLER_236_460 ();
 b15zdnd11an1n64x5 FILLER_236_465 ();
 b15zdnd11an1n64x5 FILLER_236_529 ();
 b15zdnd11an1n64x5 FILLER_236_593 ();
 b15zdnd11an1n16x5 FILLER_236_657 ();
 b15zdnd11an1n04x5 FILLER_236_676 ();
 b15zdnd11an1n32x5 FILLER_236_683 ();
 b15zdnd00an1n02x5 FILLER_236_715 ();
 b15zdnd00an1n01x5 FILLER_236_717 ();
 b15zdnd11an1n04x5 FILLER_236_726 ();
 b15zdnd11an1n04x5 FILLER_236_733 ();
 b15zdnd11an1n08x5 FILLER_236_740 ();
 b15zdnd00an1n02x5 FILLER_236_748 ();
 b15zdnd11an1n64x5 FILLER_236_792 ();
 b15zdnd11an1n64x5 FILLER_236_856 ();
 b15zdnd11an1n04x5 FILLER_236_920 ();
 b15zdnd00an1n01x5 FILLER_236_924 ();
 b15zdnd11an1n64x5 FILLER_236_977 ();
 b15zdnd11an1n32x5 FILLER_236_1041 ();
 b15zdnd11an1n08x5 FILLER_236_1073 ();
 b15zdnd00an1n02x5 FILLER_236_1081 ();
 b15zdnd00an1n01x5 FILLER_236_1083 ();
 b15zdnd11an1n64x5 FILLER_236_1108 ();
 b15zdnd11an1n64x5 FILLER_236_1172 ();
 b15zdnd11an1n64x5 FILLER_236_1236 ();
 b15zdnd11an1n64x5 FILLER_236_1300 ();
 b15zdnd11an1n64x5 FILLER_236_1364 ();
 b15zdnd11an1n64x5 FILLER_236_1428 ();
 b15zdnd11an1n64x5 FILLER_236_1492 ();
 b15zdnd11an1n64x5 FILLER_236_1556 ();
 b15zdnd11an1n64x5 FILLER_236_1620 ();
 b15zdnd11an1n64x5 FILLER_236_1684 ();
 b15zdnd11an1n64x5 FILLER_236_1748 ();
 b15zdnd11an1n64x5 FILLER_236_1812 ();
 b15zdnd11an1n64x5 FILLER_236_1876 ();
 b15zdnd11an1n64x5 FILLER_236_1940 ();
 b15zdnd11an1n32x5 FILLER_236_2004 ();
 b15zdnd11an1n16x5 FILLER_236_2036 ();
 b15zdnd11an1n08x5 FILLER_236_2052 ();
 b15zdnd11an1n04x5 FILLER_236_2060 ();
 b15zdnd00an1n01x5 FILLER_236_2064 ();
 b15zdnd11an1n16x5 FILLER_236_2068 ();
 b15zdnd11an1n08x5 FILLER_236_2084 ();
 b15zdnd11an1n16x5 FILLER_236_2134 ();
 b15zdnd11an1n04x5 FILLER_236_2150 ();
 b15zdnd11an1n16x5 FILLER_236_2162 ();
 b15zdnd11an1n08x5 FILLER_236_2178 ();
 b15zdnd11an1n04x5 FILLER_236_2228 ();
 b15zdnd00an1n02x5 FILLER_236_2274 ();
 b15zdnd11an1n64x5 FILLER_237_0 ();
 b15zdnd11an1n64x5 FILLER_237_64 ();
 b15zdnd11an1n32x5 FILLER_237_128 ();
 b15zdnd11an1n08x5 FILLER_237_160 ();
 b15zdnd00an1n01x5 FILLER_237_168 ();
 b15zdnd11an1n64x5 FILLER_237_211 ();
 b15zdnd11an1n64x5 FILLER_237_275 ();
 b15zdnd00an1n01x5 FILLER_237_339 ();
 b15zdnd11an1n64x5 FILLER_237_356 ();
 b15zdnd11an1n64x5 FILLER_237_420 ();
 b15zdnd11an1n64x5 FILLER_237_484 ();
 b15zdnd11an1n64x5 FILLER_237_548 ();
 b15zdnd11an1n64x5 FILLER_237_612 ();
 b15zdnd11an1n32x5 FILLER_237_676 ();
 b15zdnd11an1n16x5 FILLER_237_708 ();
 b15zdnd11an1n08x5 FILLER_237_724 ();
 b15zdnd00an1n02x5 FILLER_237_732 ();
 b15zdnd00an1n01x5 FILLER_237_734 ();
 b15zdnd11an1n64x5 FILLER_237_738 ();
 b15zdnd11an1n64x5 FILLER_237_802 ();
 b15zdnd11an1n64x5 FILLER_237_866 ();
 b15zdnd11an1n08x5 FILLER_237_930 ();
 b15zdnd11an1n04x5 FILLER_237_938 ();
 b15zdnd00an1n02x5 FILLER_237_942 ();
 b15zdnd00an1n01x5 FILLER_237_944 ();
 b15zdnd11an1n04x5 FILLER_237_948 ();
 b15zdnd11an1n64x5 FILLER_237_955 ();
 b15zdnd11an1n64x5 FILLER_237_1019 ();
 b15zdnd11an1n64x5 FILLER_237_1083 ();
 b15zdnd11an1n64x5 FILLER_237_1147 ();
 b15zdnd11an1n64x5 FILLER_237_1211 ();
 b15zdnd11an1n32x5 FILLER_237_1275 ();
 b15zdnd00an1n02x5 FILLER_237_1307 ();
 b15zdnd00an1n01x5 FILLER_237_1309 ();
 b15zdnd11an1n64x5 FILLER_237_1327 ();
 b15zdnd11an1n16x5 FILLER_237_1391 ();
 b15zdnd00an1n02x5 FILLER_237_1407 ();
 b15zdnd00an1n01x5 FILLER_237_1409 ();
 b15zdnd11an1n64x5 FILLER_237_1422 ();
 b15zdnd11an1n64x5 FILLER_237_1486 ();
 b15zdnd11an1n64x5 FILLER_237_1550 ();
 b15zdnd11an1n64x5 FILLER_237_1614 ();
 b15zdnd11an1n64x5 FILLER_237_1678 ();
 b15zdnd11an1n64x5 FILLER_237_1742 ();
 b15zdnd11an1n64x5 FILLER_237_1806 ();
 b15zdnd11an1n64x5 FILLER_237_1870 ();
 b15zdnd11an1n64x5 FILLER_237_1934 ();
 b15zdnd11an1n32x5 FILLER_237_1998 ();
 b15zdnd11an1n08x5 FILLER_237_2030 ();
 b15zdnd00an1n02x5 FILLER_237_2038 ();
 b15zdnd11an1n64x5 FILLER_237_2092 ();
 b15zdnd11an1n32x5 FILLER_237_2156 ();
 b15zdnd11an1n08x5 FILLER_237_2188 ();
 b15zdnd00an1n02x5 FILLER_237_2196 ();
 b15zdnd11an1n04x5 FILLER_237_2202 ();
 b15zdnd11an1n04x5 FILLER_237_2248 ();
 b15zdnd11an1n04x5 FILLER_237_2256 ();
 b15zdnd11an1n04x5 FILLER_237_2264 ();
 b15zdnd11an1n04x5 FILLER_237_2272 ();
 b15zdnd00an1n02x5 FILLER_237_2276 ();
 b15zdnd00an1n02x5 FILLER_237_2282 ();
 b15zdnd11an1n64x5 FILLER_238_8 ();
 b15zdnd11an1n64x5 FILLER_238_72 ();
 b15zdnd11an1n64x5 FILLER_238_136 ();
 b15zdnd11an1n08x5 FILLER_238_200 ();
 b15zdnd00an1n02x5 FILLER_238_208 ();
 b15zdnd11an1n04x5 FILLER_238_252 ();
 b15zdnd11an1n64x5 FILLER_238_259 ();
 b15zdnd11an1n64x5 FILLER_238_323 ();
 b15zdnd11an1n32x5 FILLER_238_387 ();
 b15zdnd11an1n16x5 FILLER_238_419 ();
 b15zdnd11an1n08x5 FILLER_238_435 ();
 b15zdnd11an1n04x5 FILLER_238_447 ();
 b15zdnd11an1n32x5 FILLER_238_458 ();
 b15zdnd11an1n16x5 FILLER_238_490 ();
 b15zdnd11an1n04x5 FILLER_238_506 ();
 b15zdnd00an1n01x5 FILLER_238_510 ();
 b15zdnd11an1n32x5 FILLER_238_532 ();
 b15zdnd11an1n16x5 FILLER_238_564 ();
 b15zdnd11an1n08x5 FILLER_238_580 ();
 b15zdnd00an1n02x5 FILLER_238_588 ();
 b15zdnd11an1n32x5 FILLER_238_593 ();
 b15zdnd11an1n04x5 FILLER_238_625 ();
 b15zdnd11an1n04x5 FILLER_238_661 ();
 b15zdnd11an1n32x5 FILLER_238_668 ();
 b15zdnd11an1n16x5 FILLER_238_700 ();
 b15zdnd00an1n02x5 FILLER_238_716 ();
 b15zdnd11an1n64x5 FILLER_238_726 ();
 b15zdnd11an1n64x5 FILLER_238_790 ();
 b15zdnd11an1n64x5 FILLER_238_854 ();
 b15zdnd11an1n64x5 FILLER_238_918 ();
 b15zdnd11an1n64x5 FILLER_238_982 ();
 b15zdnd11an1n64x5 FILLER_238_1046 ();
 b15zdnd11an1n64x5 FILLER_238_1110 ();
 b15zdnd11an1n16x5 FILLER_238_1174 ();
 b15zdnd11an1n04x5 FILLER_238_1190 ();
 b15zdnd11an1n04x5 FILLER_238_1197 ();
 b15zdnd11an1n64x5 FILLER_238_1204 ();
 b15zdnd11an1n64x5 FILLER_238_1268 ();
 b15zdnd11an1n64x5 FILLER_238_1332 ();
 b15zdnd11an1n04x5 FILLER_238_1396 ();
 b15zdnd00an1n01x5 FILLER_238_1400 ();
 b15zdnd11an1n16x5 FILLER_238_1415 ();
 b15zdnd11an1n64x5 FILLER_238_1448 ();
 b15zdnd11an1n08x5 FILLER_238_1512 ();
 b15zdnd00an1n01x5 FILLER_238_1520 ();
 b15zdnd11an1n04x5 FILLER_238_1524 ();
 b15zdnd11an1n64x5 FILLER_238_1531 ();
 b15zdnd11an1n64x5 FILLER_238_1595 ();
 b15zdnd11an1n64x5 FILLER_238_1659 ();
 b15zdnd11an1n64x5 FILLER_238_1723 ();
 b15zdnd11an1n64x5 FILLER_238_1787 ();
 b15zdnd11an1n64x5 FILLER_238_1851 ();
 b15zdnd11an1n64x5 FILLER_238_1915 ();
 b15zdnd11an1n64x5 FILLER_238_1979 ();
 b15zdnd11an1n16x5 FILLER_238_2043 ();
 b15zdnd11an1n04x5 FILLER_238_2059 ();
 b15zdnd00an1n02x5 FILLER_238_2063 ();
 b15zdnd11an1n64x5 FILLER_238_2068 ();
 b15zdnd11an1n16x5 FILLER_238_2132 ();
 b15zdnd11an1n04x5 FILLER_238_2148 ();
 b15zdnd00an1n02x5 FILLER_238_2152 ();
 b15zdnd11an1n16x5 FILLER_238_2162 ();
 b15zdnd11an1n04x5 FILLER_238_2178 ();
 b15zdnd00an1n02x5 FILLER_238_2182 ();
 b15zdnd00an1n01x5 FILLER_238_2184 ();
 b15zdnd11an1n04x5 FILLER_238_2237 ();
 b15zdnd11an1n04x5 FILLER_238_2248 ();
 b15zdnd00an1n02x5 FILLER_238_2252 ();
 b15zdnd11an1n04x5 FILLER_238_2258 ();
 b15zdnd11an1n04x5 FILLER_238_2266 ();
 b15zdnd00an1n02x5 FILLER_238_2274 ();
 b15zdnd11an1n64x5 FILLER_239_0 ();
 b15zdnd11an1n64x5 FILLER_239_64 ();
 b15zdnd11an1n32x5 FILLER_239_128 ();
 b15zdnd11an1n16x5 FILLER_239_160 ();
 b15zdnd11an1n04x5 FILLER_239_176 ();
 b15zdnd00an1n02x5 FILLER_239_180 ();
 b15zdnd00an1n01x5 FILLER_239_182 ();
 b15zdnd11an1n08x5 FILLER_239_191 ();
 b15zdnd00an1n01x5 FILLER_239_199 ();
 b15zdnd11an1n16x5 FILLER_239_220 ();
 b15zdnd11an1n64x5 FILLER_239_288 ();
 b15zdnd11an1n64x5 FILLER_239_352 ();
 b15zdnd11an1n32x5 FILLER_239_416 ();
 b15zdnd11an1n04x5 FILLER_239_448 ();
 b15zdnd11an1n32x5 FILLER_239_468 ();
 b15zdnd11an1n16x5 FILLER_239_500 ();
 b15zdnd11an1n08x5 FILLER_239_516 ();
 b15zdnd00an1n02x5 FILLER_239_524 ();
 b15zdnd11an1n32x5 FILLER_239_530 ();
 b15zdnd11an1n04x5 FILLER_239_562 ();
 b15zdnd00an1n02x5 FILLER_239_566 ();
 b15zdnd11an1n08x5 FILLER_239_600 ();
 b15zdnd11an1n04x5 FILLER_239_608 ();
 b15zdnd11an1n08x5 FILLER_239_654 ();
 b15zdnd00an1n02x5 FILLER_239_662 ();
 b15zdnd00an1n01x5 FILLER_239_664 ();
 b15zdnd11an1n64x5 FILLER_239_668 ();
 b15zdnd11an1n64x5 FILLER_239_732 ();
 b15zdnd11an1n16x5 FILLER_239_796 ();
 b15zdnd11an1n08x5 FILLER_239_812 ();
 b15zdnd00an1n01x5 FILLER_239_820 ();
 b15zdnd11an1n04x5 FILLER_239_832 ();
 b15zdnd11an1n64x5 FILLER_239_846 ();
 b15zdnd11an1n08x5 FILLER_239_910 ();
 b15zdnd11an1n04x5 FILLER_239_918 ();
 b15zdnd00an1n01x5 FILLER_239_922 ();
 b15zdnd11an1n04x5 FILLER_239_932 ();
 b15zdnd11an1n16x5 FILLER_239_939 ();
 b15zdnd11an1n04x5 FILLER_239_955 ();
 b15zdnd00an1n01x5 FILLER_239_959 ();
 b15zdnd11an1n64x5 FILLER_239_969 ();
 b15zdnd11an1n64x5 FILLER_239_1033 ();
 b15zdnd11an1n64x5 FILLER_239_1097 ();
 b15zdnd11an1n08x5 FILLER_239_1161 ();
 b15zdnd11an1n04x5 FILLER_239_1169 ();
 b15zdnd00an1n02x5 FILLER_239_1173 ();
 b15zdnd00an1n01x5 FILLER_239_1175 ();
 b15zdnd11an1n64x5 FILLER_239_1228 ();
 b15zdnd11an1n32x5 FILLER_239_1292 ();
 b15zdnd00an1n02x5 FILLER_239_1324 ();
 b15zdnd11an1n64x5 FILLER_239_1346 ();
 b15zdnd11an1n64x5 FILLER_239_1410 ();
 b15zdnd11an1n16x5 FILLER_239_1474 ();
 b15zdnd11an1n08x5 FILLER_239_1490 ();
 b15zdnd11an1n04x5 FILLER_239_1498 ();
 b15zdnd00an1n01x5 FILLER_239_1502 ();
 b15zdnd11an1n64x5 FILLER_239_1555 ();
 b15zdnd11an1n64x5 FILLER_239_1619 ();
 b15zdnd11an1n64x5 FILLER_239_1683 ();
 b15zdnd11an1n64x5 FILLER_239_1747 ();
 b15zdnd11an1n64x5 FILLER_239_1811 ();
 b15zdnd11an1n64x5 FILLER_239_1875 ();
 b15zdnd11an1n64x5 FILLER_239_1939 ();
 b15zdnd11an1n08x5 FILLER_239_2003 ();
 b15zdnd11an1n04x5 FILLER_239_2011 ();
 b15zdnd11an1n16x5 FILLER_239_2025 ();
 b15zdnd00an1n02x5 FILLER_239_2041 ();
 b15zdnd00an1n01x5 FILLER_239_2043 ();
 b15zdnd11an1n64x5 FILLER_239_2075 ();
 b15zdnd11an1n32x5 FILLER_239_2139 ();
 b15zdnd11an1n16x5 FILLER_239_2171 ();
 b15zdnd11an1n04x5 FILLER_239_2187 ();
 b15zdnd00an1n02x5 FILLER_239_2191 ();
 b15zdnd11an1n04x5 FILLER_239_2196 ();
 b15zdnd11an1n16x5 FILLER_239_2242 ();
 b15zdnd11an1n04x5 FILLER_239_2258 ();
 b15zdnd11an1n16x5 FILLER_239_2266 ();
 b15zdnd00an1n02x5 FILLER_239_2282 ();
 b15zdnd11an1n32x5 FILLER_240_8 ();
 b15zdnd11an1n08x5 FILLER_240_40 ();
 b15zdnd00an1n01x5 FILLER_240_48 ();
 b15zdnd11an1n04x5 FILLER_240_52 ();
 b15zdnd11an1n64x5 FILLER_240_59 ();
 b15zdnd11an1n32x5 FILLER_240_123 ();
 b15zdnd11an1n16x5 FILLER_240_155 ();
 b15zdnd11an1n04x5 FILLER_240_171 ();
 b15zdnd00an1n02x5 FILLER_240_175 ();
 b15zdnd11an1n08x5 FILLER_240_185 ();
 b15zdnd00an1n02x5 FILLER_240_193 ();
 b15zdnd00an1n01x5 FILLER_240_195 ();
 b15zdnd11an1n32x5 FILLER_240_208 ();
 b15zdnd11an1n16x5 FILLER_240_240 ();
 b15zdnd00an1n01x5 FILLER_240_256 ();
 b15zdnd11an1n64x5 FILLER_240_260 ();
 b15zdnd11an1n64x5 FILLER_240_324 ();
 b15zdnd11an1n08x5 FILLER_240_388 ();
 b15zdnd11an1n04x5 FILLER_240_396 ();
 b15zdnd11an1n32x5 FILLER_240_410 ();
 b15zdnd11an1n08x5 FILLER_240_442 ();
 b15zdnd11an1n04x5 FILLER_240_450 ();
 b15zdnd00an1n02x5 FILLER_240_454 ();
 b15zdnd00an1n01x5 FILLER_240_456 ();
 b15zdnd11an1n04x5 FILLER_240_469 ();
 b15zdnd11an1n08x5 FILLER_240_485 ();
 b15zdnd00an1n02x5 FILLER_240_493 ();
 b15zdnd00an1n01x5 FILLER_240_495 ();
 b15zdnd11an1n08x5 FILLER_240_510 ();
 b15zdnd00an1n01x5 FILLER_240_518 ();
 b15zdnd11an1n64x5 FILLER_240_528 ();
 b15zdnd00an1n02x5 FILLER_240_592 ();
 b15zdnd00an1n01x5 FILLER_240_594 ();
 b15zdnd11an1n64x5 FILLER_240_598 ();
 b15zdnd11an1n32x5 FILLER_240_662 ();
 b15zdnd11an1n16x5 FILLER_240_694 ();
 b15zdnd11an1n08x5 FILLER_240_710 ();
 b15zdnd11an1n64x5 FILLER_240_726 ();
 b15zdnd11an1n08x5 FILLER_240_790 ();
 b15zdnd11an1n04x5 FILLER_240_798 ();
 b15zdnd11an1n04x5 FILLER_240_816 ();
 b15zdnd00an1n01x5 FILLER_240_820 ();
 b15zdnd11an1n64x5 FILLER_240_824 ();
 b15zdnd11an1n16x5 FILLER_240_888 ();
 b15zdnd00an1n02x5 FILLER_240_904 ();
 b15zdnd11an1n04x5 FILLER_240_958 ();
 b15zdnd11an1n64x5 FILLER_240_971 ();
 b15zdnd11an1n16x5 FILLER_240_1035 ();
 b15zdnd11an1n08x5 FILLER_240_1051 ();
 b15zdnd11an1n04x5 FILLER_240_1059 ();
 b15zdnd00an1n01x5 FILLER_240_1063 ();
 b15zdnd11an1n64x5 FILLER_240_1091 ();
 b15zdnd11an1n32x5 FILLER_240_1155 ();
 b15zdnd11an1n08x5 FILLER_240_1187 ();
 b15zdnd11an1n04x5 FILLER_240_1195 ();
 b15zdnd00an1n02x5 FILLER_240_1199 ();
 b15zdnd00an1n01x5 FILLER_240_1201 ();
 b15zdnd11an1n64x5 FILLER_240_1205 ();
 b15zdnd11an1n64x5 FILLER_240_1269 ();
 b15zdnd11an1n64x5 FILLER_240_1333 ();
 b15zdnd11an1n64x5 FILLER_240_1397 ();
 b15zdnd11an1n32x5 FILLER_240_1461 ();
 b15zdnd11an1n16x5 FILLER_240_1493 ();
 b15zdnd00an1n02x5 FILLER_240_1509 ();
 b15zdnd00an1n01x5 FILLER_240_1511 ();
 b15zdnd11an1n32x5 FILLER_240_1564 ();
 b15zdnd11an1n16x5 FILLER_240_1596 ();
 b15zdnd11an1n08x5 FILLER_240_1612 ();
 b15zdnd11an1n04x5 FILLER_240_1620 ();
 b15zdnd00an1n02x5 FILLER_240_1624 ();
 b15zdnd11an1n08x5 FILLER_240_1629 ();
 b15zdnd11an1n64x5 FILLER_240_1640 ();
 b15zdnd11an1n64x5 FILLER_240_1704 ();
 b15zdnd11an1n64x5 FILLER_240_1768 ();
 b15zdnd11an1n64x5 FILLER_240_1832 ();
 b15zdnd11an1n64x5 FILLER_240_1896 ();
 b15zdnd11an1n64x5 FILLER_240_1960 ();
 b15zdnd11an1n64x5 FILLER_240_2024 ();
 b15zdnd11an1n64x5 FILLER_240_2088 ();
 b15zdnd00an1n02x5 FILLER_240_2152 ();
 b15zdnd11an1n32x5 FILLER_240_2162 ();
 b15zdnd11an1n08x5 FILLER_240_2194 ();
 b15zdnd11an1n04x5 FILLER_240_2226 ();
 b15zdnd00an1n02x5 FILLER_240_2230 ();
 b15zdnd00an1n02x5 FILLER_240_2274 ();
 b15zdnd11an1n16x5 FILLER_241_0 ();
 b15zdnd11an1n08x5 FILLER_241_16 ();
 b15zdnd00an1n02x5 FILLER_241_24 ();
 b15zdnd11an1n64x5 FILLER_241_78 ();
 b15zdnd11an1n64x5 FILLER_241_142 ();
 b15zdnd11an1n32x5 FILLER_241_206 ();
 b15zdnd11an1n16x5 FILLER_241_238 ();
 b15zdnd11an1n04x5 FILLER_241_254 ();
 b15zdnd00an1n02x5 FILLER_241_258 ();
 b15zdnd00an1n01x5 FILLER_241_260 ();
 b15zdnd11an1n64x5 FILLER_241_264 ();
 b15zdnd11an1n32x5 FILLER_241_328 ();
 b15zdnd11an1n08x5 FILLER_241_360 ();
 b15zdnd00an1n01x5 FILLER_241_368 ();
 b15zdnd11an1n64x5 FILLER_241_377 ();
 b15zdnd11an1n16x5 FILLER_241_441 ();
 b15zdnd11an1n08x5 FILLER_241_457 ();
 b15zdnd00an1n01x5 FILLER_241_465 ();
 b15zdnd11an1n64x5 FILLER_241_469 ();
 b15zdnd11an1n64x5 FILLER_241_533 ();
 b15zdnd11an1n64x5 FILLER_241_597 ();
 b15zdnd11an1n64x5 FILLER_241_661 ();
 b15zdnd11an1n04x5 FILLER_241_725 ();
 b15zdnd00an1n01x5 FILLER_241_729 ();
 b15zdnd11an1n32x5 FILLER_241_744 ();
 b15zdnd11an1n04x5 FILLER_241_794 ();
 b15zdnd11an1n64x5 FILLER_241_850 ();
 b15zdnd11an1n08x5 FILLER_241_914 ();
 b15zdnd11an1n04x5 FILLER_241_922 ();
 b15zdnd00an1n02x5 FILLER_241_926 ();
 b15zdnd00an1n01x5 FILLER_241_928 ();
 b15zdnd11an1n04x5 FILLER_241_932 ();
 b15zdnd11an1n64x5 FILLER_241_939 ();
 b15zdnd11an1n32x5 FILLER_241_1003 ();
 b15zdnd11an1n16x5 FILLER_241_1035 ();
 b15zdnd11an1n08x5 FILLER_241_1051 ();
 b15zdnd11an1n04x5 FILLER_241_1059 ();
 b15zdnd00an1n02x5 FILLER_241_1063 ();
 b15zdnd11an1n08x5 FILLER_241_1068 ();
 b15zdnd11an1n04x5 FILLER_241_1076 ();
 b15zdnd00an1n02x5 FILLER_241_1080 ();
 b15zdnd00an1n01x5 FILLER_241_1082 ();
 b15zdnd11an1n64x5 FILLER_241_1086 ();
 b15zdnd11an1n64x5 FILLER_241_1150 ();
 b15zdnd11an1n64x5 FILLER_241_1214 ();
 b15zdnd11an1n32x5 FILLER_241_1278 ();
 b15zdnd11an1n04x5 FILLER_241_1310 ();
 b15zdnd00an1n02x5 FILLER_241_1314 ();
 b15zdnd11an1n64x5 FILLER_241_1336 ();
 b15zdnd11an1n64x5 FILLER_241_1400 ();
 b15zdnd11an1n64x5 FILLER_241_1464 ();
 b15zdnd11an1n04x5 FILLER_241_1531 ();
 b15zdnd11an1n04x5 FILLER_241_1538 ();
 b15zdnd00an1n02x5 FILLER_241_1542 ();
 b15zdnd11an1n32x5 FILLER_241_1547 ();
 b15zdnd11an1n16x5 FILLER_241_1579 ();
 b15zdnd11an1n08x5 FILLER_241_1595 ();
 b15zdnd11an1n64x5 FILLER_241_1655 ();
 b15zdnd11an1n32x5 FILLER_241_1719 ();
 b15zdnd11an1n08x5 FILLER_241_1751 ();
 b15zdnd11an1n04x5 FILLER_241_1759 ();
 b15zdnd00an1n02x5 FILLER_241_1763 ();
 b15zdnd00an1n01x5 FILLER_241_1765 ();
 b15zdnd11an1n64x5 FILLER_241_1769 ();
 b15zdnd11an1n64x5 FILLER_241_1833 ();
 b15zdnd11an1n32x5 FILLER_241_1897 ();
 b15zdnd11an1n04x5 FILLER_241_1929 ();
 b15zdnd00an1n02x5 FILLER_241_1933 ();
 b15zdnd11an1n64x5 FILLER_241_1944 ();
 b15zdnd11an1n64x5 FILLER_241_2008 ();
 b15zdnd11an1n64x5 FILLER_241_2072 ();
 b15zdnd11an1n64x5 FILLER_241_2136 ();
 b15zdnd11an1n08x5 FILLER_241_2200 ();
 b15zdnd00an1n02x5 FILLER_241_2208 ();
 b15zdnd11an1n04x5 FILLER_241_2213 ();
 b15zdnd11an1n16x5 FILLER_241_2220 ();
 b15zdnd11an1n04x5 FILLER_241_2236 ();
 b15zdnd00an1n02x5 FILLER_241_2282 ();
 b15zdnd11an1n32x5 FILLER_242_8 ();
 b15zdnd11an1n04x5 FILLER_242_40 ();
 b15zdnd00an1n02x5 FILLER_242_44 ();
 b15zdnd11an1n04x5 FILLER_242_49 ();
 b15zdnd11an1n64x5 FILLER_242_56 ();
 b15zdnd11an1n64x5 FILLER_242_120 ();
 b15zdnd11an1n04x5 FILLER_242_184 ();
 b15zdnd00an1n01x5 FILLER_242_188 ();
 b15zdnd11an1n32x5 FILLER_242_231 ();
 b15zdnd00an1n02x5 FILLER_242_263 ();
 b15zdnd00an1n01x5 FILLER_242_265 ();
 b15zdnd11an1n32x5 FILLER_242_308 ();
 b15zdnd11an1n08x5 FILLER_242_340 ();
 b15zdnd11an1n04x5 FILLER_242_348 ();
 b15zdnd00an1n01x5 FILLER_242_352 ();
 b15zdnd11an1n04x5 FILLER_242_357 ();
 b15zdnd00an1n02x5 FILLER_242_361 ();
 b15zdnd00an1n01x5 FILLER_242_363 ();
 b15zdnd11an1n04x5 FILLER_242_384 ();
 b15zdnd11an1n64x5 FILLER_242_392 ();
 b15zdnd11an1n64x5 FILLER_242_456 ();
 b15zdnd11an1n64x5 FILLER_242_520 ();
 b15zdnd11an1n64x5 FILLER_242_584 ();
 b15zdnd11an1n64x5 FILLER_242_648 ();
 b15zdnd11an1n04x5 FILLER_242_712 ();
 b15zdnd00an1n02x5 FILLER_242_716 ();
 b15zdnd11an1n32x5 FILLER_242_726 ();
 b15zdnd11an1n16x5 FILLER_242_758 ();
 b15zdnd00an1n02x5 FILLER_242_774 ();
 b15zdnd00an1n01x5 FILLER_242_776 ();
 b15zdnd11an1n32x5 FILLER_242_785 ();
 b15zdnd11an1n04x5 FILLER_242_817 ();
 b15zdnd11an1n04x5 FILLER_242_824 ();
 b15zdnd11an1n04x5 FILLER_242_831 ();
 b15zdnd00an1n02x5 FILLER_242_835 ();
 b15zdnd00an1n01x5 FILLER_242_837 ();
 b15zdnd11an1n64x5 FILLER_242_880 ();
 b15zdnd11an1n64x5 FILLER_242_944 ();
 b15zdnd11an1n32x5 FILLER_242_1008 ();
 b15zdnd11an1n16x5 FILLER_242_1040 ();
 b15zdnd00an1n02x5 FILLER_242_1056 ();
 b15zdnd11an1n08x5 FILLER_242_1110 ();
 b15zdnd00an1n01x5 FILLER_242_1118 ();
 b15zdnd11an1n64x5 FILLER_242_1130 ();
 b15zdnd11an1n64x5 FILLER_242_1194 ();
 b15zdnd11an1n64x5 FILLER_242_1258 ();
 b15zdnd11an1n64x5 FILLER_242_1322 ();
 b15zdnd11an1n64x5 FILLER_242_1386 ();
 b15zdnd11an1n64x5 FILLER_242_1450 ();
 b15zdnd11an1n16x5 FILLER_242_1514 ();
 b15zdnd00an1n02x5 FILLER_242_1530 ();
 b15zdnd11an1n64x5 FILLER_242_1535 ();
 b15zdnd11an1n16x5 FILLER_242_1599 ();
 b15zdnd11an1n08x5 FILLER_242_1615 ();
 b15zdnd11an1n04x5 FILLER_242_1623 ();
 b15zdnd00an1n01x5 FILLER_242_1627 ();
 b15zdnd11an1n64x5 FILLER_242_1631 ();
 b15zdnd11an1n64x5 FILLER_242_1695 ();
 b15zdnd11an1n04x5 FILLER_242_1759 ();
 b15zdnd00an1n01x5 FILLER_242_1763 ();
 b15zdnd11an1n04x5 FILLER_242_1767 ();
 b15zdnd11an1n64x5 FILLER_242_1774 ();
 b15zdnd11an1n64x5 FILLER_242_1838 ();
 b15zdnd11an1n64x5 FILLER_242_1902 ();
 b15zdnd11an1n32x5 FILLER_242_1966 ();
 b15zdnd11an1n16x5 FILLER_242_1998 ();
 b15zdnd11an1n08x5 FILLER_242_2014 ();
 b15zdnd00an1n02x5 FILLER_242_2022 ();
 b15zdnd00an1n01x5 FILLER_242_2024 ();
 b15zdnd11an1n64x5 FILLER_242_2028 ();
 b15zdnd11an1n32x5 FILLER_242_2092 ();
 b15zdnd11an1n16x5 FILLER_242_2124 ();
 b15zdnd11an1n08x5 FILLER_242_2140 ();
 b15zdnd11an1n04x5 FILLER_242_2148 ();
 b15zdnd00an1n02x5 FILLER_242_2152 ();
 b15zdnd11an1n64x5 FILLER_242_2162 ();
 b15zdnd11an1n04x5 FILLER_242_2226 ();
 b15zdnd00an1n02x5 FILLER_242_2230 ();
 b15zdnd00an1n02x5 FILLER_242_2274 ();
 b15zdnd11an1n32x5 FILLER_243_0 ();
 b15zdnd11an1n16x5 FILLER_243_32 ();
 b15zdnd11an1n04x5 FILLER_243_48 ();
 b15zdnd00an1n02x5 FILLER_243_52 ();
 b15zdnd11an1n64x5 FILLER_243_57 ();
 b15zdnd11an1n64x5 FILLER_243_121 ();
 b15zdnd11an1n04x5 FILLER_243_185 ();
 b15zdnd00an1n01x5 FILLER_243_189 ();
 b15zdnd11an1n08x5 FILLER_243_194 ();
 b15zdnd00an1n01x5 FILLER_243_202 ();
 b15zdnd11an1n64x5 FILLER_243_224 ();
 b15zdnd11an1n04x5 FILLER_243_288 ();
 b15zdnd00an1n02x5 FILLER_243_292 ();
 b15zdnd00an1n01x5 FILLER_243_294 ();
 b15zdnd11an1n16x5 FILLER_243_337 ();
 b15zdnd11an1n08x5 FILLER_243_353 ();
 b15zdnd11an1n04x5 FILLER_243_361 ();
 b15zdnd11an1n64x5 FILLER_243_371 ();
 b15zdnd11an1n64x5 FILLER_243_435 ();
 b15zdnd11an1n64x5 FILLER_243_499 ();
 b15zdnd11an1n64x5 FILLER_243_563 ();
 b15zdnd11an1n64x5 FILLER_243_627 ();
 b15zdnd11an1n64x5 FILLER_243_691 ();
 b15zdnd11an1n16x5 FILLER_243_755 ();
 b15zdnd11an1n08x5 FILLER_243_771 ();
 b15zdnd11an1n04x5 FILLER_243_779 ();
 b15zdnd11an1n32x5 FILLER_243_790 ();
 b15zdnd11an1n08x5 FILLER_243_822 ();
 b15zdnd11an1n04x5 FILLER_243_830 ();
 b15zdnd00an1n02x5 FILLER_243_834 ();
 b15zdnd00an1n01x5 FILLER_243_836 ();
 b15zdnd11an1n64x5 FILLER_243_845 ();
 b15zdnd11an1n64x5 FILLER_243_909 ();
 b15zdnd11an1n64x5 FILLER_243_973 ();
 b15zdnd11an1n32x5 FILLER_243_1037 ();
 b15zdnd11an1n04x5 FILLER_243_1069 ();
 b15zdnd00an1n02x5 FILLER_243_1073 ();
 b15zdnd00an1n01x5 FILLER_243_1075 ();
 b15zdnd11an1n04x5 FILLER_243_1079 ();
 b15zdnd11an1n04x5 FILLER_243_1086 ();
 b15zdnd11an1n32x5 FILLER_243_1142 ();
 b15zdnd11an1n08x5 FILLER_243_1174 ();
 b15zdnd00an1n02x5 FILLER_243_1182 ();
 b15zdnd00an1n01x5 FILLER_243_1184 ();
 b15zdnd11an1n04x5 FILLER_243_1188 ();
 b15zdnd11an1n64x5 FILLER_243_1195 ();
 b15zdnd11an1n64x5 FILLER_243_1259 ();
 b15zdnd11an1n64x5 FILLER_243_1323 ();
 b15zdnd11an1n64x5 FILLER_243_1387 ();
 b15zdnd11an1n64x5 FILLER_243_1451 ();
 b15zdnd11an1n64x5 FILLER_243_1515 ();
 b15zdnd11an1n64x5 FILLER_243_1579 ();
 b15zdnd11an1n08x5 FILLER_243_1643 ();
 b15zdnd00an1n01x5 FILLER_243_1651 ();
 b15zdnd11an1n64x5 FILLER_243_1655 ();
 b15zdnd11an1n16x5 FILLER_243_1719 ();
 b15zdnd11an1n08x5 FILLER_243_1735 ();
 b15zdnd00an1n02x5 FILLER_243_1743 ();
 b15zdnd00an1n01x5 FILLER_243_1745 ();
 b15zdnd11an1n16x5 FILLER_243_1798 ();
 b15zdnd11an1n08x5 FILLER_243_1817 ();
 b15zdnd11an1n04x5 FILLER_243_1825 ();
 b15zdnd11an1n64x5 FILLER_243_1881 ();
 b15zdnd11an1n64x5 FILLER_243_1945 ();
 b15zdnd11an1n64x5 FILLER_243_2009 ();
 b15zdnd11an1n64x5 FILLER_243_2073 ();
 b15zdnd11an1n64x5 FILLER_243_2137 ();
 b15zdnd11an1n32x5 FILLER_243_2201 ();
 b15zdnd11an1n04x5 FILLER_243_2233 ();
 b15zdnd00an1n02x5 FILLER_243_2237 ();
 b15zdnd00an1n01x5 FILLER_243_2239 ();
 b15zdnd00an1n02x5 FILLER_243_2282 ();
 b15zdnd11an1n64x5 FILLER_244_8 ();
 b15zdnd11an1n64x5 FILLER_244_72 ();
 b15zdnd11an1n32x5 FILLER_244_136 ();
 b15zdnd11an1n16x5 FILLER_244_168 ();
 b15zdnd00an1n01x5 FILLER_244_184 ();
 b15zdnd11an1n64x5 FILLER_244_227 ();
 b15zdnd00an1n01x5 FILLER_244_291 ();
 b15zdnd11an1n04x5 FILLER_244_295 ();
 b15zdnd11an1n04x5 FILLER_244_302 ();
 b15zdnd11an1n64x5 FILLER_244_309 ();
 b15zdnd11an1n32x5 FILLER_244_373 ();
 b15zdnd11an1n08x5 FILLER_244_405 ();
 b15zdnd00an1n02x5 FILLER_244_413 ();
 b15zdnd00an1n01x5 FILLER_244_415 ();
 b15zdnd11an1n64x5 FILLER_244_420 ();
 b15zdnd11an1n64x5 FILLER_244_484 ();
 b15zdnd11an1n64x5 FILLER_244_548 ();
 b15zdnd11an1n64x5 FILLER_244_612 ();
 b15zdnd11an1n32x5 FILLER_244_676 ();
 b15zdnd11an1n08x5 FILLER_244_708 ();
 b15zdnd00an1n02x5 FILLER_244_716 ();
 b15zdnd11an1n64x5 FILLER_244_726 ();
 b15zdnd11an1n64x5 FILLER_244_790 ();
 b15zdnd11an1n64x5 FILLER_244_854 ();
 b15zdnd11an1n64x5 FILLER_244_918 ();
 b15zdnd11an1n64x5 FILLER_244_982 ();
 b15zdnd11an1n32x5 FILLER_244_1046 ();
 b15zdnd11an1n16x5 FILLER_244_1078 ();
 b15zdnd11an1n08x5 FILLER_244_1094 ();
 b15zdnd11an1n04x5 FILLER_244_1102 ();
 b15zdnd11an1n04x5 FILLER_244_1109 ();
 b15zdnd00an1n02x5 FILLER_244_1113 ();
 b15zdnd11an1n32x5 FILLER_244_1118 ();
 b15zdnd11an1n16x5 FILLER_244_1150 ();
 b15zdnd00an1n01x5 FILLER_244_1166 ();
 b15zdnd11an1n64x5 FILLER_244_1219 ();
 b15zdnd11an1n64x5 FILLER_244_1283 ();
 b15zdnd11an1n64x5 FILLER_244_1347 ();
 b15zdnd11an1n64x5 FILLER_244_1411 ();
 b15zdnd11an1n64x5 FILLER_244_1475 ();
 b15zdnd11an1n64x5 FILLER_244_1539 ();
 b15zdnd11an1n16x5 FILLER_244_1603 ();
 b15zdnd11an1n08x5 FILLER_244_1619 ();
 b15zdnd11an1n04x5 FILLER_244_1627 ();
 b15zdnd00an1n01x5 FILLER_244_1631 ();
 b15zdnd11an1n64x5 FILLER_244_1684 ();
 b15zdnd00an1n02x5 FILLER_244_1748 ();
 b15zdnd00an1n01x5 FILLER_244_1750 ();
 b15zdnd11an1n08x5 FILLER_244_1803 ();
 b15zdnd11an1n04x5 FILLER_244_1811 ();
 b15zdnd11an1n16x5 FILLER_244_1818 ();
 b15zdnd11an1n08x5 FILLER_244_1834 ();
 b15zdnd11an1n04x5 FILLER_244_1842 ();
 b15zdnd00an1n01x5 FILLER_244_1846 ();
 b15zdnd11an1n04x5 FILLER_244_1850 ();
 b15zdnd11an1n04x5 FILLER_244_1857 ();
 b15zdnd11an1n64x5 FILLER_244_1864 ();
 b15zdnd11an1n64x5 FILLER_244_1928 ();
 b15zdnd11an1n32x5 FILLER_244_1992 ();
 b15zdnd11an1n16x5 FILLER_244_2024 ();
 b15zdnd11an1n04x5 FILLER_244_2040 ();
 b15zdnd00an1n02x5 FILLER_244_2044 ();
 b15zdnd11an1n04x5 FILLER_244_2066 ();
 b15zdnd11an1n32x5 FILLER_244_2087 ();
 b15zdnd11an1n08x5 FILLER_244_2119 ();
 b15zdnd00an1n02x5 FILLER_244_2127 ();
 b15zdnd11an1n16x5 FILLER_244_2133 ();
 b15zdnd11an1n04x5 FILLER_244_2149 ();
 b15zdnd00an1n01x5 FILLER_244_2153 ();
 b15zdnd11an1n64x5 FILLER_244_2162 ();
 b15zdnd11an1n04x5 FILLER_244_2226 ();
 b15zdnd00an1n02x5 FILLER_244_2230 ();
 b15zdnd00an1n02x5 FILLER_244_2274 ();
 b15zdnd11an1n64x5 FILLER_245_0 ();
 b15zdnd00an1n02x5 FILLER_245_64 ();
 b15zdnd00an1n01x5 FILLER_245_66 ();
 b15zdnd11an1n04x5 FILLER_245_70 ();
 b15zdnd11an1n64x5 FILLER_245_77 ();
 b15zdnd11an1n16x5 FILLER_245_141 ();
 b15zdnd11an1n04x5 FILLER_245_157 ();
 b15zdnd00an1n01x5 FILLER_245_161 ();
 b15zdnd11an1n04x5 FILLER_245_165 ();
 b15zdnd11an1n32x5 FILLER_245_172 ();
 b15zdnd11an1n04x5 FILLER_245_204 ();
 b15zdnd00an1n02x5 FILLER_245_208 ();
 b15zdnd11an1n04x5 FILLER_245_226 ();
 b15zdnd11an1n32x5 FILLER_245_237 ();
 b15zdnd11an1n04x5 FILLER_245_269 ();
 b15zdnd11an1n32x5 FILLER_245_325 ();
 b15zdnd00an1n02x5 FILLER_245_357 ();
 b15zdnd00an1n01x5 FILLER_245_359 ();
 b15zdnd11an1n04x5 FILLER_245_368 ();
 b15zdnd00an1n02x5 FILLER_245_372 ();
 b15zdnd00an1n01x5 FILLER_245_374 ();
 b15zdnd11an1n64x5 FILLER_245_383 ();
 b15zdnd11an1n64x5 FILLER_245_447 ();
 b15zdnd11an1n32x5 FILLER_245_511 ();
 b15zdnd11an1n16x5 FILLER_245_543 ();
 b15zdnd11an1n04x5 FILLER_245_559 ();
 b15zdnd11an1n64x5 FILLER_245_572 ();
 b15zdnd11an1n64x5 FILLER_245_636 ();
 b15zdnd11an1n64x5 FILLER_245_700 ();
 b15zdnd11an1n64x5 FILLER_245_764 ();
 b15zdnd11an1n64x5 FILLER_245_828 ();
 b15zdnd11an1n32x5 FILLER_245_892 ();
 b15zdnd11an1n16x5 FILLER_245_924 ();
 b15zdnd11an1n08x5 FILLER_245_940 ();
 b15zdnd11an1n04x5 FILLER_245_948 ();
 b15zdnd00an1n02x5 FILLER_245_952 ();
 b15zdnd00an1n01x5 FILLER_245_954 ();
 b15zdnd11an1n64x5 FILLER_245_1007 ();
 b15zdnd11an1n32x5 FILLER_245_1071 ();
 b15zdnd11an1n08x5 FILLER_245_1103 ();
 b15zdnd00an1n01x5 FILLER_245_1111 ();
 b15zdnd11an1n64x5 FILLER_245_1115 ();
 b15zdnd11an1n04x5 FILLER_245_1179 ();
 b15zdnd00an1n02x5 FILLER_245_1183 ();
 b15zdnd00an1n01x5 FILLER_245_1185 ();
 b15zdnd11an1n04x5 FILLER_245_1189 ();
 b15zdnd11an1n64x5 FILLER_245_1213 ();
 b15zdnd00an1n02x5 FILLER_245_1277 ();
 b15zdnd00an1n01x5 FILLER_245_1279 ();
 b15zdnd11an1n64x5 FILLER_245_1289 ();
 b15zdnd11an1n64x5 FILLER_245_1353 ();
 b15zdnd11an1n64x5 FILLER_245_1417 ();
 b15zdnd11an1n64x5 FILLER_245_1481 ();
 b15zdnd11an1n16x5 FILLER_245_1545 ();
 b15zdnd11an1n08x5 FILLER_245_1561 ();
 b15zdnd00an1n02x5 FILLER_245_1569 ();
 b15zdnd11an1n64x5 FILLER_245_1580 ();
 b15zdnd11an1n08x5 FILLER_245_1644 ();
 b15zdnd11an1n04x5 FILLER_245_1652 ();
 b15zdnd00an1n01x5 FILLER_245_1656 ();
 b15zdnd11an1n64x5 FILLER_245_1660 ();
 b15zdnd11an1n32x5 FILLER_245_1724 ();
 b15zdnd11an1n08x5 FILLER_245_1756 ();
 b15zdnd11an1n04x5 FILLER_245_1764 ();
 b15zdnd00an1n01x5 FILLER_245_1768 ();
 b15zdnd11an1n04x5 FILLER_245_1772 ();
 b15zdnd11an1n08x5 FILLER_245_1779 ();
 b15zdnd00an1n02x5 FILLER_245_1787 ();
 b15zdnd00an1n01x5 FILLER_245_1789 ();
 b15zdnd11an1n64x5 FILLER_245_1842 ();
 b15zdnd11an1n64x5 FILLER_245_1906 ();
 b15zdnd11an1n16x5 FILLER_245_1970 ();
 b15zdnd11an1n04x5 FILLER_245_1986 ();
 b15zdnd00an1n02x5 FILLER_245_1990 ();
 b15zdnd11an1n08x5 FILLER_245_2010 ();
 b15zdnd00an1n01x5 FILLER_245_2018 ();
 b15zdnd11an1n64x5 FILLER_245_2029 ();
 b15zdnd11an1n32x5 FILLER_245_2093 ();
 b15zdnd11an1n08x5 FILLER_245_2125 ();
 b15zdnd11an1n64x5 FILLER_245_2140 ();
 b15zdnd11an1n16x5 FILLER_245_2204 ();
 b15zdnd11an1n08x5 FILLER_245_2220 ();
 b15zdnd00an1n02x5 FILLER_245_2228 ();
 b15zdnd00an1n01x5 FILLER_245_2230 ();
 b15zdnd11an1n08x5 FILLER_245_2273 ();
 b15zdnd00an1n02x5 FILLER_245_2281 ();
 b15zdnd00an1n01x5 FILLER_245_2283 ();
 b15zdnd11an1n64x5 FILLER_246_8 ();
 b15zdnd11an1n64x5 FILLER_246_72 ();
 b15zdnd11an1n04x5 FILLER_246_136 ();
 b15zdnd00an1n02x5 FILLER_246_140 ();
 b15zdnd11an1n64x5 FILLER_246_194 ();
 b15zdnd11an1n32x5 FILLER_246_258 ();
 b15zdnd11an1n16x5 FILLER_246_290 ();
 b15zdnd11an1n04x5 FILLER_246_306 ();
 b15zdnd00an1n02x5 FILLER_246_310 ();
 b15zdnd11an1n08x5 FILLER_246_343 ();
 b15zdnd11an1n04x5 FILLER_246_351 ();
 b15zdnd00an1n02x5 FILLER_246_355 ();
 b15zdnd00an1n01x5 FILLER_246_357 ();
 b15zdnd11an1n08x5 FILLER_246_365 ();
 b15zdnd11an1n64x5 FILLER_246_385 ();
 b15zdnd11an1n64x5 FILLER_246_449 ();
 b15zdnd11an1n64x5 FILLER_246_513 ();
 b15zdnd11an1n64x5 FILLER_246_577 ();
 b15zdnd11an1n64x5 FILLER_246_641 ();
 b15zdnd11an1n08x5 FILLER_246_705 ();
 b15zdnd11an1n04x5 FILLER_246_713 ();
 b15zdnd00an1n01x5 FILLER_246_717 ();
 b15zdnd11an1n64x5 FILLER_246_726 ();
 b15zdnd11an1n64x5 FILLER_246_790 ();
 b15zdnd11an1n64x5 FILLER_246_854 ();
 b15zdnd11an1n32x5 FILLER_246_918 ();
 b15zdnd11an1n16x5 FILLER_246_950 ();
 b15zdnd11an1n04x5 FILLER_246_966 ();
 b15zdnd00an1n02x5 FILLER_246_970 ();
 b15zdnd11an1n04x5 FILLER_246_975 ();
 b15zdnd00an1n02x5 FILLER_246_979 ();
 b15zdnd11an1n64x5 FILLER_246_984 ();
 b15zdnd11an1n64x5 FILLER_246_1048 ();
 b15zdnd11an1n64x5 FILLER_246_1112 ();
 b15zdnd11an1n64x5 FILLER_246_1176 ();
 b15zdnd11an1n64x5 FILLER_246_1240 ();
 b15zdnd11an1n64x5 FILLER_246_1304 ();
 b15zdnd11an1n64x5 FILLER_246_1368 ();
 b15zdnd11an1n64x5 FILLER_246_1432 ();
 b15zdnd11an1n64x5 FILLER_246_1496 ();
 b15zdnd11an1n64x5 FILLER_246_1560 ();
 b15zdnd11an1n32x5 FILLER_246_1624 ();
 b15zdnd00an1n01x5 FILLER_246_1656 ();
 b15zdnd11an1n64x5 FILLER_246_1660 ();
 b15zdnd11an1n32x5 FILLER_246_1724 ();
 b15zdnd11an1n16x5 FILLER_246_1756 ();
 b15zdnd11an1n04x5 FILLER_246_1772 ();
 b15zdnd00an1n01x5 FILLER_246_1776 ();
 b15zdnd11an1n32x5 FILLER_246_1780 ();
 b15zdnd00an1n02x5 FILLER_246_1812 ();
 b15zdnd00an1n01x5 FILLER_246_1814 ();
 b15zdnd11an1n16x5 FILLER_246_1818 ();
 b15zdnd00an1n02x5 FILLER_246_1834 ();
 b15zdnd11an1n64x5 FILLER_246_1888 ();
 b15zdnd11an1n64x5 FILLER_246_1952 ();
 b15zdnd11an1n32x5 FILLER_246_2016 ();
 b15zdnd11an1n08x5 FILLER_246_2048 ();
 b15zdnd00an1n01x5 FILLER_246_2056 ();
 b15zdnd11an1n64x5 FILLER_246_2060 ();
 b15zdnd11an1n16x5 FILLER_246_2124 ();
 b15zdnd11an1n08x5 FILLER_246_2140 ();
 b15zdnd11an1n04x5 FILLER_246_2148 ();
 b15zdnd00an1n02x5 FILLER_246_2152 ();
 b15zdnd11an1n32x5 FILLER_246_2162 ();
 b15zdnd11an1n08x5 FILLER_246_2194 ();
 b15zdnd00an1n02x5 FILLER_246_2202 ();
 b15zdnd00an1n01x5 FILLER_246_2204 ();
 b15zdnd11an1n16x5 FILLER_246_2214 ();
 b15zdnd00an1n02x5 FILLER_246_2230 ();
 b15zdnd00an1n02x5 FILLER_246_2274 ();
 b15zdnd11an1n64x5 FILLER_247_0 ();
 b15zdnd11an1n64x5 FILLER_247_64 ();
 b15zdnd11an1n32x5 FILLER_247_128 ();
 b15zdnd11an1n04x5 FILLER_247_163 ();
 b15zdnd11an1n64x5 FILLER_247_170 ();
 b15zdnd11an1n64x5 FILLER_247_234 ();
 b15zdnd11an1n64x5 FILLER_247_298 ();
 b15zdnd11an1n64x5 FILLER_247_362 ();
 b15zdnd11an1n64x5 FILLER_247_426 ();
 b15zdnd11an1n64x5 FILLER_247_490 ();
 b15zdnd11an1n64x5 FILLER_247_554 ();
 b15zdnd11an1n64x5 FILLER_247_618 ();
 b15zdnd11an1n64x5 FILLER_247_682 ();
 b15zdnd11an1n64x5 FILLER_247_746 ();
 b15zdnd11an1n64x5 FILLER_247_810 ();
 b15zdnd11an1n64x5 FILLER_247_874 ();
 b15zdnd11an1n32x5 FILLER_247_938 ();
 b15zdnd11an1n08x5 FILLER_247_970 ();
 b15zdnd11an1n04x5 FILLER_247_978 ();
 b15zdnd00an1n01x5 FILLER_247_982 ();
 b15zdnd11an1n64x5 FILLER_247_986 ();
 b15zdnd11an1n64x5 FILLER_247_1050 ();
 b15zdnd11an1n64x5 FILLER_247_1114 ();
 b15zdnd11an1n64x5 FILLER_247_1178 ();
 b15zdnd11an1n64x5 FILLER_247_1242 ();
 b15zdnd11an1n64x5 FILLER_247_1306 ();
 b15zdnd11an1n64x5 FILLER_247_1370 ();
 b15zdnd11an1n64x5 FILLER_247_1434 ();
 b15zdnd11an1n64x5 FILLER_247_1498 ();
 b15zdnd11an1n64x5 FILLER_247_1562 ();
 b15zdnd11an1n64x5 FILLER_247_1626 ();
 b15zdnd11an1n64x5 FILLER_247_1690 ();
 b15zdnd11an1n64x5 FILLER_247_1754 ();
 b15zdnd11an1n32x5 FILLER_247_1818 ();
 b15zdnd11an1n04x5 FILLER_247_1850 ();
 b15zdnd00an1n01x5 FILLER_247_1854 ();
 b15zdnd11an1n04x5 FILLER_247_1858 ();
 b15zdnd11an1n08x5 FILLER_247_1865 ();
 b15zdnd00an1n01x5 FILLER_247_1873 ();
 b15zdnd11an1n64x5 FILLER_247_1894 ();
 b15zdnd11an1n64x5 FILLER_247_1958 ();
 b15zdnd11an1n32x5 FILLER_247_2022 ();
 b15zdnd11an1n16x5 FILLER_247_2054 ();
 b15zdnd00an1n02x5 FILLER_247_2070 ();
 b15zdnd11an1n64x5 FILLER_247_2078 ();
 b15zdnd11an1n32x5 FILLER_247_2142 ();
 b15zdnd11an1n16x5 FILLER_247_2174 ();
 b15zdnd11an1n08x5 FILLER_247_2190 ();
 b15zdnd00an1n02x5 FILLER_247_2198 ();
 b15zdnd00an1n01x5 FILLER_247_2200 ();
 b15zdnd11an1n16x5 FILLER_247_2211 ();
 b15zdnd11an1n08x5 FILLER_247_2227 ();
 b15zdnd11an1n04x5 FILLER_247_2235 ();
 b15zdnd00an1n01x5 FILLER_247_2239 ();
 b15zdnd00an1n02x5 FILLER_247_2282 ();
 b15zdnd11an1n64x5 FILLER_248_8 ();
 b15zdnd11an1n64x5 FILLER_248_72 ();
 b15zdnd11an1n64x5 FILLER_248_136 ();
 b15zdnd00an1n01x5 FILLER_248_200 ();
 b15zdnd11an1n64x5 FILLER_248_243 ();
 b15zdnd11an1n32x5 FILLER_248_307 ();
 b15zdnd11an1n08x5 FILLER_248_339 ();
 b15zdnd00an1n02x5 FILLER_248_347 ();
 b15zdnd00an1n01x5 FILLER_248_349 ();
 b15zdnd11an1n64x5 FILLER_248_358 ();
 b15zdnd11an1n64x5 FILLER_248_422 ();
 b15zdnd11an1n64x5 FILLER_248_486 ();
 b15zdnd11an1n64x5 FILLER_248_550 ();
 b15zdnd11an1n64x5 FILLER_248_614 ();
 b15zdnd11an1n32x5 FILLER_248_678 ();
 b15zdnd11an1n08x5 FILLER_248_710 ();
 b15zdnd11an1n64x5 FILLER_248_726 ();
 b15zdnd11an1n64x5 FILLER_248_790 ();
 b15zdnd11an1n64x5 FILLER_248_854 ();
 b15zdnd11an1n64x5 FILLER_248_918 ();
 b15zdnd11an1n64x5 FILLER_248_982 ();
 b15zdnd11an1n64x5 FILLER_248_1046 ();
 b15zdnd11an1n64x5 FILLER_248_1110 ();
 b15zdnd11an1n64x5 FILLER_248_1174 ();
 b15zdnd11an1n16x5 FILLER_248_1238 ();
 b15zdnd11an1n08x5 FILLER_248_1254 ();
 b15zdnd11an1n04x5 FILLER_248_1262 ();
 b15zdnd11an1n64x5 FILLER_248_1275 ();
 b15zdnd11an1n64x5 FILLER_248_1339 ();
 b15zdnd11an1n64x5 FILLER_248_1403 ();
 b15zdnd11an1n64x5 FILLER_248_1467 ();
 b15zdnd11an1n64x5 FILLER_248_1531 ();
 b15zdnd11an1n64x5 FILLER_248_1595 ();
 b15zdnd11an1n64x5 FILLER_248_1659 ();
 b15zdnd11an1n64x5 FILLER_248_1723 ();
 b15zdnd11an1n64x5 FILLER_248_1787 ();
 b15zdnd11an1n08x5 FILLER_248_1851 ();
 b15zdnd00an1n02x5 FILLER_248_1859 ();
 b15zdnd11an1n64x5 FILLER_248_1864 ();
 b15zdnd11an1n64x5 FILLER_248_1928 ();
 b15zdnd11an1n32x5 FILLER_248_1992 ();
 b15zdnd11an1n16x5 FILLER_248_2024 ();
 b15zdnd11an1n08x5 FILLER_248_2040 ();
 b15zdnd11an1n04x5 FILLER_248_2048 ();
 b15zdnd00an1n02x5 FILLER_248_2052 ();
 b15zdnd11an1n08x5 FILLER_248_2071 ();
 b15zdnd00an1n02x5 FILLER_248_2079 ();
 b15zdnd00an1n01x5 FILLER_248_2081 ();
 b15zdnd11an1n64x5 FILLER_248_2090 ();
 b15zdnd11an1n32x5 FILLER_248_2162 ();
 b15zdnd11an1n04x5 FILLER_248_2194 ();
 b15zdnd11an1n32x5 FILLER_248_2213 ();
 b15zdnd11an1n16x5 FILLER_248_2245 ();
 b15zdnd11an1n08x5 FILLER_248_2261 ();
 b15zdnd11an1n04x5 FILLER_248_2269 ();
 b15zdnd00an1n02x5 FILLER_248_2273 ();
 b15zdnd00an1n01x5 FILLER_248_2275 ();
 b15zdnd11an1n64x5 FILLER_249_0 ();
 b15zdnd11an1n64x5 FILLER_249_64 ();
 b15zdnd11an1n64x5 FILLER_249_128 ();
 b15zdnd11an1n64x5 FILLER_249_192 ();
 b15zdnd11an1n64x5 FILLER_249_256 ();
 b15zdnd11an1n64x5 FILLER_249_320 ();
 b15zdnd11an1n64x5 FILLER_249_384 ();
 b15zdnd11an1n64x5 FILLER_249_448 ();
 b15zdnd11an1n64x5 FILLER_249_512 ();
 b15zdnd11an1n64x5 FILLER_249_576 ();
 b15zdnd11an1n64x5 FILLER_249_640 ();
 b15zdnd11an1n64x5 FILLER_249_704 ();
 b15zdnd11an1n64x5 FILLER_249_768 ();
 b15zdnd11an1n64x5 FILLER_249_832 ();
 b15zdnd11an1n64x5 FILLER_249_896 ();
 b15zdnd11an1n64x5 FILLER_249_960 ();
 b15zdnd11an1n64x5 FILLER_249_1024 ();
 b15zdnd11an1n64x5 FILLER_249_1088 ();
 b15zdnd11an1n64x5 FILLER_249_1152 ();
 b15zdnd11an1n16x5 FILLER_249_1216 ();
 b15zdnd11an1n08x5 FILLER_249_1232 ();
 b15zdnd11an1n04x5 FILLER_249_1240 ();
 b15zdnd00an1n01x5 FILLER_249_1244 ();
 b15zdnd11an1n64x5 FILLER_249_1248 ();
 b15zdnd11an1n64x5 FILLER_249_1312 ();
 b15zdnd11an1n64x5 FILLER_249_1376 ();
 b15zdnd11an1n64x5 FILLER_249_1440 ();
 b15zdnd11an1n64x5 FILLER_249_1504 ();
 b15zdnd11an1n16x5 FILLER_249_1568 ();
 b15zdnd11an1n08x5 FILLER_249_1584 ();
 b15zdnd11an1n04x5 FILLER_249_1592 ();
 b15zdnd00an1n02x5 FILLER_249_1596 ();
 b15zdnd00an1n01x5 FILLER_249_1598 ();
 b15zdnd11an1n64x5 FILLER_249_1608 ();
 b15zdnd11an1n64x5 FILLER_249_1672 ();
 b15zdnd11an1n32x5 FILLER_249_1736 ();
 b15zdnd11an1n16x5 FILLER_249_1768 ();
 b15zdnd11an1n08x5 FILLER_249_1784 ();
 b15zdnd00an1n02x5 FILLER_249_1792 ();
 b15zdnd11an1n64x5 FILLER_249_1803 ();
 b15zdnd11an1n64x5 FILLER_249_1867 ();
 b15zdnd11an1n64x5 FILLER_249_1931 ();
 b15zdnd11an1n16x5 FILLER_249_1995 ();
 b15zdnd00an1n01x5 FILLER_249_2011 ();
 b15zdnd11an1n64x5 FILLER_249_2030 ();
 b15zdnd11an1n64x5 FILLER_249_2094 ();
 b15zdnd11an1n08x5 FILLER_249_2158 ();
 b15zdnd11an1n64x5 FILLER_249_2208 ();
 b15zdnd11an1n08x5 FILLER_249_2272 ();
 b15zdnd11an1n04x5 FILLER_249_2280 ();
 b15zdnd11an1n64x5 FILLER_250_8 ();
 b15zdnd11an1n64x5 FILLER_250_72 ();
 b15zdnd11an1n64x5 FILLER_250_136 ();
 b15zdnd11an1n64x5 FILLER_250_200 ();
 b15zdnd11an1n64x5 FILLER_250_264 ();
 b15zdnd11an1n32x5 FILLER_250_328 ();
 b15zdnd11an1n08x5 FILLER_250_360 ();
 b15zdnd11an1n04x5 FILLER_250_368 ();
 b15zdnd00an1n02x5 FILLER_250_372 ();
 b15zdnd00an1n01x5 FILLER_250_374 ();
 b15zdnd11an1n64x5 FILLER_250_379 ();
 b15zdnd11an1n08x5 FILLER_250_443 ();
 b15zdnd11an1n04x5 FILLER_250_451 ();
 b15zdnd00an1n02x5 FILLER_250_455 ();
 b15zdnd00an1n01x5 FILLER_250_457 ();
 b15zdnd11an1n04x5 FILLER_250_465 ();
 b15zdnd11an1n04x5 FILLER_250_481 ();
 b15zdnd11an1n64x5 FILLER_250_494 ();
 b15zdnd11an1n64x5 FILLER_250_558 ();
 b15zdnd11an1n64x5 FILLER_250_622 ();
 b15zdnd11an1n32x5 FILLER_250_686 ();
 b15zdnd11an1n64x5 FILLER_250_726 ();
 b15zdnd11an1n64x5 FILLER_250_790 ();
 b15zdnd11an1n64x5 FILLER_250_854 ();
 b15zdnd11an1n64x5 FILLER_250_918 ();
 b15zdnd11an1n64x5 FILLER_250_982 ();
 b15zdnd11an1n64x5 FILLER_250_1046 ();
 b15zdnd11an1n64x5 FILLER_250_1110 ();
 b15zdnd11an1n64x5 FILLER_250_1174 ();
 b15zdnd11an1n04x5 FILLER_250_1238 ();
 b15zdnd00an1n02x5 FILLER_250_1242 ();
 b15zdnd00an1n01x5 FILLER_250_1244 ();
 b15zdnd11an1n64x5 FILLER_250_1272 ();
 b15zdnd11an1n32x5 FILLER_250_1336 ();
 b15zdnd00an1n02x5 FILLER_250_1368 ();
 b15zdnd11an1n04x5 FILLER_250_1373 ();
 b15zdnd11an1n04x5 FILLER_250_1380 ();
 b15zdnd11an1n08x5 FILLER_250_1387 ();
 b15zdnd00an1n02x5 FILLER_250_1395 ();
 b15zdnd00an1n01x5 FILLER_250_1397 ();
 b15zdnd11an1n64x5 FILLER_250_1401 ();
 b15zdnd11an1n64x5 FILLER_250_1465 ();
 b15zdnd11an1n64x5 FILLER_250_1529 ();
 b15zdnd11an1n04x5 FILLER_250_1593 ();
 b15zdnd11an1n64x5 FILLER_250_1606 ();
 b15zdnd11an1n64x5 FILLER_250_1670 ();
 b15zdnd11an1n64x5 FILLER_250_1734 ();
 b15zdnd11an1n64x5 FILLER_250_1798 ();
 b15zdnd11an1n64x5 FILLER_250_1862 ();
 b15zdnd11an1n64x5 FILLER_250_1926 ();
 b15zdnd11an1n64x5 FILLER_250_1990 ();
 b15zdnd11an1n32x5 FILLER_250_2096 ();
 b15zdnd11an1n16x5 FILLER_250_2128 ();
 b15zdnd11an1n08x5 FILLER_250_2144 ();
 b15zdnd00an1n02x5 FILLER_250_2152 ();
 b15zdnd11an1n32x5 FILLER_250_2162 ();
 b15zdnd11an1n16x5 FILLER_250_2194 ();
 b15zdnd00an1n01x5 FILLER_250_2210 ();
 b15zdnd11an1n32x5 FILLER_250_2236 ();
 b15zdnd11an1n08x5 FILLER_250_2268 ();
 b15zdnd11an1n64x5 FILLER_251_0 ();
 b15zdnd11an1n64x5 FILLER_251_64 ();
 b15zdnd11an1n64x5 FILLER_251_128 ();
 b15zdnd11an1n64x5 FILLER_251_192 ();
 b15zdnd11an1n64x5 FILLER_251_256 ();
 b15zdnd11an1n64x5 FILLER_251_320 ();
 b15zdnd11an1n64x5 FILLER_251_384 ();
 b15zdnd11an1n64x5 FILLER_251_448 ();
 b15zdnd11an1n64x5 FILLER_251_512 ();
 b15zdnd11an1n64x5 FILLER_251_576 ();
 b15zdnd11an1n32x5 FILLER_251_640 ();
 b15zdnd11an1n16x5 FILLER_251_672 ();
 b15zdnd11an1n08x5 FILLER_251_688 ();
 b15zdnd00an1n01x5 FILLER_251_696 ();
 b15zdnd11an1n64x5 FILLER_251_739 ();
 b15zdnd11an1n64x5 FILLER_251_803 ();
 b15zdnd11an1n64x5 FILLER_251_867 ();
 b15zdnd11an1n64x5 FILLER_251_931 ();
 b15zdnd11an1n64x5 FILLER_251_995 ();
 b15zdnd11an1n64x5 FILLER_251_1059 ();
 b15zdnd11an1n64x5 FILLER_251_1123 ();
 b15zdnd11an1n64x5 FILLER_251_1187 ();
 b15zdnd11an1n64x5 FILLER_251_1251 ();
 b15zdnd11an1n32x5 FILLER_251_1315 ();
 b15zdnd11an1n04x5 FILLER_251_1347 ();
 b15zdnd00an1n01x5 FILLER_251_1351 ();
 b15zdnd11an1n04x5 FILLER_251_1404 ();
 b15zdnd11an1n64x5 FILLER_251_1411 ();
 b15zdnd11an1n32x5 FILLER_251_1475 ();
 b15zdnd11an1n08x5 FILLER_251_1507 ();
 b15zdnd11an1n04x5 FILLER_251_1515 ();
 b15zdnd00an1n02x5 FILLER_251_1519 ();
 b15zdnd11an1n64x5 FILLER_251_1573 ();
 b15zdnd11an1n64x5 FILLER_251_1637 ();
 b15zdnd11an1n64x5 FILLER_251_1701 ();
 b15zdnd11an1n64x5 FILLER_251_1765 ();
 b15zdnd11an1n64x5 FILLER_251_1829 ();
 b15zdnd11an1n64x5 FILLER_251_1893 ();
 b15zdnd11an1n64x5 FILLER_251_1957 ();
 b15zdnd11an1n64x5 FILLER_251_2021 ();
 b15zdnd11an1n32x5 FILLER_251_2085 ();
 b15zdnd11an1n08x5 FILLER_251_2117 ();
 b15zdnd11an1n04x5 FILLER_251_2125 ();
 b15zdnd11an1n64x5 FILLER_251_2171 ();
 b15zdnd11an1n32x5 FILLER_251_2235 ();
 b15zdnd11an1n16x5 FILLER_251_2267 ();
 b15zdnd00an1n01x5 FILLER_251_2283 ();
 b15zdnd11an1n64x5 FILLER_252_8 ();
 b15zdnd11an1n64x5 FILLER_252_72 ();
 b15zdnd11an1n64x5 FILLER_252_136 ();
 b15zdnd11an1n64x5 FILLER_252_200 ();
 b15zdnd11an1n64x5 FILLER_252_264 ();
 b15zdnd11an1n64x5 FILLER_252_328 ();
 b15zdnd11an1n64x5 FILLER_252_392 ();
 b15zdnd11an1n16x5 FILLER_252_456 ();
 b15zdnd00an1n01x5 FILLER_252_472 ();
 b15zdnd11an1n04x5 FILLER_252_479 ();
 b15zdnd11an1n64x5 FILLER_252_495 ();
 b15zdnd11an1n64x5 FILLER_252_559 ();
 b15zdnd11an1n32x5 FILLER_252_623 ();
 b15zdnd11an1n04x5 FILLER_252_655 ();
 b15zdnd00an1n01x5 FILLER_252_659 ();
 b15zdnd11an1n32x5 FILLER_252_673 ();
 b15zdnd00an1n01x5 FILLER_252_705 ();
 b15zdnd11an1n04x5 FILLER_252_709 ();
 b15zdnd00an1n02x5 FILLER_252_716 ();
 b15zdnd11an1n64x5 FILLER_252_726 ();
 b15zdnd11an1n64x5 FILLER_252_790 ();
 b15zdnd11an1n64x5 FILLER_252_854 ();
 b15zdnd11an1n64x5 FILLER_252_918 ();
 b15zdnd11an1n64x5 FILLER_252_982 ();
 b15zdnd11an1n64x5 FILLER_252_1046 ();
 b15zdnd11an1n64x5 FILLER_252_1110 ();
 b15zdnd11an1n64x5 FILLER_252_1174 ();
 b15zdnd11an1n64x5 FILLER_252_1238 ();
 b15zdnd11an1n64x5 FILLER_252_1302 ();
 b15zdnd11an1n04x5 FILLER_252_1366 ();
 b15zdnd00an1n02x5 FILLER_252_1370 ();
 b15zdnd00an1n01x5 FILLER_252_1372 ();
 b15zdnd11an1n64x5 FILLER_252_1425 ();
 b15zdnd11an1n32x5 FILLER_252_1489 ();
 b15zdnd11an1n16x5 FILLER_252_1521 ();
 b15zdnd00an1n02x5 FILLER_252_1537 ();
 b15zdnd11an1n04x5 FILLER_252_1542 ();
 b15zdnd11an1n04x5 FILLER_252_1549 ();
 b15zdnd11an1n64x5 FILLER_252_1556 ();
 b15zdnd11an1n64x5 FILLER_252_1620 ();
 b15zdnd11an1n64x5 FILLER_252_1684 ();
 b15zdnd11an1n64x5 FILLER_252_1748 ();
 b15zdnd11an1n64x5 FILLER_252_1812 ();
 b15zdnd11an1n64x5 FILLER_252_1876 ();
 b15zdnd11an1n64x5 FILLER_252_1940 ();
 b15zdnd11an1n64x5 FILLER_252_2004 ();
 b15zdnd11an1n32x5 FILLER_252_2068 ();
 b15zdnd11an1n16x5 FILLER_252_2100 ();
 b15zdnd00an1n01x5 FILLER_252_2116 ();
 b15zdnd11an1n08x5 FILLER_252_2142 ();
 b15zdnd11an1n04x5 FILLER_252_2150 ();
 b15zdnd11an1n64x5 FILLER_252_2162 ();
 b15zdnd11an1n32x5 FILLER_252_2226 ();
 b15zdnd11an1n16x5 FILLER_252_2258 ();
 b15zdnd00an1n02x5 FILLER_252_2274 ();
 b15zdnd11an1n64x5 FILLER_253_0 ();
 b15zdnd11an1n64x5 FILLER_253_64 ();
 b15zdnd11an1n16x5 FILLER_253_128 ();
 b15zdnd11an1n08x5 FILLER_253_144 ();
 b15zdnd11an1n64x5 FILLER_253_194 ();
 b15zdnd11an1n64x5 FILLER_253_258 ();
 b15zdnd11an1n64x5 FILLER_253_322 ();
 b15zdnd11an1n64x5 FILLER_253_386 ();
 b15zdnd11an1n16x5 FILLER_253_450 ();
 b15zdnd11an1n08x5 FILLER_253_466 ();
 b15zdnd00an1n01x5 FILLER_253_474 ();
 b15zdnd11an1n64x5 FILLER_253_485 ();
 b15zdnd11an1n64x5 FILLER_253_549 ();
 b15zdnd11an1n64x5 FILLER_253_613 ();
 b15zdnd11an1n08x5 FILLER_253_677 ();
 b15zdnd00an1n01x5 FILLER_253_685 ();
 b15zdnd11an1n64x5 FILLER_253_738 ();
 b15zdnd11an1n64x5 FILLER_253_802 ();
 b15zdnd11an1n64x5 FILLER_253_866 ();
 b15zdnd11an1n64x5 FILLER_253_930 ();
 b15zdnd11an1n64x5 FILLER_253_994 ();
 b15zdnd11an1n64x5 FILLER_253_1058 ();
 b15zdnd11an1n64x5 FILLER_253_1122 ();
 b15zdnd11an1n64x5 FILLER_253_1186 ();
 b15zdnd11an1n64x5 FILLER_253_1250 ();
 b15zdnd11an1n64x5 FILLER_253_1314 ();
 b15zdnd11an1n16x5 FILLER_253_1378 ();
 b15zdnd00an1n01x5 FILLER_253_1394 ();
 b15zdnd11an1n64x5 FILLER_253_1398 ();
 b15zdnd11an1n64x5 FILLER_253_1462 ();
 b15zdnd11an1n64x5 FILLER_253_1526 ();
 b15zdnd11an1n64x5 FILLER_253_1590 ();
 b15zdnd11an1n64x5 FILLER_253_1654 ();
 b15zdnd11an1n64x5 FILLER_253_1718 ();
 b15zdnd11an1n64x5 FILLER_253_1782 ();
 b15zdnd11an1n64x5 FILLER_253_1846 ();
 b15zdnd11an1n64x5 FILLER_253_1910 ();
 b15zdnd11an1n64x5 FILLER_253_1974 ();
 b15zdnd11an1n32x5 FILLER_253_2038 ();
 b15zdnd11an1n16x5 FILLER_253_2070 ();
 b15zdnd11an1n08x5 FILLER_253_2086 ();
 b15zdnd00an1n02x5 FILLER_253_2094 ();
 b15zdnd11an1n64x5 FILLER_253_2106 ();
 b15zdnd11an1n64x5 FILLER_253_2170 ();
 b15zdnd11an1n32x5 FILLER_253_2234 ();
 b15zdnd11an1n16x5 FILLER_253_2266 ();
 b15zdnd00an1n02x5 FILLER_253_2282 ();
 b15zdnd11an1n64x5 FILLER_254_8 ();
 b15zdnd11an1n64x5 FILLER_254_72 ();
 b15zdnd11an1n64x5 FILLER_254_136 ();
 b15zdnd11an1n64x5 FILLER_254_200 ();
 b15zdnd11an1n64x5 FILLER_254_264 ();
 b15zdnd11an1n64x5 FILLER_254_328 ();
 b15zdnd11an1n64x5 FILLER_254_392 ();
 b15zdnd11an1n04x5 FILLER_254_456 ();
 b15zdnd00an1n02x5 FILLER_254_460 ();
 b15zdnd11an1n04x5 FILLER_254_467 ();
 b15zdnd00an1n02x5 FILLER_254_471 ();
 b15zdnd11an1n08x5 FILLER_254_479 ();
 b15zdnd00an1n02x5 FILLER_254_487 ();
 b15zdnd11an1n32x5 FILLER_254_492 ();
 b15zdnd11an1n08x5 FILLER_254_524 ();
 b15zdnd11an1n04x5 FILLER_254_532 ();
 b15zdnd00an1n02x5 FILLER_254_536 ();
 b15zdnd11an1n64x5 FILLER_254_541 ();
 b15zdnd11an1n64x5 FILLER_254_605 ();
 b15zdnd11an1n32x5 FILLER_254_669 ();
 b15zdnd11an1n08x5 FILLER_254_701 ();
 b15zdnd00an1n02x5 FILLER_254_709 ();
 b15zdnd11an1n04x5 FILLER_254_714 ();
 b15zdnd00an1n02x5 FILLER_254_726 ();
 b15zdnd11an1n32x5 FILLER_254_770 ();
 b15zdnd00an1n02x5 FILLER_254_802 ();
 b15zdnd11an1n64x5 FILLER_254_846 ();
 b15zdnd11an1n64x5 FILLER_254_910 ();
 b15zdnd11an1n64x5 FILLER_254_974 ();
 b15zdnd11an1n64x5 FILLER_254_1038 ();
 b15zdnd11an1n64x5 FILLER_254_1102 ();
 b15zdnd11an1n64x5 FILLER_254_1166 ();
 b15zdnd11an1n16x5 FILLER_254_1230 ();
 b15zdnd11an1n08x5 FILLER_254_1246 ();
 b15zdnd00an1n02x5 FILLER_254_1254 ();
 b15zdnd00an1n01x5 FILLER_254_1256 ();
 b15zdnd11an1n64x5 FILLER_254_1260 ();
 b15zdnd11an1n32x5 FILLER_254_1324 ();
 b15zdnd11an1n08x5 FILLER_254_1356 ();
 b15zdnd11an1n04x5 FILLER_254_1364 ();
 b15zdnd00an1n02x5 FILLER_254_1368 ();
 b15zdnd11an1n64x5 FILLER_254_1394 ();
 b15zdnd11an1n64x5 FILLER_254_1458 ();
 b15zdnd11an1n64x5 FILLER_254_1522 ();
 b15zdnd11an1n64x5 FILLER_254_1586 ();
 b15zdnd11an1n64x5 FILLER_254_1650 ();
 b15zdnd11an1n64x5 FILLER_254_1714 ();
 b15zdnd11an1n64x5 FILLER_254_1778 ();
 b15zdnd11an1n64x5 FILLER_254_1842 ();
 b15zdnd11an1n64x5 FILLER_254_1906 ();
 b15zdnd11an1n64x5 FILLER_254_1970 ();
 b15zdnd11an1n64x5 FILLER_254_2034 ();
 b15zdnd11an1n32x5 FILLER_254_2098 ();
 b15zdnd11an1n16x5 FILLER_254_2130 ();
 b15zdnd11an1n08x5 FILLER_254_2146 ();
 b15zdnd11an1n04x5 FILLER_254_2162 ();
 b15zdnd00an1n02x5 FILLER_254_2166 ();
 b15zdnd00an1n01x5 FILLER_254_2168 ();
 b15zdnd11an1n32x5 FILLER_254_2181 ();
 b15zdnd11an1n16x5 FILLER_254_2213 ();
 b15zdnd00an1n01x5 FILLER_254_2229 ();
 b15zdnd11an1n16x5 FILLER_254_2248 ();
 b15zdnd11an1n08x5 FILLER_254_2264 ();
 b15zdnd11an1n04x5 FILLER_254_2272 ();
 b15zdnd11an1n64x5 FILLER_255_0 ();
 b15zdnd11an1n64x5 FILLER_255_64 ();
 b15zdnd11an1n64x5 FILLER_255_128 ();
 b15zdnd11an1n08x5 FILLER_255_192 ();
 b15zdnd00an1n01x5 FILLER_255_200 ();
 b15zdnd11an1n64x5 FILLER_255_243 ();
 b15zdnd11an1n64x5 FILLER_255_307 ();
 b15zdnd11an1n64x5 FILLER_255_371 ();
 b15zdnd11an1n16x5 FILLER_255_435 ();
 b15zdnd11an1n04x5 FILLER_255_451 ();
 b15zdnd00an1n02x5 FILLER_255_455 ();
 b15zdnd00an1n01x5 FILLER_255_457 ();
 b15zdnd11an1n04x5 FILLER_255_465 ();
 b15zdnd11an1n04x5 FILLER_255_473 ();
 b15zdnd11an1n16x5 FILLER_255_480 ();
 b15zdnd00an1n02x5 FILLER_255_496 ();
 b15zdnd00an1n01x5 FILLER_255_498 ();
 b15zdnd11an1n04x5 FILLER_255_502 ();
 b15zdnd00an1n01x5 FILLER_255_506 ();
 b15zdnd11an1n08x5 FILLER_255_549 ();
 b15zdnd00an1n01x5 FILLER_255_557 ();
 b15zdnd11an1n64x5 FILLER_255_561 ();
 b15zdnd11an1n64x5 FILLER_255_625 ();
 b15zdnd11an1n64x5 FILLER_255_689 ();
 b15zdnd11an1n32x5 FILLER_255_753 ();
 b15zdnd11an1n08x5 FILLER_255_785 ();
 b15zdnd11an1n64x5 FILLER_255_845 ();
 b15zdnd11an1n64x5 FILLER_255_909 ();
 b15zdnd11an1n64x5 FILLER_255_973 ();
 b15zdnd11an1n64x5 FILLER_255_1037 ();
 b15zdnd11an1n64x5 FILLER_255_1101 ();
 b15zdnd11an1n64x5 FILLER_255_1165 ();
 b15zdnd11an1n16x5 FILLER_255_1229 ();
 b15zdnd11an1n08x5 FILLER_255_1245 ();
 b15zdnd11an1n04x5 FILLER_255_1253 ();
 b15zdnd11an1n64x5 FILLER_255_1260 ();
 b15zdnd11an1n64x5 FILLER_255_1324 ();
 b15zdnd11an1n64x5 FILLER_255_1388 ();
 b15zdnd11an1n64x5 FILLER_255_1452 ();
 b15zdnd11an1n64x5 FILLER_255_1516 ();
 b15zdnd11an1n64x5 FILLER_255_1580 ();
 b15zdnd11an1n64x5 FILLER_255_1644 ();
 b15zdnd11an1n64x5 FILLER_255_1708 ();
 b15zdnd11an1n64x5 FILLER_255_1772 ();
 b15zdnd11an1n64x5 FILLER_255_1836 ();
 b15zdnd11an1n64x5 FILLER_255_1900 ();
 b15zdnd11an1n64x5 FILLER_255_1964 ();
 b15zdnd11an1n64x5 FILLER_255_2028 ();
 b15zdnd11an1n32x5 FILLER_255_2092 ();
 b15zdnd11an1n16x5 FILLER_255_2124 ();
 b15zdnd11an1n04x5 FILLER_255_2140 ();
 b15zdnd11an1n64x5 FILLER_255_2186 ();
 b15zdnd11an1n32x5 FILLER_255_2250 ();
 b15zdnd00an1n02x5 FILLER_255_2282 ();
 b15zdnd11an1n64x5 FILLER_256_8 ();
 b15zdnd11an1n64x5 FILLER_256_72 ();
 b15zdnd11an1n64x5 FILLER_256_136 ();
 b15zdnd11an1n16x5 FILLER_256_200 ();
 b15zdnd11an1n04x5 FILLER_256_216 ();
 b15zdnd00an1n02x5 FILLER_256_220 ();
 b15zdnd00an1n01x5 FILLER_256_222 ();
 b15zdnd11an1n64x5 FILLER_256_226 ();
 b15zdnd11an1n64x5 FILLER_256_290 ();
 b15zdnd11an1n16x5 FILLER_256_354 ();
 b15zdnd11an1n08x5 FILLER_256_370 ();
 b15zdnd00an1n02x5 FILLER_256_378 ();
 b15zdnd11an1n32x5 FILLER_256_412 ();
 b15zdnd11an1n16x5 FILLER_256_444 ();
 b15zdnd11an1n04x5 FILLER_256_460 ();
 b15zdnd11an1n16x5 FILLER_256_485 ();
 b15zdnd11an1n08x5 FILLER_256_501 ();
 b15zdnd00an1n02x5 FILLER_256_509 ();
 b15zdnd11an1n64x5 FILLER_256_563 ();
 b15zdnd11an1n64x5 FILLER_256_627 ();
 b15zdnd11an1n16x5 FILLER_256_691 ();
 b15zdnd11an1n08x5 FILLER_256_707 ();
 b15zdnd00an1n02x5 FILLER_256_715 ();
 b15zdnd00an1n01x5 FILLER_256_717 ();
 b15zdnd11an1n64x5 FILLER_256_726 ();
 b15zdnd11an1n16x5 FILLER_256_790 ();
 b15zdnd11an1n04x5 FILLER_256_806 ();
 b15zdnd00an1n02x5 FILLER_256_810 ();
 b15zdnd00an1n01x5 FILLER_256_812 ();
 b15zdnd11an1n04x5 FILLER_256_816 ();
 b15zdnd11an1n08x5 FILLER_256_823 ();
 b15zdnd00an1n02x5 FILLER_256_831 ();
 b15zdnd11an1n64x5 FILLER_256_875 ();
 b15zdnd11an1n64x5 FILLER_256_939 ();
 b15zdnd11an1n64x5 FILLER_256_1003 ();
 b15zdnd11an1n32x5 FILLER_256_1067 ();
 b15zdnd11an1n16x5 FILLER_256_1099 ();
 b15zdnd11an1n08x5 FILLER_256_1115 ();
 b15zdnd11an1n64x5 FILLER_256_1143 ();
 b15zdnd11an1n16x5 FILLER_256_1207 ();
 b15zdnd11an1n08x5 FILLER_256_1223 ();
 b15zdnd00an1n01x5 FILLER_256_1231 ();
 b15zdnd11an1n64x5 FILLER_256_1284 ();
 b15zdnd11an1n64x5 FILLER_256_1348 ();
 b15zdnd11an1n64x5 FILLER_256_1412 ();
 b15zdnd11an1n64x5 FILLER_256_1476 ();
 b15zdnd11an1n64x5 FILLER_256_1540 ();
 b15zdnd11an1n32x5 FILLER_256_1604 ();
 b15zdnd11an1n16x5 FILLER_256_1636 ();
 b15zdnd00an1n01x5 FILLER_256_1652 ();
 b15zdnd11an1n04x5 FILLER_256_1656 ();
 b15zdnd11an1n64x5 FILLER_256_1663 ();
 b15zdnd11an1n64x5 FILLER_256_1727 ();
 b15zdnd11an1n64x5 FILLER_256_1791 ();
 b15zdnd11an1n64x5 FILLER_256_1855 ();
 b15zdnd11an1n64x5 FILLER_256_1919 ();
 b15zdnd11an1n64x5 FILLER_256_1983 ();
 b15zdnd11an1n32x5 FILLER_256_2047 ();
 b15zdnd11an1n16x5 FILLER_256_2079 ();
 b15zdnd11an1n04x5 FILLER_256_2095 ();
 b15zdnd00an1n01x5 FILLER_256_2099 ();
 b15zdnd11an1n32x5 FILLER_256_2115 ();
 b15zdnd11an1n04x5 FILLER_256_2147 ();
 b15zdnd00an1n02x5 FILLER_256_2151 ();
 b15zdnd00an1n01x5 FILLER_256_2153 ();
 b15zdnd11an1n08x5 FILLER_256_2162 ();
 b15zdnd11an1n04x5 FILLER_256_2170 ();
 b15zdnd00an1n02x5 FILLER_256_2174 ();
 b15zdnd00an1n01x5 FILLER_256_2176 ();
 b15zdnd11an1n04x5 FILLER_256_2202 ();
 b15zdnd11an1n08x5 FILLER_256_2224 ();
 b15zdnd00an1n02x5 FILLER_256_2274 ();
 b15zdnd11an1n64x5 FILLER_257_0 ();
 b15zdnd11an1n64x5 FILLER_257_64 ();
 b15zdnd11an1n64x5 FILLER_257_128 ();
 b15zdnd11an1n08x5 FILLER_257_192 ();
 b15zdnd00an1n02x5 FILLER_257_200 ();
 b15zdnd00an1n01x5 FILLER_257_202 ();
 b15zdnd11an1n04x5 FILLER_257_231 ();
 b15zdnd11an1n64x5 FILLER_257_238 ();
 b15zdnd11an1n64x5 FILLER_257_302 ();
 b15zdnd11an1n32x5 FILLER_257_366 ();
 b15zdnd11an1n04x5 FILLER_257_398 ();
 b15zdnd00an1n02x5 FILLER_257_402 ();
 b15zdnd00an1n01x5 FILLER_257_404 ();
 b15zdnd11an1n64x5 FILLER_257_408 ();
 b15zdnd11an1n04x5 FILLER_257_472 ();
 b15zdnd11an1n16x5 FILLER_257_518 ();
 b15zdnd00an1n02x5 FILLER_257_534 ();
 b15zdnd11an1n04x5 FILLER_257_539 ();
 b15zdnd11an1n32x5 FILLER_257_546 ();
 b15zdnd11an1n08x5 FILLER_257_578 ();
 b15zdnd11an1n04x5 FILLER_257_586 ();
 b15zdnd00an1n02x5 FILLER_257_590 ();
 b15zdnd00an1n01x5 FILLER_257_592 ();
 b15zdnd11an1n04x5 FILLER_257_596 ();
 b15zdnd11an1n64x5 FILLER_257_603 ();
 b15zdnd11an1n64x5 FILLER_257_667 ();
 b15zdnd11an1n64x5 FILLER_257_731 ();
 b15zdnd11an1n16x5 FILLER_257_795 ();
 b15zdnd11an1n04x5 FILLER_257_811 ();
 b15zdnd00an1n02x5 FILLER_257_815 ();
 b15zdnd00an1n01x5 FILLER_257_817 ();
 b15zdnd11an1n64x5 FILLER_257_821 ();
 b15zdnd11an1n32x5 FILLER_257_885 ();
 b15zdnd11an1n16x5 FILLER_257_917 ();
 b15zdnd11an1n04x5 FILLER_257_933 ();
 b15zdnd00an1n02x5 FILLER_257_937 ();
 b15zdnd11an1n64x5 FILLER_257_966 ();
 b15zdnd11an1n64x5 FILLER_257_1030 ();
 b15zdnd11an1n16x5 FILLER_257_1094 ();
 b15zdnd11an1n08x5 FILLER_257_1110 ();
 b15zdnd00an1n02x5 FILLER_257_1118 ();
 b15zdnd00an1n01x5 FILLER_257_1120 ();
 b15zdnd11an1n64x5 FILLER_257_1152 ();
 b15zdnd11an1n32x5 FILLER_257_1216 ();
 b15zdnd00an1n02x5 FILLER_257_1248 ();
 b15zdnd00an1n01x5 FILLER_257_1250 ();
 b15zdnd11an1n04x5 FILLER_257_1254 ();
 b15zdnd11an1n64x5 FILLER_257_1261 ();
 b15zdnd11an1n64x5 FILLER_257_1325 ();
 b15zdnd11an1n64x5 FILLER_257_1389 ();
 b15zdnd11an1n32x5 FILLER_257_1453 ();
 b15zdnd11an1n08x5 FILLER_257_1485 ();
 b15zdnd00an1n02x5 FILLER_257_1493 ();
 b15zdnd00an1n01x5 FILLER_257_1495 ();
 b15zdnd11an1n64x5 FILLER_257_1548 ();
 b15zdnd11an1n16x5 FILLER_257_1612 ();
 b15zdnd00an1n02x5 FILLER_257_1628 ();
 b15zdnd11an1n64x5 FILLER_257_1682 ();
 b15zdnd11an1n64x5 FILLER_257_1746 ();
 b15zdnd11an1n08x5 FILLER_257_1810 ();
 b15zdnd00an1n02x5 FILLER_257_1818 ();
 b15zdnd11an1n64x5 FILLER_257_1829 ();
 b15zdnd11an1n64x5 FILLER_257_1893 ();
 b15zdnd11an1n64x5 FILLER_257_1957 ();
 b15zdnd11an1n64x5 FILLER_257_2021 ();
 b15zdnd11an1n32x5 FILLER_257_2085 ();
 b15zdnd11an1n16x5 FILLER_257_2117 ();
 b15zdnd11an1n32x5 FILLER_257_2141 ();
 b15zdnd11an1n16x5 FILLER_257_2173 ();
 b15zdnd11an1n32x5 FILLER_257_2204 ();
 b15zdnd11an1n08x5 FILLER_257_2236 ();
 b15zdnd11an1n08x5 FILLER_257_2269 ();
 b15zdnd11an1n04x5 FILLER_257_2277 ();
 b15zdnd00an1n02x5 FILLER_257_2281 ();
 b15zdnd00an1n01x5 FILLER_257_2283 ();
 b15zdnd11an1n64x5 FILLER_258_8 ();
 b15zdnd00an1n02x5 FILLER_258_72 ();
 b15zdnd11an1n64x5 FILLER_258_77 ();
 b15zdnd11an1n32x5 FILLER_258_141 ();
 b15zdnd11an1n16x5 FILLER_258_173 ();
 b15zdnd11an1n08x5 FILLER_258_189 ();
 b15zdnd11an1n04x5 FILLER_258_197 ();
 b15zdnd11an1n64x5 FILLER_258_243 ();
 b15zdnd11an1n64x5 FILLER_258_307 ();
 b15zdnd11an1n32x5 FILLER_258_371 ();
 b15zdnd00an1n01x5 FILLER_258_403 ();
 b15zdnd11an1n64x5 FILLER_258_407 ();
 b15zdnd11an1n64x5 FILLER_258_471 ();
 b15zdnd11an1n16x5 FILLER_258_535 ();
 b15zdnd11an1n04x5 FILLER_258_593 ();
 b15zdnd00an1n02x5 FILLER_258_597 ();
 b15zdnd11an1n64x5 FILLER_258_602 ();
 b15zdnd11an1n32x5 FILLER_258_666 ();
 b15zdnd11an1n16x5 FILLER_258_698 ();
 b15zdnd11an1n04x5 FILLER_258_714 ();
 b15zdnd11an1n64x5 FILLER_258_726 ();
 b15zdnd11an1n64x5 FILLER_258_790 ();
 b15zdnd11an1n64x5 FILLER_258_854 ();
 b15zdnd11an1n16x5 FILLER_258_918 ();
 b15zdnd11an1n04x5 FILLER_258_934 ();
 b15zdnd00an1n01x5 FILLER_258_938 ();
 b15zdnd11an1n04x5 FILLER_258_942 ();
 b15zdnd00an1n02x5 FILLER_258_946 ();
 b15zdnd11an1n64x5 FILLER_258_1000 ();
 b15zdnd11an1n64x5 FILLER_258_1064 ();
 b15zdnd11an1n64x5 FILLER_258_1128 ();
 b15zdnd11an1n32x5 FILLER_258_1192 ();
 b15zdnd11an1n08x5 FILLER_258_1224 ();
 b15zdnd11an1n64x5 FILLER_258_1284 ();
 b15zdnd11an1n64x5 FILLER_258_1348 ();
 b15zdnd11an1n64x5 FILLER_258_1412 ();
 b15zdnd11an1n16x5 FILLER_258_1476 ();
 b15zdnd00an1n01x5 FILLER_258_1492 ();
 b15zdnd11an1n04x5 FILLER_258_1496 ();
 b15zdnd11an1n04x5 FILLER_258_1527 ();
 b15zdnd11an1n64x5 FILLER_258_1534 ();
 b15zdnd11an1n64x5 FILLER_258_1598 ();
 b15zdnd00an1n01x5 FILLER_258_1662 ();
 b15zdnd11an1n08x5 FILLER_258_1666 ();
 b15zdnd00an1n02x5 FILLER_258_1674 ();
 b15zdnd00an1n01x5 FILLER_258_1676 ();
 b15zdnd11an1n64x5 FILLER_258_1708 ();
 b15zdnd11an1n64x5 FILLER_258_1772 ();
 b15zdnd11an1n64x5 FILLER_258_1836 ();
 b15zdnd11an1n64x5 FILLER_258_1900 ();
 b15zdnd11an1n16x5 FILLER_258_1964 ();
 b15zdnd11an1n04x5 FILLER_258_1980 ();
 b15zdnd00an1n01x5 FILLER_258_1984 ();
 b15zdnd11an1n16x5 FILLER_258_2010 ();
 b15zdnd00an1n02x5 FILLER_258_2026 ();
 b15zdnd11an1n64x5 FILLER_258_2043 ();
 b15zdnd11an1n32x5 FILLER_258_2107 ();
 b15zdnd11an1n08x5 FILLER_258_2139 ();
 b15zdnd11an1n04x5 FILLER_258_2147 ();
 b15zdnd00an1n02x5 FILLER_258_2151 ();
 b15zdnd00an1n01x5 FILLER_258_2153 ();
 b15zdnd11an1n08x5 FILLER_258_2162 ();
 b15zdnd00an1n01x5 FILLER_258_2170 ();
 b15zdnd11an1n04x5 FILLER_258_2213 ();
 b15zdnd00an1n02x5 FILLER_258_2217 ();
 b15zdnd00an1n01x5 FILLER_258_2219 ();
 b15zdnd11an1n32x5 FILLER_258_2238 ();
 b15zdnd11an1n04x5 FILLER_258_2270 ();
 b15zdnd00an1n02x5 FILLER_258_2274 ();
 b15zdnd11an1n64x5 FILLER_259_0 ();
 b15zdnd11an1n04x5 FILLER_259_67 ();
 b15zdnd11an1n04x5 FILLER_259_80 ();
 b15zdnd11an1n64x5 FILLER_259_87 ();
 b15zdnd11an1n64x5 FILLER_259_151 ();
 b15zdnd11an1n64x5 FILLER_259_215 ();
 b15zdnd11an1n64x5 FILLER_259_279 ();
 b15zdnd11an1n64x5 FILLER_259_343 ();
 b15zdnd11an1n64x5 FILLER_259_407 ();
 b15zdnd11an1n64x5 FILLER_259_471 ();
 b15zdnd11an1n32x5 FILLER_259_535 ();
 b15zdnd00an1n01x5 FILLER_259_567 ();
 b15zdnd11an1n08x5 FILLER_259_620 ();
 b15zdnd11an1n64x5 FILLER_259_631 ();
 b15zdnd11an1n32x5 FILLER_259_695 ();
 b15zdnd11an1n16x5 FILLER_259_727 ();
 b15zdnd11an1n08x5 FILLER_259_743 ();
 b15zdnd11an1n04x5 FILLER_259_751 ();
 b15zdnd00an1n02x5 FILLER_259_755 ();
 b15zdnd00an1n01x5 FILLER_259_757 ();
 b15zdnd11an1n64x5 FILLER_259_761 ();
 b15zdnd11an1n64x5 FILLER_259_825 ();
 b15zdnd11an1n64x5 FILLER_259_889 ();
 b15zdnd11an1n16x5 FILLER_259_953 ();
 b15zdnd11an1n04x5 FILLER_259_969 ();
 b15zdnd00an1n01x5 FILLER_259_973 ();
 b15zdnd11an1n64x5 FILLER_259_1026 ();
 b15zdnd11an1n64x5 FILLER_259_1090 ();
 b15zdnd11an1n64x5 FILLER_259_1154 ();
 b15zdnd11an1n32x5 FILLER_259_1218 ();
 b15zdnd11an1n04x5 FILLER_259_1250 ();
 b15zdnd00an1n02x5 FILLER_259_1254 ();
 b15zdnd00an1n01x5 FILLER_259_1256 ();
 b15zdnd11an1n04x5 FILLER_259_1260 ();
 b15zdnd11an1n64x5 FILLER_259_1267 ();
 b15zdnd11an1n16x5 FILLER_259_1331 ();
 b15zdnd00an1n02x5 FILLER_259_1347 ();
 b15zdnd11an1n64x5 FILLER_259_1358 ();
 b15zdnd11an1n64x5 FILLER_259_1422 ();
 b15zdnd11an1n16x5 FILLER_259_1486 ();
 b15zdnd11an1n08x5 FILLER_259_1502 ();
 b15zdnd11an1n04x5 FILLER_259_1510 ();
 b15zdnd11an1n04x5 FILLER_259_1517 ();
 b15zdnd11an1n64x5 FILLER_259_1524 ();
 b15zdnd11an1n32x5 FILLER_259_1588 ();
 b15zdnd11an1n08x5 FILLER_259_1620 ();
 b15zdnd11an1n04x5 FILLER_259_1628 ();
 b15zdnd00an1n02x5 FILLER_259_1632 ();
 b15zdnd00an1n01x5 FILLER_259_1634 ();
 b15zdnd11an1n64x5 FILLER_259_1687 ();
 b15zdnd11an1n32x5 FILLER_259_1751 ();
 b15zdnd11an1n08x5 FILLER_259_1783 ();
 b15zdnd00an1n02x5 FILLER_259_1791 ();
 b15zdnd00an1n01x5 FILLER_259_1793 ();
 b15zdnd11an1n64x5 FILLER_259_1803 ();
 b15zdnd11an1n64x5 FILLER_259_1867 ();
 b15zdnd11an1n64x5 FILLER_259_1931 ();
 b15zdnd11an1n32x5 FILLER_259_1995 ();
 b15zdnd00an1n02x5 FILLER_259_2027 ();
 b15zdnd00an1n01x5 FILLER_259_2029 ();
 b15zdnd11an1n64x5 FILLER_259_2061 ();
 b15zdnd11an1n08x5 FILLER_259_2125 ();
 b15zdnd11an1n04x5 FILLER_259_2133 ();
 b15zdnd11an1n64x5 FILLER_259_2179 ();
 b15zdnd11an1n32x5 FILLER_259_2243 ();
 b15zdnd11an1n08x5 FILLER_259_2275 ();
 b15zdnd00an1n01x5 FILLER_259_2283 ();
 b15zdnd11an1n32x5 FILLER_260_8 ();
 b15zdnd11an1n08x5 FILLER_260_40 ();
 b15zdnd11an1n64x5 FILLER_260_100 ();
 b15zdnd11an1n64x5 FILLER_260_164 ();
 b15zdnd11an1n64x5 FILLER_260_228 ();
 b15zdnd11an1n64x5 FILLER_260_292 ();
 b15zdnd11an1n64x5 FILLER_260_356 ();
 b15zdnd11an1n64x5 FILLER_260_420 ();
 b15zdnd11an1n64x5 FILLER_260_484 ();
 b15zdnd11an1n64x5 FILLER_260_548 ();
 b15zdnd11an1n64x5 FILLER_260_654 ();
 b15zdnd11an1n16x5 FILLER_260_726 ();
 b15zdnd11an1n64x5 FILLER_260_784 ();
 b15zdnd11an1n64x5 FILLER_260_848 ();
 b15zdnd11an1n32x5 FILLER_260_912 ();
 b15zdnd11an1n16x5 FILLER_260_944 ();
 b15zdnd11an1n08x5 FILLER_260_960 ();
 b15zdnd11an1n04x5 FILLER_260_971 ();
 b15zdnd11an1n08x5 FILLER_260_978 ();
 b15zdnd11an1n04x5 FILLER_260_986 ();
 b15zdnd00an1n01x5 FILLER_260_990 ();
 b15zdnd11an1n04x5 FILLER_260_994 ();
 b15zdnd11an1n64x5 FILLER_260_1001 ();
 b15zdnd11an1n64x5 FILLER_260_1065 ();
 b15zdnd11an1n64x5 FILLER_260_1129 ();
 b15zdnd11an1n64x5 FILLER_260_1193 ();
 b15zdnd11an1n64x5 FILLER_260_1257 ();
 b15zdnd11an1n64x5 FILLER_260_1321 ();
 b15zdnd11an1n64x5 FILLER_260_1385 ();
 b15zdnd11an1n64x5 FILLER_260_1449 ();
 b15zdnd11an1n64x5 FILLER_260_1513 ();
 b15zdnd11an1n64x5 FILLER_260_1577 ();
 b15zdnd11an1n08x5 FILLER_260_1641 ();
 b15zdnd11an1n04x5 FILLER_260_1649 ();
 b15zdnd00an1n01x5 FILLER_260_1653 ();
 b15zdnd11an1n04x5 FILLER_260_1657 ();
 b15zdnd11an1n16x5 FILLER_260_1664 ();
 b15zdnd00an1n02x5 FILLER_260_1680 ();
 b15zdnd00an1n01x5 FILLER_260_1682 ();
 b15zdnd11an1n64x5 FILLER_260_1703 ();
 b15zdnd11an1n64x5 FILLER_260_1767 ();
 b15zdnd11an1n64x5 FILLER_260_1831 ();
 b15zdnd11an1n64x5 FILLER_260_1895 ();
 b15zdnd11an1n64x5 FILLER_260_1959 ();
 b15zdnd11an1n64x5 FILLER_260_2023 ();
 b15zdnd11an1n64x5 FILLER_260_2087 ();
 b15zdnd00an1n02x5 FILLER_260_2151 ();
 b15zdnd00an1n01x5 FILLER_260_2153 ();
 b15zdnd11an1n64x5 FILLER_260_2162 ();
 b15zdnd11an1n32x5 FILLER_260_2226 ();
 b15zdnd11an1n16x5 FILLER_260_2258 ();
 b15zdnd00an1n02x5 FILLER_260_2274 ();
 b15zdnd11an1n16x5 FILLER_261_0 ();
 b15zdnd11an1n08x5 FILLER_261_16 ();
 b15zdnd00an1n02x5 FILLER_261_24 ();
 b15zdnd11an1n16x5 FILLER_261_32 ();
 b15zdnd11an1n08x5 FILLER_261_48 ();
 b15zdnd11an1n04x5 FILLER_261_56 ();
 b15zdnd00an1n02x5 FILLER_261_60 ();
 b15zdnd11an1n64x5 FILLER_261_89 ();
 b15zdnd11an1n64x5 FILLER_261_153 ();
 b15zdnd11an1n64x5 FILLER_261_217 ();
 b15zdnd11an1n64x5 FILLER_261_281 ();
 b15zdnd11an1n64x5 FILLER_261_345 ();
 b15zdnd11an1n64x5 FILLER_261_409 ();
 b15zdnd11an1n64x5 FILLER_261_473 ();
 b15zdnd11an1n64x5 FILLER_261_537 ();
 b15zdnd11an1n64x5 FILLER_261_653 ();
 b15zdnd11an1n08x5 FILLER_261_717 ();
 b15zdnd11an1n04x5 FILLER_261_725 ();
 b15zdnd00an1n02x5 FILLER_261_729 ();
 b15zdnd11an1n64x5 FILLER_261_783 ();
 b15zdnd11an1n64x5 FILLER_261_847 ();
 b15zdnd11an1n32x5 FILLER_261_911 ();
 b15zdnd11an1n16x5 FILLER_261_943 ();
 b15zdnd11an1n08x5 FILLER_261_959 ();
 b15zdnd11an1n04x5 FILLER_261_967 ();
 b15zdnd00an1n01x5 FILLER_261_971 ();
 b15zdnd11an1n16x5 FILLER_261_975 ();
 b15zdnd11an1n04x5 FILLER_261_991 ();
 b15zdnd11an1n64x5 FILLER_261_998 ();
 b15zdnd11an1n64x5 FILLER_261_1062 ();
 b15zdnd11an1n64x5 FILLER_261_1126 ();
 b15zdnd11an1n64x5 FILLER_261_1190 ();
 b15zdnd11an1n64x5 FILLER_261_1254 ();
 b15zdnd11an1n64x5 FILLER_261_1318 ();
 b15zdnd11an1n64x5 FILLER_261_1382 ();
 b15zdnd11an1n64x5 FILLER_261_1446 ();
 b15zdnd11an1n64x5 FILLER_261_1510 ();
 b15zdnd11an1n64x5 FILLER_261_1574 ();
 b15zdnd00an1n01x5 FILLER_261_1638 ();
 b15zdnd11an1n04x5 FILLER_261_1659 ();
 b15zdnd11an1n16x5 FILLER_261_1666 ();
 b15zdnd11an1n08x5 FILLER_261_1682 ();
 b15zdnd11an1n04x5 FILLER_261_1690 ();
 b15zdnd11an1n64x5 FILLER_261_1714 ();
 b15zdnd11an1n64x5 FILLER_261_1778 ();
 b15zdnd11an1n64x5 FILLER_261_1842 ();
 b15zdnd11an1n64x5 FILLER_261_1906 ();
 b15zdnd11an1n64x5 FILLER_261_1970 ();
 b15zdnd11an1n32x5 FILLER_261_2034 ();
 b15zdnd11an1n16x5 FILLER_261_2066 ();
 b15zdnd00an1n02x5 FILLER_261_2082 ();
 b15zdnd11an1n64x5 FILLER_261_2099 ();
 b15zdnd11an1n16x5 FILLER_261_2163 ();
 b15zdnd11an1n08x5 FILLER_261_2179 ();
 b15zdnd11an1n04x5 FILLER_261_2187 ();
 b15zdnd11an1n32x5 FILLER_261_2233 ();
 b15zdnd11an1n16x5 FILLER_261_2265 ();
 b15zdnd00an1n02x5 FILLER_261_2281 ();
 b15zdnd00an1n01x5 FILLER_261_2283 ();
 b15zdnd11an1n32x5 FILLER_262_8 ();
 b15zdnd11an1n16x5 FILLER_262_40 ();
 b15zdnd00an1n01x5 FILLER_262_56 ();
 b15zdnd11an1n64x5 FILLER_262_109 ();
 b15zdnd11an1n64x5 FILLER_262_173 ();
 b15zdnd11an1n64x5 FILLER_262_237 ();
 b15zdnd11an1n64x5 FILLER_262_301 ();
 b15zdnd11an1n64x5 FILLER_262_365 ();
 b15zdnd11an1n64x5 FILLER_262_429 ();
 b15zdnd11an1n64x5 FILLER_262_493 ();
 b15zdnd11an1n32x5 FILLER_262_557 ();
 b15zdnd11an1n16x5 FILLER_262_589 ();
 b15zdnd11an1n08x5 FILLER_262_605 ();
 b15zdnd11an1n04x5 FILLER_262_613 ();
 b15zdnd00an1n02x5 FILLER_262_617 ();
 b15zdnd11an1n04x5 FILLER_262_622 ();
 b15zdnd11an1n08x5 FILLER_262_629 ();
 b15zdnd11an1n04x5 FILLER_262_637 ();
 b15zdnd11an1n32x5 FILLER_262_683 ();
 b15zdnd00an1n02x5 FILLER_262_715 ();
 b15zdnd00an1n01x5 FILLER_262_717 ();
 b15zdnd11an1n16x5 FILLER_262_726 ();
 b15zdnd11an1n08x5 FILLER_262_742 ();
 b15zdnd11an1n04x5 FILLER_262_750 ();
 b15zdnd00an1n02x5 FILLER_262_754 ();
 b15zdnd11an1n08x5 FILLER_262_759 ();
 b15zdnd11an1n04x5 FILLER_262_767 ();
 b15zdnd11an1n32x5 FILLER_262_813 ();
 b15zdnd11an1n16x5 FILLER_262_845 ();
 b15zdnd11an1n08x5 FILLER_262_861 ();
 b15zdnd00an1n02x5 FILLER_262_869 ();
 b15zdnd11an1n04x5 FILLER_262_903 ();
 b15zdnd11an1n64x5 FILLER_262_910 ();
 b15zdnd11an1n64x5 FILLER_262_974 ();
 b15zdnd11an1n64x5 FILLER_262_1038 ();
 b15zdnd11an1n64x5 FILLER_262_1102 ();
 b15zdnd11an1n64x5 FILLER_262_1166 ();
 b15zdnd11an1n64x5 FILLER_262_1230 ();
 b15zdnd11an1n64x5 FILLER_262_1294 ();
 b15zdnd11an1n64x5 FILLER_262_1358 ();
 b15zdnd11an1n64x5 FILLER_262_1422 ();
 b15zdnd11an1n64x5 FILLER_262_1486 ();
 b15zdnd11an1n64x5 FILLER_262_1550 ();
 b15zdnd11an1n64x5 FILLER_262_1614 ();
 b15zdnd11an1n64x5 FILLER_262_1678 ();
 b15zdnd11an1n64x5 FILLER_262_1742 ();
 b15zdnd11an1n64x5 FILLER_262_1806 ();
 b15zdnd11an1n64x5 FILLER_262_1870 ();
 b15zdnd11an1n64x5 FILLER_262_1934 ();
 b15zdnd11an1n16x5 FILLER_262_1998 ();
 b15zdnd00an1n01x5 FILLER_262_2014 ();
 b15zdnd11an1n04x5 FILLER_262_2021 ();
 b15zdnd11an1n64x5 FILLER_262_2049 ();
 b15zdnd11an1n32x5 FILLER_262_2113 ();
 b15zdnd11an1n08x5 FILLER_262_2145 ();
 b15zdnd00an1n01x5 FILLER_262_2153 ();
 b15zdnd11an1n32x5 FILLER_262_2162 ();
 b15zdnd11an1n16x5 FILLER_262_2194 ();
 b15zdnd11an1n08x5 FILLER_262_2210 ();
 b15zdnd11an1n04x5 FILLER_262_2218 ();
 b15zdnd00an1n02x5 FILLER_262_2222 ();
 b15zdnd11an1n32x5 FILLER_262_2242 ();
 b15zdnd00an1n02x5 FILLER_262_2274 ();
 b15zdnd11an1n32x5 FILLER_263_0 ();
 b15zdnd11an1n16x5 FILLER_263_32 ();
 b15zdnd11an1n08x5 FILLER_263_48 ();
 b15zdnd11an1n04x5 FILLER_263_56 ();
 b15zdnd00an1n01x5 FILLER_263_60 ();
 b15zdnd11an1n08x5 FILLER_263_64 ();
 b15zdnd11an1n04x5 FILLER_263_72 ();
 b15zdnd00an1n02x5 FILLER_263_76 ();
 b15zdnd00an1n01x5 FILLER_263_78 ();
 b15zdnd11an1n04x5 FILLER_263_82 ();
 b15zdnd11an1n64x5 FILLER_263_89 ();
 b15zdnd11an1n64x5 FILLER_263_153 ();
 b15zdnd11an1n16x5 FILLER_263_217 ();
 b15zdnd11an1n04x5 FILLER_263_233 ();
 b15zdnd00an1n01x5 FILLER_263_237 ();
 b15zdnd11an1n64x5 FILLER_263_247 ();
 b15zdnd11an1n32x5 FILLER_263_311 ();
 b15zdnd00an1n02x5 FILLER_263_343 ();
 b15zdnd00an1n01x5 FILLER_263_345 ();
 b15zdnd11an1n64x5 FILLER_263_388 ();
 b15zdnd11an1n64x5 FILLER_263_452 ();
 b15zdnd11an1n64x5 FILLER_263_516 ();
 b15zdnd11an1n64x5 FILLER_263_580 ();
 b15zdnd11an1n64x5 FILLER_263_644 ();
 b15zdnd11an1n32x5 FILLER_263_708 ();
 b15zdnd11an1n16x5 FILLER_263_740 ();
 b15zdnd11an1n64x5 FILLER_263_759 ();
 b15zdnd11an1n64x5 FILLER_263_823 ();
 b15zdnd11an1n16x5 FILLER_263_887 ();
 b15zdnd00an1n02x5 FILLER_263_903 ();
 b15zdnd11an1n64x5 FILLER_263_908 ();
 b15zdnd11an1n64x5 FILLER_263_972 ();
 b15zdnd11an1n64x5 FILLER_263_1036 ();
 b15zdnd11an1n64x5 FILLER_263_1100 ();
 b15zdnd11an1n64x5 FILLER_263_1164 ();
 b15zdnd11an1n64x5 FILLER_263_1228 ();
 b15zdnd11an1n32x5 FILLER_263_1292 ();
 b15zdnd11an1n08x5 FILLER_263_1324 ();
 b15zdnd00an1n02x5 FILLER_263_1332 ();
 b15zdnd00an1n01x5 FILLER_263_1334 ();
 b15zdnd11an1n64x5 FILLER_263_1344 ();
 b15zdnd11an1n64x5 FILLER_263_1408 ();
 b15zdnd11an1n64x5 FILLER_263_1472 ();
 b15zdnd11an1n64x5 FILLER_263_1536 ();
 b15zdnd11an1n64x5 FILLER_263_1600 ();
 b15zdnd11an1n64x5 FILLER_263_1664 ();
 b15zdnd11an1n64x5 FILLER_263_1728 ();
 b15zdnd11an1n64x5 FILLER_263_1792 ();
 b15zdnd11an1n16x5 FILLER_263_1856 ();
 b15zdnd11an1n08x5 FILLER_263_1872 ();
 b15zdnd11an1n04x5 FILLER_263_1880 ();
 b15zdnd00an1n02x5 FILLER_263_1884 ();
 b15zdnd11an1n64x5 FILLER_263_1910 ();
 b15zdnd11an1n64x5 FILLER_263_1974 ();
 b15zdnd11an1n32x5 FILLER_263_2038 ();
 b15zdnd11an1n08x5 FILLER_263_2070 ();
 b15zdnd11an1n04x5 FILLER_263_2078 ();
 b15zdnd00an1n02x5 FILLER_263_2082 ();
 b15zdnd11an1n64x5 FILLER_263_2099 ();
 b15zdnd11an1n16x5 FILLER_263_2163 ();
 b15zdnd00an1n02x5 FILLER_263_2179 ();
 b15zdnd11an1n64x5 FILLER_263_2193 ();
 b15zdnd11an1n16x5 FILLER_263_2257 ();
 b15zdnd11an1n08x5 FILLER_263_2273 ();
 b15zdnd00an1n02x5 FILLER_263_2281 ();
 b15zdnd00an1n01x5 FILLER_263_2283 ();
 b15zdnd11an1n64x5 FILLER_264_8 ();
 b15zdnd11an1n08x5 FILLER_264_72 ();
 b15zdnd11an1n64x5 FILLER_264_83 ();
 b15zdnd11an1n64x5 FILLER_264_147 ();
 b15zdnd11an1n04x5 FILLER_264_211 ();
 b15zdnd00an1n02x5 FILLER_264_215 ();
 b15zdnd11an1n04x5 FILLER_264_249 ();
 b15zdnd11an1n32x5 FILLER_264_256 ();
 b15zdnd11an1n04x5 FILLER_264_288 ();
 b15zdnd00an1n02x5 FILLER_264_292 ();
 b15zdnd11an1n64x5 FILLER_264_303 ();
 b15zdnd11an1n64x5 FILLER_264_367 ();
 b15zdnd11an1n64x5 FILLER_264_431 ();
 b15zdnd11an1n64x5 FILLER_264_495 ();
 b15zdnd11an1n64x5 FILLER_264_559 ();
 b15zdnd11an1n32x5 FILLER_264_623 ();
 b15zdnd11an1n16x5 FILLER_264_655 ();
 b15zdnd11an1n08x5 FILLER_264_671 ();
 b15zdnd11an1n04x5 FILLER_264_679 ();
 b15zdnd00an1n02x5 FILLER_264_683 ();
 b15zdnd00an1n01x5 FILLER_264_685 ();
 b15zdnd11an1n04x5 FILLER_264_701 ();
 b15zdnd00an1n02x5 FILLER_264_716 ();
 b15zdnd11an1n64x5 FILLER_264_726 ();
 b15zdnd11an1n64x5 FILLER_264_790 ();
 b15zdnd11an1n64x5 FILLER_264_854 ();
 b15zdnd11an1n32x5 FILLER_264_918 ();
 b15zdnd11an1n08x5 FILLER_264_950 ();
 b15zdnd00an1n02x5 FILLER_264_958 ();
 b15zdnd11an1n64x5 FILLER_264_969 ();
 b15zdnd11an1n64x5 FILLER_264_1033 ();
 b15zdnd11an1n64x5 FILLER_264_1097 ();
 b15zdnd11an1n64x5 FILLER_264_1161 ();
 b15zdnd11an1n64x5 FILLER_264_1225 ();
 b15zdnd11an1n04x5 FILLER_264_1289 ();
 b15zdnd00an1n01x5 FILLER_264_1293 ();
 b15zdnd11an1n64x5 FILLER_264_1303 ();
 b15zdnd11an1n64x5 FILLER_264_1367 ();
 b15zdnd11an1n64x5 FILLER_264_1431 ();
 b15zdnd11an1n64x5 FILLER_264_1495 ();
 b15zdnd11an1n64x5 FILLER_264_1559 ();
 b15zdnd11an1n64x5 FILLER_264_1623 ();
 b15zdnd11an1n64x5 FILLER_264_1687 ();
 b15zdnd11an1n64x5 FILLER_264_1751 ();
 b15zdnd11an1n64x5 FILLER_264_1815 ();
 b15zdnd11an1n64x5 FILLER_264_1879 ();
 b15zdnd11an1n64x5 FILLER_264_1943 ();
 b15zdnd11an1n32x5 FILLER_264_2007 ();
 b15zdnd11an1n16x5 FILLER_264_2039 ();
 b15zdnd11an1n64x5 FILLER_264_2065 ();
 b15zdnd11an1n16x5 FILLER_264_2129 ();
 b15zdnd11an1n08x5 FILLER_264_2145 ();
 b15zdnd00an1n01x5 FILLER_264_2153 ();
 b15zdnd11an1n64x5 FILLER_264_2162 ();
 b15zdnd11an1n32x5 FILLER_264_2226 ();
 b15zdnd11an1n16x5 FILLER_264_2258 ();
 b15zdnd00an1n02x5 FILLER_264_2274 ();
 b15zdnd11an1n64x5 FILLER_265_0 ();
 b15zdnd11an1n64x5 FILLER_265_64 ();
 b15zdnd11an1n64x5 FILLER_265_128 ();
 b15zdnd11an1n16x5 FILLER_265_192 ();
 b15zdnd11an1n08x5 FILLER_265_208 ();
 b15zdnd11an1n04x5 FILLER_265_216 ();
 b15zdnd00an1n02x5 FILLER_265_220 ();
 b15zdnd00an1n01x5 FILLER_265_222 ();
 b15zdnd11an1n64x5 FILLER_265_265 ();
 b15zdnd11an1n08x5 FILLER_265_329 ();
 b15zdnd11an1n04x5 FILLER_265_337 ();
 b15zdnd11an1n64x5 FILLER_265_344 ();
 b15zdnd11an1n64x5 FILLER_265_408 ();
 b15zdnd11an1n64x5 FILLER_265_472 ();
 b15zdnd11an1n64x5 FILLER_265_536 ();
 b15zdnd11an1n64x5 FILLER_265_600 ();
 b15zdnd11an1n64x5 FILLER_265_664 ();
 b15zdnd11an1n64x5 FILLER_265_728 ();
 b15zdnd11an1n64x5 FILLER_265_792 ();
 b15zdnd11an1n16x5 FILLER_265_856 ();
 b15zdnd11an1n64x5 FILLER_265_875 ();
 b15zdnd11an1n64x5 FILLER_265_939 ();
 b15zdnd11an1n64x5 FILLER_265_1003 ();
 b15zdnd11an1n64x5 FILLER_265_1067 ();
 b15zdnd11an1n64x5 FILLER_265_1131 ();
 b15zdnd11an1n64x5 FILLER_265_1195 ();
 b15zdnd11an1n64x5 FILLER_265_1259 ();
 b15zdnd11an1n64x5 FILLER_265_1323 ();
 b15zdnd11an1n64x5 FILLER_265_1387 ();
 b15zdnd11an1n64x5 FILLER_265_1451 ();
 b15zdnd11an1n64x5 FILLER_265_1515 ();
 b15zdnd11an1n64x5 FILLER_265_1579 ();
 b15zdnd11an1n64x5 FILLER_265_1643 ();
 b15zdnd11an1n64x5 FILLER_265_1707 ();
 b15zdnd11an1n64x5 FILLER_265_1771 ();
 b15zdnd11an1n64x5 FILLER_265_1835 ();
 b15zdnd11an1n64x5 FILLER_265_1899 ();
 b15zdnd11an1n64x5 FILLER_265_1963 ();
 b15zdnd11an1n16x5 FILLER_265_2027 ();
 b15zdnd11an1n08x5 FILLER_265_2043 ();
 b15zdnd00an1n02x5 FILLER_265_2051 ();
 b15zdnd00an1n01x5 FILLER_265_2053 ();
 b15zdnd11an1n64x5 FILLER_265_2079 ();
 b15zdnd11an1n64x5 FILLER_265_2143 ();
 b15zdnd11an1n64x5 FILLER_265_2207 ();
 b15zdnd11an1n08x5 FILLER_265_2271 ();
 b15zdnd11an1n04x5 FILLER_265_2279 ();
 b15zdnd00an1n01x5 FILLER_265_2283 ();
 b15zdnd11an1n64x5 FILLER_266_8 ();
 b15zdnd11an1n64x5 FILLER_266_72 ();
 b15zdnd11an1n64x5 FILLER_266_136 ();
 b15zdnd11an1n08x5 FILLER_266_200 ();
 b15zdnd11an1n08x5 FILLER_266_260 ();
 b15zdnd11an1n04x5 FILLER_266_275 ();
 b15zdnd11an1n16x5 FILLER_266_311 ();
 b15zdnd00an1n02x5 FILLER_266_327 ();
 b15zdnd11an1n04x5 FILLER_266_332 ();
 b15zdnd11an1n64x5 FILLER_266_378 ();
 b15zdnd11an1n64x5 FILLER_266_442 ();
 b15zdnd11an1n08x5 FILLER_266_506 ();
 b15zdnd11an1n04x5 FILLER_266_514 ();
 b15zdnd11an1n64x5 FILLER_266_560 ();
 b15zdnd11an1n64x5 FILLER_266_624 ();
 b15zdnd11an1n16x5 FILLER_266_688 ();
 b15zdnd11an1n08x5 FILLER_266_704 ();
 b15zdnd11an1n04x5 FILLER_266_712 ();
 b15zdnd00an1n02x5 FILLER_266_716 ();
 b15zdnd11an1n64x5 FILLER_266_726 ();
 b15zdnd11an1n64x5 FILLER_266_790 ();
 b15zdnd00an1n02x5 FILLER_266_854 ();
 b15zdnd11an1n64x5 FILLER_266_898 ();
 b15zdnd11an1n64x5 FILLER_266_962 ();
 b15zdnd11an1n64x5 FILLER_266_1026 ();
 b15zdnd11an1n64x5 FILLER_266_1090 ();
 b15zdnd11an1n64x5 FILLER_266_1154 ();
 b15zdnd11an1n64x5 FILLER_266_1218 ();
 b15zdnd11an1n64x5 FILLER_266_1282 ();
 b15zdnd11an1n64x5 FILLER_266_1346 ();
 b15zdnd11an1n64x5 FILLER_266_1410 ();
 b15zdnd11an1n64x5 FILLER_266_1474 ();
 b15zdnd11an1n64x5 FILLER_266_1538 ();
 b15zdnd11an1n64x5 FILLER_266_1602 ();
 b15zdnd11an1n64x5 FILLER_266_1666 ();
 b15zdnd11an1n64x5 FILLER_266_1730 ();
 b15zdnd11an1n64x5 FILLER_266_1794 ();
 b15zdnd11an1n64x5 FILLER_266_1858 ();
 b15zdnd11an1n64x5 FILLER_266_1922 ();
 b15zdnd11an1n32x5 FILLER_266_1986 ();
 b15zdnd11an1n08x5 FILLER_266_2018 ();
 b15zdnd11an1n04x5 FILLER_266_2026 ();
 b15zdnd00an1n01x5 FILLER_266_2030 ();
 b15zdnd11an1n64x5 FILLER_266_2056 ();
 b15zdnd11an1n32x5 FILLER_266_2120 ();
 b15zdnd00an1n02x5 FILLER_266_2152 ();
 b15zdnd11an1n64x5 FILLER_266_2162 ();
 b15zdnd11an1n32x5 FILLER_266_2226 ();
 b15zdnd11an1n16x5 FILLER_266_2258 ();
 b15zdnd00an1n02x5 FILLER_266_2274 ();
 b15zdnd11an1n64x5 FILLER_267_0 ();
 b15zdnd11an1n64x5 FILLER_267_64 ();
 b15zdnd11an1n64x5 FILLER_267_128 ();
 b15zdnd11an1n16x5 FILLER_267_192 ();
 b15zdnd11an1n08x5 FILLER_267_208 ();
 b15zdnd11an1n04x5 FILLER_267_216 ();
 b15zdnd00an1n01x5 FILLER_267_220 ();
 b15zdnd11an1n32x5 FILLER_267_248 ();
 b15zdnd11an1n08x5 FILLER_267_280 ();
 b15zdnd00an1n01x5 FILLER_267_288 ();
 b15zdnd11an1n04x5 FILLER_267_298 ();
 b15zdnd11an1n04x5 FILLER_267_305 ();
 b15zdnd11an1n04x5 FILLER_267_312 ();
 b15zdnd11an1n04x5 FILLER_267_368 ();
 b15zdnd11an1n64x5 FILLER_267_379 ();
 b15zdnd11an1n64x5 FILLER_267_443 ();
 b15zdnd11an1n64x5 FILLER_267_507 ();
 b15zdnd11an1n64x5 FILLER_267_571 ();
 b15zdnd11an1n64x5 FILLER_267_635 ();
 b15zdnd11an1n64x5 FILLER_267_699 ();
 b15zdnd11an1n64x5 FILLER_267_763 ();
 b15zdnd11an1n16x5 FILLER_267_827 ();
 b15zdnd00an1n02x5 FILLER_267_843 ();
 b15zdnd11an1n64x5 FILLER_267_897 ();
 b15zdnd11an1n64x5 FILLER_267_961 ();
 b15zdnd11an1n64x5 FILLER_267_1025 ();
 b15zdnd11an1n64x5 FILLER_267_1089 ();
 b15zdnd11an1n64x5 FILLER_267_1153 ();
 b15zdnd11an1n64x5 FILLER_267_1217 ();
 b15zdnd11an1n64x5 FILLER_267_1281 ();
 b15zdnd11an1n32x5 FILLER_267_1345 ();
 b15zdnd11an1n16x5 FILLER_267_1377 ();
 b15zdnd11an1n04x5 FILLER_267_1393 ();
 b15zdnd00an1n01x5 FILLER_267_1397 ();
 b15zdnd11an1n04x5 FILLER_267_1401 ();
 b15zdnd11an1n64x5 FILLER_267_1408 ();
 b15zdnd11an1n64x5 FILLER_267_1472 ();
 b15zdnd11an1n64x5 FILLER_267_1536 ();
 b15zdnd11an1n64x5 FILLER_267_1600 ();
 b15zdnd11an1n64x5 FILLER_267_1664 ();
 b15zdnd11an1n32x5 FILLER_267_1728 ();
 b15zdnd00an1n02x5 FILLER_267_1760 ();
 b15zdnd11an1n08x5 FILLER_267_1789 ();
 b15zdnd00an1n01x5 FILLER_267_1797 ();
 b15zdnd11an1n64x5 FILLER_267_1801 ();
 b15zdnd11an1n64x5 FILLER_267_1865 ();
 b15zdnd11an1n64x5 FILLER_267_1929 ();
 b15zdnd11an1n64x5 FILLER_267_1993 ();
 b15zdnd11an1n64x5 FILLER_267_2057 ();
 b15zdnd11an1n64x5 FILLER_267_2121 ();
 b15zdnd11an1n32x5 FILLER_267_2185 ();
 b15zdnd11an1n32x5 FILLER_267_2232 ();
 b15zdnd11an1n16x5 FILLER_267_2264 ();
 b15zdnd11an1n04x5 FILLER_267_2280 ();
 b15zdnd11an1n32x5 FILLER_268_8 ();
 b15zdnd11an1n16x5 FILLER_268_40 ();
 b15zdnd11an1n08x5 FILLER_268_56 ();
 b15zdnd11an1n04x5 FILLER_268_64 ();
 b15zdnd00an1n02x5 FILLER_268_68 ();
 b15zdnd00an1n01x5 FILLER_268_70 ();
 b15zdnd11an1n04x5 FILLER_268_80 ();
 b15zdnd00an1n01x5 FILLER_268_84 ();
 b15zdnd11an1n32x5 FILLER_268_94 ();
 b15zdnd11an1n16x5 FILLER_268_126 ();
 b15zdnd11an1n08x5 FILLER_268_142 ();
 b15zdnd00an1n02x5 FILLER_268_150 ();
 b15zdnd11an1n16x5 FILLER_268_194 ();
 b15zdnd11an1n08x5 FILLER_268_210 ();
 b15zdnd00an1n02x5 FILLER_268_218 ();
 b15zdnd00an1n01x5 FILLER_268_220 ();
 b15zdnd11an1n04x5 FILLER_268_224 ();
 b15zdnd11an1n04x5 FILLER_268_231 ();
 b15zdnd11an1n08x5 FILLER_268_238 ();
 b15zdnd11an1n64x5 FILLER_268_249 ();
 b15zdnd11an1n04x5 FILLER_268_313 ();
 b15zdnd11an1n64x5 FILLER_268_369 ();
 b15zdnd11an1n64x5 FILLER_268_433 ();
 b15zdnd11an1n64x5 FILLER_268_497 ();
 b15zdnd11an1n16x5 FILLER_268_561 ();
 b15zdnd11an1n04x5 FILLER_268_577 ();
 b15zdnd00an1n02x5 FILLER_268_581 ();
 b15zdnd11an1n64x5 FILLER_268_625 ();
 b15zdnd11an1n16x5 FILLER_268_689 ();
 b15zdnd11an1n08x5 FILLER_268_705 ();
 b15zdnd11an1n04x5 FILLER_268_713 ();
 b15zdnd00an1n01x5 FILLER_268_717 ();
 b15zdnd11an1n64x5 FILLER_268_726 ();
 b15zdnd11an1n64x5 FILLER_268_790 ();
 b15zdnd11an1n08x5 FILLER_268_854 ();
 b15zdnd00an1n01x5 FILLER_268_862 ();
 b15zdnd11an1n04x5 FILLER_268_866 ();
 b15zdnd11an1n08x5 FILLER_268_873 ();
 b15zdnd11an1n04x5 FILLER_268_881 ();
 b15zdnd11an1n64x5 FILLER_268_927 ();
 b15zdnd11an1n64x5 FILLER_268_991 ();
 b15zdnd11an1n16x5 FILLER_268_1055 ();
 b15zdnd11an1n08x5 FILLER_268_1071 ();
 b15zdnd00an1n02x5 FILLER_268_1079 ();
 b15zdnd00an1n01x5 FILLER_268_1081 ();
 b15zdnd11an1n04x5 FILLER_268_1109 ();
 b15zdnd00an1n02x5 FILLER_268_1113 ();
 b15zdnd11an1n64x5 FILLER_268_1118 ();
 b15zdnd11an1n64x5 FILLER_268_1182 ();
 b15zdnd11an1n64x5 FILLER_268_1246 ();
 b15zdnd11an1n64x5 FILLER_268_1310 ();
 b15zdnd11an1n04x5 FILLER_268_1374 ();
 b15zdnd00an1n02x5 FILLER_268_1378 ();
 b15zdnd11an1n32x5 FILLER_268_1432 ();
 b15zdnd11an1n08x5 FILLER_268_1464 ();
 b15zdnd00an1n02x5 FILLER_268_1472 ();
 b15zdnd00an1n01x5 FILLER_268_1474 ();
 b15zdnd11an1n64x5 FILLER_268_1495 ();
 b15zdnd11an1n64x5 FILLER_268_1559 ();
 b15zdnd11an1n32x5 FILLER_268_1623 ();
 b15zdnd11an1n08x5 FILLER_268_1655 ();
 b15zdnd00an1n02x5 FILLER_268_1663 ();
 b15zdnd11an1n64x5 FILLER_268_1689 ();
 b15zdnd11an1n08x5 FILLER_268_1753 ();
 b15zdnd00an1n01x5 FILLER_268_1761 ();
 b15zdnd11an1n08x5 FILLER_268_1765 ();
 b15zdnd11an1n16x5 FILLER_268_1825 ();
 b15zdnd11an1n04x5 FILLER_268_1841 ();
 b15zdnd00an1n01x5 FILLER_268_1845 ();
 b15zdnd11an1n04x5 FILLER_268_1849 ();
 b15zdnd11an1n64x5 FILLER_268_1856 ();
 b15zdnd11an1n64x5 FILLER_268_1920 ();
 b15zdnd11an1n64x5 FILLER_268_1984 ();
 b15zdnd11an1n64x5 FILLER_268_2048 ();
 b15zdnd11an1n32x5 FILLER_268_2112 ();
 b15zdnd11an1n08x5 FILLER_268_2144 ();
 b15zdnd00an1n02x5 FILLER_268_2152 ();
 b15zdnd11an1n64x5 FILLER_268_2162 ();
 b15zdnd11an1n32x5 FILLER_268_2226 ();
 b15zdnd11an1n16x5 FILLER_268_2258 ();
 b15zdnd00an1n02x5 FILLER_268_2274 ();
 b15zdnd11an1n64x5 FILLER_269_0 ();
 b15zdnd11an1n64x5 FILLER_269_64 ();
 b15zdnd11an1n64x5 FILLER_269_128 ();
 b15zdnd11an1n08x5 FILLER_269_192 ();
 b15zdnd11an1n04x5 FILLER_269_200 ();
 b15zdnd00an1n02x5 FILLER_269_204 ();
 b15zdnd00an1n01x5 FILLER_269_206 ();
 b15zdnd11an1n64x5 FILLER_269_249 ();
 b15zdnd11an1n16x5 FILLER_269_313 ();
 b15zdnd11an1n04x5 FILLER_269_329 ();
 b15zdnd00an1n02x5 FILLER_269_333 ();
 b15zdnd00an1n01x5 FILLER_269_335 ();
 b15zdnd11an1n64x5 FILLER_269_378 ();
 b15zdnd11an1n64x5 FILLER_269_442 ();
 b15zdnd11an1n64x5 FILLER_269_506 ();
 b15zdnd11an1n64x5 FILLER_269_570 ();
 b15zdnd11an1n32x5 FILLER_269_634 ();
 b15zdnd11an1n16x5 FILLER_269_666 ();
 b15zdnd11an1n08x5 FILLER_269_682 ();
 b15zdnd11an1n04x5 FILLER_269_690 ();
 b15zdnd00an1n02x5 FILLER_269_694 ();
 b15zdnd00an1n01x5 FILLER_269_696 ();
 b15zdnd11an1n64x5 FILLER_269_739 ();
 b15zdnd11an1n64x5 FILLER_269_803 ();
 b15zdnd11an1n64x5 FILLER_269_867 ();
 b15zdnd11an1n64x5 FILLER_269_931 ();
 b15zdnd11an1n64x5 FILLER_269_995 ();
 b15zdnd11an1n04x5 FILLER_269_1059 ();
 b15zdnd11an1n16x5 FILLER_269_1094 ();
 b15zdnd00an1n02x5 FILLER_269_1110 ();
 b15zdnd00an1n01x5 FILLER_269_1112 ();
 b15zdnd11an1n04x5 FILLER_269_1116 ();
 b15zdnd00an1n02x5 FILLER_269_1120 ();
 b15zdnd00an1n01x5 FILLER_269_1122 ();
 b15zdnd11an1n08x5 FILLER_269_1126 ();
 b15zdnd00an1n02x5 FILLER_269_1134 ();
 b15zdnd11an1n64x5 FILLER_269_1147 ();
 b15zdnd11an1n64x5 FILLER_269_1211 ();
 b15zdnd11an1n64x5 FILLER_269_1275 ();
 b15zdnd11an1n64x5 FILLER_269_1339 ();
 b15zdnd00an1n02x5 FILLER_269_1403 ();
 b15zdnd11an1n64x5 FILLER_269_1408 ();
 b15zdnd11an1n16x5 FILLER_269_1472 ();
 b15zdnd00an1n02x5 FILLER_269_1488 ();
 b15zdnd11an1n64x5 FILLER_269_1510 ();
 b15zdnd11an1n64x5 FILLER_269_1574 ();
 b15zdnd11an1n64x5 FILLER_269_1638 ();
 b15zdnd11an1n64x5 FILLER_269_1702 ();
 b15zdnd11an1n04x5 FILLER_269_1766 ();
 b15zdnd00an1n01x5 FILLER_269_1770 ();
 b15zdnd11an1n04x5 FILLER_269_1823 ();
 b15zdnd11an1n64x5 FILLER_269_1879 ();
 b15zdnd11an1n64x5 FILLER_269_1943 ();
 b15zdnd11an1n64x5 FILLER_269_2007 ();
 b15zdnd11an1n64x5 FILLER_269_2071 ();
 b15zdnd11an1n64x5 FILLER_269_2135 ();
 b15zdnd11an1n04x5 FILLER_269_2199 ();
 b15zdnd00an1n02x5 FILLER_269_2203 ();
 b15zdnd00an1n01x5 FILLER_269_2205 ();
 b15zdnd11an1n64x5 FILLER_269_2215 ();
 b15zdnd11an1n04x5 FILLER_269_2279 ();
 b15zdnd00an1n01x5 FILLER_269_2283 ();
 b15zdnd11an1n64x5 FILLER_270_8 ();
 b15zdnd11an1n64x5 FILLER_270_72 ();
 b15zdnd11an1n64x5 FILLER_270_136 ();
 b15zdnd11an1n32x5 FILLER_270_200 ();
 b15zdnd00an1n01x5 FILLER_270_232 ();
 b15zdnd11an1n64x5 FILLER_270_236 ();
 b15zdnd11an1n32x5 FILLER_270_300 ();
 b15zdnd11an1n04x5 FILLER_270_332 ();
 b15zdnd11an1n04x5 FILLER_270_339 ();
 b15zdnd11an1n04x5 FILLER_270_346 ();
 b15zdnd11an1n64x5 FILLER_270_353 ();
 b15zdnd11an1n64x5 FILLER_270_417 ();
 b15zdnd11an1n64x5 FILLER_270_481 ();
 b15zdnd11an1n64x5 FILLER_270_545 ();
 b15zdnd11an1n64x5 FILLER_270_609 ();
 b15zdnd11an1n32x5 FILLER_270_673 ();
 b15zdnd00an1n01x5 FILLER_270_705 ();
 b15zdnd11an1n04x5 FILLER_270_709 ();
 b15zdnd00an1n02x5 FILLER_270_716 ();
 b15zdnd11an1n64x5 FILLER_270_726 ();
 b15zdnd11an1n64x5 FILLER_270_790 ();
 b15zdnd11an1n64x5 FILLER_270_854 ();
 b15zdnd11an1n64x5 FILLER_270_918 ();
 b15zdnd11an1n64x5 FILLER_270_982 ();
 b15zdnd11an1n32x5 FILLER_270_1046 ();
 b15zdnd11an1n04x5 FILLER_270_1078 ();
 b15zdnd00an1n02x5 FILLER_270_1082 ();
 b15zdnd11an1n04x5 FILLER_270_1087 ();
 b15zdnd11an1n08x5 FILLER_270_1094 ();
 b15zdnd00an1n01x5 FILLER_270_1102 ();
 b15zdnd11an1n64x5 FILLER_270_1155 ();
 b15zdnd11an1n64x5 FILLER_270_1219 ();
 b15zdnd11an1n04x5 FILLER_270_1283 ();
 b15zdnd11an1n04x5 FILLER_270_1290 ();
 b15zdnd11an1n64x5 FILLER_270_1297 ();
 b15zdnd11an1n64x5 FILLER_270_1361 ();
 b15zdnd11an1n32x5 FILLER_270_1425 ();
 b15zdnd11an1n16x5 FILLER_270_1457 ();
 b15zdnd11an1n04x5 FILLER_270_1473 ();
 b15zdnd00an1n01x5 FILLER_270_1477 ();
 b15zdnd11an1n64x5 FILLER_270_1490 ();
 b15zdnd11an1n64x5 FILLER_270_1554 ();
 b15zdnd11an1n64x5 FILLER_270_1618 ();
 b15zdnd11an1n64x5 FILLER_270_1682 ();
 b15zdnd11an1n32x5 FILLER_270_1746 ();
 b15zdnd11an1n08x5 FILLER_270_1778 ();
 b15zdnd00an1n02x5 FILLER_270_1786 ();
 b15zdnd00an1n01x5 FILLER_270_1788 ();
 b15zdnd11an1n04x5 FILLER_270_1792 ();
 b15zdnd11an1n04x5 FILLER_270_1799 ();
 b15zdnd11an1n04x5 FILLER_270_1806 ();
 b15zdnd00an1n01x5 FILLER_270_1810 ();
 b15zdnd11an1n32x5 FILLER_270_1819 ();
 b15zdnd00an1n02x5 FILLER_270_1851 ();
 b15zdnd11an1n64x5 FILLER_270_1856 ();
 b15zdnd11an1n64x5 FILLER_270_1920 ();
 b15zdnd11an1n64x5 FILLER_270_1984 ();
 b15zdnd11an1n08x5 FILLER_270_2048 ();
 b15zdnd11an1n04x5 FILLER_270_2056 ();
 b15zdnd00an1n01x5 FILLER_270_2060 ();
 b15zdnd11an1n64x5 FILLER_270_2086 ();
 b15zdnd11an1n04x5 FILLER_270_2150 ();
 b15zdnd11an1n64x5 FILLER_270_2162 ();
 b15zdnd11an1n32x5 FILLER_270_2226 ();
 b15zdnd11an1n16x5 FILLER_270_2258 ();
 b15zdnd00an1n02x5 FILLER_270_2274 ();
 b15zdnd11an1n64x5 FILLER_271_0 ();
 b15zdnd11an1n64x5 FILLER_271_64 ();
 b15zdnd11an1n64x5 FILLER_271_128 ();
 b15zdnd11an1n64x5 FILLER_271_192 ();
 b15zdnd11an1n64x5 FILLER_271_256 ();
 b15zdnd11an1n16x5 FILLER_271_320 ();
 b15zdnd11an1n04x5 FILLER_271_336 ();
 b15zdnd00an1n02x5 FILLER_271_340 ();
 b15zdnd11an1n64x5 FILLER_271_345 ();
 b15zdnd11an1n64x5 FILLER_271_409 ();
 b15zdnd11an1n64x5 FILLER_271_473 ();
 b15zdnd11an1n64x5 FILLER_271_537 ();
 b15zdnd11an1n64x5 FILLER_271_601 ();
 b15zdnd11an1n16x5 FILLER_271_665 ();
 b15zdnd11an1n04x5 FILLER_271_681 ();
 b15zdnd00an1n01x5 FILLER_271_685 ();
 b15zdnd11an1n64x5 FILLER_271_738 ();
 b15zdnd11an1n64x5 FILLER_271_802 ();
 b15zdnd11an1n64x5 FILLER_271_866 ();
 b15zdnd11an1n64x5 FILLER_271_930 ();
 b15zdnd11an1n64x5 FILLER_271_994 ();
 b15zdnd11an1n16x5 FILLER_271_1058 ();
 b15zdnd11an1n08x5 FILLER_271_1074 ();
 b15zdnd11an1n04x5 FILLER_271_1082 ();
 b15zdnd00an1n01x5 FILLER_271_1086 ();
 b15zdnd11an1n04x5 FILLER_271_1139 ();
 b15zdnd11an1n64x5 FILLER_271_1169 ();
 b15zdnd11an1n32x5 FILLER_271_1233 ();
 b15zdnd11an1n04x5 FILLER_271_1265 ();
 b15zdnd11an1n64x5 FILLER_271_1321 ();
 b15zdnd11an1n64x5 FILLER_271_1385 ();
 b15zdnd11an1n64x5 FILLER_271_1449 ();
 b15zdnd11an1n64x5 FILLER_271_1513 ();
 b15zdnd11an1n64x5 FILLER_271_1577 ();
 b15zdnd11an1n64x5 FILLER_271_1641 ();
 b15zdnd11an1n64x5 FILLER_271_1705 ();
 b15zdnd11an1n16x5 FILLER_271_1769 ();
 b15zdnd11an1n08x5 FILLER_271_1785 ();
 b15zdnd00an1n01x5 FILLER_271_1793 ();
 b15zdnd11an1n04x5 FILLER_271_1797 ();
 b15zdnd11an1n64x5 FILLER_271_1804 ();
 b15zdnd11an1n64x5 FILLER_271_1868 ();
 b15zdnd11an1n64x5 FILLER_271_1932 ();
 b15zdnd11an1n32x5 FILLER_271_1996 ();
 b15zdnd11an1n04x5 FILLER_271_2028 ();
 b15zdnd00an1n01x5 FILLER_271_2032 ();
 b15zdnd11an1n16x5 FILLER_271_2051 ();
 b15zdnd00an1n02x5 FILLER_271_2067 ();
 b15zdnd11an1n64x5 FILLER_271_2084 ();
 b15zdnd11an1n64x5 FILLER_271_2148 ();
 b15zdnd11an1n64x5 FILLER_271_2212 ();
 b15zdnd11an1n08x5 FILLER_271_2276 ();
 b15zdnd11an1n64x5 FILLER_272_8 ();
 b15zdnd11an1n64x5 FILLER_272_72 ();
 b15zdnd11an1n64x5 FILLER_272_136 ();
 b15zdnd11an1n64x5 FILLER_272_200 ();
 b15zdnd11an1n64x5 FILLER_272_264 ();
 b15zdnd11an1n64x5 FILLER_272_328 ();
 b15zdnd11an1n64x5 FILLER_272_392 ();
 b15zdnd11an1n64x5 FILLER_272_456 ();
 b15zdnd11an1n64x5 FILLER_272_520 ();
 b15zdnd11an1n64x5 FILLER_272_584 ();
 b15zdnd11an1n32x5 FILLER_272_648 ();
 b15zdnd11an1n16x5 FILLER_272_680 ();
 b15zdnd11an1n08x5 FILLER_272_696 ();
 b15zdnd11an1n04x5 FILLER_272_704 ();
 b15zdnd00an1n02x5 FILLER_272_708 ();
 b15zdnd00an1n01x5 FILLER_272_710 ();
 b15zdnd11an1n04x5 FILLER_272_714 ();
 b15zdnd00an1n02x5 FILLER_272_726 ();
 b15zdnd11an1n64x5 FILLER_272_770 ();
 b15zdnd11an1n64x5 FILLER_272_834 ();
 b15zdnd11an1n64x5 FILLER_272_898 ();
 b15zdnd11an1n64x5 FILLER_272_962 ();
 b15zdnd11an1n64x5 FILLER_272_1026 ();
 b15zdnd11an1n32x5 FILLER_272_1090 ();
 b15zdnd00an1n02x5 FILLER_272_1122 ();
 b15zdnd00an1n01x5 FILLER_272_1124 ();
 b15zdnd11an1n04x5 FILLER_272_1128 ();
 b15zdnd00an1n01x5 FILLER_272_1132 ();
 b15zdnd11an1n32x5 FILLER_272_1136 ();
 b15zdnd11an1n04x5 FILLER_272_1168 ();
 b15zdnd11an1n64x5 FILLER_272_1224 ();
 b15zdnd11an1n04x5 FILLER_272_1288 ();
 b15zdnd00an1n02x5 FILLER_272_1292 ();
 b15zdnd11an1n32x5 FILLER_272_1297 ();
 b15zdnd11an1n16x5 FILLER_272_1329 ();
 b15zdnd11an1n08x5 FILLER_272_1345 ();
 b15zdnd00an1n02x5 FILLER_272_1353 ();
 b15zdnd00an1n01x5 FILLER_272_1355 ();
 b15zdnd11an1n16x5 FILLER_272_1367 ();
 b15zdnd00an1n02x5 FILLER_272_1383 ();
 b15zdnd00an1n01x5 FILLER_272_1385 ();
 b15zdnd11an1n04x5 FILLER_272_1389 ();
 b15zdnd11an1n64x5 FILLER_272_1396 ();
 b15zdnd11an1n64x5 FILLER_272_1460 ();
 b15zdnd11an1n64x5 FILLER_272_1524 ();
 b15zdnd11an1n64x5 FILLER_272_1588 ();
 b15zdnd11an1n64x5 FILLER_272_1652 ();
 b15zdnd11an1n64x5 FILLER_272_1716 ();
 b15zdnd11an1n64x5 FILLER_272_1780 ();
 b15zdnd11an1n64x5 FILLER_272_1844 ();
 b15zdnd11an1n64x5 FILLER_272_1908 ();
 b15zdnd11an1n32x5 FILLER_272_1972 ();
 b15zdnd11an1n16x5 FILLER_272_2004 ();
 b15zdnd11an1n08x5 FILLER_272_2020 ();
 b15zdnd11an1n04x5 FILLER_272_2028 ();
 b15zdnd11an1n32x5 FILLER_272_2050 ();
 b15zdnd11an1n04x5 FILLER_272_2082 ();
 b15zdnd11an1n32x5 FILLER_272_2117 ();
 b15zdnd11an1n04x5 FILLER_272_2149 ();
 b15zdnd00an1n01x5 FILLER_272_2153 ();
 b15zdnd11an1n64x5 FILLER_272_2162 ();
 b15zdnd11an1n32x5 FILLER_272_2226 ();
 b15zdnd11an1n16x5 FILLER_272_2258 ();
 b15zdnd00an1n02x5 FILLER_272_2274 ();
 b15zdnd11an1n64x5 FILLER_273_0 ();
 b15zdnd11an1n08x5 FILLER_273_64 ();
 b15zdnd11an1n04x5 FILLER_273_72 ();
 b15zdnd00an1n02x5 FILLER_273_76 ();
 b15zdnd00an1n01x5 FILLER_273_78 ();
 b15zdnd11an1n04x5 FILLER_273_82 ();
 b15zdnd11an1n64x5 FILLER_273_89 ();
 b15zdnd11an1n64x5 FILLER_273_153 ();
 b15zdnd11an1n08x5 FILLER_273_217 ();
 b15zdnd11an1n04x5 FILLER_273_225 ();
 b15zdnd00an1n02x5 FILLER_273_229 ();
 b15zdnd11an1n64x5 FILLER_273_273 ();
 b15zdnd11an1n64x5 FILLER_273_337 ();
 b15zdnd11an1n16x5 FILLER_273_401 ();
 b15zdnd11an1n08x5 FILLER_273_417 ();
 b15zdnd11an1n04x5 FILLER_273_425 ();
 b15zdnd11an1n08x5 FILLER_273_432 ();
 b15zdnd00an1n02x5 FILLER_273_440 ();
 b15zdnd11an1n64x5 FILLER_273_484 ();
 b15zdnd11an1n64x5 FILLER_273_548 ();
 b15zdnd11an1n64x5 FILLER_273_612 ();
 b15zdnd11an1n64x5 FILLER_273_676 ();
 b15zdnd11an1n64x5 FILLER_273_740 ();
 b15zdnd11an1n64x5 FILLER_273_804 ();
 b15zdnd11an1n64x5 FILLER_273_868 ();
 b15zdnd11an1n64x5 FILLER_273_932 ();
 b15zdnd11an1n64x5 FILLER_273_996 ();
 b15zdnd11an1n16x5 FILLER_273_1060 ();
 b15zdnd11an1n04x5 FILLER_273_1076 ();
 b15zdnd11an1n64x5 FILLER_273_1125 ();
 b15zdnd00an1n01x5 FILLER_273_1189 ();
 b15zdnd11an1n04x5 FILLER_273_1193 ();
 b15zdnd11an1n64x5 FILLER_273_1200 ();
 b15zdnd11an1n08x5 FILLER_273_1264 ();
 b15zdnd11an1n04x5 FILLER_273_1272 ();
 b15zdnd00an1n02x5 FILLER_273_1276 ();
 b15zdnd00an1n01x5 FILLER_273_1278 ();
 b15zdnd11an1n16x5 FILLER_273_1299 ();
 b15zdnd11an1n08x5 FILLER_273_1315 ();
 b15zdnd11an1n04x5 FILLER_273_1323 ();
 b15zdnd11an1n32x5 FILLER_273_1330 ();
 b15zdnd11an1n04x5 FILLER_273_1362 ();
 b15zdnd00an1n02x5 FILLER_273_1366 ();
 b15zdnd11an1n64x5 FILLER_273_1420 ();
 b15zdnd11an1n64x5 FILLER_273_1484 ();
 b15zdnd11an1n64x5 FILLER_273_1548 ();
 b15zdnd11an1n64x5 FILLER_273_1612 ();
 b15zdnd11an1n64x5 FILLER_273_1676 ();
 b15zdnd11an1n64x5 FILLER_273_1740 ();
 b15zdnd11an1n64x5 FILLER_273_1804 ();
 b15zdnd11an1n64x5 FILLER_273_1868 ();
 b15zdnd11an1n64x5 FILLER_273_1932 ();
 b15zdnd11an1n64x5 FILLER_273_1996 ();
 b15zdnd11an1n64x5 FILLER_273_2060 ();
 b15zdnd11an1n64x5 FILLER_273_2124 ();
 b15zdnd11an1n16x5 FILLER_273_2188 ();
 b15zdnd11an1n08x5 FILLER_273_2216 ();
 b15zdnd00an1n02x5 FILLER_273_2224 ();
 b15zdnd11an1n32x5 FILLER_273_2238 ();
 b15zdnd11an1n08x5 FILLER_273_2270 ();
 b15zdnd11an1n04x5 FILLER_273_2278 ();
 b15zdnd00an1n02x5 FILLER_273_2282 ();
 b15zdnd11an1n32x5 FILLER_274_8 ();
 b15zdnd11an1n08x5 FILLER_274_40 ();
 b15zdnd11an1n04x5 FILLER_274_48 ();
 b15zdnd00an1n01x5 FILLER_274_52 ();
 b15zdnd11an1n04x5 FILLER_274_105 ();
 b15zdnd00an1n02x5 FILLER_274_109 ();
 b15zdnd11an1n64x5 FILLER_274_153 ();
 b15zdnd11an1n64x5 FILLER_274_217 ();
 b15zdnd11an1n64x5 FILLER_274_281 ();
 b15zdnd11an1n32x5 FILLER_274_345 ();
 b15zdnd11an1n16x5 FILLER_274_377 ();
 b15zdnd11an1n08x5 FILLER_274_393 ();
 b15zdnd00an1n01x5 FILLER_274_401 ();
 b15zdnd11an1n64x5 FILLER_274_454 ();
 b15zdnd11an1n16x5 FILLER_274_518 ();
 b15zdnd11an1n08x5 FILLER_274_534 ();
 b15zdnd00an1n02x5 FILLER_274_542 ();
 b15zdnd11an1n64x5 FILLER_274_547 ();
 b15zdnd11an1n64x5 FILLER_274_611 ();
 b15zdnd11an1n32x5 FILLER_274_675 ();
 b15zdnd11an1n08x5 FILLER_274_707 ();
 b15zdnd00an1n02x5 FILLER_274_715 ();
 b15zdnd00an1n01x5 FILLER_274_717 ();
 b15zdnd11an1n64x5 FILLER_274_726 ();
 b15zdnd11an1n64x5 FILLER_274_790 ();
 b15zdnd11an1n64x5 FILLER_274_854 ();
 b15zdnd11an1n64x5 FILLER_274_918 ();
 b15zdnd11an1n64x5 FILLER_274_982 ();
 b15zdnd11an1n32x5 FILLER_274_1046 ();
 b15zdnd11an1n16x5 FILLER_274_1078 ();
 b15zdnd11an1n08x5 FILLER_274_1094 ();
 b15zdnd11an1n04x5 FILLER_274_1102 ();
 b15zdnd00an1n02x5 FILLER_274_1106 ();
 b15zdnd00an1n01x5 FILLER_274_1108 ();
 b15zdnd11an1n04x5 FILLER_274_1141 ();
 b15zdnd11an1n32x5 FILLER_274_1159 ();
 b15zdnd11an1n04x5 FILLER_274_1191 ();
 b15zdnd11an1n64x5 FILLER_274_1198 ();
 b15zdnd11an1n32x5 FILLER_274_1262 ();
 b15zdnd11an1n08x5 FILLER_274_1294 ();
 b15zdnd00an1n02x5 FILLER_274_1302 ();
 b15zdnd11an1n32x5 FILLER_274_1356 ();
 b15zdnd11an1n04x5 FILLER_274_1388 ();
 b15zdnd00an1n02x5 FILLER_274_1392 ();
 b15zdnd11an1n64x5 FILLER_274_1397 ();
 b15zdnd11an1n64x5 FILLER_274_1461 ();
 b15zdnd11an1n64x5 FILLER_274_1525 ();
 b15zdnd11an1n64x5 FILLER_274_1589 ();
 b15zdnd11an1n64x5 FILLER_274_1653 ();
 b15zdnd11an1n64x5 FILLER_274_1717 ();
 b15zdnd11an1n64x5 FILLER_274_1781 ();
 b15zdnd11an1n64x5 FILLER_274_1845 ();
 b15zdnd11an1n64x5 FILLER_274_1909 ();
 b15zdnd11an1n64x5 FILLER_274_1973 ();
 b15zdnd11an1n64x5 FILLER_274_2037 ();
 b15zdnd11an1n32x5 FILLER_274_2101 ();
 b15zdnd11an1n16x5 FILLER_274_2133 ();
 b15zdnd11an1n04x5 FILLER_274_2149 ();
 b15zdnd00an1n01x5 FILLER_274_2153 ();
 b15zdnd11an1n16x5 FILLER_274_2162 ();
 b15zdnd11an1n04x5 FILLER_274_2178 ();
 b15zdnd11an1n04x5 FILLER_274_2213 ();
 b15zdnd11an1n32x5 FILLER_274_2232 ();
 b15zdnd11an1n08x5 FILLER_274_2264 ();
 b15zdnd11an1n04x5 FILLER_274_2272 ();
 b15zdnd11an1n32x5 FILLER_275_0 ();
 b15zdnd11an1n16x5 FILLER_275_32 ();
 b15zdnd11an1n08x5 FILLER_275_48 ();
 b15zdnd11an1n64x5 FILLER_275_108 ();
 b15zdnd11an1n64x5 FILLER_275_172 ();
 b15zdnd11an1n64x5 FILLER_275_236 ();
 b15zdnd11an1n64x5 FILLER_275_300 ();
 b15zdnd11an1n32x5 FILLER_275_364 ();
 b15zdnd11an1n16x5 FILLER_275_396 ();
 b15zdnd00an1n01x5 FILLER_275_412 ();
 b15zdnd11an1n16x5 FILLER_275_455 ();
 b15zdnd00an1n01x5 FILLER_275_471 ();
 b15zdnd11an1n32x5 FILLER_275_475 ();
 b15zdnd11an1n08x5 FILLER_275_507 ();
 b15zdnd00an1n02x5 FILLER_275_515 ();
 b15zdnd11an1n64x5 FILLER_275_569 ();
 b15zdnd11an1n64x5 FILLER_275_633 ();
 b15zdnd11an1n64x5 FILLER_275_697 ();
 b15zdnd11an1n64x5 FILLER_275_761 ();
 b15zdnd00an1n01x5 FILLER_275_825 ();
 b15zdnd11an1n04x5 FILLER_275_837 ();
 b15zdnd11an1n04x5 FILLER_275_857 ();
 b15zdnd11an1n64x5 FILLER_275_864 ();
 b15zdnd11an1n64x5 FILLER_275_928 ();
 b15zdnd11an1n64x5 FILLER_275_992 ();
 b15zdnd11an1n32x5 FILLER_275_1056 ();
 b15zdnd11an1n08x5 FILLER_275_1088 ();
 b15zdnd11an1n04x5 FILLER_275_1096 ();
 b15zdnd11an1n64x5 FILLER_275_1111 ();
 b15zdnd11an1n64x5 FILLER_275_1175 ();
 b15zdnd11an1n16x5 FILLER_275_1239 ();
 b15zdnd11an1n08x5 FILLER_275_1255 ();
 b15zdnd00an1n02x5 FILLER_275_1263 ();
 b15zdnd00an1n01x5 FILLER_275_1265 ();
 b15zdnd11an1n32x5 FILLER_275_1286 ();
 b15zdnd11an1n04x5 FILLER_275_1318 ();
 b15zdnd11an1n04x5 FILLER_275_1325 ();
 b15zdnd11an1n64x5 FILLER_275_1332 ();
 b15zdnd11an1n64x5 FILLER_275_1396 ();
 b15zdnd11an1n64x5 FILLER_275_1460 ();
 b15zdnd11an1n64x5 FILLER_275_1524 ();
 b15zdnd11an1n64x5 FILLER_275_1588 ();
 b15zdnd11an1n64x5 FILLER_275_1652 ();
 b15zdnd11an1n64x5 FILLER_275_1716 ();
 b15zdnd11an1n64x5 FILLER_275_1780 ();
 b15zdnd11an1n64x5 FILLER_275_1844 ();
 b15zdnd11an1n64x5 FILLER_275_1908 ();
 b15zdnd11an1n64x5 FILLER_275_1972 ();
 b15zdnd11an1n64x5 FILLER_275_2036 ();
 b15zdnd11an1n64x5 FILLER_275_2100 ();
 b15zdnd11an1n64x5 FILLER_275_2164 ();
 b15zdnd11an1n32x5 FILLER_275_2228 ();
 b15zdnd11an1n16x5 FILLER_275_2260 ();
 b15zdnd11an1n08x5 FILLER_275_2276 ();
 b15zdnd11an1n64x5 FILLER_276_8 ();
 b15zdnd00an1n01x5 FILLER_276_72 ();
 b15zdnd11an1n04x5 FILLER_276_76 ();
 b15zdnd11an1n04x5 FILLER_276_83 ();
 b15zdnd11an1n64x5 FILLER_276_90 ();
 b15zdnd11an1n64x5 FILLER_276_154 ();
 b15zdnd11an1n64x5 FILLER_276_218 ();
 b15zdnd11an1n64x5 FILLER_276_282 ();
 b15zdnd11an1n64x5 FILLER_276_346 ();
 b15zdnd11an1n08x5 FILLER_276_410 ();
 b15zdnd00an1n02x5 FILLER_276_418 ();
 b15zdnd11an1n04x5 FILLER_276_423 ();
 b15zdnd11an1n08x5 FILLER_276_430 ();
 b15zdnd11an1n04x5 FILLER_276_438 ();
 b15zdnd00an1n02x5 FILLER_276_442 ();
 b15zdnd00an1n01x5 FILLER_276_444 ();
 b15zdnd11an1n32x5 FILLER_276_497 ();
 b15zdnd11an1n04x5 FILLER_276_529 ();
 b15zdnd00an1n02x5 FILLER_276_533 ();
 b15zdnd11an1n04x5 FILLER_276_538 ();
 b15zdnd11an1n64x5 FILLER_276_545 ();
 b15zdnd11an1n64x5 FILLER_276_609 ();
 b15zdnd11an1n32x5 FILLER_276_673 ();
 b15zdnd11an1n08x5 FILLER_276_705 ();
 b15zdnd11an1n04x5 FILLER_276_713 ();
 b15zdnd00an1n01x5 FILLER_276_717 ();
 b15zdnd11an1n64x5 FILLER_276_726 ();
 b15zdnd11an1n32x5 FILLER_276_790 ();
 b15zdnd11an1n16x5 FILLER_276_822 ();
 b15zdnd00an1n02x5 FILLER_276_838 ();
 b15zdnd11an1n64x5 FILLER_276_882 ();
 b15zdnd11an1n64x5 FILLER_276_946 ();
 b15zdnd11an1n64x5 FILLER_276_1010 ();
 b15zdnd11an1n32x5 FILLER_276_1074 ();
 b15zdnd11an1n16x5 FILLER_276_1106 ();
 b15zdnd11an1n08x5 FILLER_276_1122 ();
 b15zdnd00an1n02x5 FILLER_276_1130 ();
 b15zdnd00an1n01x5 FILLER_276_1132 ();
 b15zdnd11an1n64x5 FILLER_276_1147 ();
 b15zdnd11an1n64x5 FILLER_276_1211 ();
 b15zdnd11an1n64x5 FILLER_276_1275 ();
 b15zdnd11an1n64x5 FILLER_276_1339 ();
 b15zdnd11an1n64x5 FILLER_276_1403 ();
 b15zdnd11an1n64x5 FILLER_276_1467 ();
 b15zdnd11an1n64x5 FILLER_276_1531 ();
 b15zdnd11an1n64x5 FILLER_276_1595 ();
 b15zdnd11an1n64x5 FILLER_276_1659 ();
 b15zdnd11an1n64x5 FILLER_276_1723 ();
 b15zdnd11an1n64x5 FILLER_276_1787 ();
 b15zdnd11an1n64x5 FILLER_276_1851 ();
 b15zdnd11an1n64x5 FILLER_276_1915 ();
 b15zdnd11an1n64x5 FILLER_276_1979 ();
 b15zdnd11an1n64x5 FILLER_276_2043 ();
 b15zdnd11an1n32x5 FILLER_276_2107 ();
 b15zdnd11an1n08x5 FILLER_276_2139 ();
 b15zdnd11an1n04x5 FILLER_276_2147 ();
 b15zdnd00an1n02x5 FILLER_276_2151 ();
 b15zdnd00an1n01x5 FILLER_276_2153 ();
 b15zdnd11an1n64x5 FILLER_276_2162 ();
 b15zdnd11an1n32x5 FILLER_276_2226 ();
 b15zdnd11an1n16x5 FILLER_276_2258 ();
 b15zdnd00an1n02x5 FILLER_276_2274 ();
 b15zdnd11an1n64x5 FILLER_277_0 ();
 b15zdnd11an1n16x5 FILLER_277_64 ();
 b15zdnd00an1n01x5 FILLER_277_80 ();
 b15zdnd11an1n64x5 FILLER_277_84 ();
 b15zdnd11an1n32x5 FILLER_277_148 ();
 b15zdnd11an1n16x5 FILLER_277_180 ();
 b15zdnd11an1n08x5 FILLER_277_196 ();
 b15zdnd11an1n04x5 FILLER_277_204 ();
 b15zdnd00an1n02x5 FILLER_277_208 ();
 b15zdnd11an1n64x5 FILLER_277_219 ();
 b15zdnd11an1n64x5 FILLER_277_283 ();
 b15zdnd11an1n64x5 FILLER_277_347 ();
 b15zdnd11an1n32x5 FILLER_277_411 ();
 b15zdnd11an1n16x5 FILLER_277_443 ();
 b15zdnd11an1n04x5 FILLER_277_459 ();
 b15zdnd11an1n04x5 FILLER_277_466 ();
 b15zdnd11an1n64x5 FILLER_277_473 ();
 b15zdnd11an1n64x5 FILLER_277_537 ();
 b15zdnd11an1n04x5 FILLER_277_601 ();
 b15zdnd00an1n01x5 FILLER_277_605 ();
 b15zdnd11an1n64x5 FILLER_277_609 ();
 b15zdnd11an1n64x5 FILLER_277_673 ();
 b15zdnd11an1n64x5 FILLER_277_737 ();
 b15zdnd11an1n16x5 FILLER_277_801 ();
 b15zdnd11an1n08x5 FILLER_277_817 ();
 b15zdnd11an1n04x5 FILLER_277_825 ();
 b15zdnd11an1n64x5 FILLER_277_881 ();
 b15zdnd11an1n64x5 FILLER_277_945 ();
 b15zdnd11an1n64x5 FILLER_277_1009 ();
 b15zdnd11an1n64x5 FILLER_277_1073 ();
 b15zdnd11an1n64x5 FILLER_277_1137 ();
 b15zdnd11an1n64x5 FILLER_277_1201 ();
 b15zdnd11an1n64x5 FILLER_277_1265 ();
 b15zdnd11an1n64x5 FILLER_277_1329 ();
 b15zdnd11an1n64x5 FILLER_277_1393 ();
 b15zdnd11an1n64x5 FILLER_277_1457 ();
 b15zdnd11an1n64x5 FILLER_277_1521 ();
 b15zdnd11an1n64x5 FILLER_277_1585 ();
 b15zdnd11an1n08x5 FILLER_277_1649 ();
 b15zdnd11an1n64x5 FILLER_277_1660 ();
 b15zdnd11an1n64x5 FILLER_277_1724 ();
 b15zdnd11an1n64x5 FILLER_277_1788 ();
 b15zdnd11an1n64x5 FILLER_277_1852 ();
 b15zdnd11an1n64x5 FILLER_277_1916 ();
 b15zdnd11an1n64x5 FILLER_277_1980 ();
 b15zdnd11an1n64x5 FILLER_277_2044 ();
 b15zdnd11an1n64x5 FILLER_277_2108 ();
 b15zdnd11an1n64x5 FILLER_277_2172 ();
 b15zdnd11an1n32x5 FILLER_277_2236 ();
 b15zdnd11an1n16x5 FILLER_277_2268 ();
 b15zdnd11an1n64x5 FILLER_278_8 ();
 b15zdnd11an1n64x5 FILLER_278_72 ();
 b15zdnd11an1n64x5 FILLER_278_136 ();
 b15zdnd11an1n08x5 FILLER_278_200 ();
 b15zdnd00an1n02x5 FILLER_278_208 ();
 b15zdnd11an1n64x5 FILLER_278_252 ();
 b15zdnd11an1n64x5 FILLER_278_316 ();
 b15zdnd11an1n32x5 FILLER_278_380 ();
 b15zdnd11an1n16x5 FILLER_278_412 ();
 b15zdnd00an1n01x5 FILLER_278_428 ();
 b15zdnd11an1n64x5 FILLER_278_455 ();
 b15zdnd11an1n64x5 FILLER_278_519 ();
 b15zdnd11an1n04x5 FILLER_278_583 ();
 b15zdnd00an1n02x5 FILLER_278_587 ();
 b15zdnd00an1n01x5 FILLER_278_589 ();
 b15zdnd11an1n64x5 FILLER_278_632 ();
 b15zdnd11an1n16x5 FILLER_278_696 ();
 b15zdnd11an1n04x5 FILLER_278_712 ();
 b15zdnd00an1n02x5 FILLER_278_716 ();
 b15zdnd11an1n64x5 FILLER_278_726 ();
 b15zdnd11an1n32x5 FILLER_278_790 ();
 b15zdnd11an1n16x5 FILLER_278_822 ();
 b15zdnd11an1n08x5 FILLER_278_838 ();
 b15zdnd00an1n01x5 FILLER_278_846 ();
 b15zdnd11an1n04x5 FILLER_278_850 ();
 b15zdnd11an1n08x5 FILLER_278_857 ();
 b15zdnd11an1n04x5 FILLER_278_865 ();
 b15zdnd11an1n64x5 FILLER_278_911 ();
 b15zdnd11an1n64x5 FILLER_278_975 ();
 b15zdnd11an1n64x5 FILLER_278_1039 ();
 b15zdnd11an1n32x5 FILLER_278_1103 ();
 b15zdnd11an1n16x5 FILLER_278_1135 ();
 b15zdnd11an1n04x5 FILLER_278_1151 ();
 b15zdnd11an1n64x5 FILLER_278_1164 ();
 b15zdnd11an1n64x5 FILLER_278_1228 ();
 b15zdnd11an1n16x5 FILLER_278_1292 ();
 b15zdnd11an1n08x5 FILLER_278_1308 ();
 b15zdnd11an1n04x5 FILLER_278_1316 ();
 b15zdnd00an1n01x5 FILLER_278_1320 ();
 b15zdnd11an1n64x5 FILLER_278_1330 ();
 b15zdnd11an1n64x5 FILLER_278_1394 ();
 b15zdnd11an1n64x5 FILLER_278_1458 ();
 b15zdnd11an1n32x5 FILLER_278_1522 ();
 b15zdnd11an1n04x5 FILLER_278_1554 ();
 b15zdnd00an1n02x5 FILLER_278_1558 ();
 b15zdnd00an1n01x5 FILLER_278_1560 ();
 b15zdnd11an1n04x5 FILLER_278_1564 ();
 b15zdnd11an1n64x5 FILLER_278_1571 ();
 b15zdnd11an1n16x5 FILLER_278_1635 ();
 b15zdnd11an1n04x5 FILLER_278_1651 ();
 b15zdnd00an1n01x5 FILLER_278_1655 ();
 b15zdnd11an1n64x5 FILLER_278_1659 ();
 b15zdnd11an1n64x5 FILLER_278_1723 ();
 b15zdnd11an1n64x5 FILLER_278_1787 ();
 b15zdnd11an1n64x5 FILLER_278_1851 ();
 b15zdnd11an1n64x5 FILLER_278_1915 ();
 b15zdnd11an1n64x5 FILLER_278_1979 ();
 b15zdnd11an1n64x5 FILLER_278_2043 ();
 b15zdnd11an1n32x5 FILLER_278_2107 ();
 b15zdnd11an1n08x5 FILLER_278_2139 ();
 b15zdnd11an1n04x5 FILLER_278_2147 ();
 b15zdnd00an1n02x5 FILLER_278_2151 ();
 b15zdnd00an1n01x5 FILLER_278_2153 ();
 b15zdnd11an1n64x5 FILLER_278_2162 ();
 b15zdnd11an1n32x5 FILLER_278_2226 ();
 b15zdnd11an1n16x5 FILLER_278_2258 ();
 b15zdnd00an1n02x5 FILLER_278_2274 ();
 b15zdnd11an1n64x5 FILLER_279_0 ();
 b15zdnd11an1n64x5 FILLER_279_64 ();
 b15zdnd11an1n64x5 FILLER_279_128 ();
 b15zdnd11an1n64x5 FILLER_279_192 ();
 b15zdnd11an1n64x5 FILLER_279_256 ();
 b15zdnd11an1n64x5 FILLER_279_320 ();
 b15zdnd11an1n64x5 FILLER_279_384 ();
 b15zdnd11an1n64x5 FILLER_279_448 ();
 b15zdnd11an1n64x5 FILLER_279_512 ();
 b15zdnd00an1n02x5 FILLER_279_576 ();
 b15zdnd00an1n01x5 FILLER_279_578 ();
 b15zdnd11an1n64x5 FILLER_279_631 ();
 b15zdnd11an1n64x5 FILLER_279_695 ();
 b15zdnd11an1n64x5 FILLER_279_759 ();
 b15zdnd11an1n64x5 FILLER_279_823 ();
 b15zdnd11an1n64x5 FILLER_279_887 ();
 b15zdnd11an1n64x5 FILLER_279_951 ();
 b15zdnd11an1n64x5 FILLER_279_1015 ();
 b15zdnd11an1n64x5 FILLER_279_1079 ();
 b15zdnd11an1n64x5 FILLER_279_1143 ();
 b15zdnd11an1n64x5 FILLER_279_1207 ();
 b15zdnd11an1n64x5 FILLER_279_1271 ();
 b15zdnd11an1n64x5 FILLER_279_1335 ();
 b15zdnd11an1n64x5 FILLER_279_1399 ();
 b15zdnd11an1n64x5 FILLER_279_1463 ();
 b15zdnd11an1n04x5 FILLER_279_1530 ();
 b15zdnd11an1n04x5 FILLER_279_1537 ();
 b15zdnd00an1n02x5 FILLER_279_1541 ();
 b15zdnd11an1n32x5 FILLER_279_1595 ();
 b15zdnd11an1n04x5 FILLER_279_1627 ();
 b15zdnd11an1n64x5 FILLER_279_1683 ();
 b15zdnd11an1n64x5 FILLER_279_1747 ();
 b15zdnd11an1n64x5 FILLER_279_1811 ();
 b15zdnd11an1n64x5 FILLER_279_1875 ();
 b15zdnd11an1n64x5 FILLER_279_1939 ();
 b15zdnd11an1n64x5 FILLER_279_2003 ();
 b15zdnd11an1n64x5 FILLER_279_2067 ();
 b15zdnd11an1n64x5 FILLER_279_2131 ();
 b15zdnd11an1n64x5 FILLER_279_2195 ();
 b15zdnd11an1n16x5 FILLER_279_2259 ();
 b15zdnd11an1n08x5 FILLER_279_2275 ();
 b15zdnd00an1n01x5 FILLER_279_2283 ();
 b15zdnd11an1n32x5 FILLER_280_8 ();
 b15zdnd11an1n08x5 FILLER_280_40 ();
 b15zdnd00an1n02x5 FILLER_280_48 ();
 b15zdnd11an1n64x5 FILLER_280_92 ();
 b15zdnd11an1n64x5 FILLER_280_156 ();
 b15zdnd11an1n64x5 FILLER_280_220 ();
 b15zdnd11an1n64x5 FILLER_280_284 ();
 b15zdnd11an1n64x5 FILLER_280_348 ();
 b15zdnd11an1n16x5 FILLER_280_412 ();
 b15zdnd11an1n08x5 FILLER_280_428 ();
 b15zdnd11an1n64x5 FILLER_280_444 ();
 b15zdnd11an1n64x5 FILLER_280_508 ();
 b15zdnd11an1n32x5 FILLER_280_572 ();
 b15zdnd11an1n04x5 FILLER_280_607 ();
 b15zdnd11an1n04x5 FILLER_280_614 ();
 b15zdnd00an1n01x5 FILLER_280_618 ();
 b15zdnd11an1n32x5 FILLER_280_661 ();
 b15zdnd11an1n16x5 FILLER_280_693 ();
 b15zdnd11an1n08x5 FILLER_280_709 ();
 b15zdnd00an1n01x5 FILLER_280_717 ();
 b15zdnd11an1n64x5 FILLER_280_726 ();
 b15zdnd11an1n64x5 FILLER_280_790 ();
 b15zdnd11an1n64x5 FILLER_280_854 ();
 b15zdnd11an1n64x5 FILLER_280_918 ();
 b15zdnd11an1n64x5 FILLER_280_982 ();
 b15zdnd11an1n64x5 FILLER_280_1046 ();
 b15zdnd11an1n64x5 FILLER_280_1110 ();
 b15zdnd11an1n32x5 FILLER_280_1174 ();
 b15zdnd11an1n04x5 FILLER_280_1206 ();
 b15zdnd11an1n64x5 FILLER_280_1213 ();
 b15zdnd11an1n64x5 FILLER_280_1277 ();
 b15zdnd11an1n64x5 FILLER_280_1341 ();
 b15zdnd11an1n64x5 FILLER_280_1405 ();
 b15zdnd11an1n32x5 FILLER_280_1469 ();
 b15zdnd11an1n08x5 FILLER_280_1501 ();
 b15zdnd11an1n04x5 FILLER_280_1561 ();
 b15zdnd00an1n02x5 FILLER_280_1565 ();
 b15zdnd00an1n01x5 FILLER_280_1567 ();
 b15zdnd11an1n64x5 FILLER_280_1571 ();
 b15zdnd11an1n08x5 FILLER_280_1635 ();
 b15zdnd11an1n04x5 FILLER_280_1643 ();
 b15zdnd00an1n02x5 FILLER_280_1647 ();
 b15zdnd11an1n04x5 FILLER_280_1652 ();
 b15zdnd11an1n64x5 FILLER_280_1659 ();
 b15zdnd11an1n64x5 FILLER_280_1723 ();
 b15zdnd11an1n64x5 FILLER_280_1787 ();
 b15zdnd11an1n64x5 FILLER_280_1851 ();
 b15zdnd11an1n64x5 FILLER_280_1915 ();
 b15zdnd11an1n64x5 FILLER_280_1979 ();
 b15zdnd11an1n64x5 FILLER_280_2043 ();
 b15zdnd11an1n32x5 FILLER_280_2107 ();
 b15zdnd11an1n08x5 FILLER_280_2139 ();
 b15zdnd11an1n04x5 FILLER_280_2147 ();
 b15zdnd00an1n02x5 FILLER_280_2151 ();
 b15zdnd00an1n01x5 FILLER_280_2153 ();
 b15zdnd11an1n64x5 FILLER_280_2162 ();
 b15zdnd11an1n32x5 FILLER_280_2226 ();
 b15zdnd11an1n16x5 FILLER_280_2258 ();
 b15zdnd00an1n02x5 FILLER_280_2274 ();
 b15zdnd11an1n64x5 FILLER_281_0 ();
 b15zdnd11an1n32x5 FILLER_281_64 ();
 b15zdnd11an1n16x5 FILLER_281_96 ();
 b15zdnd11an1n08x5 FILLER_281_112 ();
 b15zdnd00an1n02x5 FILLER_281_120 ();
 b15zdnd00an1n01x5 FILLER_281_122 ();
 b15zdnd11an1n64x5 FILLER_281_165 ();
 b15zdnd11an1n64x5 FILLER_281_229 ();
 b15zdnd11an1n64x5 FILLER_281_293 ();
 b15zdnd11an1n64x5 FILLER_281_357 ();
 b15zdnd11an1n16x5 FILLER_281_421 ();
 b15zdnd00an1n02x5 FILLER_281_437 ();
 b15zdnd00an1n01x5 FILLER_281_439 ();
 b15zdnd11an1n64x5 FILLER_281_460 ();
 b15zdnd11an1n16x5 FILLER_281_524 ();
 b15zdnd11an1n08x5 FILLER_281_540 ();
 b15zdnd11an1n04x5 FILLER_281_548 ();
 b15zdnd00an1n02x5 FILLER_281_552 ();
 b15zdnd11an1n32x5 FILLER_281_558 ();
 b15zdnd11an1n08x5 FILLER_281_590 ();
 b15zdnd00an1n02x5 FILLER_281_598 ();
 b15zdnd11an1n64x5 FILLER_281_608 ();
 b15zdnd11an1n16x5 FILLER_281_672 ();
 b15zdnd00an1n02x5 FILLER_281_688 ();
 b15zdnd00an1n01x5 FILLER_281_690 ();
 b15zdnd11an1n32x5 FILLER_281_733 ();
 b15zdnd11an1n04x5 FILLER_281_765 ();
 b15zdnd11an1n64x5 FILLER_281_772 ();
 b15zdnd11an1n64x5 FILLER_281_836 ();
 b15zdnd11an1n64x5 FILLER_281_900 ();
 b15zdnd11an1n64x5 FILLER_281_964 ();
 b15zdnd11an1n64x5 FILLER_281_1028 ();
 b15zdnd11an1n64x5 FILLER_281_1092 ();
 b15zdnd11an1n32x5 FILLER_281_1156 ();
 b15zdnd11an1n16x5 FILLER_281_1188 ();
 b15zdnd11an1n04x5 FILLER_281_1204 ();
 b15zdnd00an1n02x5 FILLER_281_1208 ();
 b15zdnd11an1n64x5 FILLER_281_1213 ();
 b15zdnd11an1n64x5 FILLER_281_1277 ();
 b15zdnd11an1n64x5 FILLER_281_1341 ();
 b15zdnd11an1n64x5 FILLER_281_1405 ();
 b15zdnd11an1n16x5 FILLER_281_1469 ();
 b15zdnd11an1n08x5 FILLER_281_1485 ();
 b15zdnd11an1n04x5 FILLER_281_1493 ();
 b15zdnd00an1n02x5 FILLER_281_1497 ();
 b15zdnd00an1n01x5 FILLER_281_1499 ();
 b15zdnd11an1n04x5 FILLER_281_1503 ();
 b15zdnd11an1n04x5 FILLER_281_1534 ();
 b15zdnd11an1n64x5 FILLER_281_1541 ();
 b15zdnd11an1n16x5 FILLER_281_1605 ();
 b15zdnd00an1n02x5 FILLER_281_1621 ();
 b15zdnd00an1n01x5 FILLER_281_1623 ();
 b15zdnd11an1n64x5 FILLER_281_1676 ();
 b15zdnd11an1n64x5 FILLER_281_1740 ();
 b15zdnd11an1n64x5 FILLER_281_1804 ();
 b15zdnd11an1n64x5 FILLER_281_1868 ();
 b15zdnd11an1n64x5 FILLER_281_1932 ();
 b15zdnd11an1n64x5 FILLER_281_1996 ();
 b15zdnd11an1n64x5 FILLER_281_2060 ();
 b15zdnd11an1n64x5 FILLER_281_2124 ();
 b15zdnd11an1n64x5 FILLER_281_2188 ();
 b15zdnd11an1n32x5 FILLER_281_2252 ();
 b15zdnd11an1n64x5 FILLER_282_8 ();
 b15zdnd11an1n64x5 FILLER_282_72 ();
 b15zdnd11an1n32x5 FILLER_282_136 ();
 b15zdnd11an1n04x5 FILLER_282_168 ();
 b15zdnd00an1n02x5 FILLER_282_172 ();
 b15zdnd00an1n01x5 FILLER_282_174 ();
 b15zdnd11an1n64x5 FILLER_282_178 ();
 b15zdnd11an1n64x5 FILLER_282_242 ();
 b15zdnd11an1n64x5 FILLER_282_306 ();
 b15zdnd11an1n64x5 FILLER_282_370 ();
 b15zdnd11an1n64x5 FILLER_282_434 ();
 b15zdnd11an1n64x5 FILLER_282_498 ();
 b15zdnd11an1n64x5 FILLER_282_562 ();
 b15zdnd11an1n64x5 FILLER_282_626 ();
 b15zdnd11an1n16x5 FILLER_282_690 ();
 b15zdnd00an1n01x5 FILLER_282_706 ();
 b15zdnd11an1n08x5 FILLER_282_710 ();
 b15zdnd11an1n16x5 FILLER_282_726 ();
 b15zdnd11an1n08x5 FILLER_282_742 ();
 b15zdnd00an1n02x5 FILLER_282_750 ();
 b15zdnd00an1n01x5 FILLER_282_752 ();
 b15zdnd11an1n64x5 FILLER_282_795 ();
 b15zdnd11an1n64x5 FILLER_282_859 ();
 b15zdnd11an1n64x5 FILLER_282_923 ();
 b15zdnd11an1n64x5 FILLER_282_987 ();
 b15zdnd11an1n64x5 FILLER_282_1051 ();
 b15zdnd11an1n32x5 FILLER_282_1115 ();
 b15zdnd11an1n16x5 FILLER_282_1147 ();
 b15zdnd11an1n08x5 FILLER_282_1163 ();
 b15zdnd11an1n04x5 FILLER_282_1180 ();
 b15zdnd00an1n01x5 FILLER_282_1184 ();
 b15zdnd11an1n64x5 FILLER_282_1237 ();
 b15zdnd11an1n64x5 FILLER_282_1301 ();
 b15zdnd11an1n64x5 FILLER_282_1365 ();
 b15zdnd11an1n64x5 FILLER_282_1429 ();
 b15zdnd11an1n64x5 FILLER_282_1493 ();
 b15zdnd11an1n64x5 FILLER_282_1557 ();
 b15zdnd11an1n16x5 FILLER_282_1621 ();
 b15zdnd11an1n04x5 FILLER_282_1637 ();
 b15zdnd00an1n02x5 FILLER_282_1641 ();
 b15zdnd11an1n04x5 FILLER_282_1646 ();
 b15zdnd11an1n64x5 FILLER_282_1653 ();
 b15zdnd11an1n64x5 FILLER_282_1717 ();
 b15zdnd11an1n64x5 FILLER_282_1781 ();
 b15zdnd11an1n32x5 FILLER_282_1845 ();
 b15zdnd11an1n16x5 FILLER_282_1877 ();
 b15zdnd11an1n04x5 FILLER_282_1893 ();
 b15zdnd00an1n01x5 FILLER_282_1897 ();
 b15zdnd11an1n64x5 FILLER_282_1901 ();
 b15zdnd11an1n64x5 FILLER_282_1965 ();
 b15zdnd11an1n64x5 FILLER_282_2029 ();
 b15zdnd11an1n32x5 FILLER_282_2093 ();
 b15zdnd11an1n16x5 FILLER_282_2125 ();
 b15zdnd11an1n08x5 FILLER_282_2141 ();
 b15zdnd11an1n04x5 FILLER_282_2149 ();
 b15zdnd00an1n01x5 FILLER_282_2153 ();
 b15zdnd11an1n64x5 FILLER_282_2162 ();
 b15zdnd11an1n32x5 FILLER_282_2226 ();
 b15zdnd11an1n16x5 FILLER_282_2258 ();
 b15zdnd00an1n02x5 FILLER_282_2274 ();
 b15zdnd11an1n64x5 FILLER_283_0 ();
 b15zdnd11an1n16x5 FILLER_283_64 ();
 b15zdnd11an1n08x5 FILLER_283_80 ();
 b15zdnd11an1n04x5 FILLER_283_88 ();
 b15zdnd00an1n02x5 FILLER_283_92 ();
 b15zdnd00an1n01x5 FILLER_283_94 ();
 b15zdnd11an1n08x5 FILLER_283_137 ();
 b15zdnd00an1n02x5 FILLER_283_145 ();
 b15zdnd00an1n01x5 FILLER_283_147 ();
 b15zdnd11an1n64x5 FILLER_283_200 ();
 b15zdnd11an1n16x5 FILLER_283_264 ();
 b15zdnd11an1n04x5 FILLER_283_280 ();
 b15zdnd11an1n64x5 FILLER_283_336 ();
 b15zdnd11an1n64x5 FILLER_283_400 ();
 b15zdnd11an1n64x5 FILLER_283_464 ();
 b15zdnd11an1n64x5 FILLER_283_528 ();
 b15zdnd11an1n64x5 FILLER_283_592 ();
 b15zdnd11an1n16x5 FILLER_283_656 ();
 b15zdnd11an1n08x5 FILLER_283_672 ();
 b15zdnd11an1n08x5 FILLER_283_732 ();
 b15zdnd00an1n02x5 FILLER_283_740 ();
 b15zdnd11an1n64x5 FILLER_283_794 ();
 b15zdnd11an1n64x5 FILLER_283_858 ();
 b15zdnd11an1n64x5 FILLER_283_922 ();
 b15zdnd11an1n64x5 FILLER_283_986 ();
 b15zdnd11an1n64x5 FILLER_283_1050 ();
 b15zdnd11an1n32x5 FILLER_283_1114 ();
 b15zdnd11an1n08x5 FILLER_283_1146 ();
 b15zdnd00an1n01x5 FILLER_283_1154 ();
 b15zdnd11an1n32x5 FILLER_283_1164 ();
 b15zdnd11an1n08x5 FILLER_283_1196 ();
 b15zdnd11an1n04x5 FILLER_283_1204 ();
 b15zdnd00an1n02x5 FILLER_283_1208 ();
 b15zdnd00an1n01x5 FILLER_283_1210 ();
 b15zdnd11an1n64x5 FILLER_283_1214 ();
 b15zdnd11an1n64x5 FILLER_283_1278 ();
 b15zdnd11an1n32x5 FILLER_283_1342 ();
 b15zdnd11an1n08x5 FILLER_283_1374 ();
 b15zdnd11an1n04x5 FILLER_283_1382 ();
 b15zdnd00an1n01x5 FILLER_283_1386 ();
 b15zdnd11an1n64x5 FILLER_283_1404 ();
 b15zdnd11an1n64x5 FILLER_283_1468 ();
 b15zdnd11an1n64x5 FILLER_283_1532 ();
 b15zdnd00an1n02x5 FILLER_283_1596 ();
 b15zdnd00an1n01x5 FILLER_283_1598 ();
 b15zdnd11an1n64x5 FILLER_283_1608 ();
 b15zdnd11an1n64x5 FILLER_283_1672 ();
 b15zdnd11an1n64x5 FILLER_283_1736 ();
 b15zdnd11an1n64x5 FILLER_283_1800 ();
 b15zdnd11an1n16x5 FILLER_283_1864 ();
 b15zdnd11an1n08x5 FILLER_283_1880 ();
 b15zdnd11an1n04x5 FILLER_283_1888 ();
 b15zdnd00an1n02x5 FILLER_283_1892 ();
 b15zdnd11an1n64x5 FILLER_283_1925 ();
 b15zdnd11an1n64x5 FILLER_283_1989 ();
 b15zdnd11an1n64x5 FILLER_283_2053 ();
 b15zdnd11an1n64x5 FILLER_283_2117 ();
 b15zdnd11an1n64x5 FILLER_283_2181 ();
 b15zdnd11an1n04x5 FILLER_283_2257 ();
 b15zdnd11an1n16x5 FILLER_283_2268 ();
 b15zdnd11an1n64x5 FILLER_284_8 ();
 b15zdnd11an1n64x5 FILLER_284_72 ();
 b15zdnd11an1n16x5 FILLER_284_136 ();
 b15zdnd11an1n08x5 FILLER_284_152 ();
 b15zdnd11an1n04x5 FILLER_284_160 ();
 b15zdnd00an1n02x5 FILLER_284_164 ();
 b15zdnd11an1n04x5 FILLER_284_169 ();
 b15zdnd11an1n64x5 FILLER_284_176 ();
 b15zdnd11an1n32x5 FILLER_284_240 ();
 b15zdnd11an1n16x5 FILLER_284_272 ();
 b15zdnd11an1n08x5 FILLER_284_288 ();
 b15zdnd11an1n04x5 FILLER_284_296 ();
 b15zdnd11an1n04x5 FILLER_284_303 ();
 b15zdnd11an1n04x5 FILLER_284_310 ();
 b15zdnd11an1n64x5 FILLER_284_317 ();
 b15zdnd11an1n64x5 FILLER_284_381 ();
 b15zdnd11an1n64x5 FILLER_284_445 ();
 b15zdnd11an1n32x5 FILLER_284_509 ();
 b15zdnd11an1n64x5 FILLER_284_555 ();
 b15zdnd11an1n64x5 FILLER_284_619 ();
 b15zdnd11an1n08x5 FILLER_284_683 ();
 b15zdnd11an1n04x5 FILLER_284_691 ();
 b15zdnd00an1n02x5 FILLER_284_695 ();
 b15zdnd00an1n01x5 FILLER_284_697 ();
 b15zdnd11an1n04x5 FILLER_284_701 ();
 b15zdnd11an1n08x5 FILLER_284_708 ();
 b15zdnd00an1n02x5 FILLER_284_716 ();
 b15zdnd00an1n02x5 FILLER_284_726 ();
 b15zdnd11an1n04x5 FILLER_284_770 ();
 b15zdnd11an1n04x5 FILLER_284_777 ();
 b15zdnd00an1n01x5 FILLER_284_781 ();
 b15zdnd11an1n64x5 FILLER_284_824 ();
 b15zdnd11an1n64x5 FILLER_284_888 ();
 b15zdnd11an1n32x5 FILLER_284_952 ();
 b15zdnd11an1n16x5 FILLER_284_984 ();
 b15zdnd11an1n08x5 FILLER_284_1000 ();
 b15zdnd11an1n64x5 FILLER_284_1011 ();
 b15zdnd11an1n64x5 FILLER_284_1075 ();
 b15zdnd11an1n64x5 FILLER_284_1139 ();
 b15zdnd11an1n64x5 FILLER_284_1203 ();
 b15zdnd11an1n64x5 FILLER_284_1267 ();
 b15zdnd11an1n64x5 FILLER_284_1331 ();
 b15zdnd11an1n08x5 FILLER_284_1409 ();
 b15zdnd11an1n04x5 FILLER_284_1417 ();
 b15zdnd00an1n01x5 FILLER_284_1421 ();
 b15zdnd11an1n04x5 FILLER_284_1436 ();
 b15zdnd11an1n04x5 FILLER_284_1457 ();
 b15zdnd11an1n64x5 FILLER_284_1481 ();
 b15zdnd11an1n64x5 FILLER_284_1545 ();
 b15zdnd11an1n64x5 FILLER_284_1609 ();
 b15zdnd11an1n64x5 FILLER_284_1673 ();
 b15zdnd11an1n16x5 FILLER_284_1737 ();
 b15zdnd00an1n01x5 FILLER_284_1753 ();
 b15zdnd11an1n64x5 FILLER_284_1781 ();
 b15zdnd11an1n32x5 FILLER_284_1845 ();
 b15zdnd00an1n01x5 FILLER_284_1877 ();
 b15zdnd11an1n04x5 FILLER_284_1930 ();
 b15zdnd11an1n64x5 FILLER_284_1937 ();
 b15zdnd11an1n64x5 FILLER_284_2001 ();
 b15zdnd11an1n64x5 FILLER_284_2065 ();
 b15zdnd11an1n16x5 FILLER_284_2129 ();
 b15zdnd11an1n08x5 FILLER_284_2145 ();
 b15zdnd00an1n01x5 FILLER_284_2153 ();
 b15zdnd11an1n64x5 FILLER_284_2162 ();
 b15zdnd11an1n16x5 FILLER_284_2226 ();
 b15zdnd11an1n04x5 FILLER_284_2242 ();
 b15zdnd11an1n08x5 FILLER_284_2258 ();
 b15zdnd00an1n01x5 FILLER_284_2266 ();
 b15zdnd00an1n02x5 FILLER_284_2274 ();
 b15zdnd11an1n64x5 FILLER_285_0 ();
 b15zdnd11an1n64x5 FILLER_285_64 ();
 b15zdnd11an1n64x5 FILLER_285_128 ();
 b15zdnd11an1n64x5 FILLER_285_192 ();
 b15zdnd11an1n64x5 FILLER_285_256 ();
 b15zdnd11an1n64x5 FILLER_285_320 ();
 b15zdnd11an1n64x5 FILLER_285_384 ();
 b15zdnd11an1n64x5 FILLER_285_448 ();
 b15zdnd11an1n64x5 FILLER_285_512 ();
 b15zdnd11an1n64x5 FILLER_285_576 ();
 b15zdnd11an1n64x5 FILLER_285_640 ();
 b15zdnd11an1n32x5 FILLER_285_704 ();
 b15zdnd11an1n16x5 FILLER_285_736 ();
 b15zdnd11an1n08x5 FILLER_285_752 ();
 b15zdnd11an1n64x5 FILLER_285_763 ();
 b15zdnd11an1n64x5 FILLER_285_827 ();
 b15zdnd11an1n32x5 FILLER_285_891 ();
 b15zdnd11an1n16x5 FILLER_285_923 ();
 b15zdnd11an1n08x5 FILLER_285_939 ();
 b15zdnd00an1n02x5 FILLER_285_947 ();
 b15zdnd00an1n01x5 FILLER_285_949 ();
 b15zdnd11an1n04x5 FILLER_285_977 ();
 b15zdnd11an1n64x5 FILLER_285_1033 ();
 b15zdnd11an1n64x5 FILLER_285_1097 ();
 b15zdnd11an1n64x5 FILLER_285_1161 ();
 b15zdnd11an1n64x5 FILLER_285_1225 ();
 b15zdnd11an1n64x5 FILLER_285_1289 ();
 b15zdnd11an1n04x5 FILLER_285_1353 ();
 b15zdnd00an1n02x5 FILLER_285_1357 ();
 b15zdnd00an1n01x5 FILLER_285_1359 ();
 b15zdnd11an1n64x5 FILLER_285_1386 ();
 b15zdnd11an1n64x5 FILLER_285_1450 ();
 b15zdnd11an1n64x5 FILLER_285_1514 ();
 b15zdnd11an1n64x5 FILLER_285_1578 ();
 b15zdnd11an1n64x5 FILLER_285_1642 ();
 b15zdnd11an1n32x5 FILLER_285_1706 ();
 b15zdnd11an1n16x5 FILLER_285_1738 ();
 b15zdnd00an1n02x5 FILLER_285_1754 ();
 b15zdnd00an1n01x5 FILLER_285_1756 ();
 b15zdnd11an1n64x5 FILLER_285_1760 ();
 b15zdnd11an1n32x5 FILLER_285_1824 ();
 b15zdnd11an1n08x5 FILLER_285_1856 ();
 b15zdnd00an1n02x5 FILLER_285_1864 ();
 b15zdnd11an1n04x5 FILLER_285_1874 ();
 b15zdnd11an1n64x5 FILLER_285_1930 ();
 b15zdnd11an1n64x5 FILLER_285_1994 ();
 b15zdnd11an1n64x5 FILLER_285_2058 ();
 b15zdnd11an1n64x5 FILLER_285_2122 ();
 b15zdnd11an1n64x5 FILLER_285_2186 ();
 b15zdnd11an1n32x5 FILLER_285_2250 ();
 b15zdnd00an1n02x5 FILLER_285_2282 ();
 b15zdnd11an1n64x5 FILLER_286_8 ();
 b15zdnd11an1n64x5 FILLER_286_72 ();
 b15zdnd11an1n64x5 FILLER_286_136 ();
 b15zdnd11an1n64x5 FILLER_286_200 ();
 b15zdnd11an1n64x5 FILLER_286_264 ();
 b15zdnd11an1n64x5 FILLER_286_328 ();
 b15zdnd11an1n64x5 FILLER_286_392 ();
 b15zdnd11an1n64x5 FILLER_286_456 ();
 b15zdnd11an1n64x5 FILLER_286_520 ();
 b15zdnd11an1n64x5 FILLER_286_584 ();
 b15zdnd11an1n64x5 FILLER_286_648 ();
 b15zdnd11an1n04x5 FILLER_286_712 ();
 b15zdnd00an1n02x5 FILLER_286_716 ();
 b15zdnd11an1n64x5 FILLER_286_726 ();
 b15zdnd11an1n64x5 FILLER_286_790 ();
 b15zdnd11an1n64x5 FILLER_286_854 ();
 b15zdnd11an1n16x5 FILLER_286_918 ();
 b15zdnd11an1n08x5 FILLER_286_934 ();
 b15zdnd11an1n04x5 FILLER_286_942 ();
 b15zdnd00an1n01x5 FILLER_286_946 ();
 b15zdnd11an1n04x5 FILLER_286_950 ();
 b15zdnd11an1n32x5 FILLER_286_957 ();
 b15zdnd11an1n08x5 FILLER_286_989 ();
 b15zdnd00an1n02x5 FILLER_286_997 ();
 b15zdnd11an1n04x5 FILLER_286_1002 ();
 b15zdnd11an1n64x5 FILLER_286_1009 ();
 b15zdnd11an1n64x5 FILLER_286_1073 ();
 b15zdnd11an1n64x5 FILLER_286_1137 ();
 b15zdnd11an1n64x5 FILLER_286_1201 ();
 b15zdnd11an1n64x5 FILLER_286_1265 ();
 b15zdnd11an1n32x5 FILLER_286_1329 ();
 b15zdnd11an1n16x5 FILLER_286_1361 ();
 b15zdnd11an1n08x5 FILLER_286_1377 ();
 b15zdnd11an1n04x5 FILLER_286_1385 ();
 b15zdnd00an1n01x5 FILLER_286_1389 ();
 b15zdnd11an1n04x5 FILLER_286_1410 ();
 b15zdnd11an1n64x5 FILLER_286_1434 ();
 b15zdnd11an1n32x5 FILLER_286_1498 ();
 b15zdnd11an1n16x5 FILLER_286_1530 ();
 b15zdnd11an1n08x5 FILLER_286_1546 ();
 b15zdnd11an1n64x5 FILLER_286_1574 ();
 b15zdnd11an1n64x5 FILLER_286_1638 ();
 b15zdnd11an1n64x5 FILLER_286_1702 ();
 b15zdnd11an1n64x5 FILLER_286_1766 ();
 b15zdnd11an1n64x5 FILLER_286_1830 ();
 b15zdnd00an1n02x5 FILLER_286_1894 ();
 b15zdnd11an1n04x5 FILLER_286_1899 ();
 b15zdnd11an1n04x5 FILLER_286_1906 ();
 b15zdnd11an1n08x5 FILLER_286_1913 ();
 b15zdnd11an1n64x5 FILLER_286_1924 ();
 b15zdnd11an1n64x5 FILLER_286_1988 ();
 b15zdnd11an1n64x5 FILLER_286_2052 ();
 b15zdnd11an1n32x5 FILLER_286_2116 ();
 b15zdnd11an1n04x5 FILLER_286_2148 ();
 b15zdnd00an1n02x5 FILLER_286_2152 ();
 b15zdnd11an1n64x5 FILLER_286_2162 ();
 b15zdnd11an1n32x5 FILLER_286_2226 ();
 b15zdnd11an1n16x5 FILLER_286_2258 ();
 b15zdnd00an1n02x5 FILLER_286_2274 ();
 b15zdnd11an1n64x5 FILLER_287_0 ();
 b15zdnd11an1n64x5 FILLER_287_64 ();
 b15zdnd11an1n64x5 FILLER_287_128 ();
 b15zdnd11an1n64x5 FILLER_287_192 ();
 b15zdnd11an1n64x5 FILLER_287_256 ();
 b15zdnd11an1n64x5 FILLER_287_320 ();
 b15zdnd11an1n64x5 FILLER_287_384 ();
 b15zdnd11an1n64x5 FILLER_287_448 ();
 b15zdnd11an1n32x5 FILLER_287_512 ();
 b15zdnd11an1n16x5 FILLER_287_544 ();
 b15zdnd11an1n08x5 FILLER_287_560 ();
 b15zdnd00an1n02x5 FILLER_287_568 ();
 b15zdnd00an1n01x5 FILLER_287_570 ();
 b15zdnd11an1n64x5 FILLER_287_580 ();
 b15zdnd11an1n64x5 FILLER_287_644 ();
 b15zdnd11an1n64x5 FILLER_287_708 ();
 b15zdnd11an1n64x5 FILLER_287_772 ();
 b15zdnd11an1n64x5 FILLER_287_836 ();
 b15zdnd11an1n16x5 FILLER_287_900 ();
 b15zdnd11an1n04x5 FILLER_287_916 ();
 b15zdnd00an1n02x5 FILLER_287_920 ();
 b15zdnd11an1n64x5 FILLER_287_974 ();
 b15zdnd11an1n64x5 FILLER_287_1038 ();
 b15zdnd11an1n64x5 FILLER_287_1102 ();
 b15zdnd11an1n64x5 FILLER_287_1166 ();
 b15zdnd11an1n64x5 FILLER_287_1230 ();
 b15zdnd11an1n64x5 FILLER_287_1294 ();
 b15zdnd11an1n64x5 FILLER_287_1358 ();
 b15zdnd11an1n64x5 FILLER_287_1422 ();
 b15zdnd11an1n64x5 FILLER_287_1486 ();
 b15zdnd11an1n64x5 FILLER_287_1550 ();
 b15zdnd11an1n64x5 FILLER_287_1614 ();
 b15zdnd11an1n64x5 FILLER_287_1678 ();
 b15zdnd11an1n64x5 FILLER_287_1742 ();
 b15zdnd11an1n64x5 FILLER_287_1806 ();
 b15zdnd11an1n64x5 FILLER_287_1870 ();
 b15zdnd11an1n64x5 FILLER_287_1934 ();
 b15zdnd11an1n64x5 FILLER_287_1998 ();
 b15zdnd11an1n64x5 FILLER_287_2062 ();
 b15zdnd11an1n64x5 FILLER_287_2126 ();
 b15zdnd11an1n64x5 FILLER_287_2190 ();
 b15zdnd11an1n16x5 FILLER_287_2254 ();
 b15zdnd11an1n08x5 FILLER_287_2270 ();
 b15zdnd11an1n04x5 FILLER_287_2278 ();
 b15zdnd00an1n02x5 FILLER_287_2282 ();
 b15zdnd11an1n64x5 FILLER_288_8 ();
 b15zdnd11an1n64x5 FILLER_288_72 ();
 b15zdnd11an1n64x5 FILLER_288_136 ();
 b15zdnd11an1n16x5 FILLER_288_200 ();
 b15zdnd11an1n08x5 FILLER_288_216 ();
 b15zdnd11an1n04x5 FILLER_288_224 ();
 b15zdnd00an1n01x5 FILLER_288_228 ();
 b15zdnd11an1n04x5 FILLER_288_232 ();
 b15zdnd11an1n64x5 FILLER_288_239 ();
 b15zdnd11an1n64x5 FILLER_288_303 ();
 b15zdnd11an1n64x5 FILLER_288_367 ();
 b15zdnd11an1n64x5 FILLER_288_431 ();
 b15zdnd11an1n08x5 FILLER_288_495 ();
 b15zdnd00an1n02x5 FILLER_288_503 ();
 b15zdnd11an1n64x5 FILLER_288_521 ();
 b15zdnd11an1n16x5 FILLER_288_585 ();
 b15zdnd11an1n04x5 FILLER_288_601 ();
 b15zdnd00an1n02x5 FILLER_288_605 ();
 b15zdnd00an1n01x5 FILLER_288_607 ();
 b15zdnd11an1n64x5 FILLER_288_611 ();
 b15zdnd11an1n32x5 FILLER_288_675 ();
 b15zdnd11an1n08x5 FILLER_288_707 ();
 b15zdnd00an1n02x5 FILLER_288_715 ();
 b15zdnd00an1n01x5 FILLER_288_717 ();
 b15zdnd11an1n64x5 FILLER_288_726 ();
 b15zdnd11an1n64x5 FILLER_288_790 ();
 b15zdnd11an1n64x5 FILLER_288_854 ();
 b15zdnd11an1n08x5 FILLER_288_918 ();
 b15zdnd11an1n04x5 FILLER_288_926 ();
 b15zdnd00an1n02x5 FILLER_288_930 ();
 b15zdnd00an1n01x5 FILLER_288_932 ();
 b15zdnd11an1n08x5 FILLER_288_936 ();
 b15zdnd11an1n64x5 FILLER_288_947 ();
 b15zdnd11an1n64x5 FILLER_288_1011 ();
 b15zdnd11an1n64x5 FILLER_288_1075 ();
 b15zdnd11an1n64x5 FILLER_288_1139 ();
 b15zdnd11an1n64x5 FILLER_288_1203 ();
 b15zdnd11an1n64x5 FILLER_288_1267 ();
 b15zdnd11an1n64x5 FILLER_288_1331 ();
 b15zdnd11an1n64x5 FILLER_288_1395 ();
 b15zdnd11an1n64x5 FILLER_288_1459 ();
 b15zdnd11an1n64x5 FILLER_288_1523 ();
 b15zdnd11an1n64x5 FILLER_288_1587 ();
 b15zdnd11an1n64x5 FILLER_288_1651 ();
 b15zdnd11an1n64x5 FILLER_288_1715 ();
 b15zdnd11an1n64x5 FILLER_288_1779 ();
 b15zdnd11an1n64x5 FILLER_288_1843 ();
 b15zdnd11an1n64x5 FILLER_288_1907 ();
 b15zdnd11an1n64x5 FILLER_288_1971 ();
 b15zdnd11an1n64x5 FILLER_288_2035 ();
 b15zdnd11an1n32x5 FILLER_288_2099 ();
 b15zdnd11an1n16x5 FILLER_288_2131 ();
 b15zdnd11an1n04x5 FILLER_288_2147 ();
 b15zdnd00an1n02x5 FILLER_288_2151 ();
 b15zdnd00an1n01x5 FILLER_288_2153 ();
 b15zdnd11an1n64x5 FILLER_288_2162 ();
 b15zdnd11an1n32x5 FILLER_288_2226 ();
 b15zdnd11an1n16x5 FILLER_288_2258 ();
 b15zdnd00an1n02x5 FILLER_288_2274 ();
 b15zdnd11an1n64x5 FILLER_289_0 ();
 b15zdnd11an1n64x5 FILLER_289_64 ();
 b15zdnd11an1n64x5 FILLER_289_128 ();
 b15zdnd11an1n16x5 FILLER_289_192 ();
 b15zdnd00an1n01x5 FILLER_289_208 ();
 b15zdnd11an1n64x5 FILLER_289_261 ();
 b15zdnd11an1n64x5 FILLER_289_325 ();
 b15zdnd11an1n64x5 FILLER_289_389 ();
 b15zdnd11an1n64x5 FILLER_289_453 ();
 b15zdnd11an1n64x5 FILLER_289_517 ();
 b15zdnd11an1n64x5 FILLER_289_581 ();
 b15zdnd11an1n64x5 FILLER_289_645 ();
 b15zdnd11an1n64x5 FILLER_289_709 ();
 b15zdnd11an1n64x5 FILLER_289_773 ();
 b15zdnd11an1n16x5 FILLER_289_837 ();
 b15zdnd11an1n08x5 FILLER_289_853 ();
 b15zdnd11an1n04x5 FILLER_289_861 ();
 b15zdnd11an1n64x5 FILLER_289_907 ();
 b15zdnd11an1n64x5 FILLER_289_971 ();
 b15zdnd11an1n64x5 FILLER_289_1035 ();
 b15zdnd11an1n64x5 FILLER_289_1099 ();
 b15zdnd11an1n32x5 FILLER_289_1163 ();
 b15zdnd11an1n04x5 FILLER_289_1195 ();
 b15zdnd00an1n02x5 FILLER_289_1199 ();
 b15zdnd11an1n04x5 FILLER_289_1204 ();
 b15zdnd00an1n02x5 FILLER_289_1208 ();
 b15zdnd11an1n04x5 FILLER_289_1218 ();
 b15zdnd11an1n08x5 FILLER_289_1225 ();
 b15zdnd00an1n02x5 FILLER_289_1233 ();
 b15zdnd00an1n01x5 FILLER_289_1235 ();
 b15zdnd11an1n64x5 FILLER_289_1244 ();
 b15zdnd11an1n64x5 FILLER_289_1308 ();
 b15zdnd11an1n16x5 FILLER_289_1372 ();
 b15zdnd11an1n08x5 FILLER_289_1388 ();
 b15zdnd00an1n01x5 FILLER_289_1396 ();
 b15zdnd11an1n04x5 FILLER_289_1409 ();
 b15zdnd11an1n32x5 FILLER_289_1433 ();
 b15zdnd11an1n16x5 FILLER_289_1465 ();
 b15zdnd11an1n08x5 FILLER_289_1481 ();
 b15zdnd11an1n04x5 FILLER_289_1489 ();
 b15zdnd00an1n02x5 FILLER_289_1493 ();
 b15zdnd11an1n64x5 FILLER_289_1512 ();
 b15zdnd11an1n64x5 FILLER_289_1576 ();
 b15zdnd11an1n64x5 FILLER_289_1640 ();
 b15zdnd11an1n64x5 FILLER_289_1704 ();
 b15zdnd11an1n64x5 FILLER_289_1768 ();
 b15zdnd11an1n64x5 FILLER_289_1832 ();
 b15zdnd11an1n64x5 FILLER_289_1896 ();
 b15zdnd11an1n64x5 FILLER_289_1960 ();
 b15zdnd11an1n64x5 FILLER_289_2024 ();
 b15zdnd11an1n64x5 FILLER_289_2088 ();
 b15zdnd11an1n64x5 FILLER_289_2152 ();
 b15zdnd11an1n64x5 FILLER_289_2216 ();
 b15zdnd11an1n04x5 FILLER_289_2280 ();
 b15zdnd11an1n32x5 FILLER_290_8 ();
 b15zdnd11an1n16x5 FILLER_290_40 ();
 b15zdnd11an1n04x5 FILLER_290_56 ();
 b15zdnd00an1n02x5 FILLER_290_60 ();
 b15zdnd00an1n01x5 FILLER_290_62 ();
 b15zdnd11an1n04x5 FILLER_290_66 ();
 b15zdnd11an1n64x5 FILLER_290_81 ();
 b15zdnd11an1n64x5 FILLER_290_145 ();
 b15zdnd11an1n16x5 FILLER_290_209 ();
 b15zdnd00an1n02x5 FILLER_290_225 ();
 b15zdnd11an1n04x5 FILLER_290_230 ();
 b15zdnd11an1n64x5 FILLER_290_237 ();
 b15zdnd11an1n64x5 FILLER_290_301 ();
 b15zdnd11an1n64x5 FILLER_290_365 ();
 b15zdnd11an1n64x5 FILLER_290_429 ();
 b15zdnd11an1n32x5 FILLER_290_493 ();
 b15zdnd11an1n16x5 FILLER_290_525 ();
 b15zdnd11an1n04x5 FILLER_290_541 ();
 b15zdnd11an1n32x5 FILLER_290_561 ();
 b15zdnd11an1n08x5 FILLER_290_593 ();
 b15zdnd11an1n04x5 FILLER_290_601 ();
 b15zdnd00an1n01x5 FILLER_290_605 ();
 b15zdnd11an1n32x5 FILLER_290_615 ();
 b15zdnd11an1n08x5 FILLER_290_647 ();
 b15zdnd00an1n02x5 FILLER_290_655 ();
 b15zdnd11an1n32x5 FILLER_290_666 ();
 b15zdnd11an1n16x5 FILLER_290_698 ();
 b15zdnd11an1n04x5 FILLER_290_714 ();
 b15zdnd11an1n64x5 FILLER_290_726 ();
 b15zdnd11an1n32x5 FILLER_290_790 ();
 b15zdnd00an1n02x5 FILLER_290_822 ();
 b15zdnd00an1n01x5 FILLER_290_824 ();
 b15zdnd11an1n64x5 FILLER_290_877 ();
 b15zdnd11an1n64x5 FILLER_290_941 ();
 b15zdnd11an1n64x5 FILLER_290_1005 ();
 b15zdnd11an1n32x5 FILLER_290_1069 ();
 b15zdnd11an1n16x5 FILLER_290_1101 ();
 b15zdnd11an1n08x5 FILLER_290_1117 ();
 b15zdnd11an1n04x5 FILLER_290_1125 ();
 b15zdnd00an1n01x5 FILLER_290_1129 ();
 b15zdnd11an1n16x5 FILLER_290_1150 ();
 b15zdnd11an1n08x5 FILLER_290_1166 ();
 b15zdnd11an1n04x5 FILLER_290_1174 ();
 b15zdnd11an1n04x5 FILLER_290_1230 ();
 b15zdnd11an1n64x5 FILLER_290_1237 ();
 b15zdnd11an1n64x5 FILLER_290_1301 ();
 b15zdnd11an1n32x5 FILLER_290_1365 ();
 b15zdnd11an1n16x5 FILLER_290_1397 ();
 b15zdnd00an1n02x5 FILLER_290_1413 ();
 b15zdnd00an1n01x5 FILLER_290_1415 ();
 b15zdnd11an1n16x5 FILLER_290_1436 ();
 b15zdnd11an1n08x5 FILLER_290_1452 ();
 b15zdnd00an1n02x5 FILLER_290_1460 ();
 b15zdnd00an1n01x5 FILLER_290_1462 ();
 b15zdnd11an1n64x5 FILLER_290_1474 ();
 b15zdnd11an1n64x5 FILLER_290_1538 ();
 b15zdnd11an1n64x5 FILLER_290_1602 ();
 b15zdnd11an1n64x5 FILLER_290_1666 ();
 b15zdnd11an1n64x5 FILLER_290_1730 ();
 b15zdnd11an1n64x5 FILLER_290_1794 ();
 b15zdnd11an1n64x5 FILLER_290_1858 ();
 b15zdnd11an1n64x5 FILLER_290_1922 ();
 b15zdnd11an1n64x5 FILLER_290_1986 ();
 b15zdnd11an1n64x5 FILLER_290_2050 ();
 b15zdnd11an1n32x5 FILLER_290_2114 ();
 b15zdnd11an1n08x5 FILLER_290_2146 ();
 b15zdnd11an1n64x5 FILLER_290_2162 ();
 b15zdnd11an1n32x5 FILLER_290_2226 ();
 b15zdnd11an1n16x5 FILLER_290_2258 ();
 b15zdnd00an1n02x5 FILLER_290_2274 ();
 b15zdnd11an1n32x5 FILLER_291_0 ();
 b15zdnd11an1n16x5 FILLER_291_32 ();
 b15zdnd11an1n08x5 FILLER_291_48 ();
 b15zdnd11an1n04x5 FILLER_291_60 ();
 b15zdnd11an1n04x5 FILLER_291_80 ();
 b15zdnd11an1n64x5 FILLER_291_89 ();
 b15zdnd11an1n64x5 FILLER_291_153 ();
 b15zdnd11an1n64x5 FILLER_291_217 ();
 b15zdnd11an1n64x5 FILLER_291_281 ();
 b15zdnd11an1n64x5 FILLER_291_345 ();
 b15zdnd11an1n64x5 FILLER_291_409 ();
 b15zdnd11an1n64x5 FILLER_291_473 ();
 b15zdnd11an1n64x5 FILLER_291_537 ();
 b15zdnd11an1n08x5 FILLER_291_601 ();
 b15zdnd00an1n02x5 FILLER_291_609 ();
 b15zdnd00an1n01x5 FILLER_291_611 ();
 b15zdnd11an1n64x5 FILLER_291_616 ();
 b15zdnd11an1n64x5 FILLER_291_680 ();
 b15zdnd11an1n64x5 FILLER_291_744 ();
 b15zdnd11an1n16x5 FILLER_291_808 ();
 b15zdnd11an1n08x5 FILLER_291_824 ();
 b15zdnd11an1n04x5 FILLER_291_832 ();
 b15zdnd11an1n64x5 FILLER_291_878 ();
 b15zdnd11an1n32x5 FILLER_291_942 ();
 b15zdnd11an1n16x5 FILLER_291_974 ();
 b15zdnd11an1n04x5 FILLER_291_990 ();
 b15zdnd00an1n02x5 FILLER_291_994 ();
 b15zdnd00an1n01x5 FILLER_291_996 ();
 b15zdnd11an1n64x5 FILLER_291_1049 ();
 b15zdnd11an1n16x5 FILLER_291_1113 ();
 b15zdnd00an1n01x5 FILLER_291_1129 ();
 b15zdnd11an1n32x5 FILLER_291_1133 ();
 b15zdnd11an1n16x5 FILLER_291_1165 ();
 b15zdnd11an1n08x5 FILLER_291_1181 ();
 b15zdnd11an1n04x5 FILLER_291_1189 ();
 b15zdnd00an1n02x5 FILLER_291_1193 ();
 b15zdnd11an1n04x5 FILLER_291_1198 ();
 b15zdnd11an1n04x5 FILLER_291_1254 ();
 b15zdnd00an1n01x5 FILLER_291_1258 ();
 b15zdnd11an1n64x5 FILLER_291_1270 ();
 b15zdnd11an1n64x5 FILLER_291_1334 ();
 b15zdnd11an1n64x5 FILLER_291_1398 ();
 b15zdnd00an1n02x5 FILLER_291_1462 ();
 b15zdnd00an1n01x5 FILLER_291_1464 ();
 b15zdnd11an1n64x5 FILLER_291_1479 ();
 b15zdnd11an1n32x5 FILLER_291_1543 ();
 b15zdnd11an1n16x5 FILLER_291_1575 ();
 b15zdnd11an1n04x5 FILLER_291_1591 ();
 b15zdnd00an1n02x5 FILLER_291_1595 ();
 b15zdnd11an1n64x5 FILLER_291_1606 ();
 b15zdnd11an1n64x5 FILLER_291_1670 ();
 b15zdnd11an1n32x5 FILLER_291_1734 ();
 b15zdnd11an1n04x5 FILLER_291_1766 ();
 b15zdnd11an1n64x5 FILLER_291_1773 ();
 b15zdnd11an1n64x5 FILLER_291_1837 ();
 b15zdnd11an1n64x5 FILLER_291_1901 ();
 b15zdnd11an1n64x5 FILLER_291_1965 ();
 b15zdnd11an1n64x5 FILLER_291_2029 ();
 b15zdnd11an1n64x5 FILLER_291_2093 ();
 b15zdnd11an1n64x5 FILLER_291_2157 ();
 b15zdnd11an1n32x5 FILLER_291_2221 ();
 b15zdnd11an1n16x5 FILLER_291_2253 ();
 b15zdnd11an1n08x5 FILLER_291_2269 ();
 b15zdnd11an1n04x5 FILLER_291_2277 ();
 b15zdnd00an1n02x5 FILLER_291_2281 ();
 b15zdnd00an1n01x5 FILLER_291_2283 ();
 b15zdnd11an1n32x5 FILLER_292_8 ();
 b15zdnd11an1n08x5 FILLER_292_40 ();
 b15zdnd11an1n04x5 FILLER_292_48 ();
 b15zdnd00an1n01x5 FILLER_292_52 ();
 b15zdnd11an1n04x5 FILLER_292_71 ();
 b15zdnd11an1n04x5 FILLER_292_79 ();
 b15zdnd00an1n02x5 FILLER_292_83 ();
 b15zdnd11an1n64x5 FILLER_292_90 ();
 b15zdnd11an1n64x5 FILLER_292_154 ();
 b15zdnd11an1n64x5 FILLER_292_218 ();
 b15zdnd11an1n16x5 FILLER_292_282 ();
 b15zdnd11an1n08x5 FILLER_292_298 ();
 b15zdnd11an1n04x5 FILLER_292_306 ();
 b15zdnd11an1n08x5 FILLER_292_317 ();
 b15zdnd00an1n02x5 FILLER_292_325 ();
 b15zdnd00an1n01x5 FILLER_292_327 ();
 b15zdnd11an1n64x5 FILLER_292_335 ();
 b15zdnd11an1n32x5 FILLER_292_399 ();
 b15zdnd00an1n01x5 FILLER_292_431 ();
 b15zdnd11an1n64x5 FILLER_292_441 ();
 b15zdnd11an1n64x5 FILLER_292_505 ();
 b15zdnd11an1n64x5 FILLER_292_569 ();
 b15zdnd11an1n64x5 FILLER_292_633 ();
 b15zdnd11an1n16x5 FILLER_292_697 ();
 b15zdnd11an1n04x5 FILLER_292_713 ();
 b15zdnd00an1n01x5 FILLER_292_717 ();
 b15zdnd11an1n64x5 FILLER_292_726 ();
 b15zdnd11an1n32x5 FILLER_292_790 ();
 b15zdnd11an1n16x5 FILLER_292_822 ();
 b15zdnd11an1n04x5 FILLER_292_838 ();
 b15zdnd00an1n02x5 FILLER_292_842 ();
 b15zdnd00an1n01x5 FILLER_292_844 ();
 b15zdnd11an1n04x5 FILLER_292_848 ();
 b15zdnd11an1n04x5 FILLER_292_855 ();
 b15zdnd11an1n64x5 FILLER_292_862 ();
 b15zdnd11an1n64x5 FILLER_292_926 ();
 b15zdnd11an1n16x5 FILLER_292_990 ();
 b15zdnd11an1n08x5 FILLER_292_1006 ();
 b15zdnd11an1n04x5 FILLER_292_1014 ();
 b15zdnd00an1n01x5 FILLER_292_1018 ();
 b15zdnd11an1n04x5 FILLER_292_1022 ();
 b15zdnd11an1n16x5 FILLER_292_1029 ();
 b15zdnd00an1n01x5 FILLER_292_1045 ();
 b15zdnd11an1n04x5 FILLER_292_1066 ();
 b15zdnd11an1n08x5 FILLER_292_1090 ();
 b15zdnd11an1n04x5 FILLER_292_1098 ();
 b15zdnd11an1n08x5 FILLER_292_1113 ();
 b15zdnd00an1n02x5 FILLER_292_1121 ();
 b15zdnd00an1n01x5 FILLER_292_1123 ();
 b15zdnd11an1n04x5 FILLER_292_1127 ();
 b15zdnd11an1n64x5 FILLER_292_1134 ();
 b15zdnd11an1n04x5 FILLER_292_1198 ();
 b15zdnd00an1n01x5 FILLER_292_1202 ();
 b15zdnd11an1n16x5 FILLER_292_1206 ();
 b15zdnd00an1n02x5 FILLER_292_1222 ();
 b15zdnd00an1n01x5 FILLER_292_1224 ();
 b15zdnd11an1n64x5 FILLER_292_1228 ();
 b15zdnd11an1n64x5 FILLER_292_1292 ();
 b15zdnd11an1n64x5 FILLER_292_1356 ();
 b15zdnd11an1n64x5 FILLER_292_1420 ();
 b15zdnd11an1n64x5 FILLER_292_1484 ();
 b15zdnd11an1n32x5 FILLER_292_1548 ();
 b15zdnd11an1n16x5 FILLER_292_1580 ();
 b15zdnd00an1n02x5 FILLER_292_1596 ();
 b15zdnd00an1n01x5 FILLER_292_1598 ();
 b15zdnd11an1n64x5 FILLER_292_1608 ();
 b15zdnd11an1n64x5 FILLER_292_1672 ();
 b15zdnd11an1n32x5 FILLER_292_1736 ();
 b15zdnd00an1n01x5 FILLER_292_1768 ();
 b15zdnd11an1n32x5 FILLER_292_1772 ();
 b15zdnd11an1n16x5 FILLER_292_1804 ();
 b15zdnd00an1n01x5 FILLER_292_1820 ();
 b15zdnd11an1n16x5 FILLER_292_1830 ();
 b15zdnd00an1n02x5 FILLER_292_1846 ();
 b15zdnd00an1n01x5 FILLER_292_1848 ();
 b15zdnd11an1n32x5 FILLER_292_1858 ();
 b15zdnd11an1n04x5 FILLER_292_1890 ();
 b15zdnd00an1n02x5 FILLER_292_1894 ();
 b15zdnd11an1n64x5 FILLER_292_1938 ();
 b15zdnd11an1n64x5 FILLER_292_2002 ();
 b15zdnd11an1n64x5 FILLER_292_2066 ();
 b15zdnd11an1n16x5 FILLER_292_2130 ();
 b15zdnd11an1n08x5 FILLER_292_2146 ();
 b15zdnd11an1n64x5 FILLER_292_2162 ();
 b15zdnd11an1n32x5 FILLER_292_2226 ();
 b15zdnd11an1n16x5 FILLER_292_2258 ();
 b15zdnd00an1n02x5 FILLER_292_2274 ();
 b15zdnd11an1n32x5 FILLER_293_0 ();
 b15zdnd11an1n16x5 FILLER_293_32 ();
 b15zdnd11an1n08x5 FILLER_293_48 ();
 b15zdnd11an1n04x5 FILLER_293_56 ();
 b15zdnd11an1n64x5 FILLER_293_76 ();
 b15zdnd11an1n64x5 FILLER_293_140 ();
 b15zdnd11an1n64x5 FILLER_293_204 ();
 b15zdnd11an1n32x5 FILLER_293_268 ();
 b15zdnd11an1n16x5 FILLER_293_300 ();
 b15zdnd11an1n08x5 FILLER_293_316 ();
 b15zdnd11an1n04x5 FILLER_293_324 ();
 b15zdnd11an1n64x5 FILLER_293_344 ();
 b15zdnd11an1n64x5 FILLER_293_408 ();
 b15zdnd11an1n64x5 FILLER_293_472 ();
 b15zdnd11an1n64x5 FILLER_293_536 ();
 b15zdnd11an1n64x5 FILLER_293_600 ();
 b15zdnd11an1n64x5 FILLER_293_664 ();
 b15zdnd11an1n64x5 FILLER_293_728 ();
 b15zdnd11an1n64x5 FILLER_293_792 ();
 b15zdnd11an1n04x5 FILLER_293_856 ();
 b15zdnd00an1n01x5 FILLER_293_860 ();
 b15zdnd11an1n08x5 FILLER_293_864 ();
 b15zdnd00an1n02x5 FILLER_293_872 ();
 b15zdnd11an1n64x5 FILLER_293_916 ();
 b15zdnd11an1n32x5 FILLER_293_980 ();
 b15zdnd11an1n04x5 FILLER_293_1012 ();
 b15zdnd11an1n64x5 FILLER_293_1019 ();
 b15zdnd11an1n04x5 FILLER_293_1083 ();
 b15zdnd11an1n04x5 FILLER_293_1139 ();
 b15zdnd11an1n64x5 FILLER_293_1154 ();
 b15zdnd11an1n16x5 FILLER_293_1218 ();
 b15zdnd11an1n08x5 FILLER_293_1234 ();
 b15zdnd00an1n02x5 FILLER_293_1242 ();
 b15zdnd11an1n64x5 FILLER_293_1255 ();
 b15zdnd11an1n64x5 FILLER_293_1319 ();
 b15zdnd11an1n32x5 FILLER_293_1383 ();
 b15zdnd11an1n16x5 FILLER_293_1415 ();
 b15zdnd11an1n04x5 FILLER_293_1431 ();
 b15zdnd11an1n64x5 FILLER_293_1447 ();
 b15zdnd11an1n64x5 FILLER_293_1511 ();
 b15zdnd11an1n64x5 FILLER_293_1575 ();
 b15zdnd11an1n64x5 FILLER_293_1639 ();
 b15zdnd11an1n04x5 FILLER_293_1703 ();
 b15zdnd00an1n02x5 FILLER_293_1707 ();
 b15zdnd11an1n04x5 FILLER_293_1740 ();
 b15zdnd11an1n64x5 FILLER_293_1796 ();
 b15zdnd11an1n64x5 FILLER_293_1860 ();
 b15zdnd11an1n64x5 FILLER_293_1924 ();
 b15zdnd11an1n64x5 FILLER_293_1988 ();
 b15zdnd11an1n64x5 FILLER_293_2052 ();
 b15zdnd11an1n64x5 FILLER_293_2116 ();
 b15zdnd11an1n64x5 FILLER_293_2180 ();
 b15zdnd11an1n32x5 FILLER_293_2244 ();
 b15zdnd11an1n08x5 FILLER_293_2276 ();
 b15zdnd11an1n32x5 FILLER_294_8 ();
 b15zdnd11an1n08x5 FILLER_294_40 ();
 b15zdnd11an1n04x5 FILLER_294_48 ();
 b15zdnd00an1n02x5 FILLER_294_52 ();
 b15zdnd00an1n01x5 FILLER_294_54 ();
 b15zdnd11an1n04x5 FILLER_294_61 ();
 b15zdnd11an1n64x5 FILLER_294_73 ();
 b15zdnd11an1n64x5 FILLER_294_137 ();
 b15zdnd11an1n64x5 FILLER_294_201 ();
 b15zdnd11an1n64x5 FILLER_294_265 ();
 b15zdnd11an1n64x5 FILLER_294_329 ();
 b15zdnd11an1n32x5 FILLER_294_393 ();
 b15zdnd00an1n02x5 FILLER_294_425 ();
 b15zdnd00an1n01x5 FILLER_294_427 ();
 b15zdnd11an1n04x5 FILLER_294_431 ();
 b15zdnd11an1n64x5 FILLER_294_438 ();
 b15zdnd11an1n32x5 FILLER_294_502 ();
 b15zdnd00an1n02x5 FILLER_294_534 ();
 b15zdnd11an1n64x5 FILLER_294_540 ();
 b15zdnd11an1n64x5 FILLER_294_604 ();
 b15zdnd11an1n32x5 FILLER_294_668 ();
 b15zdnd11an1n16x5 FILLER_294_700 ();
 b15zdnd00an1n02x5 FILLER_294_716 ();
 b15zdnd11an1n64x5 FILLER_294_726 ();
 b15zdnd11an1n32x5 FILLER_294_790 ();
 b15zdnd11an1n08x5 FILLER_294_822 ();
 b15zdnd11an1n04x5 FILLER_294_830 ();
 b15zdnd11an1n64x5 FILLER_294_886 ();
 b15zdnd11an1n64x5 FILLER_294_950 ();
 b15zdnd11an1n64x5 FILLER_294_1014 ();
 b15zdnd11an1n16x5 FILLER_294_1078 ();
 b15zdnd11an1n08x5 FILLER_294_1094 ();
 b15zdnd00an1n02x5 FILLER_294_1102 ();
 b15zdnd00an1n01x5 FILLER_294_1104 ();
 b15zdnd11an1n64x5 FILLER_294_1157 ();
 b15zdnd11an1n64x5 FILLER_294_1221 ();
 b15zdnd11an1n64x5 FILLER_294_1285 ();
 b15zdnd11an1n64x5 FILLER_294_1349 ();
 b15zdnd11an1n32x5 FILLER_294_1413 ();
 b15zdnd11an1n04x5 FILLER_294_1445 ();
 b15zdnd00an1n02x5 FILLER_294_1449 ();
 b15zdnd00an1n01x5 FILLER_294_1451 ();
 b15zdnd11an1n64x5 FILLER_294_1472 ();
 b15zdnd11an1n64x5 FILLER_294_1536 ();
 b15zdnd11an1n64x5 FILLER_294_1600 ();
 b15zdnd11an1n64x5 FILLER_294_1664 ();
 b15zdnd11an1n32x5 FILLER_294_1728 ();
 b15zdnd00an1n02x5 FILLER_294_1760 ();
 b15zdnd00an1n01x5 FILLER_294_1762 ();
 b15zdnd11an1n04x5 FILLER_294_1766 ();
 b15zdnd11an1n64x5 FILLER_294_1773 ();
 b15zdnd11an1n08x5 FILLER_294_1837 ();
 b15zdnd11an1n64x5 FILLER_294_1854 ();
 b15zdnd11an1n64x5 FILLER_294_1918 ();
 b15zdnd11an1n64x5 FILLER_294_1982 ();
 b15zdnd11an1n64x5 FILLER_294_2046 ();
 b15zdnd11an1n32x5 FILLER_294_2110 ();
 b15zdnd11an1n08x5 FILLER_294_2142 ();
 b15zdnd11an1n04x5 FILLER_294_2150 ();
 b15zdnd11an1n64x5 FILLER_294_2162 ();
 b15zdnd11an1n32x5 FILLER_294_2226 ();
 b15zdnd11an1n16x5 FILLER_294_2258 ();
 b15zdnd00an1n02x5 FILLER_294_2274 ();
 b15zdnd11an1n64x5 FILLER_295_0 ();
 b15zdnd00an1n01x5 FILLER_295_64 ();
 b15zdnd11an1n64x5 FILLER_295_71 ();
 b15zdnd11an1n64x5 FILLER_295_135 ();
 b15zdnd11an1n64x5 FILLER_295_199 ();
 b15zdnd11an1n08x5 FILLER_295_263 ();
 b15zdnd11an1n04x5 FILLER_295_271 ();
 b15zdnd00an1n02x5 FILLER_295_275 ();
 b15zdnd11an1n16x5 FILLER_295_284 ();
 b15zdnd11an1n08x5 FILLER_295_300 ();
 b15zdnd11an1n64x5 FILLER_295_311 ();
 b15zdnd11an1n32x5 FILLER_295_375 ();
 b15zdnd00an1n01x5 FILLER_295_407 ();
 b15zdnd11an1n64x5 FILLER_295_460 ();
 b15zdnd11an1n64x5 FILLER_295_524 ();
 b15zdnd11an1n32x5 FILLER_295_588 ();
 b15zdnd00an1n01x5 FILLER_295_620 ();
 b15zdnd11an1n16x5 FILLER_295_637 ();
 b15zdnd11an1n08x5 FILLER_295_653 ();
 b15zdnd00an1n01x5 FILLER_295_661 ();
 b15zdnd11an1n64x5 FILLER_295_674 ();
 b15zdnd11an1n64x5 FILLER_295_738 ();
 b15zdnd11an1n32x5 FILLER_295_802 ();
 b15zdnd11an1n08x5 FILLER_295_834 ();
 b15zdnd00an1n02x5 FILLER_295_842 ();
 b15zdnd00an1n01x5 FILLER_295_844 ();
 b15zdnd11an1n64x5 FILLER_295_887 ();
 b15zdnd11an1n64x5 FILLER_295_951 ();
 b15zdnd11an1n64x5 FILLER_295_1015 ();
 b15zdnd11an1n16x5 FILLER_295_1079 ();
 b15zdnd11an1n08x5 FILLER_295_1095 ();
 b15zdnd00an1n02x5 FILLER_295_1103 ();
 b15zdnd00an1n01x5 FILLER_295_1105 ();
 b15zdnd11an1n04x5 FILLER_295_1109 ();
 b15zdnd11an1n16x5 FILLER_295_1116 ();
 b15zdnd11an1n08x5 FILLER_295_1132 ();
 b15zdnd00an1n02x5 FILLER_295_1140 ();
 b15zdnd00an1n01x5 FILLER_295_1142 ();
 b15zdnd11an1n64x5 FILLER_295_1154 ();
 b15zdnd11an1n64x5 FILLER_295_1218 ();
 b15zdnd11an1n64x5 FILLER_295_1282 ();
 b15zdnd11an1n08x5 FILLER_295_1346 ();
 b15zdnd00an1n02x5 FILLER_295_1354 ();
 b15zdnd11an1n32x5 FILLER_295_1373 ();
 b15zdnd11an1n08x5 FILLER_295_1405 ();
 b15zdnd11an1n04x5 FILLER_295_1413 ();
 b15zdnd00an1n01x5 FILLER_295_1417 ();
 b15zdnd11an1n16x5 FILLER_295_1432 ();
 b15zdnd00an1n02x5 FILLER_295_1448 ();
 b15zdnd11an1n64x5 FILLER_295_1470 ();
 b15zdnd11an1n64x5 FILLER_295_1534 ();
 b15zdnd11an1n64x5 FILLER_295_1598 ();
 b15zdnd11an1n64x5 FILLER_295_1662 ();
 b15zdnd11an1n16x5 FILLER_295_1726 ();
 b15zdnd00an1n01x5 FILLER_295_1742 ();
 b15zdnd11an1n64x5 FILLER_295_1795 ();
 b15zdnd11an1n64x5 FILLER_295_1859 ();
 b15zdnd11an1n64x5 FILLER_295_1923 ();
 b15zdnd11an1n64x5 FILLER_295_1987 ();
 b15zdnd11an1n64x5 FILLER_295_2051 ();
 b15zdnd11an1n64x5 FILLER_295_2115 ();
 b15zdnd11an1n64x5 FILLER_295_2179 ();
 b15zdnd11an1n32x5 FILLER_295_2243 ();
 b15zdnd11an1n08x5 FILLER_295_2275 ();
 b15zdnd00an1n01x5 FILLER_295_2283 ();
 b15zdnd11an1n64x5 FILLER_296_8 ();
 b15zdnd00an1n02x5 FILLER_296_72 ();
 b15zdnd00an1n01x5 FILLER_296_74 ();
 b15zdnd11an1n64x5 FILLER_296_78 ();
 b15zdnd11an1n32x5 FILLER_296_142 ();
 b15zdnd11an1n16x5 FILLER_296_174 ();
 b15zdnd00an1n02x5 FILLER_296_190 ();
 b15zdnd11an1n64x5 FILLER_296_195 ();
 b15zdnd11an1n08x5 FILLER_296_259 ();
 b15zdnd11an1n04x5 FILLER_296_267 ();
 b15zdnd00an1n01x5 FILLER_296_271 ();
 b15zdnd11an1n04x5 FILLER_296_312 ();
 b15zdnd11an1n64x5 FILLER_296_319 ();
 b15zdnd11an1n16x5 FILLER_296_383 ();
 b15zdnd11an1n08x5 FILLER_296_399 ();
 b15zdnd00an1n02x5 FILLER_296_407 ();
 b15zdnd00an1n01x5 FILLER_296_409 ();
 b15zdnd11an1n64x5 FILLER_296_462 ();
 b15zdnd11an1n64x5 FILLER_296_526 ();
 b15zdnd11an1n64x5 FILLER_296_590 ();
 b15zdnd11an1n64x5 FILLER_296_654 ();
 b15zdnd11an1n64x5 FILLER_296_726 ();
 b15zdnd11an1n32x5 FILLER_296_790 ();
 b15zdnd11an1n16x5 FILLER_296_822 ();
 b15zdnd11an1n08x5 FILLER_296_838 ();
 b15zdnd11an1n04x5 FILLER_296_846 ();
 b15zdnd00an1n02x5 FILLER_296_850 ();
 b15zdnd11an1n04x5 FILLER_296_855 ();
 b15zdnd11an1n64x5 FILLER_296_862 ();
 b15zdnd11an1n64x5 FILLER_296_926 ();
 b15zdnd11an1n64x5 FILLER_296_990 ();
 b15zdnd11an1n32x5 FILLER_296_1054 ();
 b15zdnd11an1n16x5 FILLER_296_1086 ();
 b15zdnd11an1n08x5 FILLER_296_1102 ();
 b15zdnd00an1n02x5 FILLER_296_1110 ();
 b15zdnd00an1n01x5 FILLER_296_1112 ();
 b15zdnd11an1n08x5 FILLER_296_1116 ();
 b15zdnd11an1n04x5 FILLER_296_1124 ();
 b15zdnd00an1n01x5 FILLER_296_1128 ();
 b15zdnd11an1n64x5 FILLER_296_1140 ();
 b15zdnd11an1n64x5 FILLER_296_1204 ();
 b15zdnd11an1n64x5 FILLER_296_1268 ();
 b15zdnd11an1n64x5 FILLER_296_1332 ();
 b15zdnd11an1n64x5 FILLER_296_1396 ();
 b15zdnd11an1n64x5 FILLER_296_1460 ();
 b15zdnd11an1n64x5 FILLER_296_1524 ();
 b15zdnd11an1n64x5 FILLER_296_1588 ();
 b15zdnd11an1n64x5 FILLER_296_1652 ();
 b15zdnd11an1n32x5 FILLER_296_1716 ();
 b15zdnd11an1n08x5 FILLER_296_1748 ();
 b15zdnd11an1n04x5 FILLER_296_1756 ();
 b15zdnd00an1n01x5 FILLER_296_1760 ();
 b15zdnd11an1n04x5 FILLER_296_1764 ();
 b15zdnd11an1n64x5 FILLER_296_1771 ();
 b15zdnd11an1n64x5 FILLER_296_1835 ();
 b15zdnd11an1n64x5 FILLER_296_1899 ();
 b15zdnd11an1n64x5 FILLER_296_1963 ();
 b15zdnd11an1n64x5 FILLER_296_2027 ();
 b15zdnd11an1n32x5 FILLER_296_2091 ();
 b15zdnd11an1n16x5 FILLER_296_2123 ();
 b15zdnd11an1n08x5 FILLER_296_2139 ();
 b15zdnd11an1n04x5 FILLER_296_2147 ();
 b15zdnd00an1n02x5 FILLER_296_2151 ();
 b15zdnd00an1n01x5 FILLER_296_2153 ();
 b15zdnd11an1n64x5 FILLER_296_2162 ();
 b15zdnd11an1n32x5 FILLER_296_2226 ();
 b15zdnd11an1n16x5 FILLER_296_2258 ();
 b15zdnd00an1n02x5 FILLER_296_2274 ();
 b15zdnd11an1n64x5 FILLER_297_0 ();
 b15zdnd11an1n64x5 FILLER_297_82 ();
 b15zdnd11an1n16x5 FILLER_297_146 ();
 b15zdnd11an1n04x5 FILLER_297_162 ();
 b15zdnd00an1n01x5 FILLER_297_166 ();
 b15zdnd11an1n32x5 FILLER_297_219 ();
 b15zdnd11an1n16x5 FILLER_297_251 ();
 b15zdnd11an1n04x5 FILLER_297_267 ();
 b15zdnd11an1n64x5 FILLER_297_275 ();
 b15zdnd11an1n64x5 FILLER_297_339 ();
 b15zdnd11an1n08x5 FILLER_297_403 ();
 b15zdnd11an1n04x5 FILLER_297_411 ();
 b15zdnd11an1n08x5 FILLER_297_418 ();
 b15zdnd11an1n08x5 FILLER_297_429 ();
 b15zdnd00an1n01x5 FILLER_297_437 ();
 b15zdnd11an1n04x5 FILLER_297_465 ();
 b15zdnd11an1n64x5 FILLER_297_478 ();
 b15zdnd11an1n16x5 FILLER_297_542 ();
 b15zdnd11an1n16x5 FILLER_297_574 ();
 b15zdnd11an1n04x5 FILLER_297_590 ();
 b15zdnd00an1n01x5 FILLER_297_594 ();
 b15zdnd11an1n64x5 FILLER_297_601 ();
 b15zdnd11an1n64x5 FILLER_297_665 ();
 b15zdnd11an1n64x5 FILLER_297_729 ();
 b15zdnd11an1n64x5 FILLER_297_793 ();
 b15zdnd11an1n64x5 FILLER_297_857 ();
 b15zdnd11an1n32x5 FILLER_297_921 ();
 b15zdnd11an1n04x5 FILLER_297_953 ();
 b15zdnd00an1n02x5 FILLER_297_957 ();
 b15zdnd00an1n01x5 FILLER_297_959 ();
 b15zdnd11an1n64x5 FILLER_297_969 ();
 b15zdnd11an1n32x5 FILLER_297_1033 ();
 b15zdnd11an1n16x5 FILLER_297_1065 ();
 b15zdnd11an1n04x5 FILLER_297_1081 ();
 b15zdnd00an1n02x5 FILLER_297_1085 ();
 b15zdnd11an1n64x5 FILLER_297_1118 ();
 b15zdnd11an1n64x5 FILLER_297_1182 ();
 b15zdnd11an1n64x5 FILLER_297_1246 ();
 b15zdnd11an1n64x5 FILLER_297_1310 ();
 b15zdnd11an1n64x5 FILLER_297_1374 ();
 b15zdnd11an1n08x5 FILLER_297_1438 ();
 b15zdnd00an1n02x5 FILLER_297_1446 ();
 b15zdnd11an1n64x5 FILLER_297_1480 ();
 b15zdnd11an1n64x5 FILLER_297_1544 ();
 b15zdnd11an1n64x5 FILLER_297_1608 ();
 b15zdnd11an1n64x5 FILLER_297_1672 ();
 b15zdnd11an1n64x5 FILLER_297_1736 ();
 b15zdnd11an1n64x5 FILLER_297_1800 ();
 b15zdnd11an1n64x5 FILLER_297_1864 ();
 b15zdnd11an1n64x5 FILLER_297_1928 ();
 b15zdnd11an1n64x5 FILLER_297_1992 ();
 b15zdnd11an1n64x5 FILLER_297_2056 ();
 b15zdnd11an1n64x5 FILLER_297_2120 ();
 b15zdnd11an1n64x5 FILLER_297_2184 ();
 b15zdnd11an1n32x5 FILLER_297_2248 ();
 b15zdnd11an1n04x5 FILLER_297_2280 ();
 b15zdnd11an1n64x5 FILLER_298_8 ();
 b15zdnd11an1n16x5 FILLER_298_72 ();
 b15zdnd00an1n01x5 FILLER_298_88 ();
 b15zdnd11an1n64x5 FILLER_298_92 ();
 b15zdnd11an1n16x5 FILLER_298_156 ();
 b15zdnd11an1n08x5 FILLER_298_172 ();
 b15zdnd11an1n04x5 FILLER_298_180 ();
 b15zdnd00an1n02x5 FILLER_298_184 ();
 b15zdnd11an1n04x5 FILLER_298_189 ();
 b15zdnd00an1n02x5 FILLER_298_193 ();
 b15zdnd11an1n64x5 FILLER_298_198 ();
 b15zdnd11an1n64x5 FILLER_298_262 ();
 b15zdnd11an1n32x5 FILLER_298_326 ();
 b15zdnd11an1n16x5 FILLER_298_358 ();
 b15zdnd11an1n08x5 FILLER_298_374 ();
 b15zdnd11an1n04x5 FILLER_298_382 ();
 b15zdnd11an1n04x5 FILLER_298_428 ();
 b15zdnd00an1n01x5 FILLER_298_432 ();
 b15zdnd11an1n04x5 FILLER_298_436 ();
 b15zdnd11an1n04x5 FILLER_298_443 ();
 b15zdnd00an1n02x5 FILLER_298_447 ();
 b15zdnd11an1n04x5 FILLER_298_452 ();
 b15zdnd11an1n64x5 FILLER_298_465 ();
 b15zdnd11an1n32x5 FILLER_298_529 ();
 b15zdnd11an1n08x5 FILLER_298_561 ();
 b15zdnd11an1n64x5 FILLER_298_585 ();
 b15zdnd11an1n64x5 FILLER_298_649 ();
 b15zdnd11an1n04x5 FILLER_298_713 ();
 b15zdnd00an1n01x5 FILLER_298_717 ();
 b15zdnd11an1n64x5 FILLER_298_726 ();
 b15zdnd11an1n64x5 FILLER_298_790 ();
 b15zdnd11an1n64x5 FILLER_298_854 ();
 b15zdnd11an1n64x5 FILLER_298_918 ();
 b15zdnd11an1n64x5 FILLER_298_982 ();
 b15zdnd11an1n64x5 FILLER_298_1046 ();
 b15zdnd11an1n64x5 FILLER_298_1110 ();
 b15zdnd11an1n64x5 FILLER_298_1174 ();
 b15zdnd11an1n64x5 FILLER_298_1238 ();
 b15zdnd11an1n64x5 FILLER_298_1302 ();
 b15zdnd11an1n64x5 FILLER_298_1366 ();
 b15zdnd11an1n64x5 FILLER_298_1430 ();
 b15zdnd11an1n16x5 FILLER_298_1494 ();
 b15zdnd11an1n08x5 FILLER_298_1510 ();
 b15zdnd11an1n04x5 FILLER_298_1518 ();
 b15zdnd00an1n01x5 FILLER_298_1522 ();
 b15zdnd11an1n04x5 FILLER_298_1526 ();
 b15zdnd11an1n64x5 FILLER_298_1533 ();
 b15zdnd11an1n64x5 FILLER_298_1597 ();
 b15zdnd11an1n64x5 FILLER_298_1661 ();
 b15zdnd11an1n64x5 FILLER_298_1725 ();
 b15zdnd11an1n64x5 FILLER_298_1789 ();
 b15zdnd11an1n64x5 FILLER_298_1853 ();
 b15zdnd11an1n64x5 FILLER_298_1917 ();
 b15zdnd11an1n64x5 FILLER_298_1981 ();
 b15zdnd11an1n64x5 FILLER_298_2045 ();
 b15zdnd11an1n32x5 FILLER_298_2109 ();
 b15zdnd11an1n08x5 FILLER_298_2141 ();
 b15zdnd11an1n04x5 FILLER_298_2149 ();
 b15zdnd00an1n01x5 FILLER_298_2153 ();
 b15zdnd11an1n64x5 FILLER_298_2162 ();
 b15zdnd11an1n32x5 FILLER_298_2226 ();
 b15zdnd11an1n16x5 FILLER_298_2258 ();
 b15zdnd00an1n02x5 FILLER_298_2274 ();
 b15zdnd11an1n32x5 FILLER_299_0 ();
 b15zdnd11an1n16x5 FILLER_299_32 ();
 b15zdnd11an1n08x5 FILLER_299_48 ();
 b15zdnd00an1n01x5 FILLER_299_56 ();
 b15zdnd11an1n64x5 FILLER_299_67 ();
 b15zdnd11an1n32x5 FILLER_299_131 ();
 b15zdnd11an1n16x5 FILLER_299_163 ();
 b15zdnd11an1n08x5 FILLER_299_179 ();
 b15zdnd00an1n02x5 FILLER_299_187 ();
 b15zdnd00an1n01x5 FILLER_299_189 ();
 b15zdnd11an1n16x5 FILLER_299_193 ();
 b15zdnd11an1n08x5 FILLER_299_209 ();
 b15zdnd00an1n02x5 FILLER_299_217 ();
 b15zdnd11an1n64x5 FILLER_299_239 ();
 b15zdnd11an1n64x5 FILLER_299_303 ();
 b15zdnd11an1n32x5 FILLER_299_367 ();
 b15zdnd11an1n16x5 FILLER_299_399 ();
 b15zdnd11an1n08x5 FILLER_299_415 ();
 b15zdnd11an1n04x5 FILLER_299_426 ();
 b15zdnd11an1n64x5 FILLER_299_482 ();
 b15zdnd11an1n32x5 FILLER_299_546 ();
 b15zdnd11an1n16x5 FILLER_299_578 ();
 b15zdnd11an1n08x5 FILLER_299_594 ();
 b15zdnd11an1n04x5 FILLER_299_618 ();
 b15zdnd00an1n01x5 FILLER_299_622 ();
 b15zdnd11an1n08x5 FILLER_299_626 ();
 b15zdnd00an1n02x5 FILLER_299_634 ();
 b15zdnd11an1n64x5 FILLER_299_678 ();
 b15zdnd11an1n64x5 FILLER_299_742 ();
 b15zdnd11an1n64x5 FILLER_299_806 ();
 b15zdnd11an1n64x5 FILLER_299_870 ();
 b15zdnd11an1n64x5 FILLER_299_934 ();
 b15zdnd11an1n64x5 FILLER_299_998 ();
 b15zdnd11an1n64x5 FILLER_299_1062 ();
 b15zdnd11an1n64x5 FILLER_299_1126 ();
 b15zdnd11an1n64x5 FILLER_299_1190 ();
 b15zdnd11an1n64x5 FILLER_299_1254 ();
 b15zdnd11an1n64x5 FILLER_299_1318 ();
 b15zdnd11an1n64x5 FILLER_299_1382 ();
 b15zdnd11an1n32x5 FILLER_299_1446 ();
 b15zdnd11an1n16x5 FILLER_299_1478 ();
 b15zdnd11an1n04x5 FILLER_299_1494 ();
 b15zdnd11an1n64x5 FILLER_299_1550 ();
 b15zdnd11an1n32x5 FILLER_299_1614 ();
 b15zdnd00an1n02x5 FILLER_299_1646 ();
 b15zdnd11an1n64x5 FILLER_299_1651 ();
 b15zdnd11an1n64x5 FILLER_299_1715 ();
 b15zdnd11an1n64x5 FILLER_299_1779 ();
 b15zdnd11an1n64x5 FILLER_299_1843 ();
 b15zdnd11an1n04x5 FILLER_299_1910 ();
 b15zdnd11an1n64x5 FILLER_299_1917 ();
 b15zdnd11an1n64x5 FILLER_299_1981 ();
 b15zdnd11an1n64x5 FILLER_299_2045 ();
 b15zdnd11an1n64x5 FILLER_299_2109 ();
 b15zdnd11an1n64x5 FILLER_299_2173 ();
 b15zdnd11an1n32x5 FILLER_299_2237 ();
 b15zdnd11an1n08x5 FILLER_299_2269 ();
 b15zdnd11an1n04x5 FILLER_299_2277 ();
 b15zdnd00an1n02x5 FILLER_299_2281 ();
 b15zdnd00an1n01x5 FILLER_299_2283 ();
 b15zdnd11an1n64x5 FILLER_300_8 ();
 b15zdnd11an1n16x5 FILLER_300_72 ();
 b15zdnd00an1n01x5 FILLER_300_88 ();
 b15zdnd11an1n64x5 FILLER_300_95 ();
 b15zdnd11an1n64x5 FILLER_300_159 ();
 b15zdnd11an1n64x5 FILLER_300_223 ();
 b15zdnd11an1n64x5 FILLER_300_287 ();
 b15zdnd11an1n64x5 FILLER_300_351 ();
 b15zdnd11an1n32x5 FILLER_300_415 ();
 b15zdnd00an1n01x5 FILLER_300_447 ();
 b15zdnd11an1n04x5 FILLER_300_451 ();
 b15zdnd11an1n64x5 FILLER_300_458 ();
 b15zdnd11an1n64x5 FILLER_300_522 ();
 b15zdnd11an1n08x5 FILLER_300_586 ();
 b15zdnd00an1n02x5 FILLER_300_594 ();
 b15zdnd11an1n64x5 FILLER_300_648 ();
 b15zdnd11an1n04x5 FILLER_300_712 ();
 b15zdnd00an1n02x5 FILLER_300_716 ();
 b15zdnd11an1n64x5 FILLER_300_726 ();
 b15zdnd11an1n64x5 FILLER_300_790 ();
 b15zdnd11an1n64x5 FILLER_300_854 ();
 b15zdnd11an1n64x5 FILLER_300_918 ();
 b15zdnd11an1n64x5 FILLER_300_982 ();
 b15zdnd11an1n64x5 FILLER_300_1046 ();
 b15zdnd11an1n64x5 FILLER_300_1110 ();
 b15zdnd11an1n64x5 FILLER_300_1174 ();
 b15zdnd11an1n64x5 FILLER_300_1238 ();
 b15zdnd11an1n64x5 FILLER_300_1302 ();
 b15zdnd11an1n64x5 FILLER_300_1366 ();
 b15zdnd11an1n64x5 FILLER_300_1430 ();
 b15zdnd11an1n16x5 FILLER_300_1494 ();
 b15zdnd11an1n08x5 FILLER_300_1510 ();
 b15zdnd11an1n04x5 FILLER_300_1518 ();
 b15zdnd00an1n02x5 FILLER_300_1522 ();
 b15zdnd11an1n16x5 FILLER_300_1527 ();
 b15zdnd00an1n02x5 FILLER_300_1543 ();
 b15zdnd00an1n01x5 FILLER_300_1545 ();
 b15zdnd11an1n32x5 FILLER_300_1598 ();
 b15zdnd11an1n16x5 FILLER_300_1630 ();
 b15zdnd11an1n04x5 FILLER_300_1649 ();
 b15zdnd11an1n64x5 FILLER_300_1656 ();
 b15zdnd11an1n64x5 FILLER_300_1720 ();
 b15zdnd11an1n64x5 FILLER_300_1784 ();
 b15zdnd11an1n32x5 FILLER_300_1848 ();
 b15zdnd11an1n08x5 FILLER_300_1880 ();
 b15zdnd00an1n01x5 FILLER_300_1888 ();
 b15zdnd11an1n64x5 FILLER_300_1941 ();
 b15zdnd11an1n32x5 FILLER_300_2005 ();
 b15zdnd11an1n16x5 FILLER_300_2037 ();
 b15zdnd11an1n04x5 FILLER_300_2053 ();
 b15zdnd00an1n02x5 FILLER_300_2057 ();
 b15zdnd11an1n64x5 FILLER_300_2077 ();
 b15zdnd11an1n08x5 FILLER_300_2141 ();
 b15zdnd11an1n04x5 FILLER_300_2149 ();
 b15zdnd00an1n01x5 FILLER_300_2153 ();
 b15zdnd11an1n64x5 FILLER_300_2162 ();
 b15zdnd11an1n32x5 FILLER_300_2226 ();
 b15zdnd11an1n16x5 FILLER_300_2258 ();
 b15zdnd00an1n02x5 FILLER_300_2274 ();
 b15zdnd11an1n64x5 FILLER_301_0 ();
 b15zdnd11an1n64x5 FILLER_301_64 ();
 b15zdnd11an1n64x5 FILLER_301_128 ();
 b15zdnd11an1n64x5 FILLER_301_192 ();
 b15zdnd11an1n08x5 FILLER_301_256 ();
 b15zdnd11an1n04x5 FILLER_301_264 ();
 b15zdnd00an1n02x5 FILLER_301_268 ();
 b15zdnd11an1n64x5 FILLER_301_293 ();
 b15zdnd11an1n64x5 FILLER_301_357 ();
 b15zdnd11an1n32x5 FILLER_301_421 ();
 b15zdnd11an1n04x5 FILLER_301_453 ();
 b15zdnd00an1n02x5 FILLER_301_457 ();
 b15zdnd00an1n01x5 FILLER_301_459 ();
 b15zdnd11an1n04x5 FILLER_301_463 ();
 b15zdnd11an1n64x5 FILLER_301_470 ();
 b15zdnd11an1n64x5 FILLER_301_534 ();
 b15zdnd11an1n08x5 FILLER_301_598 ();
 b15zdnd00an1n01x5 FILLER_301_606 ();
 b15zdnd11an1n64x5 FILLER_301_649 ();
 b15zdnd11an1n64x5 FILLER_301_713 ();
 b15zdnd11an1n64x5 FILLER_301_777 ();
 b15zdnd11an1n64x5 FILLER_301_841 ();
 b15zdnd11an1n64x5 FILLER_301_905 ();
 b15zdnd11an1n64x5 FILLER_301_969 ();
 b15zdnd11an1n64x5 FILLER_301_1033 ();
 b15zdnd11an1n64x5 FILLER_301_1097 ();
 b15zdnd11an1n64x5 FILLER_301_1161 ();
 b15zdnd11an1n64x5 FILLER_301_1225 ();
 b15zdnd11an1n64x5 FILLER_301_1289 ();
 b15zdnd11an1n08x5 FILLER_301_1353 ();
 b15zdnd00an1n02x5 FILLER_301_1361 ();
 b15zdnd00an1n01x5 FILLER_301_1363 ();
 b15zdnd11an1n04x5 FILLER_301_1367 ();
 b15zdnd11an1n64x5 FILLER_301_1374 ();
 b15zdnd11an1n64x5 FILLER_301_1438 ();
 b15zdnd11an1n32x5 FILLER_301_1502 ();
 b15zdnd11an1n16x5 FILLER_301_1534 ();
 b15zdnd11an1n08x5 FILLER_301_1550 ();
 b15zdnd11an1n04x5 FILLER_301_1558 ();
 b15zdnd00an1n02x5 FILLER_301_1562 ();
 b15zdnd11an1n04x5 FILLER_301_1567 ();
 b15zdnd11an1n04x5 FILLER_301_1574 ();
 b15zdnd11an1n32x5 FILLER_301_1581 ();
 b15zdnd11an1n08x5 FILLER_301_1613 ();
 b15zdnd00an1n02x5 FILLER_301_1621 ();
 b15zdnd00an1n01x5 FILLER_301_1623 ();
 b15zdnd11an1n64x5 FILLER_301_1676 ();
 b15zdnd11an1n32x5 FILLER_301_1740 ();
 b15zdnd00an1n02x5 FILLER_301_1772 ();
 b15zdnd11an1n04x5 FILLER_301_1777 ();
 b15zdnd11an1n64x5 FILLER_301_1784 ();
 b15zdnd11an1n64x5 FILLER_301_1848 ();
 b15zdnd00an1n02x5 FILLER_301_1912 ();
 b15zdnd11an1n64x5 FILLER_301_1917 ();
 b15zdnd11an1n64x5 FILLER_301_1981 ();
 b15zdnd11an1n64x5 FILLER_301_2045 ();
 b15zdnd11an1n64x5 FILLER_301_2109 ();
 b15zdnd11an1n64x5 FILLER_301_2173 ();
 b15zdnd11an1n32x5 FILLER_301_2237 ();
 b15zdnd11an1n08x5 FILLER_301_2269 ();
 b15zdnd11an1n04x5 FILLER_301_2277 ();
 b15zdnd00an1n02x5 FILLER_301_2281 ();
 b15zdnd00an1n01x5 FILLER_301_2283 ();
 b15zdnd11an1n64x5 FILLER_302_8 ();
 b15zdnd11an1n08x5 FILLER_302_72 ();
 b15zdnd00an1n02x5 FILLER_302_80 ();
 b15zdnd00an1n01x5 FILLER_302_82 ();
 b15zdnd11an1n64x5 FILLER_302_89 ();
 b15zdnd11an1n64x5 FILLER_302_153 ();
 b15zdnd11an1n64x5 FILLER_302_217 ();
 b15zdnd11an1n64x5 FILLER_302_281 ();
 b15zdnd11an1n64x5 FILLER_302_345 ();
 b15zdnd11an1n16x5 FILLER_302_409 ();
 b15zdnd11an1n08x5 FILLER_302_425 ();
 b15zdnd11an1n04x5 FILLER_302_433 ();
 b15zdnd00an1n02x5 FILLER_302_437 ();
 b15zdnd00an1n01x5 FILLER_302_439 ();
 b15zdnd11an1n64x5 FILLER_302_492 ();
 b15zdnd11an1n32x5 FILLER_302_556 ();
 b15zdnd11an1n16x5 FILLER_302_588 ();
 b15zdnd11an1n08x5 FILLER_302_604 ();
 b15zdnd11an1n04x5 FILLER_302_612 ();
 b15zdnd11an1n04x5 FILLER_302_619 ();
 b15zdnd11an1n64x5 FILLER_302_626 ();
 b15zdnd11an1n16x5 FILLER_302_690 ();
 b15zdnd11an1n08x5 FILLER_302_706 ();
 b15zdnd11an1n04x5 FILLER_302_714 ();
 b15zdnd11an1n64x5 FILLER_302_726 ();
 b15zdnd11an1n64x5 FILLER_302_790 ();
 b15zdnd11an1n64x5 FILLER_302_854 ();
 b15zdnd11an1n64x5 FILLER_302_918 ();
 b15zdnd11an1n64x5 FILLER_302_982 ();
 b15zdnd11an1n64x5 FILLER_302_1046 ();
 b15zdnd11an1n16x5 FILLER_302_1110 ();
 b15zdnd11an1n08x5 FILLER_302_1126 ();
 b15zdnd11an1n04x5 FILLER_302_1134 ();
 b15zdnd11an1n64x5 FILLER_302_1158 ();
 b15zdnd11an1n64x5 FILLER_302_1222 ();
 b15zdnd11an1n32x5 FILLER_302_1286 ();
 b15zdnd11an1n16x5 FILLER_302_1318 ();
 b15zdnd11an1n08x5 FILLER_302_1334 ();
 b15zdnd11an1n04x5 FILLER_302_1342 ();
 b15zdnd11an1n64x5 FILLER_302_1398 ();
 b15zdnd11an1n64x5 FILLER_302_1462 ();
 b15zdnd11an1n64x5 FILLER_302_1526 ();
 b15zdnd11an1n32x5 FILLER_302_1590 ();
 b15zdnd11an1n04x5 FILLER_302_1622 ();
 b15zdnd00an1n02x5 FILLER_302_1626 ();
 b15zdnd11an1n64x5 FILLER_302_1680 ();
 b15zdnd11an1n08x5 FILLER_302_1744 ();
 b15zdnd11an1n04x5 FILLER_302_1752 ();
 b15zdnd11an1n32x5 FILLER_302_1808 ();
 b15zdnd11an1n16x5 FILLER_302_1840 ();
 b15zdnd11an1n04x5 FILLER_302_1859 ();
 b15zdnd11an1n32x5 FILLER_302_1866 ();
 b15zdnd11an1n08x5 FILLER_302_1898 ();
 b15zdnd11an1n04x5 FILLER_302_1906 ();
 b15zdnd00an1n02x5 FILLER_302_1910 ();
 b15zdnd11an1n04x5 FILLER_302_1915 ();
 b15zdnd11an1n64x5 FILLER_302_1922 ();
 b15zdnd11an1n64x5 FILLER_302_1986 ();
 b15zdnd11an1n64x5 FILLER_302_2050 ();
 b15zdnd11an1n32x5 FILLER_302_2114 ();
 b15zdnd11an1n08x5 FILLER_302_2146 ();
 b15zdnd11an1n64x5 FILLER_302_2162 ();
 b15zdnd11an1n32x5 FILLER_302_2226 ();
 b15zdnd11an1n16x5 FILLER_302_2258 ();
 b15zdnd00an1n02x5 FILLER_302_2274 ();
 b15zdnd11an1n64x5 FILLER_303_0 ();
 b15zdnd11an1n08x5 FILLER_303_64 ();
 b15zdnd00an1n01x5 FILLER_303_72 ();
 b15zdnd11an1n64x5 FILLER_303_77 ();
 b15zdnd11an1n64x5 FILLER_303_141 ();
 b15zdnd11an1n64x5 FILLER_303_205 ();
 b15zdnd11an1n64x5 FILLER_303_269 ();
 b15zdnd11an1n64x5 FILLER_303_333 ();
 b15zdnd11an1n64x5 FILLER_303_397 ();
 b15zdnd11an1n04x5 FILLER_303_461 ();
 b15zdnd00an1n01x5 FILLER_303_465 ();
 b15zdnd11an1n16x5 FILLER_303_469 ();
 b15zdnd11an1n04x5 FILLER_303_485 ();
 b15zdnd00an1n01x5 FILLER_303_489 ();
 b15zdnd11an1n64x5 FILLER_303_510 ();
 b15zdnd11an1n64x5 FILLER_303_574 ();
 b15zdnd11an1n64x5 FILLER_303_638 ();
 b15zdnd11an1n64x5 FILLER_303_702 ();
 b15zdnd11an1n64x5 FILLER_303_766 ();
 b15zdnd11an1n64x5 FILLER_303_830 ();
 b15zdnd11an1n64x5 FILLER_303_894 ();
 b15zdnd11an1n08x5 FILLER_303_958 ();
 b15zdnd11an1n16x5 FILLER_303_975 ();
 b15zdnd11an1n08x5 FILLER_303_991 ();
 b15zdnd00an1n02x5 FILLER_303_999 ();
 b15zdnd11an1n04x5 FILLER_303_1004 ();
 b15zdnd11an1n64x5 FILLER_303_1011 ();
 b15zdnd11an1n64x5 FILLER_303_1075 ();
 b15zdnd11an1n08x5 FILLER_303_1139 ();
 b15zdnd11an1n04x5 FILLER_303_1147 ();
 b15zdnd00an1n02x5 FILLER_303_1151 ();
 b15zdnd00an1n01x5 FILLER_303_1153 ();
 b15zdnd11an1n64x5 FILLER_303_1174 ();
 b15zdnd11an1n32x5 FILLER_303_1238 ();
 b15zdnd11an1n16x5 FILLER_303_1270 ();
 b15zdnd11an1n08x5 FILLER_303_1286 ();
 b15zdnd11an1n04x5 FILLER_303_1294 ();
 b15zdnd11an1n04x5 FILLER_303_1301 ();
 b15zdnd11an1n32x5 FILLER_303_1308 ();
 b15zdnd11an1n16x5 FILLER_303_1340 ();
 b15zdnd11an1n08x5 FILLER_303_1356 ();
 b15zdnd11an1n04x5 FILLER_303_1364 ();
 b15zdnd00an1n02x5 FILLER_303_1368 ();
 b15zdnd00an1n01x5 FILLER_303_1370 ();
 b15zdnd11an1n64x5 FILLER_303_1374 ();
 b15zdnd11an1n64x5 FILLER_303_1438 ();
 b15zdnd11an1n64x5 FILLER_303_1502 ();
 b15zdnd11an1n32x5 FILLER_303_1566 ();
 b15zdnd11an1n16x5 FILLER_303_1598 ();
 b15zdnd11an1n04x5 FILLER_303_1614 ();
 b15zdnd00an1n02x5 FILLER_303_1618 ();
 b15zdnd00an1n01x5 FILLER_303_1620 ();
 b15zdnd11an1n04x5 FILLER_303_1641 ();
 b15zdnd11an1n08x5 FILLER_303_1648 ();
 b15zdnd11an1n64x5 FILLER_303_1659 ();
 b15zdnd11an1n32x5 FILLER_303_1723 ();
 b15zdnd11an1n16x5 FILLER_303_1755 ();
 b15zdnd11an1n08x5 FILLER_303_1771 ();
 b15zdnd00an1n02x5 FILLER_303_1779 ();
 b15zdnd00an1n01x5 FILLER_303_1781 ();
 b15zdnd11an1n32x5 FILLER_303_1785 ();
 b15zdnd11an1n16x5 FILLER_303_1817 ();
 b15zdnd11an1n04x5 FILLER_303_1833 ();
 b15zdnd00an1n01x5 FILLER_303_1837 ();
 b15zdnd11an1n04x5 FILLER_303_1890 ();
 b15zdnd11an1n64x5 FILLER_303_1946 ();
 b15zdnd11an1n64x5 FILLER_303_2010 ();
 b15zdnd11an1n64x5 FILLER_303_2074 ();
 b15zdnd11an1n64x5 FILLER_303_2138 ();
 b15zdnd11an1n64x5 FILLER_303_2202 ();
 b15zdnd11an1n16x5 FILLER_303_2266 ();
 b15zdnd00an1n02x5 FILLER_303_2282 ();
 b15zdnd11an1n64x5 FILLER_304_8 ();
 b15zdnd11an1n64x5 FILLER_304_72 ();
 b15zdnd11an1n64x5 FILLER_304_136 ();
 b15zdnd11an1n64x5 FILLER_304_200 ();
 b15zdnd11an1n64x5 FILLER_304_264 ();
 b15zdnd11an1n64x5 FILLER_304_328 ();
 b15zdnd11an1n32x5 FILLER_304_392 ();
 b15zdnd11an1n16x5 FILLER_304_424 ();
 b15zdnd11an1n08x5 FILLER_304_440 ();
 b15zdnd00an1n02x5 FILLER_304_448 ();
 b15zdnd11an1n64x5 FILLER_304_457 ();
 b15zdnd11an1n64x5 FILLER_304_521 ();
 b15zdnd11an1n64x5 FILLER_304_585 ();
 b15zdnd11an1n64x5 FILLER_304_649 ();
 b15zdnd11an1n04x5 FILLER_304_713 ();
 b15zdnd00an1n01x5 FILLER_304_717 ();
 b15zdnd00an1n02x5 FILLER_304_726 ();
 b15zdnd11an1n64x5 FILLER_304_760 ();
 b15zdnd11an1n64x5 FILLER_304_824 ();
 b15zdnd11an1n64x5 FILLER_304_888 ();
 b15zdnd11an1n16x5 FILLER_304_952 ();
 b15zdnd11an1n08x5 FILLER_304_968 ();
 b15zdnd11an1n04x5 FILLER_304_976 ();
 b15zdnd00an1n01x5 FILLER_304_980 ();
 b15zdnd11an1n04x5 FILLER_304_1033 ();
 b15zdnd00an1n02x5 FILLER_304_1037 ();
 b15zdnd11an1n64x5 FILLER_304_1053 ();
 b15zdnd11an1n64x5 FILLER_304_1117 ();
 b15zdnd11an1n64x5 FILLER_304_1181 ();
 b15zdnd11an1n04x5 FILLER_304_1245 ();
 b15zdnd11an1n04x5 FILLER_304_1276 ();
 b15zdnd11an1n32x5 FILLER_304_1332 ();
 b15zdnd11an1n04x5 FILLER_304_1364 ();
 b15zdnd00an1n02x5 FILLER_304_1368 ();
 b15zdnd11an1n04x5 FILLER_304_1373 ();
 b15zdnd11an1n64x5 FILLER_304_1380 ();
 b15zdnd11an1n64x5 FILLER_304_1444 ();
 b15zdnd11an1n64x5 FILLER_304_1508 ();
 b15zdnd11an1n64x5 FILLER_304_1572 ();
 b15zdnd11an1n16x5 FILLER_304_1636 ();
 b15zdnd11an1n04x5 FILLER_304_1652 ();
 b15zdnd11an1n64x5 FILLER_304_1659 ();
 b15zdnd11an1n64x5 FILLER_304_1723 ();
 b15zdnd11an1n64x5 FILLER_304_1787 ();
 b15zdnd11an1n08x5 FILLER_304_1851 ();
 b15zdnd11an1n04x5 FILLER_304_1859 ();
 b15zdnd00an1n01x5 FILLER_304_1863 ();
 b15zdnd11an1n32x5 FILLER_304_1867 ();
 b15zdnd11an1n08x5 FILLER_304_1899 ();
 b15zdnd11an1n04x5 FILLER_304_1907 ();
 b15zdnd00an1n02x5 FILLER_304_1911 ();
 b15zdnd11an1n64x5 FILLER_304_1916 ();
 b15zdnd11an1n64x5 FILLER_304_1980 ();
 b15zdnd11an1n64x5 FILLER_304_2044 ();
 b15zdnd11an1n32x5 FILLER_304_2108 ();
 b15zdnd11an1n08x5 FILLER_304_2140 ();
 b15zdnd11an1n04x5 FILLER_304_2148 ();
 b15zdnd00an1n02x5 FILLER_304_2152 ();
 b15zdnd11an1n64x5 FILLER_304_2162 ();
 b15zdnd11an1n32x5 FILLER_304_2226 ();
 b15zdnd11an1n16x5 FILLER_304_2258 ();
 b15zdnd00an1n02x5 FILLER_304_2274 ();
 b15zdnd11an1n64x5 FILLER_305_0 ();
 b15zdnd11an1n64x5 FILLER_305_64 ();
 b15zdnd11an1n64x5 FILLER_305_128 ();
 b15zdnd11an1n64x5 FILLER_305_192 ();
 b15zdnd11an1n64x5 FILLER_305_256 ();
 b15zdnd11an1n64x5 FILLER_305_320 ();
 b15zdnd11an1n64x5 FILLER_305_384 ();
 b15zdnd11an1n64x5 FILLER_305_448 ();
 b15zdnd11an1n64x5 FILLER_305_512 ();
 b15zdnd11an1n64x5 FILLER_305_576 ();
 b15zdnd11an1n64x5 FILLER_305_640 ();
 b15zdnd11an1n08x5 FILLER_305_704 ();
 b15zdnd00an1n01x5 FILLER_305_712 ();
 b15zdnd11an1n04x5 FILLER_305_765 ();
 b15zdnd11an1n64x5 FILLER_305_772 ();
 b15zdnd11an1n64x5 FILLER_305_836 ();
 b15zdnd11an1n64x5 FILLER_305_900 ();
 b15zdnd11an1n16x5 FILLER_305_964 ();
 b15zdnd11an1n04x5 FILLER_305_1000 ();
 b15zdnd11an1n64x5 FILLER_305_1007 ();
 b15zdnd11an1n64x5 FILLER_305_1071 ();
 b15zdnd11an1n64x5 FILLER_305_1135 ();
 b15zdnd11an1n08x5 FILLER_305_1199 ();
 b15zdnd11an1n04x5 FILLER_305_1207 ();
 b15zdnd00an1n02x5 FILLER_305_1211 ();
 b15zdnd11an1n04x5 FILLER_305_1216 ();
 b15zdnd11an1n16x5 FILLER_305_1223 ();
 b15zdnd11an1n08x5 FILLER_305_1239 ();
 b15zdnd00an1n02x5 FILLER_305_1247 ();
 b15zdnd11an1n32x5 FILLER_305_1252 ();
 b15zdnd11an1n16x5 FILLER_305_1284 ();
 b15zdnd11an1n04x5 FILLER_305_1300 ();
 b15zdnd00an1n02x5 FILLER_305_1304 ();
 b15zdnd11an1n32x5 FILLER_305_1309 ();
 b15zdnd11an1n04x5 FILLER_305_1341 ();
 b15zdnd11an1n64x5 FILLER_305_1397 ();
 b15zdnd11an1n64x5 FILLER_305_1461 ();
 b15zdnd11an1n64x5 FILLER_305_1525 ();
 b15zdnd11an1n64x5 FILLER_305_1589 ();
 b15zdnd11an1n64x5 FILLER_305_1653 ();
 b15zdnd11an1n64x5 FILLER_305_1717 ();
 b15zdnd11an1n64x5 FILLER_305_1781 ();
 b15zdnd11an1n32x5 FILLER_305_1845 ();
 b15zdnd00an1n02x5 FILLER_305_1877 ();
 b15zdnd00an1n01x5 FILLER_305_1879 ();
 b15zdnd11an1n64x5 FILLER_305_1911 ();
 b15zdnd11an1n64x5 FILLER_305_1975 ();
 b15zdnd11an1n64x5 FILLER_305_2039 ();
 b15zdnd11an1n64x5 FILLER_305_2103 ();
 b15zdnd11an1n64x5 FILLER_305_2167 ();
 b15zdnd11an1n32x5 FILLER_305_2231 ();
 b15zdnd11an1n16x5 FILLER_305_2263 ();
 b15zdnd11an1n04x5 FILLER_305_2279 ();
 b15zdnd00an1n01x5 FILLER_305_2283 ();
 b15zdnd11an1n64x5 FILLER_306_8 ();
 b15zdnd11an1n64x5 FILLER_306_72 ();
 b15zdnd11an1n64x5 FILLER_306_136 ();
 b15zdnd11an1n64x5 FILLER_306_200 ();
 b15zdnd11an1n64x5 FILLER_306_264 ();
 b15zdnd11an1n64x5 FILLER_306_328 ();
 b15zdnd11an1n64x5 FILLER_306_392 ();
 b15zdnd11an1n64x5 FILLER_306_456 ();
 b15zdnd11an1n64x5 FILLER_306_520 ();
 b15zdnd11an1n64x5 FILLER_306_584 ();
 b15zdnd11an1n64x5 FILLER_306_648 ();
 b15zdnd11an1n04x5 FILLER_306_712 ();
 b15zdnd00an1n02x5 FILLER_306_716 ();
 b15zdnd11an1n04x5 FILLER_306_726 ();
 b15zdnd11an1n04x5 FILLER_306_733 ();
 b15zdnd11an1n08x5 FILLER_306_740 ();
 b15zdnd00an1n02x5 FILLER_306_748 ();
 b15zdnd00an1n01x5 FILLER_306_750 ();
 b15zdnd11an1n64x5 FILLER_306_754 ();
 b15zdnd11an1n64x5 FILLER_306_818 ();
 b15zdnd11an1n64x5 FILLER_306_882 ();
 b15zdnd11an1n16x5 FILLER_306_946 ();
 b15zdnd00an1n01x5 FILLER_306_962 ();
 b15zdnd11an1n64x5 FILLER_306_983 ();
 b15zdnd11an1n64x5 FILLER_306_1047 ();
 b15zdnd11an1n64x5 FILLER_306_1111 ();
 b15zdnd11an1n16x5 FILLER_306_1175 ();
 b15zdnd11an1n04x5 FILLER_306_1191 ();
 b15zdnd11an1n64x5 FILLER_306_1247 ();
 b15zdnd11an1n32x5 FILLER_306_1311 ();
 b15zdnd11an1n16x5 FILLER_306_1343 ();
 b15zdnd11an1n08x5 FILLER_306_1359 ();
 b15zdnd11an1n04x5 FILLER_306_1367 ();
 b15zdnd11an1n64x5 FILLER_306_1374 ();
 b15zdnd11an1n64x5 FILLER_306_1438 ();
 b15zdnd11an1n64x5 FILLER_306_1502 ();
 b15zdnd11an1n64x5 FILLER_306_1566 ();
 b15zdnd11an1n64x5 FILLER_306_1630 ();
 b15zdnd11an1n64x5 FILLER_306_1694 ();
 b15zdnd11an1n64x5 FILLER_306_1758 ();
 b15zdnd11an1n64x5 FILLER_306_1822 ();
 b15zdnd11an1n64x5 FILLER_306_1886 ();
 b15zdnd11an1n64x5 FILLER_306_1950 ();
 b15zdnd11an1n64x5 FILLER_306_2014 ();
 b15zdnd11an1n64x5 FILLER_306_2078 ();
 b15zdnd11an1n08x5 FILLER_306_2142 ();
 b15zdnd11an1n04x5 FILLER_306_2150 ();
 b15zdnd11an1n64x5 FILLER_306_2162 ();
 b15zdnd11an1n32x5 FILLER_306_2226 ();
 b15zdnd11an1n16x5 FILLER_306_2258 ();
 b15zdnd00an1n02x5 FILLER_306_2274 ();
 b15zdnd11an1n64x5 FILLER_307_0 ();
 b15zdnd11an1n04x5 FILLER_307_64 ();
 b15zdnd00an1n02x5 FILLER_307_68 ();
 b15zdnd11an1n64x5 FILLER_307_77 ();
 b15zdnd11an1n64x5 FILLER_307_141 ();
 b15zdnd11an1n64x5 FILLER_307_205 ();
 b15zdnd11an1n64x5 FILLER_307_269 ();
 b15zdnd11an1n64x5 FILLER_307_333 ();
 b15zdnd11an1n64x5 FILLER_307_397 ();
 b15zdnd11an1n64x5 FILLER_307_461 ();
 b15zdnd11an1n64x5 FILLER_307_525 ();
 b15zdnd11an1n64x5 FILLER_307_589 ();
 b15zdnd11an1n64x5 FILLER_307_653 ();
 b15zdnd11an1n08x5 FILLER_307_717 ();
 b15zdnd11an1n04x5 FILLER_307_725 ();
 b15zdnd00an1n02x5 FILLER_307_729 ();
 b15zdnd11an1n04x5 FILLER_307_734 ();
 b15zdnd11an1n04x5 FILLER_307_747 ();
 b15zdnd00an1n02x5 FILLER_307_751 ();
 b15zdnd11an1n04x5 FILLER_307_756 ();
 b15zdnd11an1n64x5 FILLER_307_763 ();
 b15zdnd11an1n64x5 FILLER_307_827 ();
 b15zdnd11an1n32x5 FILLER_307_891 ();
 b15zdnd11an1n08x5 FILLER_307_923 ();
 b15zdnd00an1n01x5 FILLER_307_931 ();
 b15zdnd11an1n64x5 FILLER_307_941 ();
 b15zdnd11an1n16x5 FILLER_307_1005 ();
 b15zdnd11an1n08x5 FILLER_307_1021 ();
 b15zdnd00an1n01x5 FILLER_307_1029 ();
 b15zdnd11an1n64x5 FILLER_307_1044 ();
 b15zdnd11an1n64x5 FILLER_307_1108 ();
 b15zdnd11an1n32x5 FILLER_307_1172 ();
 b15zdnd11an1n16x5 FILLER_307_1204 ();
 b15zdnd00an1n01x5 FILLER_307_1220 ();
 b15zdnd11an1n64x5 FILLER_307_1224 ();
 b15zdnd11an1n64x5 FILLER_307_1288 ();
 b15zdnd11an1n64x5 FILLER_307_1352 ();
 b15zdnd11an1n64x5 FILLER_307_1416 ();
 b15zdnd11an1n64x5 FILLER_307_1480 ();
 b15zdnd11an1n64x5 FILLER_307_1544 ();
 b15zdnd11an1n64x5 FILLER_307_1608 ();
 b15zdnd11an1n64x5 FILLER_307_1672 ();
 b15zdnd11an1n64x5 FILLER_307_1736 ();
 b15zdnd11an1n64x5 FILLER_307_1800 ();
 b15zdnd11an1n64x5 FILLER_307_1864 ();
 b15zdnd11an1n64x5 FILLER_307_1928 ();
 b15zdnd11an1n64x5 FILLER_307_1992 ();
 b15zdnd11an1n64x5 FILLER_307_2056 ();
 b15zdnd11an1n64x5 FILLER_307_2120 ();
 b15zdnd11an1n64x5 FILLER_307_2184 ();
 b15zdnd11an1n32x5 FILLER_307_2248 ();
 b15zdnd11an1n04x5 FILLER_307_2280 ();
 b15zdnd11an1n64x5 FILLER_308_8 ();
 b15zdnd11an1n64x5 FILLER_308_72 ();
 b15zdnd11an1n64x5 FILLER_308_136 ();
 b15zdnd11an1n64x5 FILLER_308_200 ();
 b15zdnd11an1n64x5 FILLER_308_264 ();
 b15zdnd11an1n64x5 FILLER_308_328 ();
 b15zdnd11an1n64x5 FILLER_308_392 ();
 b15zdnd11an1n64x5 FILLER_308_456 ();
 b15zdnd11an1n64x5 FILLER_308_520 ();
 b15zdnd11an1n64x5 FILLER_308_584 ();
 b15zdnd11an1n64x5 FILLER_308_648 ();
 b15zdnd11an1n04x5 FILLER_308_712 ();
 b15zdnd00an1n02x5 FILLER_308_716 ();
 b15zdnd00an1n02x5 FILLER_308_726 ();
 b15zdnd11an1n64x5 FILLER_308_756 ();
 b15zdnd11an1n64x5 FILLER_308_820 ();
 b15zdnd11an1n08x5 FILLER_308_884 ();
 b15zdnd11an1n64x5 FILLER_308_906 ();
 b15zdnd11an1n64x5 FILLER_308_970 ();
 b15zdnd11an1n64x5 FILLER_308_1034 ();
 b15zdnd11an1n64x5 FILLER_308_1098 ();
 b15zdnd11an1n64x5 FILLER_308_1162 ();
 b15zdnd11an1n64x5 FILLER_308_1226 ();
 b15zdnd11an1n64x5 FILLER_308_1290 ();
 b15zdnd11an1n64x5 FILLER_308_1354 ();
 b15zdnd11an1n64x5 FILLER_308_1418 ();
 b15zdnd11an1n64x5 FILLER_308_1482 ();
 b15zdnd11an1n64x5 FILLER_308_1546 ();
 b15zdnd11an1n64x5 FILLER_308_1610 ();
 b15zdnd11an1n64x5 FILLER_308_1674 ();
 b15zdnd11an1n64x5 FILLER_308_1738 ();
 b15zdnd11an1n64x5 FILLER_308_1802 ();
 b15zdnd11an1n64x5 FILLER_308_1866 ();
 b15zdnd11an1n64x5 FILLER_308_1930 ();
 b15zdnd11an1n64x5 FILLER_308_1994 ();
 b15zdnd11an1n64x5 FILLER_308_2058 ();
 b15zdnd11an1n32x5 FILLER_308_2122 ();
 b15zdnd11an1n64x5 FILLER_308_2162 ();
 b15zdnd11an1n32x5 FILLER_308_2226 ();
 b15zdnd11an1n16x5 FILLER_308_2258 ();
 b15zdnd00an1n02x5 FILLER_308_2274 ();
 b15zdnd11an1n64x5 FILLER_309_0 ();
 b15zdnd11an1n04x5 FILLER_309_64 ();
 b15zdnd00an1n02x5 FILLER_309_68 ();
 b15zdnd00an1n01x5 FILLER_309_70 ();
 b15zdnd11an1n64x5 FILLER_309_78 ();
 b15zdnd11an1n64x5 FILLER_309_142 ();
 b15zdnd11an1n08x5 FILLER_309_206 ();
 b15zdnd00an1n02x5 FILLER_309_214 ();
 b15zdnd11an1n64x5 FILLER_309_219 ();
 b15zdnd11an1n64x5 FILLER_309_283 ();
 b15zdnd11an1n64x5 FILLER_309_347 ();
 b15zdnd11an1n64x5 FILLER_309_411 ();
 b15zdnd11an1n64x5 FILLER_309_475 ();
 b15zdnd11an1n64x5 FILLER_309_539 ();
 b15zdnd11an1n64x5 FILLER_309_603 ();
 b15zdnd11an1n32x5 FILLER_309_667 ();
 b15zdnd11an1n16x5 FILLER_309_699 ();
 b15zdnd11an1n08x5 FILLER_309_715 ();
 b15zdnd00an1n01x5 FILLER_309_723 ();
 b15zdnd11an1n04x5 FILLER_309_727 ();
 b15zdnd11an1n64x5 FILLER_309_758 ();
 b15zdnd11an1n64x5 FILLER_309_822 ();
 b15zdnd11an1n16x5 FILLER_309_886 ();
 b15zdnd11an1n32x5 FILLER_309_916 ();
 b15zdnd11an1n08x5 FILLER_309_948 ();
 b15zdnd00an1n02x5 FILLER_309_956 ();
 b15zdnd11an1n64x5 FILLER_309_961 ();
 b15zdnd11an1n64x5 FILLER_309_1025 ();
 b15zdnd11an1n64x5 FILLER_309_1089 ();
 b15zdnd11an1n64x5 FILLER_309_1153 ();
 b15zdnd11an1n64x5 FILLER_309_1217 ();
 b15zdnd11an1n64x5 FILLER_309_1281 ();
 b15zdnd11an1n64x5 FILLER_309_1345 ();
 b15zdnd11an1n64x5 FILLER_309_1409 ();
 b15zdnd11an1n64x5 FILLER_309_1473 ();
 b15zdnd11an1n64x5 FILLER_309_1537 ();
 b15zdnd11an1n64x5 FILLER_309_1601 ();
 b15zdnd11an1n64x5 FILLER_309_1665 ();
 b15zdnd11an1n64x5 FILLER_309_1729 ();
 b15zdnd11an1n64x5 FILLER_309_1793 ();
 b15zdnd11an1n64x5 FILLER_309_1857 ();
 b15zdnd11an1n64x5 FILLER_309_1921 ();
 b15zdnd11an1n64x5 FILLER_309_1985 ();
 b15zdnd11an1n64x5 FILLER_309_2049 ();
 b15zdnd11an1n64x5 FILLER_309_2113 ();
 b15zdnd11an1n32x5 FILLER_309_2177 ();
 b15zdnd11an1n16x5 FILLER_309_2209 ();
 b15zdnd11an1n08x5 FILLER_309_2225 ();
 b15zdnd11an1n04x5 FILLER_309_2233 ();
 b15zdnd00an1n02x5 FILLER_309_2237 ();
 b15zdnd11an1n16x5 FILLER_309_2253 ();
 b15zdnd11an1n08x5 FILLER_309_2269 ();
 b15zdnd11an1n04x5 FILLER_309_2277 ();
 b15zdnd00an1n02x5 FILLER_309_2281 ();
 b15zdnd00an1n01x5 FILLER_309_2283 ();
 b15zdnd11an1n32x5 FILLER_310_8 ();
 b15zdnd11an1n16x5 FILLER_310_40 ();
 b15zdnd00an1n01x5 FILLER_310_56 ();
 b15zdnd11an1n64x5 FILLER_310_78 ();
 b15zdnd11an1n32x5 FILLER_310_142 ();
 b15zdnd11an1n08x5 FILLER_310_174 ();
 b15zdnd11an1n04x5 FILLER_310_182 ();
 b15zdnd00an1n02x5 FILLER_310_186 ();
 b15zdnd00an1n01x5 FILLER_310_188 ();
 b15zdnd11an1n64x5 FILLER_310_241 ();
 b15zdnd11an1n64x5 FILLER_310_305 ();
 b15zdnd11an1n64x5 FILLER_310_369 ();
 b15zdnd11an1n64x5 FILLER_310_433 ();
 b15zdnd11an1n64x5 FILLER_310_497 ();
 b15zdnd11an1n64x5 FILLER_310_561 ();
 b15zdnd11an1n64x5 FILLER_310_625 ();
 b15zdnd11an1n16x5 FILLER_310_689 ();
 b15zdnd11an1n08x5 FILLER_310_705 ();
 b15zdnd11an1n04x5 FILLER_310_713 ();
 b15zdnd00an1n01x5 FILLER_310_717 ();
 b15zdnd11an1n64x5 FILLER_310_726 ();
 b15zdnd11an1n64x5 FILLER_310_790 ();
 b15zdnd11an1n32x5 FILLER_310_854 ();
 b15zdnd11an1n16x5 FILLER_310_886 ();
 b15zdnd11an1n08x5 FILLER_310_902 ();
 b15zdnd11an1n04x5 FILLER_310_910 ();
 b15zdnd00an1n01x5 FILLER_310_914 ();
 b15zdnd11an1n16x5 FILLER_310_918 ();
 b15zdnd11an1n08x5 FILLER_310_934 ();
 b15zdnd11an1n04x5 FILLER_310_942 ();
 b15zdnd00an1n02x5 FILLER_310_946 ();
 b15zdnd11an1n64x5 FILLER_310_1000 ();
 b15zdnd11an1n64x5 FILLER_310_1064 ();
 b15zdnd11an1n64x5 FILLER_310_1128 ();
 b15zdnd11an1n64x5 FILLER_310_1192 ();
 b15zdnd11an1n64x5 FILLER_310_1256 ();
 b15zdnd11an1n64x5 FILLER_310_1320 ();
 b15zdnd11an1n64x5 FILLER_310_1384 ();
 b15zdnd11an1n64x5 FILLER_310_1448 ();
 b15zdnd11an1n64x5 FILLER_310_1512 ();
 b15zdnd11an1n64x5 FILLER_310_1576 ();
 b15zdnd11an1n64x5 FILLER_310_1640 ();
 b15zdnd11an1n64x5 FILLER_310_1704 ();
 b15zdnd11an1n64x5 FILLER_310_1768 ();
 b15zdnd11an1n64x5 FILLER_310_1832 ();
 b15zdnd11an1n64x5 FILLER_310_1896 ();
 b15zdnd11an1n64x5 FILLER_310_1960 ();
 b15zdnd11an1n64x5 FILLER_310_2024 ();
 b15zdnd11an1n64x5 FILLER_310_2088 ();
 b15zdnd00an1n02x5 FILLER_310_2152 ();
 b15zdnd11an1n64x5 FILLER_310_2162 ();
 b15zdnd11an1n16x5 FILLER_310_2226 ();
 b15zdnd11an1n08x5 FILLER_310_2256 ();
 b15zdnd00an1n02x5 FILLER_310_2264 ();
 b15zdnd00an1n02x5 FILLER_310_2274 ();
 b15zdnd11an1n32x5 FILLER_311_0 ();
 b15zdnd11an1n08x5 FILLER_311_32 ();
 b15zdnd00an1n02x5 FILLER_311_40 ();
 b15zdnd11an1n04x5 FILLER_311_54 ();
 b15zdnd11an1n04x5 FILLER_311_79 ();
 b15zdnd00an1n01x5 FILLER_311_83 ();
 b15zdnd11an1n64x5 FILLER_311_87 ();
 b15zdnd11an1n32x5 FILLER_311_151 ();
 b15zdnd11an1n16x5 FILLER_311_183 ();
 b15zdnd11an1n08x5 FILLER_311_199 ();
 b15zdnd11an1n04x5 FILLER_311_210 ();
 b15zdnd11an1n08x5 FILLER_311_217 ();
 b15zdnd11an1n04x5 FILLER_311_225 ();
 b15zdnd11an1n04x5 FILLER_311_236 ();
 b15zdnd11an1n64x5 FILLER_311_282 ();
 b15zdnd11an1n64x5 FILLER_311_346 ();
 b15zdnd11an1n64x5 FILLER_311_410 ();
 b15zdnd11an1n32x5 FILLER_311_474 ();
 b15zdnd11an1n16x5 FILLER_311_506 ();
 b15zdnd11an1n08x5 FILLER_311_522 ();
 b15zdnd00an1n02x5 FILLER_311_530 ();
 b15zdnd11an1n64x5 FILLER_311_549 ();
 b15zdnd11an1n64x5 FILLER_311_613 ();
 b15zdnd11an1n32x5 FILLER_311_677 ();
 b15zdnd11an1n16x5 FILLER_311_709 ();
 b15zdnd11an1n08x5 FILLER_311_725 ();
 b15zdnd11an1n04x5 FILLER_311_733 ();
 b15zdnd11an1n04x5 FILLER_311_746 ();
 b15zdnd11an1n64x5 FILLER_311_759 ();
 b15zdnd11an1n64x5 FILLER_311_823 ();
 b15zdnd00an1n02x5 FILLER_311_887 ();
 b15zdnd00an1n01x5 FILLER_311_889 ();
 b15zdnd11an1n16x5 FILLER_311_942 ();
 b15zdnd11an1n08x5 FILLER_311_958 ();
 b15zdnd00an1n02x5 FILLER_311_966 ();
 b15zdnd00an1n01x5 FILLER_311_968 ();
 b15zdnd11an1n04x5 FILLER_311_972 ();
 b15zdnd11an1n64x5 FILLER_311_979 ();
 b15zdnd11an1n64x5 FILLER_311_1043 ();
 b15zdnd11an1n64x5 FILLER_311_1107 ();
 b15zdnd11an1n64x5 FILLER_311_1171 ();
 b15zdnd11an1n32x5 FILLER_311_1235 ();
 b15zdnd11an1n16x5 FILLER_311_1267 ();
 b15zdnd11an1n08x5 FILLER_311_1283 ();
 b15zdnd00an1n02x5 FILLER_311_1291 ();
 b15zdnd00an1n01x5 FILLER_311_1293 ();
 b15zdnd11an1n64x5 FILLER_311_1303 ();
 b15zdnd11an1n64x5 FILLER_311_1367 ();
 b15zdnd11an1n64x5 FILLER_311_1431 ();
 b15zdnd11an1n64x5 FILLER_311_1495 ();
 b15zdnd11an1n64x5 FILLER_311_1559 ();
 b15zdnd11an1n64x5 FILLER_311_1623 ();
 b15zdnd11an1n64x5 FILLER_311_1687 ();
 b15zdnd11an1n64x5 FILLER_311_1751 ();
 b15zdnd11an1n64x5 FILLER_311_1815 ();
 b15zdnd11an1n64x5 FILLER_311_1879 ();
 b15zdnd11an1n64x5 FILLER_311_1943 ();
 b15zdnd11an1n64x5 FILLER_311_2007 ();
 b15zdnd11an1n64x5 FILLER_311_2071 ();
 b15zdnd11an1n64x5 FILLER_311_2135 ();
 b15zdnd11an1n64x5 FILLER_311_2199 ();
 b15zdnd11an1n16x5 FILLER_311_2263 ();
 b15zdnd11an1n04x5 FILLER_311_2279 ();
 b15zdnd00an1n01x5 FILLER_311_2283 ();
 b15zdnd11an1n32x5 FILLER_312_8 ();
 b15zdnd11an1n16x5 FILLER_312_40 ();
 b15zdnd00an1n01x5 FILLER_312_56 ();
 b15zdnd11an1n64x5 FILLER_312_78 ();
 b15zdnd11an1n32x5 FILLER_312_142 ();
 b15zdnd11an1n08x5 FILLER_312_174 ();
 b15zdnd11an1n04x5 FILLER_312_182 ();
 b15zdnd11an1n08x5 FILLER_312_189 ();
 b15zdnd00an1n02x5 FILLER_312_197 ();
 b15zdnd00an1n01x5 FILLER_312_199 ();
 b15zdnd11an1n64x5 FILLER_312_242 ();
 b15zdnd11an1n64x5 FILLER_312_306 ();
 b15zdnd11an1n64x5 FILLER_312_370 ();
 b15zdnd11an1n64x5 FILLER_312_434 ();
 b15zdnd11an1n64x5 FILLER_312_498 ();
 b15zdnd11an1n64x5 FILLER_312_562 ();
 b15zdnd11an1n64x5 FILLER_312_626 ();
 b15zdnd11an1n16x5 FILLER_312_690 ();
 b15zdnd11an1n08x5 FILLER_312_706 ();
 b15zdnd11an1n04x5 FILLER_312_714 ();
 b15zdnd11an1n64x5 FILLER_312_726 ();
 b15zdnd11an1n64x5 FILLER_312_790 ();
 b15zdnd11an1n32x5 FILLER_312_854 ();
 b15zdnd11an1n16x5 FILLER_312_886 ();
 b15zdnd00an1n02x5 FILLER_312_902 ();
 b15zdnd00an1n01x5 FILLER_312_904 ();
 b15zdnd11an1n04x5 FILLER_312_908 ();
 b15zdnd00an1n02x5 FILLER_312_912 ();
 b15zdnd00an1n01x5 FILLER_312_914 ();
 b15zdnd11an1n64x5 FILLER_312_918 ();
 b15zdnd11an1n64x5 FILLER_312_982 ();
 b15zdnd11an1n64x5 FILLER_312_1046 ();
 b15zdnd11an1n64x5 FILLER_312_1110 ();
 b15zdnd11an1n64x5 FILLER_312_1174 ();
 b15zdnd11an1n64x5 FILLER_312_1238 ();
 b15zdnd00an1n02x5 FILLER_312_1302 ();
 b15zdnd11an1n64x5 FILLER_312_1315 ();
 b15zdnd11an1n64x5 FILLER_312_1379 ();
 b15zdnd11an1n64x5 FILLER_312_1443 ();
 b15zdnd11an1n64x5 FILLER_312_1507 ();
 b15zdnd11an1n64x5 FILLER_312_1571 ();
 b15zdnd11an1n64x5 FILLER_312_1635 ();
 b15zdnd11an1n64x5 FILLER_312_1699 ();
 b15zdnd11an1n64x5 FILLER_312_1763 ();
 b15zdnd11an1n64x5 FILLER_312_1827 ();
 b15zdnd11an1n64x5 FILLER_312_1891 ();
 b15zdnd11an1n64x5 FILLER_312_1955 ();
 b15zdnd11an1n64x5 FILLER_312_2019 ();
 b15zdnd11an1n64x5 FILLER_312_2083 ();
 b15zdnd11an1n04x5 FILLER_312_2147 ();
 b15zdnd00an1n02x5 FILLER_312_2151 ();
 b15zdnd00an1n01x5 FILLER_312_2153 ();
 b15zdnd11an1n64x5 FILLER_312_2162 ();
 b15zdnd11an1n16x5 FILLER_312_2226 ();
 b15zdnd11an1n08x5 FILLER_312_2242 ();
 b15zdnd11an1n04x5 FILLER_312_2250 ();
 b15zdnd11an1n08x5 FILLER_312_2262 ();
 b15zdnd11an1n04x5 FILLER_312_2270 ();
 b15zdnd00an1n02x5 FILLER_312_2274 ();
 b15zdnd11an1n32x5 FILLER_313_0 ();
 b15zdnd11an1n16x5 FILLER_313_32 ();
 b15zdnd11an1n08x5 FILLER_313_48 ();
 b15zdnd11an1n04x5 FILLER_313_56 ();
 b15zdnd00an1n01x5 FILLER_313_60 ();
 b15zdnd11an1n64x5 FILLER_313_87 ();
 b15zdnd11an1n08x5 FILLER_313_151 ();
 b15zdnd11an1n64x5 FILLER_313_211 ();
 b15zdnd11an1n64x5 FILLER_313_275 ();
 b15zdnd11an1n64x5 FILLER_313_339 ();
 b15zdnd11an1n64x5 FILLER_313_403 ();
 b15zdnd11an1n64x5 FILLER_313_467 ();
 b15zdnd11an1n64x5 FILLER_313_531 ();
 b15zdnd11an1n64x5 FILLER_313_595 ();
 b15zdnd11an1n64x5 FILLER_313_659 ();
 b15zdnd11an1n64x5 FILLER_313_723 ();
 b15zdnd11an1n64x5 FILLER_313_787 ();
 b15zdnd11an1n64x5 FILLER_313_851 ();
 b15zdnd11an1n64x5 FILLER_313_915 ();
 b15zdnd11an1n64x5 FILLER_313_979 ();
 b15zdnd11an1n64x5 FILLER_313_1043 ();
 b15zdnd11an1n64x5 FILLER_313_1107 ();
 b15zdnd11an1n64x5 FILLER_313_1171 ();
 b15zdnd11an1n64x5 FILLER_313_1235 ();
 b15zdnd11an1n64x5 FILLER_313_1299 ();
 b15zdnd11an1n64x5 FILLER_313_1363 ();
 b15zdnd11an1n64x5 FILLER_313_1427 ();
 b15zdnd11an1n64x5 FILLER_313_1491 ();
 b15zdnd11an1n64x5 FILLER_313_1555 ();
 b15zdnd11an1n64x5 FILLER_313_1619 ();
 b15zdnd11an1n64x5 FILLER_313_1683 ();
 b15zdnd11an1n64x5 FILLER_313_1747 ();
 b15zdnd11an1n64x5 FILLER_313_1811 ();
 b15zdnd11an1n64x5 FILLER_313_1875 ();
 b15zdnd11an1n64x5 FILLER_313_1939 ();
 b15zdnd11an1n64x5 FILLER_313_2003 ();
 b15zdnd11an1n64x5 FILLER_313_2067 ();
 b15zdnd11an1n64x5 FILLER_313_2131 ();
 b15zdnd11an1n64x5 FILLER_313_2195 ();
 b15zdnd11an1n16x5 FILLER_313_2259 ();
 b15zdnd11an1n08x5 FILLER_313_2275 ();
 b15zdnd00an1n01x5 FILLER_313_2283 ();
 b15zdnd11an1n64x5 FILLER_314_8 ();
 b15zdnd00an1n02x5 FILLER_314_72 ();
 b15zdnd00an1n01x5 FILLER_314_74 ();
 b15zdnd11an1n64x5 FILLER_314_82 ();
 b15zdnd11an1n16x5 FILLER_314_146 ();
 b15zdnd11an1n08x5 FILLER_314_162 ();
 b15zdnd11an1n04x5 FILLER_314_170 ();
 b15zdnd00an1n02x5 FILLER_314_174 ();
 b15zdnd00an1n01x5 FILLER_314_176 ();
 b15zdnd11an1n04x5 FILLER_314_180 ();
 b15zdnd11an1n16x5 FILLER_314_187 ();
 b15zdnd11an1n04x5 FILLER_314_203 ();
 b15zdnd00an1n02x5 FILLER_314_207 ();
 b15zdnd00an1n01x5 FILLER_314_209 ();
 b15zdnd11an1n64x5 FILLER_314_252 ();
 b15zdnd11an1n64x5 FILLER_314_316 ();
 b15zdnd11an1n64x5 FILLER_314_380 ();
 b15zdnd11an1n64x5 FILLER_314_444 ();
 b15zdnd11an1n64x5 FILLER_314_508 ();
 b15zdnd11an1n64x5 FILLER_314_572 ();
 b15zdnd11an1n64x5 FILLER_314_636 ();
 b15zdnd11an1n16x5 FILLER_314_700 ();
 b15zdnd00an1n02x5 FILLER_314_716 ();
 b15zdnd11an1n64x5 FILLER_314_726 ();
 b15zdnd11an1n64x5 FILLER_314_790 ();
 b15zdnd11an1n64x5 FILLER_314_854 ();
 b15zdnd11an1n64x5 FILLER_314_918 ();
 b15zdnd11an1n64x5 FILLER_314_982 ();
 b15zdnd11an1n64x5 FILLER_314_1046 ();
 b15zdnd11an1n64x5 FILLER_314_1110 ();
 b15zdnd11an1n64x5 FILLER_314_1174 ();
 b15zdnd11an1n64x5 FILLER_314_1238 ();
 b15zdnd11an1n64x5 FILLER_314_1302 ();
 b15zdnd11an1n64x5 FILLER_314_1366 ();
 b15zdnd11an1n64x5 FILLER_314_1430 ();
 b15zdnd11an1n64x5 FILLER_314_1494 ();
 b15zdnd11an1n64x5 FILLER_314_1558 ();
 b15zdnd11an1n64x5 FILLER_314_1622 ();
 b15zdnd11an1n64x5 FILLER_314_1686 ();
 b15zdnd11an1n64x5 FILLER_314_1750 ();
 b15zdnd11an1n64x5 FILLER_314_1814 ();
 b15zdnd11an1n64x5 FILLER_314_1878 ();
 b15zdnd11an1n64x5 FILLER_314_1942 ();
 b15zdnd11an1n64x5 FILLER_314_2006 ();
 b15zdnd11an1n64x5 FILLER_314_2070 ();
 b15zdnd11an1n16x5 FILLER_314_2134 ();
 b15zdnd11an1n04x5 FILLER_314_2150 ();
 b15zdnd11an1n64x5 FILLER_314_2162 ();
 b15zdnd11an1n32x5 FILLER_314_2226 ();
 b15zdnd11an1n16x5 FILLER_314_2258 ();
 b15zdnd00an1n02x5 FILLER_314_2274 ();
 b15zdnd11an1n64x5 FILLER_315_0 ();
 b15zdnd11an1n64x5 FILLER_315_64 ();
 b15zdnd11an1n64x5 FILLER_315_128 ();
 b15zdnd11an1n16x5 FILLER_315_192 ();
 b15zdnd00an1n02x5 FILLER_315_208 ();
 b15zdnd11an1n64x5 FILLER_315_217 ();
 b15zdnd11an1n64x5 FILLER_315_281 ();
 b15zdnd11an1n64x5 FILLER_315_345 ();
 b15zdnd11an1n64x5 FILLER_315_409 ();
 b15zdnd11an1n64x5 FILLER_315_473 ();
 b15zdnd11an1n64x5 FILLER_315_537 ();
 b15zdnd11an1n64x5 FILLER_315_601 ();
 b15zdnd11an1n64x5 FILLER_315_665 ();
 b15zdnd11an1n16x5 FILLER_315_729 ();
 b15zdnd00an1n02x5 FILLER_315_745 ();
 b15zdnd00an1n01x5 FILLER_315_747 ();
 b15zdnd11an1n64x5 FILLER_315_751 ();
 b15zdnd11an1n64x5 FILLER_315_815 ();
 b15zdnd11an1n64x5 FILLER_315_879 ();
 b15zdnd11an1n64x5 FILLER_315_943 ();
 b15zdnd11an1n64x5 FILLER_315_1007 ();
 b15zdnd11an1n64x5 FILLER_315_1071 ();
 b15zdnd11an1n64x5 FILLER_315_1135 ();
 b15zdnd11an1n64x5 FILLER_315_1199 ();
 b15zdnd11an1n32x5 FILLER_315_1263 ();
 b15zdnd11an1n08x5 FILLER_315_1295 ();
 b15zdnd11an1n64x5 FILLER_315_1312 ();
 b15zdnd11an1n64x5 FILLER_315_1376 ();
 b15zdnd11an1n64x5 FILLER_315_1440 ();
 b15zdnd11an1n08x5 FILLER_315_1504 ();
 b15zdnd00an1n02x5 FILLER_315_1512 ();
 b15zdnd00an1n01x5 FILLER_315_1514 ();
 b15zdnd11an1n64x5 FILLER_315_1518 ();
 b15zdnd11an1n64x5 FILLER_315_1582 ();
 b15zdnd11an1n64x5 FILLER_315_1646 ();
 b15zdnd11an1n64x5 FILLER_315_1710 ();
 b15zdnd11an1n64x5 FILLER_315_1774 ();
 b15zdnd11an1n64x5 FILLER_315_1838 ();
 b15zdnd11an1n64x5 FILLER_315_1902 ();
 b15zdnd11an1n64x5 FILLER_315_1966 ();
 b15zdnd11an1n64x5 FILLER_315_2030 ();
 b15zdnd11an1n64x5 FILLER_315_2094 ();
 b15zdnd11an1n64x5 FILLER_315_2158 ();
 b15zdnd11an1n32x5 FILLER_315_2222 ();
 b15zdnd11an1n16x5 FILLER_315_2254 ();
 b15zdnd11an1n08x5 FILLER_315_2270 ();
 b15zdnd11an1n04x5 FILLER_315_2278 ();
 b15zdnd00an1n02x5 FILLER_315_2282 ();
 b15zdnd11an1n64x5 FILLER_316_8 ();
 b15zdnd11an1n64x5 FILLER_316_72 ();
 b15zdnd11an1n64x5 FILLER_316_136 ();
 b15zdnd11an1n64x5 FILLER_316_200 ();
 b15zdnd11an1n64x5 FILLER_316_264 ();
 b15zdnd11an1n16x5 FILLER_316_328 ();
 b15zdnd11an1n04x5 FILLER_316_344 ();
 b15zdnd00an1n01x5 FILLER_316_348 ();
 b15zdnd11an1n64x5 FILLER_316_358 ();
 b15zdnd11an1n64x5 FILLER_316_422 ();
 b15zdnd11an1n64x5 FILLER_316_486 ();
 b15zdnd11an1n64x5 FILLER_316_550 ();
 b15zdnd11an1n64x5 FILLER_316_614 ();
 b15zdnd11an1n32x5 FILLER_316_678 ();
 b15zdnd11an1n08x5 FILLER_316_710 ();
 b15zdnd00an1n02x5 FILLER_316_726 ();
 b15zdnd11an1n08x5 FILLER_316_780 ();
 b15zdnd11an1n04x5 FILLER_316_805 ();
 b15zdnd00an1n01x5 FILLER_316_809 ();
 b15zdnd11an1n64x5 FILLER_316_827 ();
 b15zdnd11an1n64x5 FILLER_316_891 ();
 b15zdnd11an1n64x5 FILLER_316_955 ();
 b15zdnd11an1n64x5 FILLER_316_1019 ();
 b15zdnd11an1n64x5 FILLER_316_1083 ();
 b15zdnd11an1n16x5 FILLER_316_1147 ();
 b15zdnd11an1n64x5 FILLER_316_1194 ();
 b15zdnd11an1n08x5 FILLER_316_1258 ();
 b15zdnd11an1n64x5 FILLER_316_1275 ();
 b15zdnd11an1n64x5 FILLER_316_1339 ();
 b15zdnd11an1n64x5 FILLER_316_1403 ();
 b15zdnd11an1n16x5 FILLER_316_1467 ();
 b15zdnd11an1n04x5 FILLER_316_1483 ();
 b15zdnd00an1n01x5 FILLER_316_1487 ();
 b15zdnd11an1n64x5 FILLER_316_1540 ();
 b15zdnd11an1n64x5 FILLER_316_1604 ();
 b15zdnd11an1n64x5 FILLER_316_1668 ();
 b15zdnd11an1n64x5 FILLER_316_1732 ();
 b15zdnd11an1n64x5 FILLER_316_1796 ();
 b15zdnd11an1n64x5 FILLER_316_1860 ();
 b15zdnd11an1n64x5 FILLER_316_1924 ();
 b15zdnd11an1n64x5 FILLER_316_1988 ();
 b15zdnd11an1n64x5 FILLER_316_2052 ();
 b15zdnd11an1n32x5 FILLER_316_2116 ();
 b15zdnd11an1n04x5 FILLER_316_2148 ();
 b15zdnd00an1n02x5 FILLER_316_2152 ();
 b15zdnd11an1n64x5 FILLER_316_2162 ();
 b15zdnd11an1n32x5 FILLER_316_2226 ();
 b15zdnd11an1n16x5 FILLER_316_2258 ();
 b15zdnd00an1n02x5 FILLER_316_2274 ();
 b15zdnd11an1n64x5 FILLER_317_0 ();
 b15zdnd11an1n64x5 FILLER_317_64 ();
 b15zdnd11an1n64x5 FILLER_317_128 ();
 b15zdnd11an1n64x5 FILLER_317_192 ();
 b15zdnd11an1n64x5 FILLER_317_256 ();
 b15zdnd11an1n16x5 FILLER_317_320 ();
 b15zdnd11an1n08x5 FILLER_317_336 ();
 b15zdnd00an1n02x5 FILLER_317_344 ();
 b15zdnd11an1n64x5 FILLER_317_349 ();
 b15zdnd11an1n64x5 FILLER_317_413 ();
 b15zdnd11an1n64x5 FILLER_317_477 ();
 b15zdnd11an1n64x5 FILLER_317_541 ();
 b15zdnd11an1n64x5 FILLER_317_605 ();
 b15zdnd11an1n32x5 FILLER_317_669 ();
 b15zdnd11an1n16x5 FILLER_317_701 ();
 b15zdnd11an1n04x5 FILLER_317_717 ();
 b15zdnd00an1n01x5 FILLER_317_721 ();
 b15zdnd11an1n64x5 FILLER_317_774 ();
 b15zdnd11an1n64x5 FILLER_317_838 ();
 b15zdnd11an1n64x5 FILLER_317_902 ();
 b15zdnd11an1n64x5 FILLER_317_966 ();
 b15zdnd11an1n64x5 FILLER_317_1030 ();
 b15zdnd11an1n64x5 FILLER_317_1094 ();
 b15zdnd11an1n64x5 FILLER_317_1158 ();
 b15zdnd11an1n64x5 FILLER_317_1222 ();
 b15zdnd11an1n64x5 FILLER_317_1286 ();
 b15zdnd11an1n64x5 FILLER_317_1350 ();
 b15zdnd11an1n64x5 FILLER_317_1414 ();
 b15zdnd11an1n08x5 FILLER_317_1478 ();
 b15zdnd00an1n01x5 FILLER_317_1486 ();
 b15zdnd11an1n64x5 FILLER_317_1539 ();
 b15zdnd11an1n64x5 FILLER_317_1603 ();
 b15zdnd11an1n64x5 FILLER_317_1667 ();
 b15zdnd11an1n64x5 FILLER_317_1731 ();
 b15zdnd11an1n64x5 FILLER_317_1798 ();
 b15zdnd11an1n64x5 FILLER_317_1862 ();
 b15zdnd11an1n64x5 FILLER_317_1926 ();
 b15zdnd11an1n64x5 FILLER_317_1990 ();
 b15zdnd11an1n64x5 FILLER_317_2054 ();
 b15zdnd11an1n64x5 FILLER_317_2118 ();
 b15zdnd11an1n64x5 FILLER_317_2182 ();
 b15zdnd11an1n32x5 FILLER_317_2246 ();
 b15zdnd11an1n04x5 FILLER_317_2278 ();
 b15zdnd00an1n02x5 FILLER_317_2282 ();
 b15zdnd11an1n64x5 FILLER_318_8 ();
 b15zdnd11an1n64x5 FILLER_318_72 ();
 b15zdnd11an1n64x5 FILLER_318_136 ();
 b15zdnd11an1n64x5 FILLER_318_200 ();
 b15zdnd11an1n32x5 FILLER_318_264 ();
 b15zdnd11an1n16x5 FILLER_318_296 ();
 b15zdnd11an1n04x5 FILLER_318_315 ();
 b15zdnd11an1n64x5 FILLER_318_371 ();
 b15zdnd11an1n64x5 FILLER_318_435 ();
 b15zdnd11an1n64x5 FILLER_318_499 ();
 b15zdnd11an1n64x5 FILLER_318_563 ();
 b15zdnd11an1n64x5 FILLER_318_627 ();
 b15zdnd11an1n16x5 FILLER_318_691 ();
 b15zdnd11an1n08x5 FILLER_318_707 ();
 b15zdnd00an1n02x5 FILLER_318_715 ();
 b15zdnd00an1n01x5 FILLER_318_717 ();
 b15zdnd11an1n16x5 FILLER_318_726 ();
 b15zdnd00an1n02x5 FILLER_318_742 ();
 b15zdnd00an1n01x5 FILLER_318_744 ();
 b15zdnd11an1n04x5 FILLER_318_748 ();
 b15zdnd11an1n04x5 FILLER_318_755 ();
 b15zdnd11an1n64x5 FILLER_318_762 ();
 b15zdnd11an1n32x5 FILLER_318_826 ();
 b15zdnd11an1n16x5 FILLER_318_858 ();
 b15zdnd11an1n08x5 FILLER_318_874 ();
 b15zdnd11an1n64x5 FILLER_318_934 ();
 b15zdnd11an1n16x5 FILLER_318_998 ();
 b15zdnd11an1n08x5 FILLER_318_1014 ();
 b15zdnd00an1n01x5 FILLER_318_1022 ();
 b15zdnd11an1n16x5 FILLER_318_1054 ();
 b15zdnd00an1n01x5 FILLER_318_1070 ();
 b15zdnd11an1n64x5 FILLER_318_1074 ();
 b15zdnd11an1n64x5 FILLER_318_1138 ();
 b15zdnd11an1n64x5 FILLER_318_1202 ();
 b15zdnd11an1n64x5 FILLER_318_1266 ();
 b15zdnd11an1n32x5 FILLER_318_1330 ();
 b15zdnd11an1n16x5 FILLER_318_1362 ();
 b15zdnd11an1n08x5 FILLER_318_1378 ();
 b15zdnd00an1n02x5 FILLER_318_1386 ();
 b15zdnd00an1n01x5 FILLER_318_1388 ();
 b15zdnd11an1n04x5 FILLER_318_1397 ();
 b15zdnd11an1n64x5 FILLER_318_1413 ();
 b15zdnd11an1n16x5 FILLER_318_1477 ();
 b15zdnd11an1n08x5 FILLER_318_1493 ();
 b15zdnd11an1n04x5 FILLER_318_1501 ();
 b15zdnd00an1n01x5 FILLER_318_1505 ();
 b15zdnd11an1n04x5 FILLER_318_1509 ();
 b15zdnd11an1n04x5 FILLER_318_1516 ();
 b15zdnd11an1n64x5 FILLER_318_1523 ();
 b15zdnd11an1n16x5 FILLER_318_1587 ();
 b15zdnd11an1n04x5 FILLER_318_1603 ();
 b15zdnd11an1n64x5 FILLER_318_1634 ();
 b15zdnd11an1n64x5 FILLER_318_1698 ();
 b15zdnd11an1n32x5 FILLER_318_1762 ();
 b15zdnd00an1n01x5 FILLER_318_1794 ();
 b15zdnd11an1n64x5 FILLER_318_1798 ();
 b15zdnd11an1n64x5 FILLER_318_1862 ();
 b15zdnd11an1n64x5 FILLER_318_1926 ();
 b15zdnd11an1n64x5 FILLER_318_1990 ();
 b15zdnd11an1n64x5 FILLER_318_2054 ();
 b15zdnd11an1n32x5 FILLER_318_2118 ();
 b15zdnd11an1n04x5 FILLER_318_2150 ();
 b15zdnd11an1n64x5 FILLER_318_2162 ();
 b15zdnd11an1n32x5 FILLER_318_2226 ();
 b15zdnd11an1n16x5 FILLER_318_2258 ();
 b15zdnd00an1n02x5 FILLER_318_2274 ();
 b15zdnd11an1n64x5 FILLER_319_0 ();
 b15zdnd11an1n64x5 FILLER_319_64 ();
 b15zdnd11an1n64x5 FILLER_319_128 ();
 b15zdnd11an1n64x5 FILLER_319_192 ();
 b15zdnd11an1n16x5 FILLER_319_256 ();
 b15zdnd00an1n02x5 FILLER_319_272 ();
 b15zdnd11an1n08x5 FILLER_319_301 ();
 b15zdnd11an1n04x5 FILLER_319_309 ();
 b15zdnd11an1n04x5 FILLER_319_316 ();
 b15zdnd11an1n08x5 FILLER_319_323 ();
 b15zdnd00an1n01x5 FILLER_319_331 ();
 b15zdnd11an1n64x5 FILLER_319_384 ();
 b15zdnd11an1n08x5 FILLER_319_448 ();
 b15zdnd11an1n04x5 FILLER_319_456 ();
 b15zdnd00an1n02x5 FILLER_319_460 ();
 b15zdnd11an1n08x5 FILLER_319_465 ();
 b15zdnd00an1n02x5 FILLER_319_473 ();
 b15zdnd11an1n64x5 FILLER_319_517 ();
 b15zdnd11an1n64x5 FILLER_319_581 ();
 b15zdnd11an1n64x5 FILLER_319_645 ();
 b15zdnd11an1n32x5 FILLER_319_709 ();
 b15zdnd11an1n04x5 FILLER_319_741 ();
 b15zdnd00an1n02x5 FILLER_319_745 ();
 b15zdnd00an1n01x5 FILLER_319_747 ();
 b15zdnd11an1n04x5 FILLER_319_751 ();
 b15zdnd11an1n64x5 FILLER_319_758 ();
 b15zdnd11an1n64x5 FILLER_319_822 ();
 b15zdnd11an1n08x5 FILLER_319_886 ();
 b15zdnd00an1n02x5 FILLER_319_894 ();
 b15zdnd00an1n01x5 FILLER_319_896 ();
 b15zdnd11an1n04x5 FILLER_319_900 ();
 b15zdnd00an1n02x5 FILLER_319_904 ();
 b15zdnd00an1n01x5 FILLER_319_906 ();
 b15zdnd11an1n16x5 FILLER_319_910 ();
 b15zdnd11an1n04x5 FILLER_319_926 ();
 b15zdnd00an1n02x5 FILLER_319_930 ();
 b15zdnd00an1n01x5 FILLER_319_932 ();
 b15zdnd11an1n04x5 FILLER_319_950 ();
 b15zdnd11an1n64x5 FILLER_319_971 ();
 b15zdnd11an1n08x5 FILLER_319_1035 ();
 b15zdnd00an1n01x5 FILLER_319_1043 ();
 b15zdnd11an1n16x5 FILLER_319_1096 ();
 b15zdnd11an1n08x5 FILLER_319_1112 ();
 b15zdnd11an1n04x5 FILLER_319_1120 ();
 b15zdnd11an1n04x5 FILLER_319_1127 ();
 b15zdnd11an1n04x5 FILLER_319_1134 ();
 b15zdnd11an1n64x5 FILLER_319_1141 ();
 b15zdnd11an1n64x5 FILLER_319_1205 ();
 b15zdnd11an1n64x5 FILLER_319_1269 ();
 b15zdnd11an1n32x5 FILLER_319_1333 ();
 b15zdnd11an1n04x5 FILLER_319_1365 ();
 b15zdnd00an1n01x5 FILLER_319_1369 ();
 b15zdnd11an1n04x5 FILLER_319_1378 ();
 b15zdnd11an1n04x5 FILLER_319_1402 ();
 b15zdnd00an1n02x5 FILLER_319_1406 ();
 b15zdnd11an1n64x5 FILLER_319_1428 ();
 b15zdnd11an1n08x5 FILLER_319_1492 ();
 b15zdnd11an1n04x5 FILLER_319_1500 ();
 b15zdnd00an1n01x5 FILLER_319_1504 ();
 b15zdnd11an1n04x5 FILLER_319_1508 ();
 b15zdnd11an1n64x5 FILLER_319_1515 ();
 b15zdnd11an1n16x5 FILLER_319_1579 ();
 b15zdnd11an1n08x5 FILLER_319_1595 ();
 b15zdnd11an1n04x5 FILLER_319_1603 ();
 b15zdnd11an1n08x5 FILLER_319_1610 ();
 b15zdnd00an1n01x5 FILLER_319_1618 ();
 b15zdnd11an1n64x5 FILLER_319_1622 ();
 b15zdnd11an1n64x5 FILLER_319_1686 ();
 b15zdnd11an1n16x5 FILLER_319_1750 ();
 b15zdnd11an1n04x5 FILLER_319_1766 ();
 b15zdnd11an1n64x5 FILLER_319_1822 ();
 b15zdnd11an1n64x5 FILLER_319_1886 ();
 b15zdnd11an1n64x5 FILLER_319_1950 ();
 b15zdnd11an1n64x5 FILLER_319_2014 ();
 b15zdnd11an1n64x5 FILLER_319_2078 ();
 b15zdnd11an1n64x5 FILLER_319_2142 ();
 b15zdnd11an1n64x5 FILLER_319_2206 ();
 b15zdnd11an1n08x5 FILLER_319_2270 ();
 b15zdnd11an1n04x5 FILLER_319_2278 ();
 b15zdnd00an1n02x5 FILLER_319_2282 ();
 b15zdnd11an1n64x5 FILLER_320_8 ();
 b15zdnd11an1n64x5 FILLER_320_72 ();
 b15zdnd11an1n64x5 FILLER_320_136 ();
 b15zdnd11an1n64x5 FILLER_320_200 ();
 b15zdnd11an1n08x5 FILLER_320_264 ();
 b15zdnd00an1n01x5 FILLER_320_272 ();
 b15zdnd11an1n16x5 FILLER_320_276 ();
 b15zdnd00an1n01x5 FILLER_320_292 ();
 b15zdnd11an1n04x5 FILLER_320_345 ();
 b15zdnd11an1n04x5 FILLER_320_358 ();
 b15zdnd00an1n01x5 FILLER_320_362 ();
 b15zdnd11an1n64x5 FILLER_320_366 ();
 b15zdnd11an1n04x5 FILLER_320_430 ();
 b15zdnd00an1n01x5 FILLER_320_434 ();
 b15zdnd11an1n32x5 FILLER_320_487 ();
 b15zdnd11an1n16x5 FILLER_320_519 ();
 b15zdnd11an1n08x5 FILLER_320_535 ();
 b15zdnd00an1n01x5 FILLER_320_543 ();
 b15zdnd11an1n04x5 FILLER_320_553 ();
 b15zdnd00an1n02x5 FILLER_320_557 ();
 b15zdnd00an1n01x5 FILLER_320_559 ();
 b15zdnd11an1n04x5 FILLER_320_587 ();
 b15zdnd11an1n64x5 FILLER_320_594 ();
 b15zdnd11an1n32x5 FILLER_320_658 ();
 b15zdnd11an1n16x5 FILLER_320_690 ();
 b15zdnd11an1n08x5 FILLER_320_706 ();
 b15zdnd11an1n04x5 FILLER_320_714 ();
 b15zdnd11an1n64x5 FILLER_320_726 ();
 b15zdnd11an1n64x5 FILLER_320_790 ();
 b15zdnd11an1n32x5 FILLER_320_854 ();
 b15zdnd11an1n16x5 FILLER_320_886 ();
 b15zdnd11an1n32x5 FILLER_320_905 ();
 b15zdnd11an1n04x5 FILLER_320_937 ();
 b15zdnd00an1n02x5 FILLER_320_941 ();
 b15zdnd11an1n32x5 FILLER_320_995 ();
 b15zdnd11an1n16x5 FILLER_320_1027 ();
 b15zdnd11an1n16x5 FILLER_320_1046 ();
 b15zdnd11an1n04x5 FILLER_320_1065 ();
 b15zdnd11an1n32x5 FILLER_320_1072 ();
 b15zdnd11an1n64x5 FILLER_320_1156 ();
 b15zdnd11an1n64x5 FILLER_320_1220 ();
 b15zdnd11an1n64x5 FILLER_320_1284 ();
 b15zdnd11an1n16x5 FILLER_320_1348 ();
 b15zdnd11an1n04x5 FILLER_320_1364 ();
 b15zdnd00an1n02x5 FILLER_320_1368 ();
 b15zdnd11an1n04x5 FILLER_320_1373 ();
 b15zdnd00an1n01x5 FILLER_320_1377 ();
 b15zdnd11an1n08x5 FILLER_320_1392 ();
 b15zdnd11an1n04x5 FILLER_320_1400 ();
 b15zdnd00an1n02x5 FILLER_320_1404 ();
 b15zdnd11an1n64x5 FILLER_320_1426 ();
 b15zdnd11an1n64x5 FILLER_320_1490 ();
 b15zdnd11an1n64x5 FILLER_320_1554 ();
 b15zdnd00an1n02x5 FILLER_320_1618 ();
 b15zdnd00an1n01x5 FILLER_320_1620 ();
 b15zdnd11an1n04x5 FILLER_320_1624 ();
 b15zdnd00an1n01x5 FILLER_320_1628 ();
 b15zdnd11an1n04x5 FILLER_320_1632 ();
 b15zdnd11an1n64x5 FILLER_320_1656 ();
 b15zdnd11an1n32x5 FILLER_320_1720 ();
 b15zdnd11an1n08x5 FILLER_320_1752 ();
 b15zdnd00an1n02x5 FILLER_320_1760 ();
 b15zdnd00an1n01x5 FILLER_320_1762 ();
 b15zdnd11an1n16x5 FILLER_320_1774 ();
 b15zdnd11an1n04x5 FILLER_320_1790 ();
 b15zdnd00an1n02x5 FILLER_320_1794 ();
 b15zdnd11an1n64x5 FILLER_320_1799 ();
 b15zdnd11an1n16x5 FILLER_320_1863 ();
 b15zdnd11an1n08x5 FILLER_320_1879 ();
 b15zdnd00an1n01x5 FILLER_320_1887 ();
 b15zdnd11an1n64x5 FILLER_320_1940 ();
 b15zdnd11an1n64x5 FILLER_320_2004 ();
 b15zdnd11an1n64x5 FILLER_320_2068 ();
 b15zdnd11an1n16x5 FILLER_320_2132 ();
 b15zdnd11an1n04x5 FILLER_320_2148 ();
 b15zdnd00an1n02x5 FILLER_320_2152 ();
 b15zdnd11an1n64x5 FILLER_320_2162 ();
 b15zdnd11an1n32x5 FILLER_320_2226 ();
 b15zdnd11an1n16x5 FILLER_320_2258 ();
 b15zdnd00an1n02x5 FILLER_320_2274 ();
 b15zdnd11an1n64x5 FILLER_321_0 ();
 b15zdnd11an1n64x5 FILLER_321_64 ();
 b15zdnd11an1n64x5 FILLER_321_128 ();
 b15zdnd11an1n64x5 FILLER_321_192 ();
 b15zdnd11an1n32x5 FILLER_321_256 ();
 b15zdnd11an1n08x5 FILLER_321_340 ();
 b15zdnd00an1n01x5 FILLER_321_348 ();
 b15zdnd11an1n04x5 FILLER_321_352 ();
 b15zdnd11an1n04x5 FILLER_321_359 ();
 b15zdnd11an1n64x5 FILLER_321_366 ();
 b15zdnd11an1n16x5 FILLER_321_430 ();
 b15zdnd11an1n32x5 FILLER_321_488 ();
 b15zdnd11an1n16x5 FILLER_321_520 ();
 b15zdnd11an1n08x5 FILLER_321_536 ();
 b15zdnd11an1n04x5 FILLER_321_544 ();
 b15zdnd11an1n04x5 FILLER_321_600 ();
 b15zdnd11an1n64x5 FILLER_321_613 ();
 b15zdnd11an1n64x5 FILLER_321_677 ();
 b15zdnd11an1n64x5 FILLER_321_741 ();
 b15zdnd11an1n64x5 FILLER_321_805 ();
 b15zdnd11an1n64x5 FILLER_321_869 ();
 b15zdnd11an1n16x5 FILLER_321_933 ();
 b15zdnd11an1n04x5 FILLER_321_949 ();
 b15zdnd11an1n04x5 FILLER_321_956 ();
 b15zdnd11an1n04x5 FILLER_321_963 ();
 b15zdnd11an1n32x5 FILLER_321_970 ();
 b15zdnd11an1n08x5 FILLER_321_1002 ();
 b15zdnd11an1n04x5 FILLER_321_1010 ();
 b15zdnd00an1n02x5 FILLER_321_1014 ();
 b15zdnd11an1n32x5 FILLER_321_1068 ();
 b15zdnd00an1n02x5 FILLER_321_1100 ();
 b15zdnd00an1n01x5 FILLER_321_1102 ();
 b15zdnd11an1n04x5 FILLER_321_1106 ();
 b15zdnd11an1n64x5 FILLER_321_1137 ();
 b15zdnd11an1n32x5 FILLER_321_1201 ();
 b15zdnd11an1n08x5 FILLER_321_1233 ();
 b15zdnd00an1n01x5 FILLER_321_1241 ();
 b15zdnd11an1n64x5 FILLER_321_1245 ();
 b15zdnd11an1n32x5 FILLER_321_1309 ();
 b15zdnd00an1n02x5 FILLER_321_1341 ();
 b15zdnd00an1n01x5 FILLER_321_1343 ();
 b15zdnd11an1n16x5 FILLER_321_1396 ();
 b15zdnd11an1n04x5 FILLER_321_1412 ();
 b15zdnd00an1n02x5 FILLER_321_1416 ();
 b15zdnd00an1n01x5 FILLER_321_1418 ();
 b15zdnd11an1n64x5 FILLER_321_1433 ();
 b15zdnd11an1n64x5 FILLER_321_1497 ();
 b15zdnd11an1n32x5 FILLER_321_1561 ();
 b15zdnd11an1n04x5 FILLER_321_1593 ();
 b15zdnd11an1n64x5 FILLER_321_1649 ();
 b15zdnd11an1n64x5 FILLER_321_1713 ();
 b15zdnd11an1n64x5 FILLER_321_1777 ();
 b15zdnd11an1n64x5 FILLER_321_1841 ();
 b15zdnd11an1n04x5 FILLER_321_1905 ();
 b15zdnd00an1n02x5 FILLER_321_1909 ();
 b15zdnd11an1n04x5 FILLER_321_1914 ();
 b15zdnd11an1n64x5 FILLER_321_1921 ();
 b15zdnd11an1n64x5 FILLER_321_1985 ();
 b15zdnd11an1n64x5 FILLER_321_2049 ();
 b15zdnd11an1n64x5 FILLER_321_2113 ();
 b15zdnd11an1n64x5 FILLER_321_2177 ();
 b15zdnd11an1n32x5 FILLER_321_2241 ();
 b15zdnd11an1n08x5 FILLER_321_2273 ();
 b15zdnd00an1n02x5 FILLER_321_2281 ();
 b15zdnd00an1n01x5 FILLER_321_2283 ();
 b15zdnd11an1n64x5 FILLER_322_8 ();
 b15zdnd11an1n08x5 FILLER_322_72 ();
 b15zdnd00an1n02x5 FILLER_322_80 ();
 b15zdnd11an1n64x5 FILLER_322_85 ();
 b15zdnd11an1n64x5 FILLER_322_149 ();
 b15zdnd11an1n64x5 FILLER_322_213 ();
 b15zdnd11an1n16x5 FILLER_322_277 ();
 b15zdnd00an1n01x5 FILLER_322_293 ();
 b15zdnd11an1n04x5 FILLER_322_303 ();
 b15zdnd00an1n02x5 FILLER_322_307 ();
 b15zdnd11an1n04x5 FILLER_322_312 ();
 b15zdnd11an1n16x5 FILLER_322_319 ();
 b15zdnd11an1n08x5 FILLER_322_335 ();
 b15zdnd00an1n01x5 FILLER_322_343 ();
 b15zdnd11an1n64x5 FILLER_322_347 ();
 b15zdnd11an1n32x5 FILLER_322_411 ();
 b15zdnd11an1n08x5 FILLER_322_443 ();
 b15zdnd00an1n01x5 FILLER_322_451 ();
 b15zdnd11an1n04x5 FILLER_322_455 ();
 b15zdnd00an1n01x5 FILLER_322_459 ();
 b15zdnd11an1n64x5 FILLER_322_463 ();
 b15zdnd11an1n16x5 FILLER_322_527 ();
 b15zdnd11an1n08x5 FILLER_322_543 ();
 b15zdnd11an1n04x5 FILLER_322_551 ();
 b15zdnd11an1n04x5 FILLER_322_558 ();
 b15zdnd11an1n64x5 FILLER_322_614 ();
 b15zdnd11an1n32x5 FILLER_322_678 ();
 b15zdnd11an1n08x5 FILLER_322_710 ();
 b15zdnd11an1n64x5 FILLER_322_726 ();
 b15zdnd11an1n64x5 FILLER_322_790 ();
 b15zdnd11an1n64x5 FILLER_322_854 ();
 b15zdnd11an1n64x5 FILLER_322_918 ();
 b15zdnd11an1n32x5 FILLER_322_982 ();
 b15zdnd11an1n16x5 FILLER_322_1014 ();
 b15zdnd11an1n04x5 FILLER_322_1030 ();
 b15zdnd11an1n04x5 FILLER_322_1037 ();
 b15zdnd11an1n64x5 FILLER_322_1044 ();
 b15zdnd11an1n64x5 FILLER_322_1108 ();
 b15zdnd11an1n64x5 FILLER_322_1172 ();
 b15zdnd11an1n04x5 FILLER_322_1236 ();
 b15zdnd00an1n01x5 FILLER_322_1240 ();
 b15zdnd11an1n64x5 FILLER_322_1244 ();
 b15zdnd11an1n32x5 FILLER_322_1308 ();
 b15zdnd11an1n16x5 FILLER_322_1340 ();
 b15zdnd11an1n04x5 FILLER_322_1356 ();
 b15zdnd00an1n02x5 FILLER_322_1360 ();
 b15zdnd11an1n04x5 FILLER_322_1365 ();
 b15zdnd11an1n08x5 FILLER_322_1372 ();
 b15zdnd00an1n01x5 FILLER_322_1380 ();
 b15zdnd11an1n64x5 FILLER_322_1398 ();
 b15zdnd11an1n64x5 FILLER_322_1462 ();
 b15zdnd11an1n64x5 FILLER_322_1526 ();
 b15zdnd11an1n64x5 FILLER_322_1590 ();
 b15zdnd11an1n64x5 FILLER_322_1654 ();
 b15zdnd11an1n32x5 FILLER_322_1718 ();
 b15zdnd11an1n16x5 FILLER_322_1750 ();
 b15zdnd11an1n08x5 FILLER_322_1766 ();
 b15zdnd11an1n64x5 FILLER_322_1777 ();
 b15zdnd11an1n64x5 FILLER_322_1841 ();
 b15zdnd11an1n04x5 FILLER_322_1905 ();
 b15zdnd00an1n02x5 FILLER_322_1909 ();
 b15zdnd11an1n64x5 FILLER_322_1914 ();
 b15zdnd11an1n64x5 FILLER_322_1978 ();
 b15zdnd11an1n64x5 FILLER_322_2042 ();
 b15zdnd11an1n32x5 FILLER_322_2106 ();
 b15zdnd11an1n16x5 FILLER_322_2138 ();
 b15zdnd11an1n64x5 FILLER_322_2162 ();
 b15zdnd11an1n32x5 FILLER_322_2226 ();
 b15zdnd11an1n16x5 FILLER_322_2258 ();
 b15zdnd00an1n02x5 FILLER_322_2274 ();
 b15zdnd11an1n32x5 FILLER_323_0 ();
 b15zdnd11an1n16x5 FILLER_323_32 ();
 b15zdnd11an1n08x5 FILLER_323_48 ();
 b15zdnd11an1n04x5 FILLER_323_56 ();
 b15zdnd00an1n01x5 FILLER_323_60 ();
 b15zdnd11an1n64x5 FILLER_323_115 ();
 b15zdnd11an1n64x5 FILLER_323_179 ();
 b15zdnd11an1n32x5 FILLER_323_243 ();
 b15zdnd11an1n16x5 FILLER_323_275 ();
 b15zdnd11an1n08x5 FILLER_323_291 ();
 b15zdnd00an1n02x5 FILLER_323_299 ();
 b15zdnd00an1n01x5 FILLER_323_301 ();
 b15zdnd11an1n64x5 FILLER_323_305 ();
 b15zdnd11an1n64x5 FILLER_323_369 ();
 b15zdnd11an1n64x5 FILLER_323_433 ();
 b15zdnd11an1n64x5 FILLER_323_497 ();
 b15zdnd11an1n04x5 FILLER_323_564 ();
 b15zdnd11an1n64x5 FILLER_323_620 ();
 b15zdnd11an1n32x5 FILLER_323_684 ();
 b15zdnd00an1n02x5 FILLER_323_716 ();
 b15zdnd11an1n64x5 FILLER_323_760 ();
 b15zdnd11an1n64x5 FILLER_323_824 ();
 b15zdnd11an1n64x5 FILLER_323_888 ();
 b15zdnd11an1n64x5 FILLER_323_952 ();
 b15zdnd11an1n64x5 FILLER_323_1016 ();
 b15zdnd11an1n64x5 FILLER_323_1080 ();
 b15zdnd11an1n64x5 FILLER_323_1144 ();
 b15zdnd11an1n08x5 FILLER_323_1208 ();
 b15zdnd11an1n64x5 FILLER_323_1268 ();
 b15zdnd11an1n64x5 FILLER_323_1332 ();
 b15zdnd11an1n64x5 FILLER_323_1396 ();
 b15zdnd11an1n64x5 FILLER_323_1460 ();
 b15zdnd11an1n64x5 FILLER_323_1524 ();
 b15zdnd11an1n64x5 FILLER_323_1588 ();
 b15zdnd11an1n64x5 FILLER_323_1652 ();
 b15zdnd11an1n32x5 FILLER_323_1716 ();
 b15zdnd11an1n16x5 FILLER_323_1748 ();
 b15zdnd11an1n04x5 FILLER_323_1764 ();
 b15zdnd00an1n01x5 FILLER_323_1768 ();
 b15zdnd11an1n04x5 FILLER_323_1772 ();
 b15zdnd11an1n64x5 FILLER_323_1779 ();
 b15zdnd11an1n64x5 FILLER_323_1843 ();
 b15zdnd11an1n64x5 FILLER_323_1907 ();
 b15zdnd11an1n64x5 FILLER_323_1971 ();
 b15zdnd11an1n64x5 FILLER_323_2035 ();
 b15zdnd11an1n64x5 FILLER_323_2099 ();
 b15zdnd11an1n64x5 FILLER_323_2163 ();
 b15zdnd11an1n32x5 FILLER_323_2227 ();
 b15zdnd11an1n16x5 FILLER_323_2259 ();
 b15zdnd11an1n08x5 FILLER_323_2275 ();
 b15zdnd00an1n01x5 FILLER_323_2283 ();
 b15zdnd11an1n64x5 FILLER_324_8 ();
 b15zdnd11an1n08x5 FILLER_324_72 ();
 b15zdnd11an1n04x5 FILLER_324_80 ();
 b15zdnd00an1n01x5 FILLER_324_84 ();
 b15zdnd11an1n64x5 FILLER_324_88 ();
 b15zdnd11an1n64x5 FILLER_324_152 ();
 b15zdnd11an1n64x5 FILLER_324_216 ();
 b15zdnd11an1n64x5 FILLER_324_280 ();
 b15zdnd11an1n64x5 FILLER_324_344 ();
 b15zdnd11an1n64x5 FILLER_324_408 ();
 b15zdnd11an1n64x5 FILLER_324_472 ();
 b15zdnd11an1n16x5 FILLER_324_536 ();
 b15zdnd00an1n02x5 FILLER_324_552 ();
 b15zdnd00an1n01x5 FILLER_324_554 ();
 b15zdnd11an1n08x5 FILLER_324_558 ();
 b15zdnd11an1n04x5 FILLER_324_569 ();
 b15zdnd00an1n02x5 FILLER_324_573 ();
 b15zdnd11an1n64x5 FILLER_324_627 ();
 b15zdnd11an1n16x5 FILLER_324_691 ();
 b15zdnd11an1n08x5 FILLER_324_707 ();
 b15zdnd00an1n02x5 FILLER_324_715 ();
 b15zdnd00an1n01x5 FILLER_324_717 ();
 b15zdnd11an1n64x5 FILLER_324_726 ();
 b15zdnd11an1n64x5 FILLER_324_790 ();
 b15zdnd11an1n64x5 FILLER_324_854 ();
 b15zdnd11an1n64x5 FILLER_324_918 ();
 b15zdnd11an1n64x5 FILLER_324_982 ();
 b15zdnd11an1n64x5 FILLER_324_1046 ();
 b15zdnd11an1n64x5 FILLER_324_1110 ();
 b15zdnd11an1n64x5 FILLER_324_1174 ();
 b15zdnd00an1n02x5 FILLER_324_1238 ();
 b15zdnd00an1n01x5 FILLER_324_1240 ();
 b15zdnd11an1n04x5 FILLER_324_1244 ();
 b15zdnd00an1n01x5 FILLER_324_1248 ();
 b15zdnd11an1n64x5 FILLER_324_1252 ();
 b15zdnd11an1n64x5 FILLER_324_1316 ();
 b15zdnd11an1n64x5 FILLER_324_1380 ();
 b15zdnd11an1n64x5 FILLER_324_1444 ();
 b15zdnd11an1n64x5 FILLER_324_1508 ();
 b15zdnd11an1n64x5 FILLER_324_1572 ();
 b15zdnd11an1n64x5 FILLER_324_1636 ();
 b15zdnd11an1n32x5 FILLER_324_1700 ();
 b15zdnd11an1n16x5 FILLER_324_1732 ();
 b15zdnd00an1n02x5 FILLER_324_1748 ();
 b15zdnd00an1n01x5 FILLER_324_1750 ();
 b15zdnd11an1n64x5 FILLER_324_1803 ();
 b15zdnd11an1n64x5 FILLER_324_1867 ();
 b15zdnd11an1n64x5 FILLER_324_1931 ();
 b15zdnd11an1n64x5 FILLER_324_1995 ();
 b15zdnd11an1n64x5 FILLER_324_2059 ();
 b15zdnd11an1n16x5 FILLER_324_2123 ();
 b15zdnd11an1n08x5 FILLER_324_2139 ();
 b15zdnd11an1n04x5 FILLER_324_2147 ();
 b15zdnd00an1n02x5 FILLER_324_2151 ();
 b15zdnd00an1n01x5 FILLER_324_2153 ();
 b15zdnd11an1n64x5 FILLER_324_2162 ();
 b15zdnd11an1n32x5 FILLER_324_2226 ();
 b15zdnd11an1n16x5 FILLER_324_2258 ();
 b15zdnd00an1n02x5 FILLER_324_2274 ();
 b15zdnd11an1n64x5 FILLER_325_0 ();
 b15zdnd11an1n16x5 FILLER_325_64 ();
 b15zdnd11an1n04x5 FILLER_325_80 ();
 b15zdnd00an1n02x5 FILLER_325_84 ();
 b15zdnd00an1n01x5 FILLER_325_86 ();
 b15zdnd11an1n64x5 FILLER_325_90 ();
 b15zdnd11an1n64x5 FILLER_325_154 ();
 b15zdnd11an1n64x5 FILLER_325_218 ();
 b15zdnd11an1n64x5 FILLER_325_282 ();
 b15zdnd11an1n64x5 FILLER_325_346 ();
 b15zdnd11an1n64x5 FILLER_325_410 ();
 b15zdnd11an1n64x5 FILLER_325_474 ();
 b15zdnd11an1n32x5 FILLER_325_538 ();
 b15zdnd11an1n04x5 FILLER_325_570 ();
 b15zdnd11an1n04x5 FILLER_325_577 ();
 b15zdnd11an1n04x5 FILLER_325_584 ();
 b15zdnd11an1n04x5 FILLER_325_597 ();
 b15zdnd00an1n01x5 FILLER_325_601 ();
 b15zdnd11an1n64x5 FILLER_325_605 ();
 b15zdnd11an1n64x5 FILLER_325_669 ();
 b15zdnd11an1n64x5 FILLER_325_733 ();
 b15zdnd11an1n64x5 FILLER_325_797 ();
 b15zdnd11an1n64x5 FILLER_325_861 ();
 b15zdnd11an1n64x5 FILLER_325_925 ();
 b15zdnd11an1n64x5 FILLER_325_989 ();
 b15zdnd11an1n64x5 FILLER_325_1053 ();
 b15zdnd11an1n64x5 FILLER_325_1117 ();
 b15zdnd11an1n64x5 FILLER_325_1181 ();
 b15zdnd00an1n01x5 FILLER_325_1245 ();
 b15zdnd11an1n04x5 FILLER_325_1249 ();
 b15zdnd11an1n04x5 FILLER_325_1256 ();
 b15zdnd11an1n64x5 FILLER_325_1263 ();
 b15zdnd11an1n64x5 FILLER_325_1327 ();
 b15zdnd11an1n64x5 FILLER_325_1391 ();
 b15zdnd11an1n64x5 FILLER_325_1455 ();
 b15zdnd11an1n64x5 FILLER_325_1519 ();
 b15zdnd11an1n64x5 FILLER_325_1583 ();
 b15zdnd11an1n64x5 FILLER_325_1647 ();
 b15zdnd11an1n64x5 FILLER_325_1711 ();
 b15zdnd00an1n02x5 FILLER_325_1775 ();
 b15zdnd11an1n64x5 FILLER_325_1804 ();
 b15zdnd11an1n64x5 FILLER_325_1868 ();
 b15zdnd11an1n64x5 FILLER_325_1932 ();
 b15zdnd11an1n64x5 FILLER_325_1996 ();
 b15zdnd11an1n64x5 FILLER_325_2060 ();
 b15zdnd11an1n64x5 FILLER_325_2124 ();
 b15zdnd11an1n64x5 FILLER_325_2188 ();
 b15zdnd11an1n32x5 FILLER_325_2252 ();
 b15zdnd11an1n64x5 FILLER_326_8 ();
 b15zdnd11an1n08x5 FILLER_326_72 ();
 b15zdnd00an1n02x5 FILLER_326_80 ();
 b15zdnd00an1n01x5 FILLER_326_82 ();
 b15zdnd11an1n64x5 FILLER_326_91 ();
 b15zdnd11an1n64x5 FILLER_326_155 ();
 b15zdnd11an1n64x5 FILLER_326_219 ();
 b15zdnd11an1n64x5 FILLER_326_283 ();
 b15zdnd11an1n64x5 FILLER_326_347 ();
 b15zdnd11an1n64x5 FILLER_326_411 ();
 b15zdnd11an1n64x5 FILLER_326_475 ();
 b15zdnd11an1n32x5 FILLER_326_539 ();
 b15zdnd11an1n08x5 FILLER_326_571 ();
 b15zdnd00an1n02x5 FILLER_326_579 ();
 b15zdnd11an1n04x5 FILLER_326_584 ();
 b15zdnd11an1n04x5 FILLER_326_591 ();
 b15zdnd11an1n04x5 FILLER_326_598 ();
 b15zdnd11an1n64x5 FILLER_326_605 ();
 b15zdnd11an1n32x5 FILLER_326_669 ();
 b15zdnd11an1n16x5 FILLER_326_701 ();
 b15zdnd00an1n01x5 FILLER_326_717 ();
 b15zdnd11an1n64x5 FILLER_326_726 ();
 b15zdnd11an1n64x5 FILLER_326_790 ();
 b15zdnd11an1n64x5 FILLER_326_854 ();
 b15zdnd11an1n64x5 FILLER_326_918 ();
 b15zdnd11an1n64x5 FILLER_326_982 ();
 b15zdnd11an1n16x5 FILLER_326_1046 ();
 b15zdnd11an1n08x5 FILLER_326_1062 ();
 b15zdnd00an1n01x5 FILLER_326_1070 ();
 b15zdnd11an1n64x5 FILLER_326_1080 ();
 b15zdnd11an1n64x5 FILLER_326_1144 ();
 b15zdnd11an1n16x5 FILLER_326_1208 ();
 b15zdnd11an1n04x5 FILLER_326_1224 ();
 b15zdnd11an1n64x5 FILLER_326_1280 ();
 b15zdnd11an1n64x5 FILLER_326_1344 ();
 b15zdnd11an1n64x5 FILLER_326_1408 ();
 b15zdnd11an1n64x5 FILLER_326_1472 ();
 b15zdnd11an1n08x5 FILLER_326_1536 ();
 b15zdnd11an1n64x5 FILLER_326_1553 ();
 b15zdnd11an1n64x5 FILLER_326_1617 ();
 b15zdnd11an1n64x5 FILLER_326_1681 ();
 b15zdnd11an1n32x5 FILLER_326_1745 ();
 b15zdnd11an1n64x5 FILLER_326_1780 ();
 b15zdnd11an1n04x5 FILLER_326_1844 ();
 b15zdnd00an1n01x5 FILLER_326_1848 ();
 b15zdnd11an1n64x5 FILLER_326_1858 ();
 b15zdnd11an1n64x5 FILLER_326_1922 ();
 b15zdnd11an1n32x5 FILLER_326_1986 ();
 b15zdnd11an1n16x5 FILLER_326_2018 ();
 b15zdnd11an1n04x5 FILLER_326_2034 ();
 b15zdnd00an1n01x5 FILLER_326_2038 ();
 b15zdnd11an1n64x5 FILLER_326_2059 ();
 b15zdnd11an1n16x5 FILLER_326_2123 ();
 b15zdnd11an1n08x5 FILLER_326_2139 ();
 b15zdnd11an1n04x5 FILLER_326_2147 ();
 b15zdnd00an1n02x5 FILLER_326_2151 ();
 b15zdnd00an1n01x5 FILLER_326_2153 ();
 b15zdnd11an1n64x5 FILLER_326_2162 ();
 b15zdnd11an1n32x5 FILLER_326_2226 ();
 b15zdnd11an1n16x5 FILLER_326_2258 ();
 b15zdnd00an1n02x5 FILLER_326_2274 ();
 b15zdnd11an1n64x5 FILLER_327_0 ();
 b15zdnd11an1n64x5 FILLER_327_64 ();
 b15zdnd11an1n64x5 FILLER_327_128 ();
 b15zdnd11an1n64x5 FILLER_327_192 ();
 b15zdnd11an1n64x5 FILLER_327_256 ();
 b15zdnd11an1n64x5 FILLER_327_320 ();
 b15zdnd11an1n64x5 FILLER_327_384 ();
 b15zdnd11an1n64x5 FILLER_327_448 ();
 b15zdnd11an1n64x5 FILLER_327_512 ();
 b15zdnd11an1n08x5 FILLER_327_576 ();
 b15zdnd11an1n04x5 FILLER_327_584 ();
 b15zdnd00an1n01x5 FILLER_327_588 ();
 b15zdnd11an1n64x5 FILLER_327_592 ();
 b15zdnd11an1n08x5 FILLER_327_656 ();
 b15zdnd11an1n04x5 FILLER_327_664 ();
 b15zdnd11an1n64x5 FILLER_327_676 ();
 b15zdnd11an1n64x5 FILLER_327_740 ();
 b15zdnd11an1n64x5 FILLER_327_804 ();
 b15zdnd11an1n64x5 FILLER_327_868 ();
 b15zdnd11an1n64x5 FILLER_327_932 ();
 b15zdnd11an1n64x5 FILLER_327_996 ();
 b15zdnd11an1n64x5 FILLER_327_1060 ();
 b15zdnd11an1n64x5 FILLER_327_1124 ();
 b15zdnd11an1n32x5 FILLER_327_1188 ();
 b15zdnd11an1n16x5 FILLER_327_1220 ();
 b15zdnd00an1n01x5 FILLER_327_1236 ();
 b15zdnd11an1n64x5 FILLER_327_1289 ();
 b15zdnd11an1n32x5 FILLER_327_1353 ();
 b15zdnd11an1n08x5 FILLER_327_1385 ();
 b15zdnd11an1n04x5 FILLER_327_1393 ();
 b15zdnd00an1n02x5 FILLER_327_1397 ();
 b15zdnd00an1n01x5 FILLER_327_1399 ();
 b15zdnd11an1n64x5 FILLER_327_1420 ();
 b15zdnd11an1n64x5 FILLER_327_1484 ();
 b15zdnd11an1n64x5 FILLER_327_1548 ();
 b15zdnd11an1n08x5 FILLER_327_1612 ();
 b15zdnd11an1n04x5 FILLER_327_1620 ();
 b15zdnd00an1n01x5 FILLER_327_1624 ();
 b15zdnd11an1n64x5 FILLER_327_1642 ();
 b15zdnd11an1n64x5 FILLER_327_1706 ();
 b15zdnd11an1n64x5 FILLER_327_1770 ();
 b15zdnd11an1n64x5 FILLER_327_1834 ();
 b15zdnd11an1n64x5 FILLER_327_1898 ();
 b15zdnd11an1n64x5 FILLER_327_1962 ();
 b15zdnd11an1n64x5 FILLER_327_2026 ();
 b15zdnd11an1n64x5 FILLER_327_2090 ();
 b15zdnd11an1n64x5 FILLER_327_2154 ();
 b15zdnd11an1n64x5 FILLER_327_2218 ();
 b15zdnd00an1n02x5 FILLER_327_2282 ();
 b15zdnd11an1n64x5 FILLER_328_8 ();
 b15zdnd11an1n64x5 FILLER_328_72 ();
 b15zdnd11an1n64x5 FILLER_328_136 ();
 b15zdnd11an1n64x5 FILLER_328_200 ();
 b15zdnd11an1n64x5 FILLER_328_264 ();
 b15zdnd11an1n64x5 FILLER_328_328 ();
 b15zdnd11an1n64x5 FILLER_328_392 ();
 b15zdnd11an1n64x5 FILLER_328_456 ();
 b15zdnd11an1n64x5 FILLER_328_520 ();
 b15zdnd11an1n64x5 FILLER_328_584 ();
 b15zdnd11an1n64x5 FILLER_328_648 ();
 b15zdnd11an1n04x5 FILLER_328_712 ();
 b15zdnd00an1n02x5 FILLER_328_716 ();
 b15zdnd00an1n02x5 FILLER_328_726 ();
 b15zdnd11an1n64x5 FILLER_328_770 ();
 b15zdnd11an1n64x5 FILLER_328_834 ();
 b15zdnd11an1n64x5 FILLER_328_898 ();
 b15zdnd11an1n64x5 FILLER_328_962 ();
 b15zdnd11an1n64x5 FILLER_328_1026 ();
 b15zdnd11an1n64x5 FILLER_328_1090 ();
 b15zdnd11an1n64x5 FILLER_328_1154 ();
 b15zdnd11an1n32x5 FILLER_328_1218 ();
 b15zdnd11an1n08x5 FILLER_328_1250 ();
 b15zdnd00an1n02x5 FILLER_328_1258 ();
 b15zdnd11an1n04x5 FILLER_328_1263 ();
 b15zdnd11an1n16x5 FILLER_328_1270 ();
 b15zdnd11an1n08x5 FILLER_328_1286 ();
 b15zdnd00an1n01x5 FILLER_328_1294 ();
 b15zdnd11an1n64x5 FILLER_328_1306 ();
 b15zdnd11an1n64x5 FILLER_328_1370 ();
 b15zdnd11an1n64x5 FILLER_328_1434 ();
 b15zdnd11an1n64x5 FILLER_328_1498 ();
 b15zdnd11an1n64x5 FILLER_328_1562 ();
 b15zdnd11an1n64x5 FILLER_328_1626 ();
 b15zdnd11an1n64x5 FILLER_328_1690 ();
 b15zdnd11an1n04x5 FILLER_328_1754 ();
 b15zdnd00an1n01x5 FILLER_328_1758 ();
 b15zdnd11an1n04x5 FILLER_328_1762 ();
 b15zdnd11an1n64x5 FILLER_328_1769 ();
 b15zdnd11an1n64x5 FILLER_328_1833 ();
 b15zdnd11an1n64x5 FILLER_328_1897 ();
 b15zdnd11an1n64x5 FILLER_328_1961 ();
 b15zdnd11an1n64x5 FILLER_328_2025 ();
 b15zdnd11an1n64x5 FILLER_328_2089 ();
 b15zdnd00an1n01x5 FILLER_328_2153 ();
 b15zdnd11an1n64x5 FILLER_328_2162 ();
 b15zdnd11an1n32x5 FILLER_328_2226 ();
 b15zdnd11an1n16x5 FILLER_328_2258 ();
 b15zdnd00an1n02x5 FILLER_328_2274 ();
 b15zdnd11an1n64x5 FILLER_329_0 ();
 b15zdnd11an1n64x5 FILLER_329_64 ();
 b15zdnd11an1n64x5 FILLER_329_128 ();
 b15zdnd11an1n64x5 FILLER_329_192 ();
 b15zdnd11an1n64x5 FILLER_329_256 ();
 b15zdnd11an1n64x5 FILLER_329_320 ();
 b15zdnd11an1n64x5 FILLER_329_384 ();
 b15zdnd11an1n64x5 FILLER_329_448 ();
 b15zdnd11an1n64x5 FILLER_329_512 ();
 b15zdnd11an1n64x5 FILLER_329_576 ();
 b15zdnd11an1n16x5 FILLER_329_640 ();
 b15zdnd11an1n08x5 FILLER_329_656 ();
 b15zdnd11an1n04x5 FILLER_329_664 ();
 b15zdnd00an1n02x5 FILLER_329_668 ();
 b15zdnd00an1n01x5 FILLER_329_670 ();
 b15zdnd11an1n64x5 FILLER_329_677 ();
 b15zdnd11an1n64x5 FILLER_329_741 ();
 b15zdnd11an1n64x5 FILLER_329_805 ();
 b15zdnd11an1n64x5 FILLER_329_869 ();
 b15zdnd11an1n64x5 FILLER_329_933 ();
 b15zdnd11an1n64x5 FILLER_329_997 ();
 b15zdnd11an1n64x5 FILLER_329_1061 ();
 b15zdnd11an1n64x5 FILLER_329_1125 ();
 b15zdnd11an1n64x5 FILLER_329_1189 ();
 b15zdnd11an1n08x5 FILLER_329_1253 ();
 b15zdnd00an1n02x5 FILLER_329_1261 ();
 b15zdnd11an1n64x5 FILLER_329_1274 ();
 b15zdnd11an1n64x5 FILLER_329_1338 ();
 b15zdnd11an1n64x5 FILLER_329_1402 ();
 b15zdnd11an1n32x5 FILLER_329_1466 ();
 b15zdnd11an1n16x5 FILLER_329_1498 ();
 b15zdnd11an1n08x5 FILLER_329_1514 ();
 b15zdnd11an1n64x5 FILLER_329_1536 ();
 b15zdnd11an1n64x5 FILLER_329_1600 ();
 b15zdnd11an1n64x5 FILLER_329_1664 ();
 b15zdnd11an1n08x5 FILLER_329_1728 ();
 b15zdnd11an1n04x5 FILLER_329_1736 ();
 b15zdnd00an1n01x5 FILLER_329_1740 ();
 b15zdnd11an1n64x5 FILLER_329_1793 ();
 b15zdnd11an1n32x5 FILLER_329_1857 ();
 b15zdnd11an1n08x5 FILLER_329_1889 ();
 b15zdnd11an1n04x5 FILLER_329_1897 ();
 b15zdnd00an1n02x5 FILLER_329_1901 ();
 b15zdnd11an1n04x5 FILLER_329_1906 ();
 b15zdnd11an1n64x5 FILLER_329_1913 ();
 b15zdnd11an1n64x5 FILLER_329_1977 ();
 b15zdnd11an1n64x5 FILLER_329_2041 ();
 b15zdnd11an1n64x5 FILLER_329_2105 ();
 b15zdnd11an1n64x5 FILLER_329_2169 ();
 b15zdnd11an1n32x5 FILLER_329_2233 ();
 b15zdnd11an1n16x5 FILLER_329_2265 ();
 b15zdnd00an1n02x5 FILLER_329_2281 ();
 b15zdnd00an1n01x5 FILLER_329_2283 ();
 b15zdnd11an1n64x5 FILLER_330_8 ();
 b15zdnd11an1n04x5 FILLER_330_72 ();
 b15zdnd00an1n02x5 FILLER_330_76 ();
 b15zdnd11an1n64x5 FILLER_330_81 ();
 b15zdnd11an1n64x5 FILLER_330_145 ();
 b15zdnd11an1n64x5 FILLER_330_209 ();
 b15zdnd11an1n64x5 FILLER_330_273 ();
 b15zdnd11an1n64x5 FILLER_330_337 ();
 b15zdnd11an1n64x5 FILLER_330_401 ();
 b15zdnd11an1n64x5 FILLER_330_465 ();
 b15zdnd11an1n64x5 FILLER_330_529 ();
 b15zdnd11an1n64x5 FILLER_330_593 ();
 b15zdnd11an1n32x5 FILLER_330_657 ();
 b15zdnd11an1n16x5 FILLER_330_689 ();
 b15zdnd11an1n08x5 FILLER_330_705 ();
 b15zdnd11an1n04x5 FILLER_330_713 ();
 b15zdnd00an1n01x5 FILLER_330_717 ();
 b15zdnd11an1n16x5 FILLER_330_726 ();
 b15zdnd11an1n08x5 FILLER_330_742 ();
 b15zdnd00an1n02x5 FILLER_330_750 ();
 b15zdnd11an1n64x5 FILLER_330_772 ();
 b15zdnd11an1n64x5 FILLER_330_836 ();
 b15zdnd11an1n64x5 FILLER_330_900 ();
 b15zdnd11an1n64x5 FILLER_330_964 ();
 b15zdnd11an1n64x5 FILLER_330_1028 ();
 b15zdnd11an1n64x5 FILLER_330_1092 ();
 b15zdnd11an1n64x5 FILLER_330_1156 ();
 b15zdnd11an1n64x5 FILLER_330_1220 ();
 b15zdnd11an1n64x5 FILLER_330_1284 ();
 b15zdnd11an1n64x5 FILLER_330_1348 ();
 b15zdnd11an1n64x5 FILLER_330_1412 ();
 b15zdnd11an1n16x5 FILLER_330_1476 ();
 b15zdnd00an1n01x5 FILLER_330_1492 ();
 b15zdnd11an1n16x5 FILLER_330_1545 ();
 b15zdnd11an1n08x5 FILLER_330_1561 ();
 b15zdnd00an1n02x5 FILLER_330_1569 ();
 b15zdnd11an1n04x5 FILLER_330_1580 ();
 b15zdnd11an1n64x5 FILLER_330_1593 ();
 b15zdnd11an1n64x5 FILLER_330_1657 ();
 b15zdnd11an1n32x5 FILLER_330_1721 ();
 b15zdnd11an1n08x5 FILLER_330_1753 ();
 b15zdnd11an1n04x5 FILLER_330_1761 ();
 b15zdnd00an1n02x5 FILLER_330_1765 ();
 b15zdnd11an1n32x5 FILLER_330_1770 ();
 b15zdnd11an1n16x5 FILLER_330_1802 ();
 b15zdnd00an1n02x5 FILLER_330_1818 ();
 b15zdnd00an1n01x5 FILLER_330_1820 ();
 b15zdnd11an1n32x5 FILLER_330_1830 ();
 b15zdnd11an1n16x5 FILLER_330_1862 ();
 b15zdnd11an1n04x5 FILLER_330_1878 ();
 b15zdnd00an1n02x5 FILLER_330_1882 ();
 b15zdnd00an1n01x5 FILLER_330_1884 ();
 b15zdnd11an1n64x5 FILLER_330_1937 ();
 b15zdnd11an1n64x5 FILLER_330_2001 ();
 b15zdnd11an1n64x5 FILLER_330_2065 ();
 b15zdnd11an1n16x5 FILLER_330_2129 ();
 b15zdnd11an1n08x5 FILLER_330_2145 ();
 b15zdnd00an1n01x5 FILLER_330_2153 ();
 b15zdnd11an1n64x5 FILLER_330_2162 ();
 b15zdnd11an1n32x5 FILLER_330_2226 ();
 b15zdnd11an1n16x5 FILLER_330_2258 ();
 b15zdnd00an1n02x5 FILLER_330_2274 ();
 b15zdnd11an1n64x5 FILLER_331_0 ();
 b15zdnd11an1n64x5 FILLER_331_64 ();
 b15zdnd11an1n32x5 FILLER_331_128 ();
 b15zdnd11an1n08x5 FILLER_331_160 ();
 b15zdnd11an1n04x5 FILLER_331_168 ();
 b15zdnd11an1n64x5 FILLER_331_175 ();
 b15zdnd11an1n64x5 FILLER_331_239 ();
 b15zdnd11an1n64x5 FILLER_331_303 ();
 b15zdnd11an1n64x5 FILLER_331_367 ();
 b15zdnd11an1n64x5 FILLER_331_431 ();
 b15zdnd11an1n64x5 FILLER_331_495 ();
 b15zdnd11an1n64x5 FILLER_331_559 ();
 b15zdnd11an1n64x5 FILLER_331_623 ();
 b15zdnd11an1n64x5 FILLER_331_687 ();
 b15zdnd11an1n64x5 FILLER_331_751 ();
 b15zdnd11an1n64x5 FILLER_331_815 ();
 b15zdnd11an1n64x5 FILLER_331_879 ();
 b15zdnd11an1n64x5 FILLER_331_943 ();
 b15zdnd11an1n64x5 FILLER_331_1007 ();
 b15zdnd11an1n64x5 FILLER_331_1071 ();
 b15zdnd11an1n64x5 FILLER_331_1135 ();
 b15zdnd11an1n64x5 FILLER_331_1199 ();
 b15zdnd11an1n64x5 FILLER_331_1263 ();
 b15zdnd11an1n64x5 FILLER_331_1327 ();
 b15zdnd11an1n64x5 FILLER_331_1391 ();
 b15zdnd11an1n32x5 FILLER_331_1455 ();
 b15zdnd11an1n16x5 FILLER_331_1487 ();
 b15zdnd11an1n08x5 FILLER_331_1503 ();
 b15zdnd11an1n04x5 FILLER_331_1511 ();
 b15zdnd00an1n01x5 FILLER_331_1515 ();
 b15zdnd11an1n64x5 FILLER_331_1519 ();
 b15zdnd11an1n64x5 FILLER_331_1583 ();
 b15zdnd11an1n64x5 FILLER_331_1647 ();
 b15zdnd11an1n64x5 FILLER_331_1711 ();
 b15zdnd11an1n16x5 FILLER_331_1775 ();
 b15zdnd11an1n04x5 FILLER_331_1791 ();
 b15zdnd00an1n02x5 FILLER_331_1795 ();
 b15zdnd11an1n64x5 FILLER_331_1839 ();
 b15zdnd11an1n04x5 FILLER_331_1903 ();
 b15zdnd00an1n02x5 FILLER_331_1907 ();
 b15zdnd00an1n01x5 FILLER_331_1909 ();
 b15zdnd11an1n64x5 FILLER_331_1913 ();
 b15zdnd11an1n64x5 FILLER_331_1977 ();
 b15zdnd11an1n64x5 FILLER_331_2041 ();
 b15zdnd11an1n64x5 FILLER_331_2105 ();
 b15zdnd11an1n64x5 FILLER_331_2169 ();
 b15zdnd11an1n32x5 FILLER_331_2233 ();
 b15zdnd11an1n16x5 FILLER_331_2265 ();
 b15zdnd00an1n02x5 FILLER_331_2281 ();
 b15zdnd00an1n01x5 FILLER_331_2283 ();
 b15zdnd11an1n64x5 FILLER_332_8 ();
 b15zdnd11an1n04x5 FILLER_332_72 ();
 b15zdnd00an1n02x5 FILLER_332_76 ();
 b15zdnd11an1n64x5 FILLER_332_81 ();
 b15zdnd11an1n64x5 FILLER_332_197 ();
 b15zdnd11an1n64x5 FILLER_332_261 ();
 b15zdnd11an1n64x5 FILLER_332_325 ();
 b15zdnd11an1n64x5 FILLER_332_389 ();
 b15zdnd11an1n64x5 FILLER_332_453 ();
 b15zdnd11an1n64x5 FILLER_332_517 ();
 b15zdnd11an1n64x5 FILLER_332_581 ();
 b15zdnd11an1n32x5 FILLER_332_645 ();
 b15zdnd11an1n16x5 FILLER_332_694 ();
 b15zdnd11an1n08x5 FILLER_332_710 ();
 b15zdnd11an1n32x5 FILLER_332_726 ();
 b15zdnd11an1n16x5 FILLER_332_758 ();
 b15zdnd11an1n04x5 FILLER_332_774 ();
 b15zdnd00an1n02x5 FILLER_332_778 ();
 b15zdnd11an1n64x5 FILLER_332_800 ();
 b15zdnd11an1n64x5 FILLER_332_864 ();
 b15zdnd11an1n64x5 FILLER_332_928 ();
 b15zdnd11an1n64x5 FILLER_332_992 ();
 b15zdnd11an1n16x5 FILLER_332_1056 ();
 b15zdnd11an1n04x5 FILLER_332_1072 ();
 b15zdnd00an1n02x5 FILLER_332_1076 ();
 b15zdnd00an1n01x5 FILLER_332_1078 ();
 b15zdnd11an1n64x5 FILLER_332_1088 ();
 b15zdnd11an1n64x5 FILLER_332_1152 ();
 b15zdnd11an1n64x5 FILLER_332_1216 ();
 b15zdnd11an1n64x5 FILLER_332_1280 ();
 b15zdnd11an1n64x5 FILLER_332_1344 ();
 b15zdnd11an1n64x5 FILLER_332_1408 ();
 b15zdnd11an1n32x5 FILLER_332_1472 ();
 b15zdnd11an1n08x5 FILLER_332_1504 ();
 b15zdnd11an1n04x5 FILLER_332_1512 ();
 b15zdnd11an1n04x5 FILLER_332_1519 ();
 b15zdnd11an1n64x5 FILLER_332_1526 ();
 b15zdnd11an1n64x5 FILLER_332_1590 ();
 b15zdnd11an1n64x5 FILLER_332_1654 ();
 b15zdnd11an1n64x5 FILLER_332_1718 ();
 b15zdnd11an1n64x5 FILLER_332_1782 ();
 b15zdnd11an1n64x5 FILLER_332_1855 ();
 b15zdnd11an1n64x5 FILLER_332_1919 ();
 b15zdnd11an1n64x5 FILLER_332_1983 ();
 b15zdnd11an1n64x5 FILLER_332_2047 ();
 b15zdnd11an1n32x5 FILLER_332_2111 ();
 b15zdnd11an1n08x5 FILLER_332_2143 ();
 b15zdnd00an1n02x5 FILLER_332_2151 ();
 b15zdnd00an1n01x5 FILLER_332_2153 ();
 b15zdnd11an1n64x5 FILLER_332_2162 ();
 b15zdnd11an1n32x5 FILLER_332_2226 ();
 b15zdnd11an1n16x5 FILLER_332_2258 ();
 b15zdnd00an1n02x5 FILLER_332_2274 ();
 b15zdnd11an1n64x5 FILLER_333_0 ();
 b15zdnd11an1n08x5 FILLER_333_64 ();
 b15zdnd00an1n02x5 FILLER_333_72 ();
 b15zdnd11an1n64x5 FILLER_333_78 ();
 b15zdnd11an1n16x5 FILLER_333_142 ();
 b15zdnd11an1n04x5 FILLER_333_158 ();
 b15zdnd00an1n01x5 FILLER_333_162 ();
 b15zdnd11an1n04x5 FILLER_333_166 ();
 b15zdnd11an1n64x5 FILLER_333_173 ();
 b15zdnd11an1n08x5 FILLER_333_237 ();
 b15zdnd11an1n64x5 FILLER_333_287 ();
 b15zdnd11an1n64x5 FILLER_333_351 ();
 b15zdnd11an1n64x5 FILLER_333_415 ();
 b15zdnd11an1n64x5 FILLER_333_479 ();
 b15zdnd11an1n64x5 FILLER_333_543 ();
 b15zdnd11an1n64x5 FILLER_333_607 ();
 b15zdnd11an1n16x5 FILLER_333_671 ();
 b15zdnd00an1n01x5 FILLER_333_687 ();
 b15zdnd11an1n64x5 FILLER_333_696 ();
 b15zdnd11an1n64x5 FILLER_333_760 ();
 b15zdnd11an1n64x5 FILLER_333_824 ();
 b15zdnd11an1n64x5 FILLER_333_888 ();
 b15zdnd11an1n64x5 FILLER_333_952 ();
 b15zdnd11an1n64x5 FILLER_333_1016 ();
 b15zdnd11an1n64x5 FILLER_333_1080 ();
 b15zdnd11an1n64x5 FILLER_333_1144 ();
 b15zdnd11an1n64x5 FILLER_333_1208 ();
 b15zdnd11an1n32x5 FILLER_333_1272 ();
 b15zdnd11an1n08x5 FILLER_333_1304 ();
 b15zdnd11an1n04x5 FILLER_333_1312 ();
 b15zdnd00an1n02x5 FILLER_333_1316 ();
 b15zdnd11an1n32x5 FILLER_333_1332 ();
 b15zdnd11an1n16x5 FILLER_333_1364 ();
 b15zdnd11an1n08x5 FILLER_333_1380 ();
 b15zdnd11an1n04x5 FILLER_333_1388 ();
 b15zdnd11an1n04x5 FILLER_333_1406 ();
 b15zdnd11an1n32x5 FILLER_333_1424 ();
 b15zdnd00an1n01x5 FILLER_333_1456 ();
 b15zdnd11an1n64x5 FILLER_333_1474 ();
 b15zdnd11an1n64x5 FILLER_333_1538 ();
 b15zdnd11an1n16x5 FILLER_333_1602 ();
 b15zdnd11an1n08x5 FILLER_333_1618 ();
 b15zdnd11an1n04x5 FILLER_333_1626 ();
 b15zdnd11an1n04x5 FILLER_333_1633 ();
 b15zdnd11an1n64x5 FILLER_333_1640 ();
 b15zdnd11an1n64x5 FILLER_333_1704 ();
 b15zdnd11an1n64x5 FILLER_333_1768 ();
 b15zdnd11an1n64x5 FILLER_333_1832 ();
 b15zdnd11an1n64x5 FILLER_333_1896 ();
 b15zdnd11an1n64x5 FILLER_333_1960 ();
 b15zdnd11an1n64x5 FILLER_333_2024 ();
 b15zdnd11an1n64x5 FILLER_333_2088 ();
 b15zdnd11an1n64x5 FILLER_333_2152 ();
 b15zdnd11an1n64x5 FILLER_333_2216 ();
 b15zdnd11an1n04x5 FILLER_333_2280 ();
 b15zdnd11an1n64x5 FILLER_334_8 ();
 b15zdnd11an1n32x5 FILLER_334_72 ();
 b15zdnd11an1n16x5 FILLER_334_104 ();
 b15zdnd11an1n08x5 FILLER_334_120 ();
 b15zdnd11an1n04x5 FILLER_334_128 ();
 b15zdnd11an1n64x5 FILLER_334_159 ();
 b15zdnd11an1n64x5 FILLER_334_223 ();
 b15zdnd11an1n64x5 FILLER_334_287 ();
 b15zdnd11an1n64x5 FILLER_334_351 ();
 b15zdnd11an1n64x5 FILLER_334_415 ();
 b15zdnd11an1n64x5 FILLER_334_479 ();
 b15zdnd11an1n64x5 FILLER_334_543 ();
 b15zdnd11an1n64x5 FILLER_334_607 ();
 b15zdnd11an1n08x5 FILLER_334_671 ();
 b15zdnd11an1n04x5 FILLER_334_679 ();
 b15zdnd11an1n16x5 FILLER_334_688 ();
 b15zdnd11an1n08x5 FILLER_334_704 ();
 b15zdnd11an1n04x5 FILLER_334_712 ();
 b15zdnd00an1n02x5 FILLER_334_716 ();
 b15zdnd11an1n64x5 FILLER_334_726 ();
 b15zdnd11an1n16x5 FILLER_334_790 ();
 b15zdnd11an1n64x5 FILLER_334_833 ();
 b15zdnd11an1n64x5 FILLER_334_897 ();
 b15zdnd11an1n64x5 FILLER_334_961 ();
 b15zdnd11an1n64x5 FILLER_334_1025 ();
 b15zdnd11an1n64x5 FILLER_334_1089 ();
 b15zdnd11an1n64x5 FILLER_334_1153 ();
 b15zdnd11an1n64x5 FILLER_334_1217 ();
 b15zdnd11an1n64x5 FILLER_334_1281 ();
 b15zdnd11an1n64x5 FILLER_334_1345 ();
 b15zdnd11an1n64x5 FILLER_334_1409 ();
 b15zdnd11an1n64x5 FILLER_334_1473 ();
 b15zdnd11an1n64x5 FILLER_334_1537 ();
 b15zdnd11an1n04x5 FILLER_334_1601 ();
 b15zdnd11an1n64x5 FILLER_334_1657 ();
 b15zdnd11an1n64x5 FILLER_334_1721 ();
 b15zdnd11an1n64x5 FILLER_334_1785 ();
 b15zdnd11an1n64x5 FILLER_334_1849 ();
 b15zdnd11an1n64x5 FILLER_334_1913 ();
 b15zdnd11an1n64x5 FILLER_334_1977 ();
 b15zdnd11an1n64x5 FILLER_334_2041 ();
 b15zdnd11an1n32x5 FILLER_334_2105 ();
 b15zdnd11an1n16x5 FILLER_334_2137 ();
 b15zdnd00an1n01x5 FILLER_334_2153 ();
 b15zdnd11an1n64x5 FILLER_334_2162 ();
 b15zdnd11an1n32x5 FILLER_334_2226 ();
 b15zdnd11an1n16x5 FILLER_334_2258 ();
 b15zdnd00an1n02x5 FILLER_334_2274 ();
 b15zdnd11an1n64x5 FILLER_335_0 ();
 b15zdnd11an1n08x5 FILLER_335_64 ();
 b15zdnd11an1n04x5 FILLER_335_72 ();
 b15zdnd11an1n32x5 FILLER_335_79 ();
 b15zdnd11an1n16x5 FILLER_335_111 ();
 b15zdnd11an1n04x5 FILLER_335_127 ();
 b15zdnd00an1n01x5 FILLER_335_131 ();
 b15zdnd11an1n04x5 FILLER_335_135 ();
 b15zdnd11an1n04x5 FILLER_335_167 ();
 b15zdnd11an1n64x5 FILLER_335_174 ();
 b15zdnd11an1n64x5 FILLER_335_238 ();
 b15zdnd11an1n64x5 FILLER_335_302 ();
 b15zdnd11an1n64x5 FILLER_335_366 ();
 b15zdnd11an1n64x5 FILLER_335_430 ();
 b15zdnd11an1n64x5 FILLER_335_494 ();
 b15zdnd11an1n64x5 FILLER_335_558 ();
 b15zdnd11an1n64x5 FILLER_335_622 ();
 b15zdnd11an1n64x5 FILLER_335_686 ();
 b15zdnd11an1n32x5 FILLER_335_750 ();
 b15zdnd11an1n16x5 FILLER_335_782 ();
 b15zdnd11an1n08x5 FILLER_335_798 ();
 b15zdnd00an1n02x5 FILLER_335_806 ();
 b15zdnd11an1n08x5 FILLER_335_811 ();
 b15zdnd00an1n02x5 FILLER_335_819 ();
 b15zdnd11an1n64x5 FILLER_335_830 ();
 b15zdnd11an1n64x5 FILLER_335_894 ();
 b15zdnd11an1n64x5 FILLER_335_958 ();
 b15zdnd11an1n32x5 FILLER_335_1022 ();
 b15zdnd11an1n16x5 FILLER_335_1054 ();
 b15zdnd00an1n01x5 FILLER_335_1070 ();
 b15zdnd11an1n64x5 FILLER_335_1080 ();
 b15zdnd11an1n64x5 FILLER_335_1144 ();
 b15zdnd11an1n64x5 FILLER_335_1208 ();
 b15zdnd11an1n64x5 FILLER_335_1272 ();
 b15zdnd11an1n64x5 FILLER_335_1336 ();
 b15zdnd11an1n64x5 FILLER_335_1400 ();
 b15zdnd11an1n08x5 FILLER_335_1464 ();
 b15zdnd11an1n04x5 FILLER_335_1472 ();
 b15zdnd00an1n02x5 FILLER_335_1476 ();
 b15zdnd11an1n64x5 FILLER_335_1498 ();
 b15zdnd11an1n64x5 FILLER_335_1562 ();
 b15zdnd11an1n04x5 FILLER_335_1626 ();
 b15zdnd11an1n64x5 FILLER_335_1633 ();
 b15zdnd11an1n64x5 FILLER_335_1697 ();
 b15zdnd11an1n64x5 FILLER_335_1761 ();
 b15zdnd11an1n64x5 FILLER_335_1825 ();
 b15zdnd11an1n64x5 FILLER_335_1889 ();
 b15zdnd11an1n64x5 FILLER_335_1953 ();
 b15zdnd11an1n64x5 FILLER_335_2017 ();
 b15zdnd11an1n64x5 FILLER_335_2081 ();
 b15zdnd11an1n64x5 FILLER_335_2145 ();
 b15zdnd11an1n64x5 FILLER_335_2209 ();
 b15zdnd11an1n08x5 FILLER_335_2273 ();
 b15zdnd00an1n02x5 FILLER_335_2281 ();
 b15zdnd00an1n01x5 FILLER_335_2283 ();
 b15zdnd11an1n32x5 FILLER_336_8 ();
 b15zdnd11an1n04x5 FILLER_336_40 ();
 b15zdnd00an1n02x5 FILLER_336_44 ();
 b15zdnd11an1n04x5 FILLER_336_72 ();
 b15zdnd11an1n64x5 FILLER_336_88 ();
 b15zdnd00an1n02x5 FILLER_336_152 ();
 b15zdnd00an1n01x5 FILLER_336_154 ();
 b15zdnd11an1n64x5 FILLER_336_164 ();
 b15zdnd11an1n64x5 FILLER_336_228 ();
 b15zdnd11an1n64x5 FILLER_336_292 ();
 b15zdnd11an1n64x5 FILLER_336_356 ();
 b15zdnd11an1n64x5 FILLER_336_420 ();
 b15zdnd11an1n64x5 FILLER_336_484 ();
 b15zdnd11an1n64x5 FILLER_336_548 ();
 b15zdnd11an1n64x5 FILLER_336_612 ();
 b15zdnd11an1n32x5 FILLER_336_676 ();
 b15zdnd11an1n08x5 FILLER_336_708 ();
 b15zdnd00an1n02x5 FILLER_336_716 ();
 b15zdnd11an1n64x5 FILLER_336_726 ();
 b15zdnd11an1n64x5 FILLER_336_790 ();
 b15zdnd11an1n64x5 FILLER_336_854 ();
 b15zdnd11an1n64x5 FILLER_336_918 ();
 b15zdnd11an1n64x5 FILLER_336_982 ();
 b15zdnd11an1n64x5 FILLER_336_1046 ();
 b15zdnd11an1n64x5 FILLER_336_1110 ();
 b15zdnd11an1n64x5 FILLER_336_1174 ();
 b15zdnd11an1n64x5 FILLER_336_1238 ();
 b15zdnd11an1n32x5 FILLER_336_1302 ();
 b15zdnd00an1n02x5 FILLER_336_1334 ();
 b15zdnd00an1n01x5 FILLER_336_1336 ();
 b15zdnd11an1n64x5 FILLER_336_1351 ();
 b15zdnd11an1n64x5 FILLER_336_1415 ();
 b15zdnd11an1n64x5 FILLER_336_1479 ();
 b15zdnd11an1n64x5 FILLER_336_1543 ();
 b15zdnd11an1n64x5 FILLER_336_1607 ();
 b15zdnd11an1n64x5 FILLER_336_1671 ();
 b15zdnd11an1n64x5 FILLER_336_1735 ();
 b15zdnd11an1n32x5 FILLER_336_1799 ();
 b15zdnd11an1n16x5 FILLER_336_1831 ();
 b15zdnd11an1n08x5 FILLER_336_1847 ();
 b15zdnd11an1n04x5 FILLER_336_1855 ();
 b15zdnd00an1n01x5 FILLER_336_1859 ();
 b15zdnd11an1n08x5 FILLER_336_1863 ();
 b15zdnd11an1n64x5 FILLER_336_1874 ();
 b15zdnd11an1n64x5 FILLER_336_1938 ();
 b15zdnd11an1n64x5 FILLER_336_2002 ();
 b15zdnd11an1n64x5 FILLER_336_2066 ();
 b15zdnd11an1n16x5 FILLER_336_2130 ();
 b15zdnd11an1n08x5 FILLER_336_2146 ();
 b15zdnd11an1n64x5 FILLER_336_2162 ();
 b15zdnd11an1n32x5 FILLER_336_2226 ();
 b15zdnd11an1n16x5 FILLER_336_2258 ();
 b15zdnd00an1n02x5 FILLER_336_2274 ();
 b15zdnd11an1n64x5 FILLER_337_0 ();
 b15zdnd11an1n08x5 FILLER_337_64 ();
 b15zdnd00an1n02x5 FILLER_337_72 ();
 b15zdnd00an1n01x5 FILLER_337_74 ();
 b15zdnd11an1n64x5 FILLER_337_87 ();
 b15zdnd11an1n04x5 FILLER_337_151 ();
 b15zdnd00an1n02x5 FILLER_337_155 ();
 b15zdnd11an1n64x5 FILLER_337_160 ();
 b15zdnd11an1n64x5 FILLER_337_224 ();
 b15zdnd11an1n64x5 FILLER_337_288 ();
 b15zdnd11an1n04x5 FILLER_337_352 ();
 b15zdnd00an1n02x5 FILLER_337_356 ();
 b15zdnd11an1n64x5 FILLER_337_370 ();
 b15zdnd11an1n64x5 FILLER_337_434 ();
 b15zdnd11an1n64x5 FILLER_337_498 ();
 b15zdnd11an1n64x5 FILLER_337_562 ();
 b15zdnd11an1n64x5 FILLER_337_626 ();
 b15zdnd11an1n64x5 FILLER_337_690 ();
 b15zdnd11an1n64x5 FILLER_337_754 ();
 b15zdnd11an1n64x5 FILLER_337_818 ();
 b15zdnd11an1n64x5 FILLER_337_882 ();
 b15zdnd11an1n64x5 FILLER_337_946 ();
 b15zdnd11an1n64x5 FILLER_337_1010 ();
 b15zdnd11an1n64x5 FILLER_337_1074 ();
 b15zdnd11an1n64x5 FILLER_337_1138 ();
 b15zdnd11an1n64x5 FILLER_337_1202 ();
 b15zdnd11an1n64x5 FILLER_337_1266 ();
 b15zdnd11an1n64x5 FILLER_337_1330 ();
 b15zdnd11an1n64x5 FILLER_337_1394 ();
 b15zdnd11an1n16x5 FILLER_337_1458 ();
 b15zdnd11an1n08x5 FILLER_337_1474 ();
 b15zdnd11an1n04x5 FILLER_337_1482 ();
 b15zdnd00an1n01x5 FILLER_337_1486 ();
 b15zdnd11an1n64x5 FILLER_337_1501 ();
 b15zdnd11an1n64x5 FILLER_337_1565 ();
 b15zdnd11an1n64x5 FILLER_337_1629 ();
 b15zdnd11an1n64x5 FILLER_337_1693 ();
 b15zdnd11an1n64x5 FILLER_337_1757 ();
 b15zdnd11an1n16x5 FILLER_337_1821 ();
 b15zdnd11an1n64x5 FILLER_337_1889 ();
 b15zdnd11an1n64x5 FILLER_337_1953 ();
 b15zdnd11an1n64x5 FILLER_337_2017 ();
 b15zdnd11an1n64x5 FILLER_337_2081 ();
 b15zdnd11an1n64x5 FILLER_337_2145 ();
 b15zdnd11an1n64x5 FILLER_337_2209 ();
 b15zdnd11an1n08x5 FILLER_337_2273 ();
 b15zdnd00an1n02x5 FILLER_337_2281 ();
 b15zdnd00an1n01x5 FILLER_337_2283 ();
 b15zdnd11an1n64x5 FILLER_338_8 ();
 b15zdnd11an1n64x5 FILLER_338_72 ();
 b15zdnd11an1n32x5 FILLER_338_136 ();
 b15zdnd11an1n04x5 FILLER_338_168 ();
 b15zdnd00an1n02x5 FILLER_338_172 ();
 b15zdnd00an1n01x5 FILLER_338_174 ();
 b15zdnd11an1n64x5 FILLER_338_178 ();
 b15zdnd11an1n64x5 FILLER_338_242 ();
 b15zdnd11an1n64x5 FILLER_338_306 ();
 b15zdnd11an1n64x5 FILLER_338_370 ();
 b15zdnd11an1n08x5 FILLER_338_434 ();
 b15zdnd00an1n02x5 FILLER_338_442 ();
 b15zdnd00an1n01x5 FILLER_338_444 ();
 b15zdnd11an1n64x5 FILLER_338_461 ();
 b15zdnd11an1n64x5 FILLER_338_525 ();
 b15zdnd11an1n64x5 FILLER_338_589 ();
 b15zdnd11an1n32x5 FILLER_338_653 ();
 b15zdnd11an1n16x5 FILLER_338_685 ();
 b15zdnd11an1n04x5 FILLER_338_701 ();
 b15zdnd00an1n02x5 FILLER_338_705 ();
 b15zdnd11an1n04x5 FILLER_338_711 ();
 b15zdnd00an1n02x5 FILLER_338_715 ();
 b15zdnd00an1n01x5 FILLER_338_717 ();
 b15zdnd11an1n64x5 FILLER_338_726 ();
 b15zdnd11an1n64x5 FILLER_338_790 ();
 b15zdnd11an1n64x5 FILLER_338_854 ();
 b15zdnd11an1n64x5 FILLER_338_918 ();
 b15zdnd11an1n32x5 FILLER_338_982 ();
 b15zdnd11an1n64x5 FILLER_338_1017 ();
 b15zdnd11an1n64x5 FILLER_338_1081 ();
 b15zdnd00an1n01x5 FILLER_338_1145 ();
 b15zdnd11an1n64x5 FILLER_338_1166 ();
 b15zdnd11an1n64x5 FILLER_338_1230 ();
 b15zdnd11an1n64x5 FILLER_338_1294 ();
 b15zdnd11an1n32x5 FILLER_338_1358 ();
 b15zdnd11an1n08x5 FILLER_338_1390 ();
 b15zdnd11an1n04x5 FILLER_338_1398 ();
 b15zdnd00an1n02x5 FILLER_338_1402 ();
 b15zdnd00an1n01x5 FILLER_338_1404 ();
 b15zdnd11an1n64x5 FILLER_338_1425 ();
 b15zdnd11an1n64x5 FILLER_338_1489 ();
 b15zdnd11an1n64x5 FILLER_338_1553 ();
 b15zdnd11an1n64x5 FILLER_338_1617 ();
 b15zdnd11an1n64x5 FILLER_338_1681 ();
 b15zdnd11an1n64x5 FILLER_338_1745 ();
 b15zdnd11an1n32x5 FILLER_338_1809 ();
 b15zdnd11an1n16x5 FILLER_338_1841 ();
 b15zdnd00an1n02x5 FILLER_338_1857 ();
 b15zdnd00an1n01x5 FILLER_338_1859 ();
 b15zdnd11an1n04x5 FILLER_338_1863 ();
 b15zdnd00an1n02x5 FILLER_338_1867 ();
 b15zdnd11an1n64x5 FILLER_338_1889 ();
 b15zdnd11an1n64x5 FILLER_338_1953 ();
 b15zdnd11an1n64x5 FILLER_338_2017 ();
 b15zdnd11an1n64x5 FILLER_338_2081 ();
 b15zdnd11an1n08x5 FILLER_338_2145 ();
 b15zdnd00an1n01x5 FILLER_338_2153 ();
 b15zdnd11an1n64x5 FILLER_338_2162 ();
 b15zdnd11an1n32x5 FILLER_338_2226 ();
 b15zdnd11an1n16x5 FILLER_338_2258 ();
 b15zdnd00an1n02x5 FILLER_338_2274 ();
 b15zdnd11an1n64x5 FILLER_339_0 ();
 b15zdnd11an1n64x5 FILLER_339_64 ();
 b15zdnd11an1n16x5 FILLER_339_128 ();
 b15zdnd11an1n04x5 FILLER_339_144 ();
 b15zdnd11an1n64x5 FILLER_339_200 ();
 b15zdnd11an1n64x5 FILLER_339_264 ();
 b15zdnd11an1n32x5 FILLER_339_328 ();
 b15zdnd11an1n08x5 FILLER_339_360 ();
 b15zdnd11an1n04x5 FILLER_339_368 ();
 b15zdnd00an1n01x5 FILLER_339_372 ();
 b15zdnd11an1n64x5 FILLER_339_397 ();
 b15zdnd11an1n64x5 FILLER_339_461 ();
 b15zdnd11an1n64x5 FILLER_339_525 ();
 b15zdnd11an1n64x5 FILLER_339_589 ();
 b15zdnd11an1n32x5 FILLER_339_653 ();
 b15zdnd00an1n01x5 FILLER_339_685 ();
 b15zdnd11an1n64x5 FILLER_339_697 ();
 b15zdnd11an1n64x5 FILLER_339_761 ();
 b15zdnd11an1n64x5 FILLER_339_825 ();
 b15zdnd11an1n64x5 FILLER_339_889 ();
 b15zdnd11an1n32x5 FILLER_339_953 ();
 b15zdnd11an1n16x5 FILLER_339_985 ();
 b15zdnd00an1n02x5 FILLER_339_1001 ();
 b15zdnd00an1n01x5 FILLER_339_1003 ();
 b15zdnd11an1n08x5 FILLER_339_1007 ();
 b15zdnd11an1n04x5 FILLER_339_1018 ();
 b15zdnd00an1n02x5 FILLER_339_1022 ();
 b15zdnd11an1n64x5 FILLER_339_1027 ();
 b15zdnd11an1n08x5 FILLER_339_1091 ();
 b15zdnd11an1n04x5 FILLER_339_1099 ();
 b15zdnd11an1n64x5 FILLER_339_1123 ();
 b15zdnd11an1n32x5 FILLER_339_1187 ();
 b15zdnd11an1n16x5 FILLER_339_1219 ();
 b15zdnd11an1n64x5 FILLER_339_1255 ();
 b15zdnd11an1n64x5 FILLER_339_1319 ();
 b15zdnd11an1n08x5 FILLER_339_1383 ();
 b15zdnd00an1n02x5 FILLER_339_1391 ();
 b15zdnd11an1n32x5 FILLER_339_1407 ();
 b15zdnd11an1n16x5 FILLER_339_1439 ();
 b15zdnd11an1n08x5 FILLER_339_1455 ();
 b15zdnd11an1n04x5 FILLER_339_1463 ();
 b15zdnd00an1n02x5 FILLER_339_1467 ();
 b15zdnd11an1n64x5 FILLER_339_1483 ();
 b15zdnd11an1n64x5 FILLER_339_1547 ();
 b15zdnd11an1n64x5 FILLER_339_1611 ();
 b15zdnd11an1n64x5 FILLER_339_1675 ();
 b15zdnd11an1n64x5 FILLER_339_1739 ();
 b15zdnd11an1n64x5 FILLER_339_1803 ();
 b15zdnd11an1n64x5 FILLER_339_1867 ();
 b15zdnd11an1n64x5 FILLER_339_1931 ();
 b15zdnd11an1n32x5 FILLER_339_1995 ();
 b15zdnd11an1n08x5 FILLER_339_2027 ();
 b15zdnd11an1n04x5 FILLER_339_2035 ();
 b15zdnd11an1n64x5 FILLER_339_2047 ();
 b15zdnd11an1n64x5 FILLER_339_2111 ();
 b15zdnd11an1n64x5 FILLER_339_2175 ();
 b15zdnd11an1n32x5 FILLER_339_2239 ();
 b15zdnd11an1n08x5 FILLER_339_2271 ();
 b15zdnd11an1n04x5 FILLER_339_2279 ();
 b15zdnd00an1n01x5 FILLER_339_2283 ();
 b15zdnd11an1n64x5 FILLER_340_8 ();
 b15zdnd11an1n32x5 FILLER_340_72 ();
 b15zdnd11an1n16x5 FILLER_340_104 ();
 b15zdnd11an1n04x5 FILLER_340_120 ();
 b15zdnd00an1n02x5 FILLER_340_124 ();
 b15zdnd00an1n01x5 FILLER_340_126 ();
 b15zdnd11an1n16x5 FILLER_340_136 ();
 b15zdnd11an1n04x5 FILLER_340_152 ();
 b15zdnd00an1n01x5 FILLER_340_156 ();
 b15zdnd11an1n04x5 FILLER_340_166 ();
 b15zdnd00an1n02x5 FILLER_340_170 ();
 b15zdnd00an1n01x5 FILLER_340_172 ();
 b15zdnd11an1n64x5 FILLER_340_176 ();
 b15zdnd11an1n64x5 FILLER_340_240 ();
 b15zdnd11an1n16x5 FILLER_340_304 ();
 b15zdnd11an1n04x5 FILLER_340_320 ();
 b15zdnd00an1n02x5 FILLER_340_324 ();
 b15zdnd11an1n32x5 FILLER_340_347 ();
 b15zdnd11an1n08x5 FILLER_340_379 ();
 b15zdnd11an1n04x5 FILLER_340_387 ();
 b15zdnd00an1n01x5 FILLER_340_391 ();
 b15zdnd11an1n64x5 FILLER_340_396 ();
 b15zdnd11an1n64x5 FILLER_340_460 ();
 b15zdnd11an1n64x5 FILLER_340_524 ();
 b15zdnd11an1n64x5 FILLER_340_588 ();
 b15zdnd11an1n64x5 FILLER_340_652 ();
 b15zdnd00an1n02x5 FILLER_340_716 ();
 b15zdnd11an1n64x5 FILLER_340_726 ();
 b15zdnd11an1n04x5 FILLER_340_790 ();
 b15zdnd00an1n02x5 FILLER_340_794 ();
 b15zdnd00an1n01x5 FILLER_340_796 ();
 b15zdnd11an1n64x5 FILLER_340_849 ();
 b15zdnd11an1n64x5 FILLER_340_913 ();
 b15zdnd11an1n16x5 FILLER_340_977 ();
 b15zdnd11an1n04x5 FILLER_340_993 ();
 b15zdnd00an1n02x5 FILLER_340_997 ();
 b15zdnd00an1n01x5 FILLER_340_999 ();
 b15zdnd11an1n64x5 FILLER_340_1052 ();
 b15zdnd11an1n04x5 FILLER_340_1116 ();
 b15zdnd00an1n02x5 FILLER_340_1120 ();
 b15zdnd11an1n04x5 FILLER_340_1125 ();
 b15zdnd11an1n64x5 FILLER_340_1132 ();
 b15zdnd11an1n64x5 FILLER_340_1196 ();
 b15zdnd11an1n64x5 FILLER_340_1260 ();
 b15zdnd11an1n08x5 FILLER_340_1324 ();
 b15zdnd11an1n04x5 FILLER_340_1332 ();
 b15zdnd00an1n02x5 FILLER_340_1336 ();
 b15zdnd11an1n64x5 FILLER_340_1358 ();
 b15zdnd11an1n16x5 FILLER_340_1422 ();
 b15zdnd11an1n08x5 FILLER_340_1438 ();
 b15zdnd11an1n04x5 FILLER_340_1446 ();
 b15zdnd11an1n64x5 FILLER_340_1470 ();
 b15zdnd11an1n64x5 FILLER_340_1534 ();
 b15zdnd11an1n64x5 FILLER_340_1598 ();
 b15zdnd11an1n64x5 FILLER_340_1662 ();
 b15zdnd11an1n64x5 FILLER_340_1726 ();
 b15zdnd11an1n08x5 FILLER_340_1790 ();
 b15zdnd00an1n01x5 FILLER_340_1798 ();
 b15zdnd11an1n64x5 FILLER_340_1802 ();
 b15zdnd11an1n64x5 FILLER_340_1866 ();
 b15zdnd11an1n64x5 FILLER_340_1930 ();
 b15zdnd11an1n64x5 FILLER_340_1994 ();
 b15zdnd11an1n64x5 FILLER_340_2058 ();
 b15zdnd11an1n32x5 FILLER_340_2122 ();
 b15zdnd11an1n64x5 FILLER_340_2162 ();
 b15zdnd11an1n32x5 FILLER_340_2226 ();
 b15zdnd11an1n16x5 FILLER_340_2258 ();
 b15zdnd00an1n02x5 FILLER_340_2274 ();
 b15zdnd11an1n64x5 FILLER_341_0 ();
 b15zdnd11an1n64x5 FILLER_341_64 ();
 b15zdnd11an1n32x5 FILLER_341_128 ();
 b15zdnd11an1n04x5 FILLER_341_160 ();
 b15zdnd00an1n02x5 FILLER_341_164 ();
 b15zdnd11an1n64x5 FILLER_341_169 ();
 b15zdnd11an1n64x5 FILLER_341_233 ();
 b15zdnd11an1n08x5 FILLER_341_297 ();
 b15zdnd11an1n04x5 FILLER_341_305 ();
 b15zdnd11an1n32x5 FILLER_341_333 ();
 b15zdnd11an1n08x5 FILLER_341_365 ();
 b15zdnd11an1n04x5 FILLER_341_373 ();
 b15zdnd00an1n01x5 FILLER_341_377 ();
 b15zdnd11an1n04x5 FILLER_341_383 ();
 b15zdnd00an1n01x5 FILLER_341_387 ();
 b15zdnd11an1n04x5 FILLER_341_394 ();
 b15zdnd00an1n01x5 FILLER_341_398 ();
 b15zdnd11an1n04x5 FILLER_341_415 ();
 b15zdnd00an1n01x5 FILLER_341_419 ();
 b15zdnd11an1n04x5 FILLER_341_439 ();
 b15zdnd00an1n02x5 FILLER_341_443 ();
 b15zdnd11an1n04x5 FILLER_341_451 ();
 b15zdnd00an1n02x5 FILLER_341_455 ();
 b15zdnd11an1n64x5 FILLER_341_481 ();
 b15zdnd11an1n08x5 FILLER_341_545 ();
 b15zdnd11an1n04x5 FILLER_341_553 ();
 b15zdnd00an1n02x5 FILLER_341_557 ();
 b15zdnd11an1n04x5 FILLER_341_574 ();
 b15zdnd00an1n02x5 FILLER_341_578 ();
 b15zdnd11an1n32x5 FILLER_341_611 ();
 b15zdnd11an1n16x5 FILLER_341_643 ();
 b15zdnd11an1n08x5 FILLER_341_659 ();
 b15zdnd00an1n02x5 FILLER_341_667 ();
 b15zdnd00an1n01x5 FILLER_341_669 ();
 b15zdnd11an1n04x5 FILLER_341_684 ();
 b15zdnd11an1n08x5 FILLER_341_695 ();
 b15zdnd00an1n02x5 FILLER_341_703 ();
 b15zdnd11an1n64x5 FILLER_341_709 ();
 b15zdnd11an1n32x5 FILLER_341_773 ();
 b15zdnd00an1n01x5 FILLER_341_805 ();
 b15zdnd11an1n64x5 FILLER_341_858 ();
 b15zdnd11an1n64x5 FILLER_341_922 ();
 b15zdnd11an1n04x5 FILLER_341_986 ();
 b15zdnd00an1n01x5 FILLER_341_990 ();
 b15zdnd11an1n32x5 FILLER_341_1043 ();
 b15zdnd11an1n16x5 FILLER_341_1075 ();
 b15zdnd11an1n08x5 FILLER_341_1091 ();
 b15zdnd00an1n02x5 FILLER_341_1099 ();
 b15zdnd11an1n64x5 FILLER_341_1153 ();
 b15zdnd11an1n64x5 FILLER_341_1217 ();
 b15zdnd11an1n32x5 FILLER_341_1281 ();
 b15zdnd11an1n16x5 FILLER_341_1313 ();
 b15zdnd11an1n04x5 FILLER_341_1329 ();
 b15zdnd11an1n64x5 FILLER_341_1345 ();
 b15zdnd11an1n64x5 FILLER_341_1409 ();
 b15zdnd11an1n32x5 FILLER_341_1473 ();
 b15zdnd00an1n02x5 FILLER_341_1505 ();
 b15zdnd11an1n32x5 FILLER_341_1510 ();
 b15zdnd11an1n16x5 FILLER_341_1542 ();
 b15zdnd11an1n04x5 FILLER_341_1558 ();
 b15zdnd00an1n01x5 FILLER_341_1562 ();
 b15zdnd11an1n64x5 FILLER_341_1583 ();
 b15zdnd11an1n64x5 FILLER_341_1647 ();
 b15zdnd11an1n64x5 FILLER_341_1711 ();
 b15zdnd11an1n16x5 FILLER_341_1775 ();
 b15zdnd00an1n02x5 FILLER_341_1791 ();
 b15zdnd11an1n04x5 FILLER_341_1796 ();
 b15zdnd11an1n04x5 FILLER_341_1803 ();
 b15zdnd11an1n32x5 FILLER_341_1810 ();
 b15zdnd11an1n16x5 FILLER_341_1842 ();
 b15zdnd11an1n08x5 FILLER_341_1858 ();
 b15zdnd00an1n01x5 FILLER_341_1866 ();
 b15zdnd11an1n64x5 FILLER_341_1887 ();
 b15zdnd11an1n64x5 FILLER_341_1951 ();
 b15zdnd11an1n64x5 FILLER_341_2015 ();
 b15zdnd11an1n64x5 FILLER_341_2079 ();
 b15zdnd11an1n64x5 FILLER_341_2143 ();
 b15zdnd11an1n64x5 FILLER_341_2207 ();
 b15zdnd11an1n08x5 FILLER_341_2271 ();
 b15zdnd11an1n04x5 FILLER_341_2279 ();
 b15zdnd00an1n01x5 FILLER_341_2283 ();
 b15zdnd11an1n64x5 FILLER_342_8 ();
 b15zdnd11an1n64x5 FILLER_342_72 ();
 b15zdnd11an1n64x5 FILLER_342_136 ();
 b15zdnd11an1n64x5 FILLER_342_200 ();
 b15zdnd11an1n16x5 FILLER_342_264 ();
 b15zdnd11an1n08x5 FILLER_342_280 ();
 b15zdnd00an1n01x5 FILLER_342_288 ();
 b15zdnd11an1n32x5 FILLER_342_292 ();
 b15zdnd00an1n01x5 FILLER_342_324 ();
 b15zdnd11an1n04x5 FILLER_342_333 ();
 b15zdnd11an1n32x5 FILLER_342_343 ();
 b15zdnd11an1n08x5 FILLER_342_375 ();
 b15zdnd00an1n01x5 FILLER_342_383 ();
 b15zdnd11an1n04x5 FILLER_342_395 ();
 b15zdnd11an1n04x5 FILLER_342_405 ();
 b15zdnd11an1n08x5 FILLER_342_429 ();
 b15zdnd11an1n04x5 FILLER_342_437 ();
 b15zdnd11an1n32x5 FILLER_342_452 ();
 b15zdnd11an1n08x5 FILLER_342_484 ();
 b15zdnd00an1n02x5 FILLER_342_492 ();
 b15zdnd00an1n01x5 FILLER_342_494 ();
 b15zdnd11an1n16x5 FILLER_342_505 ();
 b15zdnd11an1n64x5 FILLER_342_531 ();
 b15zdnd11an1n64x5 FILLER_342_595 ();
 b15zdnd11an1n32x5 FILLER_342_659 ();
 b15zdnd11an1n16x5 FILLER_342_691 ();
 b15zdnd11an1n08x5 FILLER_342_707 ();
 b15zdnd00an1n02x5 FILLER_342_715 ();
 b15zdnd00an1n01x5 FILLER_342_717 ();
 b15zdnd11an1n64x5 FILLER_342_726 ();
 b15zdnd11an1n08x5 FILLER_342_790 ();
 b15zdnd00an1n02x5 FILLER_342_798 ();
 b15zdnd00an1n01x5 FILLER_342_800 ();
 b15zdnd11an1n04x5 FILLER_342_804 ();
 b15zdnd11an1n04x5 FILLER_342_811 ();
 b15zdnd11an1n04x5 FILLER_342_818 ();
 b15zdnd11an1n04x5 FILLER_342_825 ();
 b15zdnd11an1n08x5 FILLER_342_838 ();
 b15zdnd00an1n01x5 FILLER_342_846 ();
 b15zdnd11an1n04x5 FILLER_342_850 ();
 b15zdnd11an1n64x5 FILLER_342_857 ();
 b15zdnd11an1n32x5 FILLER_342_921 ();
 b15zdnd11an1n08x5 FILLER_342_953 ();
 b15zdnd11an1n04x5 FILLER_342_961 ();
 b15zdnd00an1n02x5 FILLER_342_965 ();
 b15zdnd11an1n04x5 FILLER_342_1012 ();
 b15zdnd00an1n02x5 FILLER_342_1016 ();
 b15zdnd11an1n04x5 FILLER_342_1021 ();
 b15zdnd11an1n16x5 FILLER_342_1028 ();
 b15zdnd11an1n04x5 FILLER_342_1044 ();
 b15zdnd00an1n01x5 FILLER_342_1048 ();
 b15zdnd11an1n32x5 FILLER_342_1052 ();
 b15zdnd11an1n16x5 FILLER_342_1084 ();
 b15zdnd11an1n08x5 FILLER_342_1100 ();
 b15zdnd11an1n04x5 FILLER_342_1108 ();
 b15zdnd11an1n04x5 FILLER_342_1115 ();
 b15zdnd00an1n01x5 FILLER_342_1119 ();
 b15zdnd11an1n04x5 FILLER_342_1123 ();
 b15zdnd11an1n04x5 FILLER_342_1147 ();
 b15zdnd11an1n32x5 FILLER_342_1175 ();
 b15zdnd11an1n16x5 FILLER_342_1207 ();
 b15zdnd11an1n08x5 FILLER_342_1223 ();
 b15zdnd11an1n16x5 FILLER_342_1245 ();
 b15zdnd00an1n02x5 FILLER_342_1261 ();
 b15zdnd00an1n01x5 FILLER_342_1263 ();
 b15zdnd11an1n16x5 FILLER_342_1276 ();
 b15zdnd11an1n08x5 FILLER_342_1292 ();
 b15zdnd11an1n64x5 FILLER_342_1314 ();
 b15zdnd11an1n64x5 FILLER_342_1378 ();
 b15zdnd11an1n64x5 FILLER_342_1442 ();
 b15zdnd00an1n02x5 FILLER_342_1506 ();
 b15zdnd11an1n64x5 FILLER_342_1511 ();
 b15zdnd11an1n32x5 FILLER_342_1575 ();
 b15zdnd11an1n08x5 FILLER_342_1607 ();
 b15zdnd00an1n02x5 FILLER_342_1615 ();
 b15zdnd11an1n04x5 FILLER_342_1620 ();
 b15zdnd11an1n64x5 FILLER_342_1627 ();
 b15zdnd11an1n64x5 FILLER_342_1691 ();
 b15zdnd11an1n16x5 FILLER_342_1755 ();
 b15zdnd11an1n08x5 FILLER_342_1771 ();
 b15zdnd11an1n32x5 FILLER_342_1831 ();
 b15zdnd11an1n04x5 FILLER_342_1863 ();
 b15zdnd00an1n01x5 FILLER_342_1867 ();
 b15zdnd11an1n64x5 FILLER_342_1882 ();
 b15zdnd11an1n64x5 FILLER_342_1946 ();
 b15zdnd11an1n64x5 FILLER_342_2010 ();
 b15zdnd11an1n64x5 FILLER_342_2074 ();
 b15zdnd11an1n16x5 FILLER_342_2138 ();
 b15zdnd11an1n64x5 FILLER_342_2162 ();
 b15zdnd11an1n32x5 FILLER_342_2226 ();
 b15zdnd11an1n16x5 FILLER_342_2258 ();
 b15zdnd00an1n02x5 FILLER_342_2274 ();
 b15zdnd11an1n64x5 FILLER_343_0 ();
 b15zdnd11an1n64x5 FILLER_343_64 ();
 b15zdnd11an1n64x5 FILLER_343_128 ();
 b15zdnd11an1n64x5 FILLER_343_192 ();
 b15zdnd11an1n32x5 FILLER_343_256 ();
 b15zdnd11an1n16x5 FILLER_343_300 ();
 b15zdnd00an1n02x5 FILLER_343_316 ();
 b15zdnd11an1n08x5 FILLER_343_322 ();
 b15zdnd11an1n04x5 FILLER_343_330 ();
 b15zdnd00an1n02x5 FILLER_343_334 ();
 b15zdnd11an1n16x5 FILLER_343_355 ();
 b15zdnd11an1n08x5 FILLER_343_371 ();
 b15zdnd00an1n01x5 FILLER_343_379 ();
 b15zdnd11an1n08x5 FILLER_343_391 ();
 b15zdnd00an1n01x5 FILLER_343_399 ();
 b15zdnd11an1n32x5 FILLER_343_419 ();
 b15zdnd11an1n08x5 FILLER_343_451 ();
 b15zdnd11an1n04x5 FILLER_343_459 ();
 b15zdnd00an1n02x5 FILLER_343_463 ();
 b15zdnd11an1n64x5 FILLER_343_468 ();
 b15zdnd11an1n16x5 FILLER_343_532 ();
 b15zdnd11an1n08x5 FILLER_343_548 ();
 b15zdnd00an1n01x5 FILLER_343_556 ();
 b15zdnd11an1n04x5 FILLER_343_562 ();
 b15zdnd00an1n02x5 FILLER_343_566 ();
 b15zdnd00an1n01x5 FILLER_343_568 ();
 b15zdnd11an1n04x5 FILLER_343_588 ();
 b15zdnd00an1n01x5 FILLER_343_592 ();
 b15zdnd11an1n64x5 FILLER_343_605 ();
 b15zdnd11an1n08x5 FILLER_343_669 ();
 b15zdnd11an1n04x5 FILLER_343_677 ();
 b15zdnd00an1n02x5 FILLER_343_681 ();
 b15zdnd00an1n01x5 FILLER_343_683 ();
 b15zdnd11an1n64x5 FILLER_343_695 ();
 b15zdnd11an1n32x5 FILLER_343_759 ();
 b15zdnd11an1n04x5 FILLER_343_791 ();
 b15zdnd00an1n02x5 FILLER_343_795 ();
 b15zdnd00an1n01x5 FILLER_343_797 ();
 b15zdnd11an1n64x5 FILLER_343_850 ();
 b15zdnd11an1n64x5 FILLER_343_914 ();
 b15zdnd11an1n32x5 FILLER_343_978 ();
 b15zdnd11an1n08x5 FILLER_343_1010 ();
 b15zdnd11an1n04x5 FILLER_343_1018 ();
 b15zdnd11an1n08x5 FILLER_343_1074 ();
 b15zdnd11an1n04x5 FILLER_343_1082 ();
 b15zdnd00an1n01x5 FILLER_343_1086 ();
 b15zdnd11an1n16x5 FILLER_343_1139 ();
 b15zdnd11an1n04x5 FILLER_343_1155 ();
 b15zdnd00an1n02x5 FILLER_343_1159 ();
 b15zdnd11an1n32x5 FILLER_343_1181 ();
 b15zdnd11an1n08x5 FILLER_343_1213 ();
 b15zdnd00an1n01x5 FILLER_343_1221 ();
 b15zdnd11an1n64x5 FILLER_343_1236 ();
 b15zdnd00an1n02x5 FILLER_343_1300 ();
 b15zdnd11an1n32x5 FILLER_343_1322 ();
 b15zdnd11an1n08x5 FILLER_343_1354 ();
 b15zdnd11an1n32x5 FILLER_343_1374 ();
 b15zdnd00an1n01x5 FILLER_343_1406 ();
 b15zdnd11an1n32x5 FILLER_343_1424 ();
 b15zdnd00an1n02x5 FILLER_343_1456 ();
 b15zdnd11an1n04x5 FILLER_343_1478 ();
 b15zdnd00an1n01x5 FILLER_343_1482 ();
 b15zdnd11an1n64x5 FILLER_343_1535 ();
 b15zdnd11an1n04x5 FILLER_343_1651 ();
 b15zdnd00an1n02x5 FILLER_343_1655 ();
 b15zdnd11an1n64x5 FILLER_343_1681 ();
 b15zdnd11an1n16x5 FILLER_343_1745 ();
 b15zdnd11an1n04x5 FILLER_343_1761 ();
 b15zdnd00an1n01x5 FILLER_343_1765 ();
 b15zdnd11an1n64x5 FILLER_343_1818 ();
 b15zdnd11an1n64x5 FILLER_343_1882 ();
 b15zdnd11an1n64x5 FILLER_343_1946 ();
 b15zdnd11an1n64x5 FILLER_343_2010 ();
 b15zdnd11an1n64x5 FILLER_343_2074 ();
 b15zdnd11an1n64x5 FILLER_343_2138 ();
 b15zdnd11an1n64x5 FILLER_343_2202 ();
 b15zdnd11an1n16x5 FILLER_343_2266 ();
 b15zdnd00an1n02x5 FILLER_343_2282 ();
 b15zdnd11an1n64x5 FILLER_344_8 ();
 b15zdnd11an1n64x5 FILLER_344_72 ();
 b15zdnd11an1n64x5 FILLER_344_136 ();
 b15zdnd11an1n64x5 FILLER_344_200 ();
 b15zdnd11an1n64x5 FILLER_344_264 ();
 b15zdnd11an1n64x5 FILLER_344_328 ();
 b15zdnd11an1n08x5 FILLER_344_392 ();
 b15zdnd11an1n04x5 FILLER_344_400 ();
 b15zdnd11an1n64x5 FILLER_344_420 ();
 b15zdnd11an1n64x5 FILLER_344_484 ();
 b15zdnd11an1n32x5 FILLER_344_548 ();
 b15zdnd11an1n16x5 FILLER_344_580 ();
 b15zdnd11an1n08x5 FILLER_344_596 ();
 b15zdnd00an1n02x5 FILLER_344_604 ();
 b15zdnd00an1n01x5 FILLER_344_606 ();
 b15zdnd11an1n16x5 FILLER_344_613 ();
 b15zdnd11an1n08x5 FILLER_344_629 ();
 b15zdnd00an1n02x5 FILLER_344_637 ();
 b15zdnd11an1n32x5 FILLER_344_651 ();
 b15zdnd00an1n01x5 FILLER_344_683 ();
 b15zdnd11an1n16x5 FILLER_344_698 ();
 b15zdnd11an1n04x5 FILLER_344_714 ();
 b15zdnd11an1n64x5 FILLER_344_726 ();
 b15zdnd11an1n08x5 FILLER_344_790 ();
 b15zdnd00an1n01x5 FILLER_344_798 ();
 b15zdnd11an1n64x5 FILLER_344_851 ();
 b15zdnd11an1n64x5 FILLER_344_915 ();
 b15zdnd11an1n32x5 FILLER_344_979 ();
 b15zdnd11an1n16x5 FILLER_344_1011 ();
 b15zdnd11an1n08x5 FILLER_344_1027 ();
 b15zdnd11an1n04x5 FILLER_344_1035 ();
 b15zdnd00an1n01x5 FILLER_344_1039 ();
 b15zdnd11an1n04x5 FILLER_344_1043 ();
 b15zdnd11an1n32x5 FILLER_344_1050 ();
 b15zdnd11an1n16x5 FILLER_344_1082 ();
 b15zdnd11an1n08x5 FILLER_344_1098 ();
 b15zdnd00an1n01x5 FILLER_344_1106 ();
 b15zdnd11an1n04x5 FILLER_344_1110 ();
 b15zdnd11an1n16x5 FILLER_344_1117 ();
 b15zdnd11an1n04x5 FILLER_344_1157 ();
 b15zdnd11an1n64x5 FILLER_344_1175 ();
 b15zdnd11an1n64x5 FILLER_344_1239 ();
 b15zdnd11an1n32x5 FILLER_344_1303 ();
 b15zdnd11an1n16x5 FILLER_344_1335 ();
 b15zdnd11an1n08x5 FILLER_344_1351 ();
 b15zdnd11an1n04x5 FILLER_344_1359 ();
 b15zdnd00an1n01x5 FILLER_344_1363 ();
 b15zdnd11an1n32x5 FILLER_344_1370 ();
 b15zdnd11an1n16x5 FILLER_344_1402 ();
 b15zdnd11an1n04x5 FILLER_344_1418 ();
 b15zdnd00an1n02x5 FILLER_344_1422 ();
 b15zdnd11an1n04x5 FILLER_344_1444 ();
 b15zdnd11an1n32x5 FILLER_344_1460 ();
 b15zdnd11an1n16x5 FILLER_344_1492 ();
 b15zdnd00an1n01x5 FILLER_344_1508 ();
 b15zdnd11an1n64x5 FILLER_344_1512 ();
 b15zdnd11an1n04x5 FILLER_344_1576 ();
 b15zdnd00an1n02x5 FILLER_344_1580 ();
 b15zdnd00an1n01x5 FILLER_344_1582 ();
 b15zdnd11an1n04x5 FILLER_344_1635 ();
 b15zdnd11an1n04x5 FILLER_344_1659 ();
 b15zdnd11an1n64x5 FILLER_344_1683 ();
 b15zdnd11an1n32x5 FILLER_344_1747 ();
 b15zdnd11an1n04x5 FILLER_344_1779 ();
 b15zdnd00an1n01x5 FILLER_344_1783 ();
 b15zdnd11an1n04x5 FILLER_344_1787 ();
 b15zdnd11an1n64x5 FILLER_344_1794 ();
 b15zdnd11an1n64x5 FILLER_344_1858 ();
 b15zdnd11an1n64x5 FILLER_344_1922 ();
 b15zdnd11an1n64x5 FILLER_344_1986 ();
 b15zdnd11an1n64x5 FILLER_344_2050 ();
 b15zdnd11an1n32x5 FILLER_344_2114 ();
 b15zdnd11an1n08x5 FILLER_344_2146 ();
 b15zdnd11an1n64x5 FILLER_344_2162 ();
 b15zdnd11an1n32x5 FILLER_344_2226 ();
 b15zdnd11an1n16x5 FILLER_344_2258 ();
 b15zdnd00an1n02x5 FILLER_344_2274 ();
 b15zdnd11an1n64x5 FILLER_345_0 ();
 b15zdnd11an1n64x5 FILLER_345_64 ();
 b15zdnd11an1n16x5 FILLER_345_128 ();
 b15zdnd11an1n04x5 FILLER_345_144 ();
 b15zdnd00an1n02x5 FILLER_345_148 ();
 b15zdnd11an1n64x5 FILLER_345_153 ();
 b15zdnd11an1n64x5 FILLER_345_217 ();
 b15zdnd11an1n64x5 FILLER_345_281 ();
 b15zdnd11an1n32x5 FILLER_345_345 ();
 b15zdnd11an1n16x5 FILLER_345_377 ();
 b15zdnd11an1n08x5 FILLER_345_393 ();
 b15zdnd11an1n04x5 FILLER_345_401 ();
 b15zdnd00an1n02x5 FILLER_345_405 ();
 b15zdnd00an1n01x5 FILLER_345_407 ();
 b15zdnd11an1n64x5 FILLER_345_424 ();
 b15zdnd11an1n08x5 FILLER_345_488 ();
 b15zdnd11an1n08x5 FILLER_345_506 ();
 b15zdnd11an1n04x5 FILLER_345_514 ();
 b15zdnd00an1n02x5 FILLER_345_518 ();
 b15zdnd11an1n04x5 FILLER_345_534 ();
 b15zdnd11an1n32x5 FILLER_345_552 ();
 b15zdnd11an1n08x5 FILLER_345_584 ();
 b15zdnd00an1n02x5 FILLER_345_592 ();
 b15zdnd00an1n01x5 FILLER_345_594 ();
 b15zdnd11an1n16x5 FILLER_345_598 ();
 b15zdnd11an1n08x5 FILLER_345_614 ();
 b15zdnd11an1n64x5 FILLER_345_637 ();
 b15zdnd11an1n64x5 FILLER_345_701 ();
 b15zdnd11an1n32x5 FILLER_345_765 ();
 b15zdnd11an1n16x5 FILLER_345_797 ();
 b15zdnd00an1n01x5 FILLER_345_813 ();
 b15zdnd11an1n04x5 FILLER_345_817 ();
 b15zdnd11an1n04x5 FILLER_345_830 ();
 b15zdnd00an1n02x5 FILLER_345_834 ();
 b15zdnd00an1n01x5 FILLER_345_836 ();
 b15zdnd11an1n64x5 FILLER_345_840 ();
 b15zdnd11an1n64x5 FILLER_345_904 ();
 b15zdnd11an1n64x5 FILLER_345_968 ();
 b15zdnd11an1n64x5 FILLER_345_1032 ();
 b15zdnd11an1n64x5 FILLER_345_1096 ();
 b15zdnd11an1n32x5 FILLER_345_1160 ();
 b15zdnd11an1n08x5 FILLER_345_1192 ();
 b15zdnd00an1n02x5 FILLER_345_1200 ();
 b15zdnd11an1n64x5 FILLER_345_1226 ();
 b15zdnd11an1n64x5 FILLER_345_1290 ();
 b15zdnd11an1n64x5 FILLER_345_1354 ();
 b15zdnd11an1n64x5 FILLER_345_1418 ();
 b15zdnd11an1n64x5 FILLER_345_1482 ();
 b15zdnd11an1n32x5 FILLER_345_1546 ();
 b15zdnd11an1n16x5 FILLER_345_1578 ();
 b15zdnd11an1n04x5 FILLER_345_1594 ();
 b15zdnd00an1n02x5 FILLER_345_1598 ();
 b15zdnd00an1n01x5 FILLER_345_1600 ();
 b15zdnd11an1n04x5 FILLER_345_1604 ();
 b15zdnd11an1n04x5 FILLER_345_1611 ();
 b15zdnd11an1n04x5 FILLER_345_1618 ();
 b15zdnd00an1n02x5 FILLER_345_1622 ();
 b15zdnd00an1n01x5 FILLER_345_1624 ();
 b15zdnd11an1n16x5 FILLER_345_1628 ();
 b15zdnd11an1n04x5 FILLER_345_1644 ();
 b15zdnd00an1n02x5 FILLER_345_1648 ();
 b15zdnd11an1n64x5 FILLER_345_1670 ();
 b15zdnd11an1n64x5 FILLER_345_1734 ();
 b15zdnd11an1n64x5 FILLER_345_1798 ();
 b15zdnd11an1n64x5 FILLER_345_1862 ();
 b15zdnd11an1n64x5 FILLER_345_1926 ();
 b15zdnd11an1n64x5 FILLER_345_1990 ();
 b15zdnd11an1n64x5 FILLER_345_2054 ();
 b15zdnd11an1n64x5 FILLER_345_2118 ();
 b15zdnd11an1n64x5 FILLER_345_2182 ();
 b15zdnd11an1n32x5 FILLER_345_2246 ();
 b15zdnd11an1n04x5 FILLER_345_2278 ();
 b15zdnd00an1n02x5 FILLER_345_2282 ();
 b15zdnd11an1n64x5 FILLER_346_8 ();
 b15zdnd11an1n32x5 FILLER_346_72 ();
 b15zdnd11an1n16x5 FILLER_346_104 ();
 b15zdnd00an1n02x5 FILLER_346_120 ();
 b15zdnd11an1n04x5 FILLER_346_154 ();
 b15zdnd11an1n64x5 FILLER_346_161 ();
 b15zdnd11an1n32x5 FILLER_346_225 ();
 b15zdnd11an1n16x5 FILLER_346_257 ();
 b15zdnd11an1n08x5 FILLER_346_273 ();
 b15zdnd00an1n02x5 FILLER_346_281 ();
 b15zdnd00an1n01x5 FILLER_346_283 ();
 b15zdnd11an1n64x5 FILLER_346_296 ();
 b15zdnd11an1n64x5 FILLER_346_360 ();
 b15zdnd11an1n08x5 FILLER_346_424 ();
 b15zdnd00an1n01x5 FILLER_346_432 ();
 b15zdnd11an1n16x5 FILLER_346_442 ();
 b15zdnd00an1n01x5 FILLER_346_458 ();
 b15zdnd11an1n64x5 FILLER_346_473 ();
 b15zdnd11an1n64x5 FILLER_346_537 ();
 b15zdnd11an1n64x5 FILLER_346_601 ();
 b15zdnd11an1n32x5 FILLER_346_665 ();
 b15zdnd11an1n16x5 FILLER_346_697 ();
 b15zdnd11an1n04x5 FILLER_346_713 ();
 b15zdnd00an1n01x5 FILLER_346_717 ();
 b15zdnd11an1n64x5 FILLER_346_726 ();
 b15zdnd11an1n16x5 FILLER_346_790 ();
 b15zdnd11an1n08x5 FILLER_346_806 ();
 b15zdnd00an1n02x5 FILLER_346_814 ();
 b15zdnd11an1n04x5 FILLER_346_819 ();
 b15zdnd11an1n04x5 FILLER_346_826 ();
 b15zdnd11an1n64x5 FILLER_346_833 ();
 b15zdnd11an1n64x5 FILLER_346_897 ();
 b15zdnd11an1n64x5 FILLER_346_961 ();
 b15zdnd11an1n64x5 FILLER_346_1025 ();
 b15zdnd11an1n64x5 FILLER_346_1089 ();
 b15zdnd11an1n64x5 FILLER_346_1153 ();
 b15zdnd11an1n32x5 FILLER_346_1217 ();
 b15zdnd11an1n04x5 FILLER_346_1249 ();
 b15zdnd11an1n64x5 FILLER_346_1270 ();
 b15zdnd11an1n08x5 FILLER_346_1334 ();
 b15zdnd11an1n04x5 FILLER_346_1342 ();
 b15zdnd11an1n64x5 FILLER_346_1358 ();
 b15zdnd11an1n64x5 FILLER_346_1422 ();
 b15zdnd11an1n64x5 FILLER_346_1486 ();
 b15zdnd11an1n64x5 FILLER_346_1550 ();
 b15zdnd11an1n64x5 FILLER_346_1614 ();
 b15zdnd11an1n32x5 FILLER_346_1678 ();
 b15zdnd11an1n08x5 FILLER_346_1710 ();
 b15zdnd00an1n01x5 FILLER_346_1718 ();
 b15zdnd11an1n32x5 FILLER_346_1743 ();
 b15zdnd11an1n08x5 FILLER_346_1775 ();
 b15zdnd11an1n64x5 FILLER_346_1814 ();
 b15zdnd11an1n64x5 FILLER_346_1878 ();
 b15zdnd11an1n64x5 FILLER_346_1942 ();
 b15zdnd11an1n64x5 FILLER_346_2006 ();
 b15zdnd11an1n64x5 FILLER_346_2070 ();
 b15zdnd11an1n16x5 FILLER_346_2134 ();
 b15zdnd11an1n04x5 FILLER_346_2150 ();
 b15zdnd11an1n64x5 FILLER_346_2162 ();
 b15zdnd11an1n32x5 FILLER_346_2226 ();
 b15zdnd11an1n16x5 FILLER_346_2258 ();
 b15zdnd00an1n02x5 FILLER_346_2274 ();
 b15zdnd11an1n64x5 FILLER_347_0 ();
 b15zdnd11an1n08x5 FILLER_347_64 ();
 b15zdnd11an1n04x5 FILLER_347_72 ();
 b15zdnd00an1n01x5 FILLER_347_76 ();
 b15zdnd11an1n16x5 FILLER_347_89 ();
 b15zdnd11an1n08x5 FILLER_347_105 ();
 b15zdnd00an1n01x5 FILLER_347_113 ();
 b15zdnd11an1n64x5 FILLER_347_166 ();
 b15zdnd11an1n32x5 FILLER_347_230 ();
 b15zdnd11an1n16x5 FILLER_347_262 ();
 b15zdnd11an1n08x5 FILLER_347_278 ();
 b15zdnd00an1n01x5 FILLER_347_286 ();
 b15zdnd11an1n64x5 FILLER_347_290 ();
 b15zdnd11an1n64x5 FILLER_347_354 ();
 b15zdnd11an1n64x5 FILLER_347_418 ();
 b15zdnd11an1n32x5 FILLER_347_482 ();
 b15zdnd11an1n08x5 FILLER_347_514 ();
 b15zdnd11an1n04x5 FILLER_347_522 ();
 b15zdnd11an1n64x5 FILLER_347_530 ();
 b15zdnd11an1n64x5 FILLER_347_594 ();
 b15zdnd11an1n64x5 FILLER_347_658 ();
 b15zdnd11an1n64x5 FILLER_347_722 ();
 b15zdnd11an1n32x5 FILLER_347_786 ();
 b15zdnd11an1n04x5 FILLER_347_818 ();
 b15zdnd00an1n02x5 FILLER_347_822 ();
 b15zdnd11an1n64x5 FILLER_347_827 ();
 b15zdnd11an1n64x5 FILLER_347_891 ();
 b15zdnd11an1n64x5 FILLER_347_955 ();
 b15zdnd11an1n64x5 FILLER_347_1019 ();
 b15zdnd11an1n64x5 FILLER_347_1083 ();
 b15zdnd11an1n64x5 FILLER_347_1147 ();
 b15zdnd11an1n64x5 FILLER_347_1211 ();
 b15zdnd11an1n64x5 FILLER_347_1275 ();
 b15zdnd11an1n08x5 FILLER_347_1339 ();
 b15zdnd11an1n04x5 FILLER_347_1347 ();
 b15zdnd11an1n64x5 FILLER_347_1365 ();
 b15zdnd11an1n64x5 FILLER_347_1429 ();
 b15zdnd11an1n64x5 FILLER_347_1493 ();
 b15zdnd11an1n64x5 FILLER_347_1557 ();
 b15zdnd11an1n32x5 FILLER_347_1621 ();
 b15zdnd11an1n08x5 FILLER_347_1653 ();
 b15zdnd11an1n04x5 FILLER_347_1661 ();
 b15zdnd00an1n02x5 FILLER_347_1665 ();
 b15zdnd11an1n64x5 FILLER_347_1687 ();
 b15zdnd11an1n64x5 FILLER_347_1751 ();
 b15zdnd11an1n64x5 FILLER_347_1815 ();
 b15zdnd11an1n64x5 FILLER_347_1879 ();
 b15zdnd11an1n64x5 FILLER_347_1943 ();
 b15zdnd11an1n64x5 FILLER_347_2007 ();
 b15zdnd11an1n64x5 FILLER_347_2071 ();
 b15zdnd11an1n64x5 FILLER_347_2135 ();
 b15zdnd11an1n64x5 FILLER_347_2199 ();
 b15zdnd11an1n16x5 FILLER_347_2263 ();
 b15zdnd11an1n04x5 FILLER_347_2279 ();
 b15zdnd00an1n01x5 FILLER_347_2283 ();
 b15zdnd11an1n64x5 FILLER_348_8 ();
 b15zdnd00an1n01x5 FILLER_348_72 ();
 b15zdnd11an1n32x5 FILLER_348_85 ();
 b15zdnd11an1n16x5 FILLER_348_117 ();
 b15zdnd00an1n01x5 FILLER_348_133 ();
 b15zdnd11an1n04x5 FILLER_348_137 ();
 b15zdnd11an1n64x5 FILLER_348_144 ();
 b15zdnd11an1n08x5 FILLER_348_208 ();
 b15zdnd11an1n04x5 FILLER_348_216 ();
 b15zdnd11an1n32x5 FILLER_348_262 ();
 b15zdnd11an1n16x5 FILLER_348_294 ();
 b15zdnd11an1n04x5 FILLER_348_310 ();
 b15zdnd00an1n02x5 FILLER_348_314 ();
 b15zdnd00an1n01x5 FILLER_348_316 ();
 b15zdnd11an1n64x5 FILLER_348_321 ();
 b15zdnd11an1n64x5 FILLER_348_385 ();
 b15zdnd11an1n64x5 FILLER_348_449 ();
 b15zdnd11an1n64x5 FILLER_348_513 ();
 b15zdnd11an1n64x5 FILLER_348_577 ();
 b15zdnd11an1n64x5 FILLER_348_641 ();
 b15zdnd11an1n08x5 FILLER_348_705 ();
 b15zdnd11an1n04x5 FILLER_348_713 ();
 b15zdnd00an1n01x5 FILLER_348_717 ();
 b15zdnd11an1n64x5 FILLER_348_726 ();
 b15zdnd11an1n64x5 FILLER_348_790 ();
 b15zdnd11an1n64x5 FILLER_348_854 ();
 b15zdnd11an1n64x5 FILLER_348_918 ();
 b15zdnd11an1n64x5 FILLER_348_982 ();
 b15zdnd11an1n64x5 FILLER_348_1046 ();
 b15zdnd11an1n64x5 FILLER_348_1110 ();
 b15zdnd11an1n64x5 FILLER_348_1174 ();
 b15zdnd11an1n64x5 FILLER_348_1238 ();
 b15zdnd11an1n32x5 FILLER_348_1302 ();
 b15zdnd11an1n04x5 FILLER_348_1334 ();
 b15zdnd00an1n02x5 FILLER_348_1338 ();
 b15zdnd11an1n64x5 FILLER_348_1360 ();
 b15zdnd11an1n64x5 FILLER_348_1424 ();
 b15zdnd11an1n64x5 FILLER_348_1488 ();
 b15zdnd11an1n64x5 FILLER_348_1552 ();
 b15zdnd11an1n64x5 FILLER_348_1616 ();
 b15zdnd11an1n64x5 FILLER_348_1680 ();
 b15zdnd11an1n64x5 FILLER_348_1744 ();
 b15zdnd11an1n64x5 FILLER_348_1808 ();
 b15zdnd11an1n64x5 FILLER_348_1872 ();
 b15zdnd11an1n64x5 FILLER_348_1936 ();
 b15zdnd11an1n64x5 FILLER_348_2000 ();
 b15zdnd11an1n64x5 FILLER_348_2064 ();
 b15zdnd11an1n16x5 FILLER_348_2128 ();
 b15zdnd11an1n08x5 FILLER_348_2144 ();
 b15zdnd00an1n02x5 FILLER_348_2152 ();
 b15zdnd11an1n64x5 FILLER_348_2162 ();
 b15zdnd11an1n32x5 FILLER_348_2226 ();
 b15zdnd11an1n16x5 FILLER_348_2258 ();
 b15zdnd00an1n02x5 FILLER_348_2274 ();
 b15zdnd11an1n64x5 FILLER_349_0 ();
 b15zdnd11an1n64x5 FILLER_349_64 ();
 b15zdnd11an1n04x5 FILLER_349_128 ();
 b15zdnd00an1n02x5 FILLER_349_132 ();
 b15zdnd11an1n64x5 FILLER_349_137 ();
 b15zdnd11an1n64x5 FILLER_349_201 ();
 b15zdnd11an1n64x5 FILLER_349_265 ();
 b15zdnd11an1n16x5 FILLER_349_329 ();
 b15zdnd11an1n08x5 FILLER_349_345 ();
 b15zdnd00an1n02x5 FILLER_349_353 ();
 b15zdnd00an1n01x5 FILLER_349_355 ();
 b15zdnd11an1n64x5 FILLER_349_375 ();
 b15zdnd11an1n64x5 FILLER_349_439 ();
 b15zdnd11an1n64x5 FILLER_349_503 ();
 b15zdnd11an1n64x5 FILLER_349_567 ();
 b15zdnd11an1n64x5 FILLER_349_631 ();
 b15zdnd11an1n64x5 FILLER_349_695 ();
 b15zdnd11an1n64x5 FILLER_349_759 ();
 b15zdnd11an1n64x5 FILLER_349_823 ();
 b15zdnd11an1n64x5 FILLER_349_887 ();
 b15zdnd11an1n64x5 FILLER_349_951 ();
 b15zdnd11an1n64x5 FILLER_349_1015 ();
 b15zdnd11an1n64x5 FILLER_349_1079 ();
 b15zdnd11an1n64x5 FILLER_349_1143 ();
 b15zdnd11an1n64x5 FILLER_349_1207 ();
 b15zdnd11an1n64x5 FILLER_349_1271 ();
 b15zdnd11an1n64x5 FILLER_349_1335 ();
 b15zdnd11an1n64x5 FILLER_349_1399 ();
 b15zdnd11an1n64x5 FILLER_349_1463 ();
 b15zdnd11an1n64x5 FILLER_349_1527 ();
 b15zdnd11an1n64x5 FILLER_349_1591 ();
 b15zdnd11an1n32x5 FILLER_349_1655 ();
 b15zdnd11an1n64x5 FILLER_349_1718 ();
 b15zdnd11an1n64x5 FILLER_349_1782 ();
 b15zdnd11an1n64x5 FILLER_349_1846 ();
 b15zdnd11an1n64x5 FILLER_349_1910 ();
 b15zdnd11an1n64x5 FILLER_349_1974 ();
 b15zdnd11an1n64x5 FILLER_349_2038 ();
 b15zdnd11an1n64x5 FILLER_349_2102 ();
 b15zdnd11an1n64x5 FILLER_349_2166 ();
 b15zdnd11an1n32x5 FILLER_349_2230 ();
 b15zdnd11an1n16x5 FILLER_349_2262 ();
 b15zdnd11an1n04x5 FILLER_349_2278 ();
 b15zdnd00an1n02x5 FILLER_349_2282 ();
 b15zdnd11an1n64x5 FILLER_350_8 ();
 b15zdnd11an1n04x5 FILLER_350_72 ();
 b15zdnd00an1n01x5 FILLER_350_76 ();
 b15zdnd11an1n04x5 FILLER_350_81 ();
 b15zdnd11an1n64x5 FILLER_350_89 ();
 b15zdnd11an1n64x5 FILLER_350_153 ();
 b15zdnd11an1n64x5 FILLER_350_217 ();
 b15zdnd11an1n64x5 FILLER_350_281 ();
 b15zdnd11an1n64x5 FILLER_350_345 ();
 b15zdnd11an1n32x5 FILLER_350_409 ();
 b15zdnd11an1n16x5 FILLER_350_441 ();
 b15zdnd11an1n64x5 FILLER_350_494 ();
 b15zdnd11an1n64x5 FILLER_350_558 ();
 b15zdnd11an1n64x5 FILLER_350_622 ();
 b15zdnd11an1n32x5 FILLER_350_686 ();
 b15zdnd11an1n64x5 FILLER_350_726 ();
 b15zdnd11an1n64x5 FILLER_350_790 ();
 b15zdnd11an1n64x5 FILLER_350_854 ();
 b15zdnd11an1n64x5 FILLER_350_918 ();
 b15zdnd11an1n64x5 FILLER_350_982 ();
 b15zdnd11an1n64x5 FILLER_350_1046 ();
 b15zdnd11an1n64x5 FILLER_350_1110 ();
 b15zdnd11an1n64x5 FILLER_350_1174 ();
 b15zdnd11an1n64x5 FILLER_350_1238 ();
 b15zdnd11an1n64x5 FILLER_350_1302 ();
 b15zdnd11an1n64x5 FILLER_350_1366 ();
 b15zdnd11an1n64x5 FILLER_350_1430 ();
 b15zdnd11an1n64x5 FILLER_350_1494 ();
 b15zdnd11an1n64x5 FILLER_350_1558 ();
 b15zdnd11an1n64x5 FILLER_350_1622 ();
 b15zdnd11an1n64x5 FILLER_350_1686 ();
 b15zdnd11an1n64x5 FILLER_350_1750 ();
 b15zdnd11an1n64x5 FILLER_350_1814 ();
 b15zdnd11an1n64x5 FILLER_350_1878 ();
 b15zdnd11an1n64x5 FILLER_350_1942 ();
 b15zdnd11an1n64x5 FILLER_350_2006 ();
 b15zdnd11an1n64x5 FILLER_350_2070 ();
 b15zdnd11an1n16x5 FILLER_350_2134 ();
 b15zdnd11an1n04x5 FILLER_350_2150 ();
 b15zdnd11an1n64x5 FILLER_350_2162 ();
 b15zdnd11an1n32x5 FILLER_350_2226 ();
 b15zdnd11an1n16x5 FILLER_350_2258 ();
 b15zdnd00an1n02x5 FILLER_350_2274 ();
 b15zdnd11an1n64x5 FILLER_351_0 ();
 b15zdnd11an1n64x5 FILLER_351_64 ();
 b15zdnd11an1n64x5 FILLER_351_128 ();
 b15zdnd11an1n32x5 FILLER_351_192 ();
 b15zdnd11an1n16x5 FILLER_351_224 ();
 b15zdnd11an1n08x5 FILLER_351_240 ();
 b15zdnd00an1n02x5 FILLER_351_248 ();
 b15zdnd11an1n64x5 FILLER_351_273 ();
 b15zdnd11an1n64x5 FILLER_351_337 ();
 b15zdnd11an1n64x5 FILLER_351_401 ();
 b15zdnd11an1n64x5 FILLER_351_465 ();
 b15zdnd00an1n01x5 FILLER_351_529 ();
 b15zdnd11an1n04x5 FILLER_351_541 ();
 b15zdnd11an1n64x5 FILLER_351_556 ();
 b15zdnd11an1n32x5 FILLER_351_620 ();
 b15zdnd11an1n16x5 FILLER_351_652 ();
 b15zdnd11an1n08x5 FILLER_351_668 ();
 b15zdnd11an1n04x5 FILLER_351_676 ();
 b15zdnd00an1n02x5 FILLER_351_680 ();
 b15zdnd11an1n64x5 FILLER_351_686 ();
 b15zdnd11an1n64x5 FILLER_351_750 ();
 b15zdnd11an1n64x5 FILLER_351_814 ();
 b15zdnd11an1n64x5 FILLER_351_878 ();
 b15zdnd11an1n64x5 FILLER_351_942 ();
 b15zdnd11an1n64x5 FILLER_351_1006 ();
 b15zdnd11an1n64x5 FILLER_351_1070 ();
 b15zdnd11an1n64x5 FILLER_351_1134 ();
 b15zdnd11an1n64x5 FILLER_351_1198 ();
 b15zdnd11an1n64x5 FILLER_351_1262 ();
 b15zdnd11an1n64x5 FILLER_351_1326 ();
 b15zdnd11an1n64x5 FILLER_351_1390 ();
 b15zdnd11an1n64x5 FILLER_351_1454 ();
 b15zdnd11an1n64x5 FILLER_351_1518 ();
 b15zdnd11an1n64x5 FILLER_351_1582 ();
 b15zdnd11an1n64x5 FILLER_351_1646 ();
 b15zdnd11an1n64x5 FILLER_351_1710 ();
 b15zdnd11an1n64x5 FILLER_351_1774 ();
 b15zdnd11an1n64x5 FILLER_351_1838 ();
 b15zdnd11an1n64x5 FILLER_351_1902 ();
 b15zdnd11an1n64x5 FILLER_351_1966 ();
 b15zdnd11an1n64x5 FILLER_351_2030 ();
 b15zdnd11an1n64x5 FILLER_351_2094 ();
 b15zdnd11an1n64x5 FILLER_351_2158 ();
 b15zdnd11an1n32x5 FILLER_351_2222 ();
 b15zdnd11an1n16x5 FILLER_351_2254 ();
 b15zdnd11an1n08x5 FILLER_351_2270 ();
 b15zdnd11an1n04x5 FILLER_351_2278 ();
 b15zdnd00an1n02x5 FILLER_351_2282 ();
 b15zdnd11an1n64x5 FILLER_352_8 ();
 b15zdnd11an1n64x5 FILLER_352_72 ();
 b15zdnd11an1n64x5 FILLER_352_136 ();
 b15zdnd11an1n64x5 FILLER_352_200 ();
 b15zdnd11an1n64x5 FILLER_352_264 ();
 b15zdnd11an1n64x5 FILLER_352_328 ();
 b15zdnd11an1n32x5 FILLER_352_392 ();
 b15zdnd11an1n16x5 FILLER_352_424 ();
 b15zdnd11an1n08x5 FILLER_352_440 ();
 b15zdnd11an1n04x5 FILLER_352_448 ();
 b15zdnd00an1n02x5 FILLER_352_452 ();
 b15zdnd00an1n01x5 FILLER_352_454 ();
 b15zdnd11an1n32x5 FILLER_352_471 ();
 b15zdnd11an1n16x5 FILLER_352_503 ();
 b15zdnd11an1n08x5 FILLER_352_519 ();
 b15zdnd11an1n04x5 FILLER_352_527 ();
 b15zdnd00an1n01x5 FILLER_352_531 ();
 b15zdnd11an1n64x5 FILLER_352_538 ();
 b15zdnd11an1n64x5 FILLER_352_602 ();
 b15zdnd11an1n32x5 FILLER_352_666 ();
 b15zdnd11an1n16x5 FILLER_352_698 ();
 b15zdnd11an1n04x5 FILLER_352_714 ();
 b15zdnd11an1n64x5 FILLER_352_726 ();
 b15zdnd11an1n64x5 FILLER_352_790 ();
 b15zdnd11an1n64x5 FILLER_352_854 ();
 b15zdnd11an1n64x5 FILLER_352_918 ();
 b15zdnd11an1n64x5 FILLER_352_982 ();
 b15zdnd11an1n64x5 FILLER_352_1046 ();
 b15zdnd11an1n64x5 FILLER_352_1110 ();
 b15zdnd11an1n64x5 FILLER_352_1174 ();
 b15zdnd11an1n64x5 FILLER_352_1238 ();
 b15zdnd11an1n64x5 FILLER_352_1302 ();
 b15zdnd11an1n64x5 FILLER_352_1366 ();
 b15zdnd11an1n64x5 FILLER_352_1430 ();
 b15zdnd11an1n64x5 FILLER_352_1494 ();
 b15zdnd11an1n64x5 FILLER_352_1558 ();
 b15zdnd11an1n64x5 FILLER_352_1622 ();
 b15zdnd11an1n64x5 FILLER_352_1686 ();
 b15zdnd11an1n64x5 FILLER_352_1750 ();
 b15zdnd11an1n64x5 FILLER_352_1814 ();
 b15zdnd11an1n64x5 FILLER_352_1878 ();
 b15zdnd11an1n64x5 FILLER_352_1942 ();
 b15zdnd11an1n64x5 FILLER_352_2006 ();
 b15zdnd11an1n64x5 FILLER_352_2070 ();
 b15zdnd11an1n16x5 FILLER_352_2134 ();
 b15zdnd11an1n04x5 FILLER_352_2150 ();
 b15zdnd11an1n64x5 FILLER_352_2162 ();
 b15zdnd11an1n32x5 FILLER_352_2226 ();
 b15zdnd11an1n16x5 FILLER_352_2258 ();
 b15zdnd00an1n02x5 FILLER_352_2274 ();
 b15zdnd11an1n64x5 FILLER_353_0 ();
 b15zdnd11an1n16x5 FILLER_353_64 ();
 b15zdnd11an1n04x5 FILLER_353_80 ();
 b15zdnd00an1n02x5 FILLER_353_84 ();
 b15zdnd11an1n64x5 FILLER_353_95 ();
 b15zdnd11an1n64x5 FILLER_353_159 ();
 b15zdnd11an1n64x5 FILLER_353_223 ();
 b15zdnd11an1n64x5 FILLER_353_287 ();
 b15zdnd11an1n64x5 FILLER_353_351 ();
 b15zdnd11an1n64x5 FILLER_353_415 ();
 b15zdnd11an1n64x5 FILLER_353_479 ();
 b15zdnd11an1n64x5 FILLER_353_543 ();
 b15zdnd11an1n64x5 FILLER_353_607 ();
 b15zdnd11an1n64x5 FILLER_353_671 ();
 b15zdnd11an1n64x5 FILLER_353_735 ();
 b15zdnd11an1n64x5 FILLER_353_799 ();
 b15zdnd11an1n64x5 FILLER_353_863 ();
 b15zdnd11an1n64x5 FILLER_353_927 ();
 b15zdnd11an1n64x5 FILLER_353_991 ();
 b15zdnd11an1n64x5 FILLER_353_1055 ();
 b15zdnd11an1n64x5 FILLER_353_1119 ();
 b15zdnd11an1n64x5 FILLER_353_1183 ();
 b15zdnd11an1n64x5 FILLER_353_1247 ();
 b15zdnd11an1n64x5 FILLER_353_1311 ();
 b15zdnd11an1n64x5 FILLER_353_1375 ();
 b15zdnd11an1n64x5 FILLER_353_1439 ();
 b15zdnd11an1n64x5 FILLER_353_1503 ();
 b15zdnd11an1n64x5 FILLER_353_1567 ();
 b15zdnd11an1n32x5 FILLER_353_1631 ();
 b15zdnd11an1n04x5 FILLER_353_1663 ();
 b15zdnd11an1n64x5 FILLER_353_1681 ();
 b15zdnd11an1n64x5 FILLER_353_1745 ();
 b15zdnd11an1n64x5 FILLER_353_1809 ();
 b15zdnd11an1n64x5 FILLER_353_1873 ();
 b15zdnd11an1n64x5 FILLER_353_1937 ();
 b15zdnd11an1n64x5 FILLER_353_2001 ();
 b15zdnd11an1n64x5 FILLER_353_2065 ();
 b15zdnd11an1n64x5 FILLER_353_2129 ();
 b15zdnd11an1n64x5 FILLER_353_2193 ();
 b15zdnd11an1n16x5 FILLER_353_2257 ();
 b15zdnd11an1n08x5 FILLER_353_2273 ();
 b15zdnd00an1n02x5 FILLER_353_2281 ();
 b15zdnd00an1n01x5 FILLER_353_2283 ();
 b15zdnd11an1n64x5 FILLER_354_8 ();
 b15zdnd11an1n64x5 FILLER_354_72 ();
 b15zdnd11an1n64x5 FILLER_354_136 ();
 b15zdnd11an1n32x5 FILLER_354_200 ();
 b15zdnd11an1n08x5 FILLER_354_232 ();
 b15zdnd11an1n04x5 FILLER_354_240 ();
 b15zdnd11an1n64x5 FILLER_354_251 ();
 b15zdnd11an1n64x5 FILLER_354_315 ();
 b15zdnd11an1n64x5 FILLER_354_379 ();
 b15zdnd11an1n64x5 FILLER_354_443 ();
 b15zdnd11an1n64x5 FILLER_354_507 ();
 b15zdnd11an1n64x5 FILLER_354_571 ();
 b15zdnd11an1n64x5 FILLER_354_635 ();
 b15zdnd11an1n16x5 FILLER_354_699 ();
 b15zdnd00an1n02x5 FILLER_354_715 ();
 b15zdnd00an1n01x5 FILLER_354_717 ();
 b15zdnd11an1n64x5 FILLER_354_726 ();
 b15zdnd11an1n64x5 FILLER_354_790 ();
 b15zdnd11an1n64x5 FILLER_354_854 ();
 b15zdnd11an1n64x5 FILLER_354_918 ();
 b15zdnd11an1n64x5 FILLER_354_982 ();
 b15zdnd11an1n64x5 FILLER_354_1046 ();
 b15zdnd11an1n64x5 FILLER_354_1110 ();
 b15zdnd11an1n64x5 FILLER_354_1174 ();
 b15zdnd11an1n64x5 FILLER_354_1238 ();
 b15zdnd11an1n64x5 FILLER_354_1302 ();
 b15zdnd11an1n64x5 FILLER_354_1366 ();
 b15zdnd11an1n64x5 FILLER_354_1430 ();
 b15zdnd11an1n64x5 FILLER_354_1494 ();
 b15zdnd11an1n32x5 FILLER_354_1558 ();
 b15zdnd11an1n08x5 FILLER_354_1590 ();
 b15zdnd11an1n04x5 FILLER_354_1598 ();
 b15zdnd11an1n04x5 FILLER_354_1616 ();
 b15zdnd11an1n08x5 FILLER_354_1634 ();
 b15zdnd00an1n02x5 FILLER_354_1642 ();
 b15zdnd00an1n01x5 FILLER_354_1644 ();
 b15zdnd11an1n64x5 FILLER_354_1659 ();
 b15zdnd11an1n64x5 FILLER_354_1723 ();
 b15zdnd11an1n64x5 FILLER_354_1787 ();
 b15zdnd11an1n64x5 FILLER_354_1851 ();
 b15zdnd11an1n64x5 FILLER_354_1915 ();
 b15zdnd11an1n64x5 FILLER_354_1979 ();
 b15zdnd11an1n64x5 FILLER_354_2043 ();
 b15zdnd11an1n32x5 FILLER_354_2107 ();
 b15zdnd11an1n08x5 FILLER_354_2139 ();
 b15zdnd11an1n04x5 FILLER_354_2147 ();
 b15zdnd00an1n02x5 FILLER_354_2151 ();
 b15zdnd00an1n01x5 FILLER_354_2153 ();
 b15zdnd11an1n64x5 FILLER_354_2162 ();
 b15zdnd11an1n32x5 FILLER_354_2226 ();
 b15zdnd11an1n16x5 FILLER_354_2258 ();
 b15zdnd00an1n02x5 FILLER_354_2274 ();
 b15zdnd11an1n64x5 FILLER_355_0 ();
 b15zdnd11an1n08x5 FILLER_355_64 ();
 b15zdnd11an1n04x5 FILLER_355_72 ();
 b15zdnd00an1n01x5 FILLER_355_76 ();
 b15zdnd11an1n64x5 FILLER_355_96 ();
 b15zdnd11an1n64x5 FILLER_355_160 ();
 b15zdnd11an1n64x5 FILLER_355_224 ();
 b15zdnd11an1n64x5 FILLER_355_288 ();
 b15zdnd11an1n64x5 FILLER_355_352 ();
 b15zdnd11an1n64x5 FILLER_355_416 ();
 b15zdnd11an1n64x5 FILLER_355_480 ();
 b15zdnd11an1n64x5 FILLER_355_544 ();
 b15zdnd11an1n64x5 FILLER_355_608 ();
 b15zdnd11an1n64x5 FILLER_355_672 ();
 b15zdnd11an1n64x5 FILLER_355_736 ();
 b15zdnd11an1n64x5 FILLER_355_800 ();
 b15zdnd11an1n64x5 FILLER_355_864 ();
 b15zdnd11an1n64x5 FILLER_355_928 ();
 b15zdnd11an1n64x5 FILLER_355_992 ();
 b15zdnd11an1n64x5 FILLER_355_1056 ();
 b15zdnd11an1n64x5 FILLER_355_1120 ();
 b15zdnd11an1n64x5 FILLER_355_1184 ();
 b15zdnd11an1n64x5 FILLER_355_1248 ();
 b15zdnd11an1n64x5 FILLER_355_1312 ();
 b15zdnd11an1n64x5 FILLER_355_1376 ();
 b15zdnd11an1n64x5 FILLER_355_1440 ();
 b15zdnd11an1n64x5 FILLER_355_1504 ();
 b15zdnd11an1n32x5 FILLER_355_1568 ();
 b15zdnd11an1n16x5 FILLER_355_1600 ();
 b15zdnd11an1n04x5 FILLER_355_1616 ();
 b15zdnd11an1n64x5 FILLER_355_1662 ();
 b15zdnd11an1n64x5 FILLER_355_1726 ();
 b15zdnd11an1n64x5 FILLER_355_1790 ();
 b15zdnd11an1n64x5 FILLER_355_1854 ();
 b15zdnd11an1n64x5 FILLER_355_1918 ();
 b15zdnd11an1n64x5 FILLER_355_1982 ();
 b15zdnd11an1n64x5 FILLER_355_2046 ();
 b15zdnd11an1n64x5 FILLER_355_2110 ();
 b15zdnd11an1n64x5 FILLER_355_2174 ();
 b15zdnd11an1n32x5 FILLER_355_2238 ();
 b15zdnd11an1n08x5 FILLER_355_2270 ();
 b15zdnd11an1n04x5 FILLER_355_2278 ();
 b15zdnd00an1n02x5 FILLER_355_2282 ();
 b15zdnd11an1n64x5 FILLER_356_8 ();
 b15zdnd11an1n64x5 FILLER_356_72 ();
 b15zdnd11an1n64x5 FILLER_356_136 ();
 b15zdnd11an1n16x5 FILLER_356_200 ();
 b15zdnd11an1n08x5 FILLER_356_216 ();
 b15zdnd11an1n04x5 FILLER_356_224 ();
 b15zdnd11an1n16x5 FILLER_356_234 ();
 b15zdnd11an1n08x5 FILLER_356_250 ();
 b15zdnd00an1n02x5 FILLER_356_258 ();
 b15zdnd00an1n01x5 FILLER_356_260 ();
 b15zdnd11an1n64x5 FILLER_356_303 ();
 b15zdnd11an1n32x5 FILLER_356_367 ();
 b15zdnd11an1n08x5 FILLER_356_399 ();
 b15zdnd11an1n04x5 FILLER_356_407 ();
 b15zdnd00an1n02x5 FILLER_356_411 ();
 b15zdnd00an1n01x5 FILLER_356_413 ();
 b15zdnd11an1n64x5 FILLER_356_426 ();
 b15zdnd11an1n64x5 FILLER_356_490 ();
 b15zdnd11an1n64x5 FILLER_356_554 ();
 b15zdnd11an1n64x5 FILLER_356_618 ();
 b15zdnd11an1n32x5 FILLER_356_682 ();
 b15zdnd11an1n04x5 FILLER_356_714 ();
 b15zdnd11an1n64x5 FILLER_356_726 ();
 b15zdnd11an1n64x5 FILLER_356_790 ();
 b15zdnd11an1n64x5 FILLER_356_854 ();
 b15zdnd11an1n64x5 FILLER_356_918 ();
 b15zdnd11an1n64x5 FILLER_356_982 ();
 b15zdnd11an1n64x5 FILLER_356_1046 ();
 b15zdnd11an1n64x5 FILLER_356_1110 ();
 b15zdnd11an1n64x5 FILLER_356_1174 ();
 b15zdnd11an1n64x5 FILLER_356_1238 ();
 b15zdnd11an1n64x5 FILLER_356_1302 ();
 b15zdnd11an1n64x5 FILLER_356_1366 ();
 b15zdnd11an1n64x5 FILLER_356_1430 ();
 b15zdnd11an1n64x5 FILLER_356_1494 ();
 b15zdnd11an1n64x5 FILLER_356_1558 ();
 b15zdnd11an1n64x5 FILLER_356_1622 ();
 b15zdnd11an1n64x5 FILLER_356_1686 ();
 b15zdnd11an1n64x5 FILLER_356_1750 ();
 b15zdnd11an1n64x5 FILLER_356_1814 ();
 b15zdnd11an1n64x5 FILLER_356_1878 ();
 b15zdnd11an1n64x5 FILLER_356_1942 ();
 b15zdnd11an1n32x5 FILLER_356_2006 ();
 b15zdnd11an1n08x5 FILLER_356_2038 ();
 b15zdnd11an1n04x5 FILLER_356_2046 ();
 b15zdnd00an1n01x5 FILLER_356_2050 ();
 b15zdnd11an1n64x5 FILLER_356_2061 ();
 b15zdnd11an1n16x5 FILLER_356_2125 ();
 b15zdnd11an1n08x5 FILLER_356_2141 ();
 b15zdnd11an1n04x5 FILLER_356_2149 ();
 b15zdnd00an1n01x5 FILLER_356_2153 ();
 b15zdnd11an1n64x5 FILLER_356_2162 ();
 b15zdnd11an1n32x5 FILLER_356_2226 ();
 b15zdnd11an1n16x5 FILLER_356_2258 ();
 b15zdnd00an1n02x5 FILLER_356_2274 ();
 b15zdnd11an1n64x5 FILLER_357_0 ();
 b15zdnd11an1n04x5 FILLER_357_64 ();
 b15zdnd00an1n01x5 FILLER_357_68 ();
 b15zdnd11an1n64x5 FILLER_357_73 ();
 b15zdnd11an1n64x5 FILLER_357_137 ();
 b15zdnd11an1n64x5 FILLER_357_201 ();
 b15zdnd11an1n08x5 FILLER_357_265 ();
 b15zdnd11an1n64x5 FILLER_357_277 ();
 b15zdnd11an1n64x5 FILLER_357_341 ();
 b15zdnd11an1n64x5 FILLER_357_405 ();
 b15zdnd11an1n64x5 FILLER_357_469 ();
 b15zdnd11an1n64x5 FILLER_357_533 ();
 b15zdnd11an1n64x5 FILLER_357_597 ();
 b15zdnd11an1n64x5 FILLER_357_661 ();
 b15zdnd11an1n64x5 FILLER_357_725 ();
 b15zdnd11an1n64x5 FILLER_357_789 ();
 b15zdnd11an1n64x5 FILLER_357_853 ();
 b15zdnd11an1n64x5 FILLER_357_917 ();
 b15zdnd11an1n64x5 FILLER_357_981 ();
 b15zdnd11an1n64x5 FILLER_357_1045 ();
 b15zdnd11an1n64x5 FILLER_357_1109 ();
 b15zdnd11an1n64x5 FILLER_357_1173 ();
 b15zdnd11an1n64x5 FILLER_357_1237 ();
 b15zdnd11an1n64x5 FILLER_357_1301 ();
 b15zdnd11an1n64x5 FILLER_357_1365 ();
 b15zdnd11an1n64x5 FILLER_357_1429 ();
 b15zdnd11an1n64x5 FILLER_357_1493 ();
 b15zdnd11an1n64x5 FILLER_357_1557 ();
 b15zdnd11an1n64x5 FILLER_357_1621 ();
 b15zdnd11an1n64x5 FILLER_357_1685 ();
 b15zdnd11an1n64x5 FILLER_357_1749 ();
 b15zdnd11an1n64x5 FILLER_357_1813 ();
 b15zdnd11an1n64x5 FILLER_357_1877 ();
 b15zdnd11an1n64x5 FILLER_357_1941 ();
 b15zdnd11an1n64x5 FILLER_357_2005 ();
 b15zdnd11an1n64x5 FILLER_357_2069 ();
 b15zdnd11an1n64x5 FILLER_357_2133 ();
 b15zdnd11an1n64x5 FILLER_357_2197 ();
 b15zdnd11an1n16x5 FILLER_357_2261 ();
 b15zdnd11an1n04x5 FILLER_357_2277 ();
 b15zdnd00an1n02x5 FILLER_357_2281 ();
 b15zdnd00an1n01x5 FILLER_357_2283 ();
 b15zdnd11an1n64x5 FILLER_358_8 ();
 b15zdnd11an1n64x5 FILLER_358_72 ();
 b15zdnd11an1n64x5 FILLER_358_136 ();
 b15zdnd11an1n64x5 FILLER_358_200 ();
 b15zdnd11an1n08x5 FILLER_358_264 ();
 b15zdnd11an1n64x5 FILLER_358_283 ();
 b15zdnd11an1n64x5 FILLER_358_347 ();
 b15zdnd11an1n64x5 FILLER_358_411 ();
 b15zdnd11an1n64x5 FILLER_358_475 ();
 b15zdnd11an1n64x5 FILLER_358_539 ();
 b15zdnd11an1n64x5 FILLER_358_603 ();
 b15zdnd11an1n32x5 FILLER_358_667 ();
 b15zdnd11an1n16x5 FILLER_358_699 ();
 b15zdnd00an1n02x5 FILLER_358_715 ();
 b15zdnd00an1n01x5 FILLER_358_717 ();
 b15zdnd11an1n64x5 FILLER_358_726 ();
 b15zdnd11an1n64x5 FILLER_358_790 ();
 b15zdnd11an1n64x5 FILLER_358_854 ();
 b15zdnd11an1n64x5 FILLER_358_918 ();
 b15zdnd11an1n64x5 FILLER_358_982 ();
 b15zdnd11an1n64x5 FILLER_358_1046 ();
 b15zdnd11an1n64x5 FILLER_358_1110 ();
 b15zdnd11an1n64x5 FILLER_358_1174 ();
 b15zdnd11an1n64x5 FILLER_358_1238 ();
 b15zdnd11an1n64x5 FILLER_358_1302 ();
 b15zdnd11an1n64x5 FILLER_358_1366 ();
 b15zdnd11an1n64x5 FILLER_358_1430 ();
 b15zdnd11an1n64x5 FILLER_358_1494 ();
 b15zdnd11an1n64x5 FILLER_358_1558 ();
 b15zdnd11an1n64x5 FILLER_358_1622 ();
 b15zdnd11an1n64x5 FILLER_358_1686 ();
 b15zdnd11an1n64x5 FILLER_358_1750 ();
 b15zdnd11an1n64x5 FILLER_358_1814 ();
 b15zdnd11an1n64x5 FILLER_358_1878 ();
 b15zdnd11an1n64x5 FILLER_358_1942 ();
 b15zdnd11an1n64x5 FILLER_358_2006 ();
 b15zdnd11an1n16x5 FILLER_358_2070 ();
 b15zdnd00an1n01x5 FILLER_358_2086 ();
 b15zdnd11an1n32x5 FILLER_358_2101 ();
 b15zdnd11an1n16x5 FILLER_358_2133 ();
 b15zdnd11an1n04x5 FILLER_358_2149 ();
 b15zdnd00an1n01x5 FILLER_358_2153 ();
 b15zdnd11an1n64x5 FILLER_358_2162 ();
 b15zdnd11an1n32x5 FILLER_358_2226 ();
 b15zdnd11an1n16x5 FILLER_358_2258 ();
 b15zdnd00an1n02x5 FILLER_358_2274 ();
 b15zdnd11an1n64x5 FILLER_359_0 ();
 b15zdnd11an1n64x5 FILLER_359_64 ();
 b15zdnd11an1n64x5 FILLER_359_128 ();
 b15zdnd11an1n32x5 FILLER_359_192 ();
 b15zdnd00an1n01x5 FILLER_359_224 ();
 b15zdnd11an1n64x5 FILLER_359_241 ();
 b15zdnd11an1n64x5 FILLER_359_305 ();
 b15zdnd11an1n08x5 FILLER_359_369 ();
 b15zdnd11an1n64x5 FILLER_359_398 ();
 b15zdnd11an1n64x5 FILLER_359_462 ();
 b15zdnd11an1n64x5 FILLER_359_526 ();
 b15zdnd11an1n64x5 FILLER_359_590 ();
 b15zdnd11an1n64x5 FILLER_359_654 ();
 b15zdnd11an1n64x5 FILLER_359_718 ();
 b15zdnd11an1n64x5 FILLER_359_782 ();
 b15zdnd11an1n64x5 FILLER_359_846 ();
 b15zdnd11an1n64x5 FILLER_359_910 ();
 b15zdnd11an1n64x5 FILLER_359_974 ();
 b15zdnd11an1n64x5 FILLER_359_1038 ();
 b15zdnd11an1n64x5 FILLER_359_1102 ();
 b15zdnd11an1n64x5 FILLER_359_1166 ();
 b15zdnd11an1n64x5 FILLER_359_1230 ();
 b15zdnd11an1n64x5 FILLER_359_1294 ();
 b15zdnd11an1n64x5 FILLER_359_1358 ();
 b15zdnd11an1n64x5 FILLER_359_1422 ();
 b15zdnd11an1n64x5 FILLER_359_1486 ();
 b15zdnd11an1n64x5 FILLER_359_1550 ();
 b15zdnd11an1n64x5 FILLER_359_1614 ();
 b15zdnd11an1n64x5 FILLER_359_1678 ();
 b15zdnd11an1n64x5 FILLER_359_1742 ();
 b15zdnd11an1n32x5 FILLER_359_1806 ();
 b15zdnd11an1n08x5 FILLER_359_1838 ();
 b15zdnd00an1n02x5 FILLER_359_1846 ();
 b15zdnd00an1n01x5 FILLER_359_1848 ();
 b15zdnd11an1n04x5 FILLER_359_1863 ();
 b15zdnd11an1n64x5 FILLER_359_1881 ();
 b15zdnd11an1n64x5 FILLER_359_1945 ();
 b15zdnd11an1n64x5 FILLER_359_2009 ();
 b15zdnd11an1n16x5 FILLER_359_2073 ();
 b15zdnd11an1n64x5 FILLER_359_2103 ();
 b15zdnd11an1n64x5 FILLER_359_2167 ();
 b15zdnd11an1n32x5 FILLER_359_2231 ();
 b15zdnd11an1n16x5 FILLER_359_2263 ();
 b15zdnd11an1n04x5 FILLER_359_2279 ();
 b15zdnd00an1n01x5 FILLER_359_2283 ();
 b15zdnd11an1n64x5 FILLER_360_8 ();
 b15zdnd11an1n64x5 FILLER_360_72 ();
 b15zdnd11an1n64x5 FILLER_360_136 ();
 b15zdnd11an1n16x5 FILLER_360_200 ();
 b15zdnd11an1n08x5 FILLER_360_216 ();
 b15zdnd11an1n04x5 FILLER_360_224 ();
 b15zdnd00an1n01x5 FILLER_360_228 ();
 b15zdnd11an1n64x5 FILLER_360_271 ();
 b15zdnd11an1n64x5 FILLER_360_335 ();
 b15zdnd11an1n32x5 FILLER_360_399 ();
 b15zdnd11an1n08x5 FILLER_360_431 ();
 b15zdnd11an1n04x5 FILLER_360_439 ();
 b15zdnd00an1n02x5 FILLER_360_443 ();
 b15zdnd11an1n64x5 FILLER_360_449 ();
 b15zdnd11an1n64x5 FILLER_360_513 ();
 b15zdnd11an1n64x5 FILLER_360_577 ();
 b15zdnd11an1n64x5 FILLER_360_641 ();
 b15zdnd11an1n08x5 FILLER_360_705 ();
 b15zdnd11an1n04x5 FILLER_360_713 ();
 b15zdnd00an1n01x5 FILLER_360_717 ();
 b15zdnd11an1n64x5 FILLER_360_726 ();
 b15zdnd11an1n64x5 FILLER_360_790 ();
 b15zdnd11an1n64x5 FILLER_360_854 ();
 b15zdnd11an1n64x5 FILLER_360_918 ();
 b15zdnd11an1n64x5 FILLER_360_982 ();
 b15zdnd11an1n64x5 FILLER_360_1046 ();
 b15zdnd11an1n64x5 FILLER_360_1110 ();
 b15zdnd11an1n64x5 FILLER_360_1174 ();
 b15zdnd11an1n64x5 FILLER_360_1238 ();
 b15zdnd11an1n64x5 FILLER_360_1302 ();
 b15zdnd11an1n64x5 FILLER_360_1366 ();
 b15zdnd11an1n64x5 FILLER_360_1430 ();
 b15zdnd11an1n64x5 FILLER_360_1494 ();
 b15zdnd11an1n64x5 FILLER_360_1558 ();
 b15zdnd11an1n64x5 FILLER_360_1622 ();
 b15zdnd11an1n64x5 FILLER_360_1686 ();
 b15zdnd11an1n64x5 FILLER_360_1750 ();
 b15zdnd11an1n64x5 FILLER_360_1814 ();
 b15zdnd11an1n64x5 FILLER_360_1878 ();
 b15zdnd11an1n64x5 FILLER_360_1942 ();
 b15zdnd11an1n64x5 FILLER_360_2006 ();
 b15zdnd11an1n64x5 FILLER_360_2070 ();
 b15zdnd11an1n16x5 FILLER_360_2134 ();
 b15zdnd11an1n04x5 FILLER_360_2150 ();
 b15zdnd11an1n64x5 FILLER_360_2162 ();
 b15zdnd11an1n32x5 FILLER_360_2226 ();
 b15zdnd11an1n16x5 FILLER_360_2258 ();
 b15zdnd00an1n02x5 FILLER_360_2274 ();
 b15zdnd11an1n64x5 FILLER_361_0 ();
 b15zdnd11an1n32x5 FILLER_361_64 ();
 b15zdnd11an1n08x5 FILLER_361_96 ();
 b15zdnd11an1n04x5 FILLER_361_104 ();
 b15zdnd00an1n02x5 FILLER_361_108 ();
 b15zdnd00an1n01x5 FILLER_361_110 ();
 b15zdnd11an1n32x5 FILLER_361_129 ();
 b15zdnd11an1n16x5 FILLER_361_161 ();
 b15zdnd00an1n02x5 FILLER_361_177 ();
 b15zdnd00an1n01x5 FILLER_361_179 ();
 b15zdnd11an1n08x5 FILLER_361_196 ();
 b15zdnd00an1n01x5 FILLER_361_204 ();
 b15zdnd11an1n64x5 FILLER_361_217 ();
 b15zdnd11an1n16x5 FILLER_361_281 ();
 b15zdnd11an1n04x5 FILLER_361_297 ();
 b15zdnd00an1n02x5 FILLER_361_301 ();
 b15zdnd11an1n64x5 FILLER_361_311 ();
 b15zdnd00an1n02x5 FILLER_361_375 ();
 b15zdnd00an1n01x5 FILLER_361_377 ();
 b15zdnd11an1n08x5 FILLER_361_398 ();
 b15zdnd00an1n02x5 FILLER_361_406 ();
 b15zdnd11an1n16x5 FILLER_361_422 ();
 b15zdnd11an1n64x5 FILLER_361_454 ();
 b15zdnd11an1n64x5 FILLER_361_518 ();
 b15zdnd11an1n64x5 FILLER_361_582 ();
 b15zdnd11an1n64x5 FILLER_361_646 ();
 b15zdnd11an1n64x5 FILLER_361_710 ();
 b15zdnd11an1n64x5 FILLER_361_774 ();
 b15zdnd11an1n64x5 FILLER_361_838 ();
 b15zdnd11an1n64x5 FILLER_361_902 ();
 b15zdnd11an1n64x5 FILLER_361_966 ();
 b15zdnd11an1n64x5 FILLER_361_1030 ();
 b15zdnd11an1n64x5 FILLER_361_1094 ();
 b15zdnd11an1n64x5 FILLER_361_1158 ();
 b15zdnd11an1n64x5 FILLER_361_1222 ();
 b15zdnd11an1n64x5 FILLER_361_1286 ();
 b15zdnd11an1n64x5 FILLER_361_1350 ();
 b15zdnd11an1n64x5 FILLER_361_1414 ();
 b15zdnd11an1n64x5 FILLER_361_1478 ();
 b15zdnd11an1n64x5 FILLER_361_1542 ();
 b15zdnd11an1n64x5 FILLER_361_1606 ();
 b15zdnd11an1n64x5 FILLER_361_1670 ();
 b15zdnd11an1n64x5 FILLER_361_1734 ();
 b15zdnd11an1n64x5 FILLER_361_1798 ();
 b15zdnd11an1n08x5 FILLER_361_1862 ();
 b15zdnd11an1n04x5 FILLER_361_1870 ();
 b15zdnd00an1n01x5 FILLER_361_1874 ();
 b15zdnd11an1n64x5 FILLER_361_1889 ();
 b15zdnd11an1n64x5 FILLER_361_1953 ();
 b15zdnd11an1n64x5 FILLER_361_2017 ();
 b15zdnd11an1n64x5 FILLER_361_2081 ();
 b15zdnd11an1n64x5 FILLER_361_2145 ();
 b15zdnd11an1n64x5 FILLER_361_2209 ();
 b15zdnd11an1n08x5 FILLER_361_2273 ();
 b15zdnd00an1n02x5 FILLER_361_2281 ();
 b15zdnd00an1n01x5 FILLER_361_2283 ();
 b15zdnd11an1n64x5 FILLER_362_8 ();
 b15zdnd11an1n32x5 FILLER_362_72 ();
 b15zdnd11an1n04x5 FILLER_362_104 ();
 b15zdnd11an1n64x5 FILLER_362_112 ();
 b15zdnd11an1n16x5 FILLER_362_176 ();
 b15zdnd11an1n04x5 FILLER_362_192 ();
 b15zdnd11an1n32x5 FILLER_362_204 ();
 b15zdnd00an1n02x5 FILLER_362_236 ();
 b15zdnd11an1n04x5 FILLER_362_245 ();
 b15zdnd11an1n16x5 FILLER_362_267 ();
 b15zdnd11an1n04x5 FILLER_362_283 ();
 b15zdnd00an1n02x5 FILLER_362_287 ();
 b15zdnd11an1n64x5 FILLER_362_296 ();
 b15zdnd11an1n32x5 FILLER_362_360 ();
 b15zdnd11an1n04x5 FILLER_362_392 ();
 b15zdnd00an1n02x5 FILLER_362_396 ();
 b15zdnd00an1n01x5 FILLER_362_398 ();
 b15zdnd11an1n16x5 FILLER_362_409 ();
 b15zdnd11an1n08x5 FILLER_362_425 ();
 b15zdnd00an1n02x5 FILLER_362_433 ();
 b15zdnd11an1n04x5 FILLER_362_451 ();
 b15zdnd11an1n04x5 FILLER_362_458 ();
 b15zdnd11an1n08x5 FILLER_362_474 ();
 b15zdnd00an1n02x5 FILLER_362_482 ();
 b15zdnd00an1n01x5 FILLER_362_484 ();
 b15zdnd11an1n64x5 FILLER_362_497 ();
 b15zdnd11an1n64x5 FILLER_362_561 ();
 b15zdnd11an1n64x5 FILLER_362_625 ();
 b15zdnd11an1n16x5 FILLER_362_689 ();
 b15zdnd11an1n08x5 FILLER_362_705 ();
 b15zdnd11an1n04x5 FILLER_362_713 ();
 b15zdnd00an1n01x5 FILLER_362_717 ();
 b15zdnd11an1n64x5 FILLER_362_726 ();
 b15zdnd11an1n64x5 FILLER_362_790 ();
 b15zdnd11an1n64x5 FILLER_362_854 ();
 b15zdnd11an1n64x5 FILLER_362_918 ();
 b15zdnd11an1n64x5 FILLER_362_982 ();
 b15zdnd11an1n64x5 FILLER_362_1046 ();
 b15zdnd11an1n64x5 FILLER_362_1110 ();
 b15zdnd11an1n64x5 FILLER_362_1174 ();
 b15zdnd11an1n64x5 FILLER_362_1238 ();
 b15zdnd11an1n64x5 FILLER_362_1302 ();
 b15zdnd11an1n64x5 FILLER_362_1366 ();
 b15zdnd11an1n64x5 FILLER_362_1430 ();
 b15zdnd11an1n64x5 FILLER_362_1494 ();
 b15zdnd11an1n64x5 FILLER_362_1558 ();
 b15zdnd11an1n64x5 FILLER_362_1622 ();
 b15zdnd11an1n64x5 FILLER_362_1686 ();
 b15zdnd11an1n64x5 FILLER_362_1750 ();
 b15zdnd11an1n64x5 FILLER_362_1814 ();
 b15zdnd11an1n64x5 FILLER_362_1878 ();
 b15zdnd11an1n64x5 FILLER_362_1942 ();
 b15zdnd11an1n64x5 FILLER_362_2006 ();
 b15zdnd11an1n64x5 FILLER_362_2070 ();
 b15zdnd11an1n16x5 FILLER_362_2134 ();
 b15zdnd11an1n04x5 FILLER_362_2150 ();
 b15zdnd11an1n64x5 FILLER_362_2162 ();
 b15zdnd11an1n32x5 FILLER_362_2226 ();
 b15zdnd11an1n16x5 FILLER_362_2258 ();
 b15zdnd00an1n02x5 FILLER_362_2274 ();
 b15zdnd11an1n64x5 FILLER_363_0 ();
 b15zdnd11an1n64x5 FILLER_363_64 ();
 b15zdnd11an1n32x5 FILLER_363_128 ();
 b15zdnd11an1n32x5 FILLER_363_176 ();
 b15zdnd11an1n16x5 FILLER_363_208 ();
 b15zdnd11an1n08x5 FILLER_363_224 ();
 b15zdnd11an1n04x5 FILLER_363_232 ();
 b15zdnd00an1n02x5 FILLER_363_236 ();
 b15zdnd00an1n01x5 FILLER_363_238 ();
 b15zdnd11an1n04x5 FILLER_363_257 ();
 b15zdnd11an1n64x5 FILLER_363_279 ();
 b15zdnd11an1n64x5 FILLER_363_343 ();
 b15zdnd11an1n64x5 FILLER_363_407 ();
 b15zdnd11an1n08x5 FILLER_363_471 ();
 b15zdnd11an1n04x5 FILLER_363_479 ();
 b15zdnd00an1n02x5 FILLER_363_483 ();
 b15zdnd00an1n01x5 FILLER_363_485 ();
 b15zdnd11an1n32x5 FILLER_363_490 ();
 b15zdnd11an1n16x5 FILLER_363_522 ();
 b15zdnd11an1n04x5 FILLER_363_538 ();
 b15zdnd00an1n02x5 FILLER_363_542 ();
 b15zdnd00an1n01x5 FILLER_363_544 ();
 b15zdnd11an1n64x5 FILLER_363_559 ();
 b15zdnd11an1n64x5 FILLER_363_623 ();
 b15zdnd11an1n64x5 FILLER_363_687 ();
 b15zdnd11an1n64x5 FILLER_363_751 ();
 b15zdnd11an1n64x5 FILLER_363_815 ();
 b15zdnd11an1n64x5 FILLER_363_879 ();
 b15zdnd11an1n64x5 FILLER_363_943 ();
 b15zdnd11an1n64x5 FILLER_363_1007 ();
 b15zdnd11an1n64x5 FILLER_363_1071 ();
 b15zdnd11an1n64x5 FILLER_363_1135 ();
 b15zdnd11an1n64x5 FILLER_363_1199 ();
 b15zdnd11an1n64x5 FILLER_363_1263 ();
 b15zdnd11an1n64x5 FILLER_363_1327 ();
 b15zdnd11an1n64x5 FILLER_363_1391 ();
 b15zdnd11an1n64x5 FILLER_363_1455 ();
 b15zdnd11an1n64x5 FILLER_363_1519 ();
 b15zdnd11an1n64x5 FILLER_363_1583 ();
 b15zdnd11an1n64x5 FILLER_363_1647 ();
 b15zdnd11an1n64x5 FILLER_363_1711 ();
 b15zdnd11an1n64x5 FILLER_363_1775 ();
 b15zdnd11an1n32x5 FILLER_363_1839 ();
 b15zdnd11an1n16x5 FILLER_363_1871 ();
 b15zdnd00an1n02x5 FILLER_363_1887 ();
 b15zdnd00an1n01x5 FILLER_363_1889 ();
 b15zdnd11an1n64x5 FILLER_363_1904 ();
 b15zdnd11an1n64x5 FILLER_363_1968 ();
 b15zdnd11an1n64x5 FILLER_363_2032 ();
 b15zdnd11an1n64x5 FILLER_363_2096 ();
 b15zdnd11an1n64x5 FILLER_363_2160 ();
 b15zdnd11an1n32x5 FILLER_363_2224 ();
 b15zdnd11an1n16x5 FILLER_363_2256 ();
 b15zdnd11an1n08x5 FILLER_363_2272 ();
 b15zdnd11an1n04x5 FILLER_363_2280 ();
 b15zdnd11an1n64x5 FILLER_364_8 ();
 b15zdnd11an1n64x5 FILLER_364_72 ();
 b15zdnd11an1n32x5 FILLER_364_136 ();
 b15zdnd00an1n02x5 FILLER_364_168 ();
 b15zdnd11an1n32x5 FILLER_364_186 ();
 b15zdnd11an1n04x5 FILLER_364_218 ();
 b15zdnd00an1n02x5 FILLER_364_222 ();
 b15zdnd11an1n04x5 FILLER_364_240 ();
 b15zdnd11an1n16x5 FILLER_364_261 ();
 b15zdnd11an1n08x5 FILLER_364_277 ();
 b15zdnd11an1n04x5 FILLER_364_285 ();
 b15zdnd00an1n01x5 FILLER_364_289 ();
 b15zdnd11an1n64x5 FILLER_364_306 ();
 b15zdnd11an1n64x5 FILLER_364_370 ();
 b15zdnd11an1n16x5 FILLER_364_434 ();
 b15zdnd11an1n04x5 FILLER_364_450 ();
 b15zdnd00an1n01x5 FILLER_364_454 ();
 b15zdnd11an1n64x5 FILLER_364_476 ();
 b15zdnd11an1n08x5 FILLER_364_540 ();
 b15zdnd00an1n02x5 FILLER_364_548 ();
 b15zdnd11an1n04x5 FILLER_364_564 ();
 b15zdnd00an1n02x5 FILLER_364_568 ();
 b15zdnd00an1n01x5 FILLER_364_570 ();
 b15zdnd11an1n64x5 FILLER_364_575 ();
 b15zdnd11an1n64x5 FILLER_364_639 ();
 b15zdnd11an1n08x5 FILLER_364_703 ();
 b15zdnd11an1n04x5 FILLER_364_711 ();
 b15zdnd00an1n02x5 FILLER_364_715 ();
 b15zdnd00an1n01x5 FILLER_364_717 ();
 b15zdnd11an1n64x5 FILLER_364_726 ();
 b15zdnd11an1n64x5 FILLER_364_790 ();
 b15zdnd11an1n64x5 FILLER_364_854 ();
 b15zdnd11an1n64x5 FILLER_364_918 ();
 b15zdnd11an1n64x5 FILLER_364_982 ();
 b15zdnd11an1n64x5 FILLER_364_1046 ();
 b15zdnd11an1n64x5 FILLER_364_1110 ();
 b15zdnd11an1n64x5 FILLER_364_1174 ();
 b15zdnd11an1n64x5 FILLER_364_1238 ();
 b15zdnd11an1n64x5 FILLER_364_1302 ();
 b15zdnd11an1n64x5 FILLER_364_1366 ();
 b15zdnd11an1n64x5 FILLER_364_1430 ();
 b15zdnd11an1n64x5 FILLER_364_1494 ();
 b15zdnd11an1n64x5 FILLER_364_1558 ();
 b15zdnd11an1n64x5 FILLER_364_1622 ();
 b15zdnd11an1n64x5 FILLER_364_1686 ();
 b15zdnd11an1n64x5 FILLER_364_1750 ();
 b15zdnd11an1n64x5 FILLER_364_1814 ();
 b15zdnd11an1n64x5 FILLER_364_1878 ();
 b15zdnd11an1n64x5 FILLER_364_1942 ();
 b15zdnd11an1n64x5 FILLER_364_2006 ();
 b15zdnd11an1n64x5 FILLER_364_2070 ();
 b15zdnd11an1n16x5 FILLER_364_2134 ();
 b15zdnd11an1n04x5 FILLER_364_2150 ();
 b15zdnd11an1n64x5 FILLER_364_2162 ();
 b15zdnd11an1n32x5 FILLER_364_2226 ();
 b15zdnd11an1n16x5 FILLER_364_2258 ();
 b15zdnd00an1n02x5 FILLER_364_2274 ();
 b15zdnd11an1n64x5 FILLER_365_0 ();
 b15zdnd11an1n64x5 FILLER_365_64 ();
 b15zdnd11an1n08x5 FILLER_365_128 ();
 b15zdnd11an1n04x5 FILLER_365_136 ();
 b15zdnd00an1n01x5 FILLER_365_140 ();
 b15zdnd11an1n32x5 FILLER_365_183 ();
 b15zdnd11an1n08x5 FILLER_365_215 ();
 b15zdnd00an1n02x5 FILLER_365_223 ();
 b15zdnd11an1n04x5 FILLER_365_239 ();
 b15zdnd11an1n08x5 FILLER_365_250 ();
 b15zdnd00an1n02x5 FILLER_365_258 ();
 b15zdnd00an1n01x5 FILLER_365_260 ();
 b15zdnd11an1n64x5 FILLER_365_274 ();
 b15zdnd11an1n64x5 FILLER_365_338 ();
 b15zdnd11an1n64x5 FILLER_365_402 ();
 b15zdnd11an1n64x5 FILLER_365_466 ();
 b15zdnd11an1n64x5 FILLER_365_530 ();
 b15zdnd11an1n64x5 FILLER_365_594 ();
 b15zdnd11an1n64x5 FILLER_365_658 ();
 b15zdnd11an1n64x5 FILLER_365_722 ();
 b15zdnd11an1n64x5 FILLER_365_786 ();
 b15zdnd11an1n64x5 FILLER_365_850 ();
 b15zdnd11an1n64x5 FILLER_365_914 ();
 b15zdnd11an1n64x5 FILLER_365_978 ();
 b15zdnd11an1n64x5 FILLER_365_1042 ();
 b15zdnd11an1n64x5 FILLER_365_1106 ();
 b15zdnd11an1n64x5 FILLER_365_1170 ();
 b15zdnd11an1n64x5 FILLER_365_1234 ();
 b15zdnd11an1n64x5 FILLER_365_1298 ();
 b15zdnd11an1n64x5 FILLER_365_1362 ();
 b15zdnd11an1n64x5 FILLER_365_1426 ();
 b15zdnd11an1n64x5 FILLER_365_1490 ();
 b15zdnd11an1n64x5 FILLER_365_1554 ();
 b15zdnd11an1n64x5 FILLER_365_1618 ();
 b15zdnd11an1n64x5 FILLER_365_1682 ();
 b15zdnd11an1n64x5 FILLER_365_1746 ();
 b15zdnd11an1n64x5 FILLER_365_1810 ();
 b15zdnd11an1n64x5 FILLER_365_1874 ();
 b15zdnd11an1n64x5 FILLER_365_1938 ();
 b15zdnd11an1n64x5 FILLER_365_2002 ();
 b15zdnd11an1n64x5 FILLER_365_2066 ();
 b15zdnd11an1n64x5 FILLER_365_2130 ();
 b15zdnd11an1n64x5 FILLER_365_2194 ();
 b15zdnd11an1n16x5 FILLER_365_2258 ();
 b15zdnd11an1n08x5 FILLER_365_2274 ();
 b15zdnd00an1n02x5 FILLER_365_2282 ();
 b15zdnd11an1n64x5 FILLER_366_8 ();
 b15zdnd11an1n64x5 FILLER_366_72 ();
 b15zdnd11an1n64x5 FILLER_366_136 ();
 b15zdnd11an1n64x5 FILLER_366_200 ();
 b15zdnd11an1n64x5 FILLER_366_264 ();
 b15zdnd11an1n64x5 FILLER_366_328 ();
 b15zdnd11an1n64x5 FILLER_366_392 ();
 b15zdnd00an1n02x5 FILLER_366_456 ();
 b15zdnd11an1n64x5 FILLER_366_463 ();
 b15zdnd11an1n64x5 FILLER_366_527 ();
 b15zdnd11an1n64x5 FILLER_366_591 ();
 b15zdnd11an1n32x5 FILLER_366_655 ();
 b15zdnd11an1n16x5 FILLER_366_687 ();
 b15zdnd11an1n08x5 FILLER_366_703 ();
 b15zdnd11an1n04x5 FILLER_366_711 ();
 b15zdnd00an1n02x5 FILLER_366_715 ();
 b15zdnd00an1n01x5 FILLER_366_717 ();
 b15zdnd11an1n64x5 FILLER_366_726 ();
 b15zdnd11an1n64x5 FILLER_366_790 ();
 b15zdnd11an1n64x5 FILLER_366_854 ();
 b15zdnd11an1n64x5 FILLER_366_918 ();
 b15zdnd11an1n64x5 FILLER_366_982 ();
 b15zdnd11an1n64x5 FILLER_366_1046 ();
 b15zdnd11an1n64x5 FILLER_366_1110 ();
 b15zdnd11an1n64x5 FILLER_366_1174 ();
 b15zdnd11an1n64x5 FILLER_366_1238 ();
 b15zdnd11an1n64x5 FILLER_366_1302 ();
 b15zdnd11an1n64x5 FILLER_366_1366 ();
 b15zdnd11an1n64x5 FILLER_366_1430 ();
 b15zdnd11an1n64x5 FILLER_366_1494 ();
 b15zdnd11an1n64x5 FILLER_366_1558 ();
 b15zdnd11an1n64x5 FILLER_366_1622 ();
 b15zdnd11an1n64x5 FILLER_366_1686 ();
 b15zdnd11an1n64x5 FILLER_366_1750 ();
 b15zdnd11an1n64x5 FILLER_366_1814 ();
 b15zdnd11an1n64x5 FILLER_366_1878 ();
 b15zdnd11an1n64x5 FILLER_366_1942 ();
 b15zdnd11an1n64x5 FILLER_366_2006 ();
 b15zdnd11an1n64x5 FILLER_366_2070 ();
 b15zdnd11an1n16x5 FILLER_366_2134 ();
 b15zdnd11an1n04x5 FILLER_366_2150 ();
 b15zdnd11an1n64x5 FILLER_366_2162 ();
 b15zdnd11an1n32x5 FILLER_366_2226 ();
 b15zdnd11an1n16x5 FILLER_366_2258 ();
 b15zdnd00an1n02x5 FILLER_366_2274 ();
 b15zdnd11an1n64x5 FILLER_367_0 ();
 b15zdnd11an1n64x5 FILLER_367_64 ();
 b15zdnd11an1n64x5 FILLER_367_128 ();
 b15zdnd11an1n64x5 FILLER_367_192 ();
 b15zdnd11an1n64x5 FILLER_367_256 ();
 b15zdnd11an1n64x5 FILLER_367_320 ();
 b15zdnd11an1n64x5 FILLER_367_384 ();
 b15zdnd11an1n64x5 FILLER_367_448 ();
 b15zdnd11an1n64x5 FILLER_367_512 ();
 b15zdnd11an1n64x5 FILLER_367_576 ();
 b15zdnd11an1n64x5 FILLER_367_640 ();
 b15zdnd11an1n64x5 FILLER_367_704 ();
 b15zdnd11an1n64x5 FILLER_367_768 ();
 b15zdnd11an1n64x5 FILLER_367_832 ();
 b15zdnd11an1n64x5 FILLER_367_896 ();
 b15zdnd11an1n64x5 FILLER_367_960 ();
 b15zdnd11an1n64x5 FILLER_367_1024 ();
 b15zdnd11an1n64x5 FILLER_367_1088 ();
 b15zdnd11an1n64x5 FILLER_367_1152 ();
 b15zdnd11an1n64x5 FILLER_367_1216 ();
 b15zdnd11an1n64x5 FILLER_367_1280 ();
 b15zdnd11an1n64x5 FILLER_367_1344 ();
 b15zdnd11an1n64x5 FILLER_367_1408 ();
 b15zdnd11an1n64x5 FILLER_367_1472 ();
 b15zdnd11an1n64x5 FILLER_367_1536 ();
 b15zdnd11an1n64x5 FILLER_367_1600 ();
 b15zdnd11an1n64x5 FILLER_367_1664 ();
 b15zdnd11an1n64x5 FILLER_367_1728 ();
 b15zdnd11an1n64x5 FILLER_367_1792 ();
 b15zdnd11an1n64x5 FILLER_367_1856 ();
 b15zdnd11an1n64x5 FILLER_367_1920 ();
 b15zdnd11an1n64x5 FILLER_367_1984 ();
 b15zdnd11an1n64x5 FILLER_367_2048 ();
 b15zdnd11an1n64x5 FILLER_367_2112 ();
 b15zdnd11an1n64x5 FILLER_367_2176 ();
 b15zdnd11an1n32x5 FILLER_367_2240 ();
 b15zdnd11an1n08x5 FILLER_367_2272 ();
 b15zdnd11an1n04x5 FILLER_367_2280 ();
 b15zdnd11an1n64x5 FILLER_368_8 ();
 b15zdnd11an1n64x5 FILLER_368_72 ();
 b15zdnd11an1n64x5 FILLER_368_136 ();
 b15zdnd11an1n64x5 FILLER_368_200 ();
 b15zdnd11an1n64x5 FILLER_368_264 ();
 b15zdnd11an1n08x5 FILLER_368_328 ();
 b15zdnd00an1n02x5 FILLER_368_336 ();
 b15zdnd11an1n64x5 FILLER_368_347 ();
 b15zdnd11an1n08x5 FILLER_368_411 ();
 b15zdnd11an1n04x5 FILLER_368_419 ();
 b15zdnd11an1n64x5 FILLER_368_427 ();
 b15zdnd11an1n64x5 FILLER_368_491 ();
 b15zdnd11an1n64x5 FILLER_368_555 ();
 b15zdnd11an1n64x5 FILLER_368_619 ();
 b15zdnd11an1n32x5 FILLER_368_683 ();
 b15zdnd00an1n02x5 FILLER_368_715 ();
 b15zdnd00an1n01x5 FILLER_368_717 ();
 b15zdnd11an1n64x5 FILLER_368_726 ();
 b15zdnd11an1n64x5 FILLER_368_790 ();
 b15zdnd11an1n64x5 FILLER_368_854 ();
 b15zdnd11an1n64x5 FILLER_368_918 ();
 b15zdnd11an1n64x5 FILLER_368_982 ();
 b15zdnd11an1n64x5 FILLER_368_1046 ();
 b15zdnd11an1n64x5 FILLER_368_1110 ();
 b15zdnd11an1n64x5 FILLER_368_1174 ();
 b15zdnd11an1n64x5 FILLER_368_1238 ();
 b15zdnd11an1n64x5 FILLER_368_1302 ();
 b15zdnd11an1n64x5 FILLER_368_1366 ();
 b15zdnd11an1n64x5 FILLER_368_1430 ();
 b15zdnd11an1n64x5 FILLER_368_1494 ();
 b15zdnd11an1n64x5 FILLER_368_1558 ();
 b15zdnd11an1n64x5 FILLER_368_1622 ();
 b15zdnd11an1n64x5 FILLER_368_1686 ();
 b15zdnd11an1n64x5 FILLER_368_1750 ();
 b15zdnd11an1n64x5 FILLER_368_1814 ();
 b15zdnd11an1n64x5 FILLER_368_1878 ();
 b15zdnd11an1n64x5 FILLER_368_1942 ();
 b15zdnd11an1n64x5 FILLER_368_2006 ();
 b15zdnd11an1n64x5 FILLER_368_2070 ();
 b15zdnd11an1n16x5 FILLER_368_2134 ();
 b15zdnd11an1n04x5 FILLER_368_2150 ();
 b15zdnd11an1n64x5 FILLER_368_2162 ();
 b15zdnd11an1n32x5 FILLER_368_2226 ();
 b15zdnd11an1n16x5 FILLER_368_2258 ();
 b15zdnd00an1n02x5 FILLER_368_2274 ();
 b15zdnd11an1n64x5 FILLER_369_0 ();
 b15zdnd11an1n64x5 FILLER_369_64 ();
 b15zdnd11an1n64x5 FILLER_369_128 ();
 b15zdnd11an1n64x5 FILLER_369_192 ();
 b15zdnd11an1n64x5 FILLER_369_256 ();
 b15zdnd11an1n08x5 FILLER_369_320 ();
 b15zdnd11an1n04x5 FILLER_369_328 ();
 b15zdnd00an1n02x5 FILLER_369_332 ();
 b15zdnd11an1n64x5 FILLER_369_348 ();
 b15zdnd11an1n32x5 FILLER_369_412 ();
 b15zdnd11an1n08x5 FILLER_369_444 ();
 b15zdnd00an1n02x5 FILLER_369_452 ();
 b15zdnd00an1n01x5 FILLER_369_454 ();
 b15zdnd11an1n04x5 FILLER_369_464 ();
 b15zdnd11an1n16x5 FILLER_369_475 ();
 b15zdnd00an1n01x5 FILLER_369_491 ();
 b15zdnd11an1n64x5 FILLER_369_510 ();
 b15zdnd11an1n64x5 FILLER_369_574 ();
 b15zdnd11an1n64x5 FILLER_369_638 ();
 b15zdnd11an1n64x5 FILLER_369_702 ();
 b15zdnd11an1n64x5 FILLER_369_766 ();
 b15zdnd11an1n64x5 FILLER_369_830 ();
 b15zdnd11an1n64x5 FILLER_369_894 ();
 b15zdnd11an1n64x5 FILLER_369_958 ();
 b15zdnd11an1n64x5 FILLER_369_1022 ();
 b15zdnd11an1n64x5 FILLER_369_1086 ();
 b15zdnd11an1n64x5 FILLER_369_1150 ();
 b15zdnd11an1n64x5 FILLER_369_1214 ();
 b15zdnd11an1n64x5 FILLER_369_1278 ();
 b15zdnd11an1n64x5 FILLER_369_1342 ();
 b15zdnd11an1n64x5 FILLER_369_1406 ();
 b15zdnd11an1n64x5 FILLER_369_1470 ();
 b15zdnd11an1n64x5 FILLER_369_1534 ();
 b15zdnd11an1n64x5 FILLER_369_1598 ();
 b15zdnd11an1n64x5 FILLER_369_1662 ();
 b15zdnd11an1n64x5 FILLER_369_1726 ();
 b15zdnd11an1n64x5 FILLER_369_1790 ();
 b15zdnd11an1n64x5 FILLER_369_1854 ();
 b15zdnd11an1n64x5 FILLER_369_1918 ();
 b15zdnd11an1n64x5 FILLER_369_1982 ();
 b15zdnd11an1n64x5 FILLER_369_2046 ();
 b15zdnd11an1n64x5 FILLER_369_2110 ();
 b15zdnd11an1n64x5 FILLER_369_2174 ();
 b15zdnd11an1n32x5 FILLER_369_2238 ();
 b15zdnd11an1n08x5 FILLER_369_2270 ();
 b15zdnd11an1n04x5 FILLER_369_2278 ();
 b15zdnd00an1n02x5 FILLER_369_2282 ();
 b15zdnd11an1n64x5 FILLER_370_8 ();
 b15zdnd11an1n64x5 FILLER_370_72 ();
 b15zdnd11an1n64x5 FILLER_370_136 ();
 b15zdnd11an1n64x5 FILLER_370_200 ();
 b15zdnd11an1n16x5 FILLER_370_264 ();
 b15zdnd00an1n01x5 FILLER_370_280 ();
 b15zdnd11an1n08x5 FILLER_370_293 ();
 b15zdnd11an1n04x5 FILLER_370_301 ();
 b15zdnd00an1n02x5 FILLER_370_305 ();
 b15zdnd00an1n01x5 FILLER_370_307 ();
 b15zdnd11an1n64x5 FILLER_370_315 ();
 b15zdnd11an1n64x5 FILLER_370_379 ();
 b15zdnd11an1n04x5 FILLER_370_443 ();
 b15zdnd00an1n02x5 FILLER_370_447 ();
 b15zdnd11an1n64x5 FILLER_370_462 ();
 b15zdnd11an1n64x5 FILLER_370_526 ();
 b15zdnd11an1n64x5 FILLER_370_590 ();
 b15zdnd11an1n64x5 FILLER_370_654 ();
 b15zdnd11an1n64x5 FILLER_370_726 ();
 b15zdnd11an1n64x5 FILLER_370_790 ();
 b15zdnd11an1n64x5 FILLER_370_854 ();
 b15zdnd11an1n64x5 FILLER_370_918 ();
 b15zdnd11an1n64x5 FILLER_370_982 ();
 b15zdnd11an1n64x5 FILLER_370_1046 ();
 b15zdnd11an1n64x5 FILLER_370_1110 ();
 b15zdnd11an1n64x5 FILLER_370_1174 ();
 b15zdnd11an1n64x5 FILLER_370_1238 ();
 b15zdnd11an1n64x5 FILLER_370_1302 ();
 b15zdnd11an1n64x5 FILLER_370_1366 ();
 b15zdnd11an1n64x5 FILLER_370_1430 ();
 b15zdnd11an1n64x5 FILLER_370_1494 ();
 b15zdnd11an1n64x5 FILLER_370_1558 ();
 b15zdnd11an1n64x5 FILLER_370_1622 ();
 b15zdnd11an1n64x5 FILLER_370_1686 ();
 b15zdnd11an1n64x5 FILLER_370_1750 ();
 b15zdnd11an1n64x5 FILLER_370_1814 ();
 b15zdnd11an1n64x5 FILLER_370_1878 ();
 b15zdnd11an1n64x5 FILLER_370_1942 ();
 b15zdnd11an1n64x5 FILLER_370_2006 ();
 b15zdnd11an1n64x5 FILLER_370_2070 ();
 b15zdnd11an1n16x5 FILLER_370_2134 ();
 b15zdnd11an1n04x5 FILLER_370_2150 ();
 b15zdnd11an1n64x5 FILLER_370_2162 ();
 b15zdnd11an1n32x5 FILLER_370_2226 ();
 b15zdnd11an1n16x5 FILLER_370_2258 ();
 b15zdnd00an1n02x5 FILLER_370_2274 ();
 b15zdnd11an1n64x5 FILLER_371_0 ();
 b15zdnd11an1n64x5 FILLER_371_64 ();
 b15zdnd11an1n64x5 FILLER_371_128 ();
 b15zdnd11an1n64x5 FILLER_371_192 ();
 b15zdnd11an1n64x5 FILLER_371_256 ();
 b15zdnd11an1n16x5 FILLER_371_320 ();
 b15zdnd00an1n02x5 FILLER_371_336 ();
 b15zdnd11an1n32x5 FILLER_371_354 ();
 b15zdnd11an1n16x5 FILLER_371_386 ();
 b15zdnd11an1n08x5 FILLER_371_402 ();
 b15zdnd00an1n02x5 FILLER_371_410 ();
 b15zdnd00an1n01x5 FILLER_371_412 ();
 b15zdnd11an1n16x5 FILLER_371_425 ();
 b15zdnd11an1n08x5 FILLER_371_441 ();
 b15zdnd11an1n64x5 FILLER_371_465 ();
 b15zdnd11an1n64x5 FILLER_371_529 ();
 b15zdnd11an1n64x5 FILLER_371_593 ();
 b15zdnd11an1n64x5 FILLER_371_657 ();
 b15zdnd11an1n64x5 FILLER_371_721 ();
 b15zdnd11an1n64x5 FILLER_371_785 ();
 b15zdnd11an1n64x5 FILLER_371_849 ();
 b15zdnd11an1n64x5 FILLER_371_913 ();
 b15zdnd11an1n64x5 FILLER_371_977 ();
 b15zdnd11an1n64x5 FILLER_371_1041 ();
 b15zdnd11an1n64x5 FILLER_371_1105 ();
 b15zdnd11an1n64x5 FILLER_371_1169 ();
 b15zdnd11an1n64x5 FILLER_371_1233 ();
 b15zdnd11an1n64x5 FILLER_371_1297 ();
 b15zdnd11an1n64x5 FILLER_371_1361 ();
 b15zdnd11an1n64x5 FILLER_371_1425 ();
 b15zdnd11an1n64x5 FILLER_371_1489 ();
 b15zdnd11an1n64x5 FILLER_371_1553 ();
 b15zdnd11an1n64x5 FILLER_371_1617 ();
 b15zdnd11an1n16x5 FILLER_371_1681 ();
 b15zdnd11an1n04x5 FILLER_371_1697 ();
 b15zdnd00an1n02x5 FILLER_371_1701 ();
 b15zdnd00an1n01x5 FILLER_371_1703 ();
 b15zdnd11an1n04x5 FILLER_371_1718 ();
 b15zdnd11an1n64x5 FILLER_371_1736 ();
 b15zdnd11an1n64x5 FILLER_371_1800 ();
 b15zdnd11an1n64x5 FILLER_371_1864 ();
 b15zdnd11an1n64x5 FILLER_371_1928 ();
 b15zdnd11an1n64x5 FILLER_371_1992 ();
 b15zdnd11an1n64x5 FILLER_371_2056 ();
 b15zdnd11an1n64x5 FILLER_371_2120 ();
 b15zdnd11an1n64x5 FILLER_371_2184 ();
 b15zdnd11an1n32x5 FILLER_371_2248 ();
 b15zdnd11an1n04x5 FILLER_371_2280 ();
 b15zdnd11an1n64x5 FILLER_372_8 ();
 b15zdnd11an1n64x5 FILLER_372_72 ();
 b15zdnd11an1n32x5 FILLER_372_136 ();
 b15zdnd00an1n02x5 FILLER_372_168 ();
 b15zdnd11an1n32x5 FILLER_372_187 ();
 b15zdnd11an1n08x5 FILLER_372_219 ();
 b15zdnd11an1n04x5 FILLER_372_227 ();
 b15zdnd00an1n02x5 FILLER_372_231 ();
 b15zdnd11an1n64x5 FILLER_372_239 ();
 b15zdnd11an1n64x5 FILLER_372_303 ();
 b15zdnd11an1n64x5 FILLER_372_367 ();
 b15zdnd11an1n64x5 FILLER_372_431 ();
 b15zdnd11an1n64x5 FILLER_372_495 ();
 b15zdnd11an1n64x5 FILLER_372_559 ();
 b15zdnd11an1n64x5 FILLER_372_623 ();
 b15zdnd11an1n16x5 FILLER_372_687 ();
 b15zdnd11an1n08x5 FILLER_372_703 ();
 b15zdnd11an1n04x5 FILLER_372_711 ();
 b15zdnd00an1n02x5 FILLER_372_715 ();
 b15zdnd00an1n01x5 FILLER_372_717 ();
 b15zdnd11an1n64x5 FILLER_372_726 ();
 b15zdnd11an1n64x5 FILLER_372_790 ();
 b15zdnd11an1n64x5 FILLER_372_854 ();
 b15zdnd11an1n64x5 FILLER_372_918 ();
 b15zdnd11an1n64x5 FILLER_372_982 ();
 b15zdnd11an1n64x5 FILLER_372_1046 ();
 b15zdnd11an1n64x5 FILLER_372_1110 ();
 b15zdnd11an1n64x5 FILLER_372_1174 ();
 b15zdnd11an1n64x5 FILLER_372_1238 ();
 b15zdnd11an1n64x5 FILLER_372_1302 ();
 b15zdnd11an1n64x5 FILLER_372_1366 ();
 b15zdnd11an1n64x5 FILLER_372_1430 ();
 b15zdnd11an1n64x5 FILLER_372_1494 ();
 b15zdnd11an1n64x5 FILLER_372_1558 ();
 b15zdnd11an1n64x5 FILLER_372_1622 ();
 b15zdnd11an1n64x5 FILLER_372_1686 ();
 b15zdnd11an1n64x5 FILLER_372_1750 ();
 b15zdnd11an1n64x5 FILLER_372_1814 ();
 b15zdnd11an1n64x5 FILLER_372_1878 ();
 b15zdnd11an1n64x5 FILLER_372_1942 ();
 b15zdnd11an1n64x5 FILLER_372_2006 ();
 b15zdnd11an1n64x5 FILLER_372_2070 ();
 b15zdnd11an1n16x5 FILLER_372_2134 ();
 b15zdnd11an1n04x5 FILLER_372_2150 ();
 b15zdnd11an1n64x5 FILLER_372_2162 ();
 b15zdnd11an1n32x5 FILLER_372_2226 ();
 b15zdnd11an1n16x5 FILLER_372_2258 ();
 b15zdnd00an1n02x5 FILLER_372_2274 ();
 b15zdnd11an1n64x5 FILLER_373_0 ();
 b15zdnd11an1n64x5 FILLER_373_64 ();
 b15zdnd11an1n64x5 FILLER_373_128 ();
 b15zdnd11an1n64x5 FILLER_373_192 ();
 b15zdnd11an1n64x5 FILLER_373_256 ();
 b15zdnd11an1n64x5 FILLER_373_320 ();
 b15zdnd11an1n64x5 FILLER_373_384 ();
 b15zdnd11an1n64x5 FILLER_373_448 ();
 b15zdnd11an1n64x5 FILLER_373_512 ();
 b15zdnd11an1n64x5 FILLER_373_576 ();
 b15zdnd11an1n64x5 FILLER_373_640 ();
 b15zdnd11an1n64x5 FILLER_373_704 ();
 b15zdnd11an1n64x5 FILLER_373_768 ();
 b15zdnd11an1n64x5 FILLER_373_832 ();
 b15zdnd11an1n64x5 FILLER_373_896 ();
 b15zdnd11an1n64x5 FILLER_373_960 ();
 b15zdnd11an1n64x5 FILLER_373_1024 ();
 b15zdnd11an1n64x5 FILLER_373_1088 ();
 b15zdnd11an1n64x5 FILLER_373_1152 ();
 b15zdnd11an1n64x5 FILLER_373_1216 ();
 b15zdnd11an1n64x5 FILLER_373_1280 ();
 b15zdnd11an1n64x5 FILLER_373_1344 ();
 b15zdnd11an1n64x5 FILLER_373_1408 ();
 b15zdnd11an1n64x5 FILLER_373_1472 ();
 b15zdnd11an1n64x5 FILLER_373_1536 ();
 b15zdnd11an1n64x5 FILLER_373_1600 ();
 b15zdnd11an1n64x5 FILLER_373_1664 ();
 b15zdnd11an1n64x5 FILLER_373_1728 ();
 b15zdnd11an1n64x5 FILLER_373_1792 ();
 b15zdnd11an1n64x5 FILLER_373_1856 ();
 b15zdnd11an1n64x5 FILLER_373_1920 ();
 b15zdnd11an1n64x5 FILLER_373_1984 ();
 b15zdnd11an1n64x5 FILLER_373_2048 ();
 b15zdnd11an1n64x5 FILLER_373_2112 ();
 b15zdnd11an1n64x5 FILLER_373_2176 ();
 b15zdnd11an1n32x5 FILLER_373_2240 ();
 b15zdnd11an1n08x5 FILLER_373_2272 ();
 b15zdnd11an1n04x5 FILLER_373_2280 ();
 b15zdnd11an1n64x5 FILLER_374_8 ();
 b15zdnd11an1n64x5 FILLER_374_72 ();
 b15zdnd11an1n64x5 FILLER_374_136 ();
 b15zdnd11an1n04x5 FILLER_374_200 ();
 b15zdnd00an1n01x5 FILLER_374_204 ();
 b15zdnd11an1n08x5 FILLER_374_221 ();
 b15zdnd00an1n01x5 FILLER_374_229 ();
 b15zdnd11an1n04x5 FILLER_374_245 ();
 b15zdnd11an1n16x5 FILLER_374_257 ();
 b15zdnd00an1n02x5 FILLER_374_273 ();
 b15zdnd11an1n64x5 FILLER_374_293 ();
 b15zdnd11an1n64x5 FILLER_374_357 ();
 b15zdnd11an1n64x5 FILLER_374_421 ();
 b15zdnd11an1n64x5 FILLER_374_485 ();
 b15zdnd11an1n64x5 FILLER_374_549 ();
 b15zdnd11an1n64x5 FILLER_374_613 ();
 b15zdnd11an1n32x5 FILLER_374_677 ();
 b15zdnd11an1n08x5 FILLER_374_709 ();
 b15zdnd00an1n01x5 FILLER_374_717 ();
 b15zdnd11an1n64x5 FILLER_374_726 ();
 b15zdnd11an1n64x5 FILLER_374_790 ();
 b15zdnd11an1n64x5 FILLER_374_854 ();
 b15zdnd11an1n64x5 FILLER_374_918 ();
 b15zdnd11an1n64x5 FILLER_374_982 ();
 b15zdnd11an1n64x5 FILLER_374_1046 ();
 b15zdnd11an1n64x5 FILLER_374_1110 ();
 b15zdnd11an1n64x5 FILLER_374_1174 ();
 b15zdnd11an1n64x5 FILLER_374_1238 ();
 b15zdnd11an1n64x5 FILLER_374_1302 ();
 b15zdnd11an1n64x5 FILLER_374_1366 ();
 b15zdnd11an1n64x5 FILLER_374_1430 ();
 b15zdnd11an1n64x5 FILLER_374_1494 ();
 b15zdnd11an1n64x5 FILLER_374_1558 ();
 b15zdnd11an1n64x5 FILLER_374_1622 ();
 b15zdnd11an1n64x5 FILLER_374_1686 ();
 b15zdnd11an1n64x5 FILLER_374_1750 ();
 b15zdnd11an1n64x5 FILLER_374_1814 ();
 b15zdnd11an1n64x5 FILLER_374_1878 ();
 b15zdnd11an1n64x5 FILLER_374_1942 ();
 b15zdnd11an1n64x5 FILLER_374_2006 ();
 b15zdnd11an1n64x5 FILLER_374_2070 ();
 b15zdnd11an1n16x5 FILLER_374_2134 ();
 b15zdnd11an1n04x5 FILLER_374_2150 ();
 b15zdnd11an1n64x5 FILLER_374_2162 ();
 b15zdnd11an1n32x5 FILLER_374_2226 ();
 b15zdnd11an1n16x5 FILLER_374_2258 ();
 b15zdnd00an1n02x5 FILLER_374_2274 ();
 b15zdnd11an1n64x5 FILLER_375_0 ();
 b15zdnd11an1n64x5 FILLER_375_64 ();
 b15zdnd11an1n64x5 FILLER_375_128 ();
 b15zdnd00an1n02x5 FILLER_375_192 ();
 b15zdnd00an1n01x5 FILLER_375_194 ();
 b15zdnd11an1n04x5 FILLER_375_199 ();
 b15zdnd11an1n04x5 FILLER_375_224 ();
 b15zdnd00an1n02x5 FILLER_375_228 ();
 b15zdnd11an1n32x5 FILLER_375_242 ();
 b15zdnd11an1n04x5 FILLER_375_274 ();
 b15zdnd00an1n01x5 FILLER_375_278 ();
 b15zdnd11an1n16x5 FILLER_375_289 ();
 b15zdnd11an1n08x5 FILLER_375_305 ();
 b15zdnd00an1n01x5 FILLER_375_313 ();
 b15zdnd11an1n04x5 FILLER_375_330 ();
 b15zdnd11an1n08x5 FILLER_375_346 ();
 b15zdnd11an1n04x5 FILLER_375_354 ();
 b15zdnd11an1n64x5 FILLER_375_370 ();
 b15zdnd11an1n64x5 FILLER_375_434 ();
 b15zdnd11an1n64x5 FILLER_375_498 ();
 b15zdnd11an1n64x5 FILLER_375_562 ();
 b15zdnd11an1n64x5 FILLER_375_626 ();
 b15zdnd11an1n64x5 FILLER_375_690 ();
 b15zdnd11an1n64x5 FILLER_375_754 ();
 b15zdnd11an1n64x5 FILLER_375_818 ();
 b15zdnd11an1n64x5 FILLER_375_882 ();
 b15zdnd11an1n64x5 FILLER_375_946 ();
 b15zdnd11an1n64x5 FILLER_375_1010 ();
 b15zdnd11an1n64x5 FILLER_375_1074 ();
 b15zdnd11an1n64x5 FILLER_375_1138 ();
 b15zdnd11an1n64x5 FILLER_375_1202 ();
 b15zdnd11an1n64x5 FILLER_375_1266 ();
 b15zdnd11an1n64x5 FILLER_375_1330 ();
 b15zdnd11an1n64x5 FILLER_375_1394 ();
 b15zdnd11an1n64x5 FILLER_375_1458 ();
 b15zdnd11an1n64x5 FILLER_375_1522 ();
 b15zdnd11an1n64x5 FILLER_375_1586 ();
 b15zdnd11an1n64x5 FILLER_375_1650 ();
 b15zdnd11an1n64x5 FILLER_375_1714 ();
 b15zdnd11an1n64x5 FILLER_375_1778 ();
 b15zdnd11an1n64x5 FILLER_375_1842 ();
 b15zdnd11an1n64x5 FILLER_375_1906 ();
 b15zdnd11an1n64x5 FILLER_375_1970 ();
 b15zdnd11an1n64x5 FILLER_375_2034 ();
 b15zdnd11an1n64x5 FILLER_375_2098 ();
 b15zdnd11an1n64x5 FILLER_375_2162 ();
 b15zdnd11an1n32x5 FILLER_375_2226 ();
 b15zdnd11an1n16x5 FILLER_375_2258 ();
 b15zdnd11an1n08x5 FILLER_375_2274 ();
 b15zdnd00an1n02x5 FILLER_375_2282 ();
 b15zdnd11an1n64x5 FILLER_376_8 ();
 b15zdnd11an1n64x5 FILLER_376_72 ();
 b15zdnd11an1n64x5 FILLER_376_136 ();
 b15zdnd11an1n64x5 FILLER_376_200 ();
 b15zdnd11an1n32x5 FILLER_376_264 ();
 b15zdnd11an1n08x5 FILLER_376_296 ();
 b15zdnd00an1n02x5 FILLER_376_304 ();
 b15zdnd00an1n01x5 FILLER_376_306 ();
 b15zdnd11an1n08x5 FILLER_376_313 ();
 b15zdnd00an1n02x5 FILLER_376_321 ();
 b15zdnd00an1n01x5 FILLER_376_323 ();
 b15zdnd11an1n64x5 FILLER_376_333 ();
 b15zdnd11an1n64x5 FILLER_376_397 ();
 b15zdnd11an1n64x5 FILLER_376_461 ();
 b15zdnd11an1n64x5 FILLER_376_525 ();
 b15zdnd11an1n64x5 FILLER_376_589 ();
 b15zdnd11an1n64x5 FILLER_376_653 ();
 b15zdnd00an1n01x5 FILLER_376_717 ();
 b15zdnd11an1n64x5 FILLER_376_726 ();
 b15zdnd11an1n64x5 FILLER_376_790 ();
 b15zdnd11an1n64x5 FILLER_376_854 ();
 b15zdnd11an1n64x5 FILLER_376_918 ();
 b15zdnd11an1n64x5 FILLER_376_982 ();
 b15zdnd11an1n64x5 FILLER_376_1046 ();
 b15zdnd11an1n64x5 FILLER_376_1110 ();
 b15zdnd11an1n64x5 FILLER_376_1174 ();
 b15zdnd11an1n64x5 FILLER_376_1238 ();
 b15zdnd11an1n64x5 FILLER_376_1302 ();
 b15zdnd11an1n64x5 FILLER_376_1366 ();
 b15zdnd11an1n64x5 FILLER_376_1430 ();
 b15zdnd11an1n64x5 FILLER_376_1494 ();
 b15zdnd11an1n64x5 FILLER_376_1558 ();
 b15zdnd11an1n64x5 FILLER_376_1622 ();
 b15zdnd11an1n64x5 FILLER_376_1686 ();
 b15zdnd11an1n64x5 FILLER_376_1750 ();
 b15zdnd11an1n64x5 FILLER_376_1814 ();
 b15zdnd11an1n64x5 FILLER_376_1878 ();
 b15zdnd11an1n64x5 FILLER_376_1942 ();
 b15zdnd11an1n64x5 FILLER_376_2006 ();
 b15zdnd11an1n64x5 FILLER_376_2070 ();
 b15zdnd11an1n16x5 FILLER_376_2134 ();
 b15zdnd11an1n04x5 FILLER_376_2150 ();
 b15zdnd11an1n64x5 FILLER_376_2162 ();
 b15zdnd11an1n32x5 FILLER_376_2226 ();
 b15zdnd11an1n16x5 FILLER_376_2258 ();
 b15zdnd00an1n02x5 FILLER_376_2274 ();
 b15zdnd11an1n64x5 FILLER_377_0 ();
 b15zdnd11an1n64x5 FILLER_377_64 ();
 b15zdnd11an1n64x5 FILLER_377_128 ();
 b15zdnd11an1n32x5 FILLER_377_192 ();
 b15zdnd11an1n08x5 FILLER_377_224 ();
 b15zdnd11an1n64x5 FILLER_377_250 ();
 b15zdnd11an1n04x5 FILLER_377_314 ();
 b15zdnd00an1n01x5 FILLER_377_318 ();
 b15zdnd11an1n64x5 FILLER_377_340 ();
 b15zdnd11an1n64x5 FILLER_377_404 ();
 b15zdnd11an1n64x5 FILLER_377_468 ();
 b15zdnd11an1n64x5 FILLER_377_532 ();
 b15zdnd11an1n64x5 FILLER_377_596 ();
 b15zdnd11an1n64x5 FILLER_377_660 ();
 b15zdnd11an1n64x5 FILLER_377_724 ();
 b15zdnd11an1n64x5 FILLER_377_788 ();
 b15zdnd11an1n64x5 FILLER_377_852 ();
 b15zdnd11an1n64x5 FILLER_377_916 ();
 b15zdnd11an1n64x5 FILLER_377_980 ();
 b15zdnd11an1n64x5 FILLER_377_1044 ();
 b15zdnd11an1n64x5 FILLER_377_1108 ();
 b15zdnd11an1n64x5 FILLER_377_1172 ();
 b15zdnd11an1n64x5 FILLER_377_1236 ();
 b15zdnd11an1n64x5 FILLER_377_1300 ();
 b15zdnd11an1n64x5 FILLER_377_1364 ();
 b15zdnd11an1n64x5 FILLER_377_1428 ();
 b15zdnd11an1n64x5 FILLER_377_1492 ();
 b15zdnd11an1n64x5 FILLER_377_1556 ();
 b15zdnd11an1n64x5 FILLER_377_1620 ();
 b15zdnd11an1n64x5 FILLER_377_1684 ();
 b15zdnd11an1n64x5 FILLER_377_1748 ();
 b15zdnd11an1n64x5 FILLER_377_1812 ();
 b15zdnd11an1n64x5 FILLER_377_1876 ();
 b15zdnd11an1n64x5 FILLER_377_1940 ();
 b15zdnd11an1n64x5 FILLER_377_2004 ();
 b15zdnd11an1n64x5 FILLER_377_2068 ();
 b15zdnd11an1n64x5 FILLER_377_2132 ();
 b15zdnd11an1n64x5 FILLER_377_2196 ();
 b15zdnd11an1n16x5 FILLER_377_2260 ();
 b15zdnd11an1n08x5 FILLER_377_2276 ();
 b15zdnd11an1n64x5 FILLER_378_8 ();
 b15zdnd11an1n64x5 FILLER_378_72 ();
 b15zdnd11an1n64x5 FILLER_378_136 ();
 b15zdnd11an1n16x5 FILLER_378_200 ();
 b15zdnd11an1n08x5 FILLER_378_216 ();
 b15zdnd11an1n04x5 FILLER_378_224 ();
 b15zdnd00an1n01x5 FILLER_378_228 ();
 b15zdnd11an1n64x5 FILLER_378_235 ();
 b15zdnd11an1n64x5 FILLER_378_299 ();
 b15zdnd11an1n64x5 FILLER_378_363 ();
 b15zdnd11an1n64x5 FILLER_378_427 ();
 b15zdnd11an1n64x5 FILLER_378_491 ();
 b15zdnd11an1n64x5 FILLER_378_555 ();
 b15zdnd11an1n64x5 FILLER_378_619 ();
 b15zdnd11an1n32x5 FILLER_378_683 ();
 b15zdnd00an1n02x5 FILLER_378_715 ();
 b15zdnd00an1n01x5 FILLER_378_717 ();
 b15zdnd11an1n64x5 FILLER_378_726 ();
 b15zdnd11an1n64x5 FILLER_378_790 ();
 b15zdnd11an1n64x5 FILLER_378_854 ();
 b15zdnd11an1n64x5 FILLER_378_918 ();
 b15zdnd11an1n64x5 FILLER_378_982 ();
 b15zdnd11an1n64x5 FILLER_378_1046 ();
 b15zdnd11an1n64x5 FILLER_378_1110 ();
 b15zdnd11an1n64x5 FILLER_378_1174 ();
 b15zdnd11an1n64x5 FILLER_378_1238 ();
 b15zdnd11an1n64x5 FILLER_378_1302 ();
 b15zdnd11an1n64x5 FILLER_378_1366 ();
 b15zdnd11an1n64x5 FILLER_378_1430 ();
 b15zdnd11an1n64x5 FILLER_378_1494 ();
 b15zdnd11an1n64x5 FILLER_378_1558 ();
 b15zdnd11an1n64x5 FILLER_378_1622 ();
 b15zdnd11an1n64x5 FILLER_378_1686 ();
 b15zdnd11an1n64x5 FILLER_378_1750 ();
 b15zdnd11an1n64x5 FILLER_378_1814 ();
 b15zdnd11an1n64x5 FILLER_378_1878 ();
 b15zdnd11an1n64x5 FILLER_378_1942 ();
 b15zdnd11an1n64x5 FILLER_378_2006 ();
 b15zdnd11an1n64x5 FILLER_378_2070 ();
 b15zdnd11an1n16x5 FILLER_378_2134 ();
 b15zdnd11an1n04x5 FILLER_378_2150 ();
 b15zdnd11an1n64x5 FILLER_378_2162 ();
 b15zdnd11an1n32x5 FILLER_378_2226 ();
 b15zdnd11an1n16x5 FILLER_378_2258 ();
 b15zdnd00an1n02x5 FILLER_378_2274 ();
 b15zdnd11an1n64x5 FILLER_379_0 ();
 b15zdnd11an1n64x5 FILLER_379_64 ();
 b15zdnd11an1n64x5 FILLER_379_128 ();
 b15zdnd11an1n16x5 FILLER_379_192 ();
 b15zdnd11an1n08x5 FILLER_379_208 ();
 b15zdnd00an1n02x5 FILLER_379_216 ();
 b15zdnd00an1n01x5 FILLER_379_218 ();
 b15zdnd11an1n08x5 FILLER_379_235 ();
 b15zdnd11an1n04x5 FILLER_379_243 ();
 b15zdnd00an1n02x5 FILLER_379_247 ();
 b15zdnd00an1n01x5 FILLER_379_249 ();
 b15zdnd11an1n64x5 FILLER_379_260 ();
 b15zdnd11an1n32x5 FILLER_379_324 ();
 b15zdnd11an1n04x5 FILLER_379_356 ();
 b15zdnd00an1n02x5 FILLER_379_360 ();
 b15zdnd11an1n64x5 FILLER_379_367 ();
 b15zdnd11an1n64x5 FILLER_379_431 ();
 b15zdnd11an1n64x5 FILLER_379_495 ();
 b15zdnd11an1n64x5 FILLER_379_559 ();
 b15zdnd11an1n64x5 FILLER_379_623 ();
 b15zdnd11an1n64x5 FILLER_379_687 ();
 b15zdnd11an1n64x5 FILLER_379_751 ();
 b15zdnd11an1n64x5 FILLER_379_815 ();
 b15zdnd11an1n64x5 FILLER_379_879 ();
 b15zdnd11an1n64x5 FILLER_379_943 ();
 b15zdnd11an1n64x5 FILLER_379_1007 ();
 b15zdnd11an1n64x5 FILLER_379_1071 ();
 b15zdnd11an1n64x5 FILLER_379_1135 ();
 b15zdnd11an1n64x5 FILLER_379_1199 ();
 b15zdnd11an1n64x5 FILLER_379_1263 ();
 b15zdnd11an1n64x5 FILLER_379_1327 ();
 b15zdnd11an1n64x5 FILLER_379_1391 ();
 b15zdnd11an1n64x5 FILLER_379_1455 ();
 b15zdnd11an1n64x5 FILLER_379_1519 ();
 b15zdnd11an1n64x5 FILLER_379_1583 ();
 b15zdnd11an1n64x5 FILLER_379_1647 ();
 b15zdnd11an1n64x5 FILLER_379_1711 ();
 b15zdnd11an1n64x5 FILLER_379_1775 ();
 b15zdnd11an1n64x5 FILLER_379_1839 ();
 b15zdnd11an1n64x5 FILLER_379_1903 ();
 b15zdnd11an1n64x5 FILLER_379_1967 ();
 b15zdnd11an1n64x5 FILLER_379_2031 ();
 b15zdnd11an1n64x5 FILLER_379_2095 ();
 b15zdnd11an1n64x5 FILLER_379_2159 ();
 b15zdnd11an1n32x5 FILLER_379_2223 ();
 b15zdnd11an1n16x5 FILLER_379_2255 ();
 b15zdnd11an1n08x5 FILLER_379_2271 ();
 b15zdnd11an1n04x5 FILLER_379_2279 ();
 b15zdnd00an1n01x5 FILLER_379_2283 ();
 b15zdnd11an1n64x5 FILLER_380_8 ();
 b15zdnd11an1n64x5 FILLER_380_72 ();
 b15zdnd11an1n32x5 FILLER_380_136 ();
 b15zdnd11an1n16x5 FILLER_380_168 ();
 b15zdnd00an1n02x5 FILLER_380_184 ();
 b15zdnd00an1n01x5 FILLER_380_186 ();
 b15zdnd11an1n04x5 FILLER_380_206 ();
 b15zdnd11an1n04x5 FILLER_380_252 ();
 b15zdnd11an1n04x5 FILLER_380_278 ();
 b15zdnd11an1n08x5 FILLER_380_288 ();
 b15zdnd11an1n04x5 FILLER_380_296 ();
 b15zdnd11an1n16x5 FILLER_380_304 ();
 b15zdnd11an1n04x5 FILLER_380_320 ();
 b15zdnd11an1n04x5 FILLER_380_330 ();
 b15zdnd11an1n04x5 FILLER_380_342 ();
 b15zdnd11an1n64x5 FILLER_380_351 ();
 b15zdnd00an1n01x5 FILLER_380_415 ();
 b15zdnd11an1n04x5 FILLER_380_432 ();
 b15zdnd11an1n08x5 FILLER_380_442 ();
 b15zdnd00an1n01x5 FILLER_380_450 ();
 b15zdnd11an1n64x5 FILLER_380_470 ();
 b15zdnd11an1n64x5 FILLER_380_534 ();
 b15zdnd11an1n64x5 FILLER_380_598 ();
 b15zdnd11an1n32x5 FILLER_380_662 ();
 b15zdnd11an1n16x5 FILLER_380_694 ();
 b15zdnd11an1n08x5 FILLER_380_710 ();
 b15zdnd11an1n64x5 FILLER_380_726 ();
 b15zdnd11an1n64x5 FILLER_380_790 ();
 b15zdnd11an1n64x5 FILLER_380_854 ();
 b15zdnd11an1n64x5 FILLER_380_918 ();
 b15zdnd11an1n64x5 FILLER_380_982 ();
 b15zdnd11an1n64x5 FILLER_380_1046 ();
 b15zdnd11an1n64x5 FILLER_380_1110 ();
 b15zdnd11an1n64x5 FILLER_380_1174 ();
 b15zdnd11an1n64x5 FILLER_380_1238 ();
 b15zdnd11an1n64x5 FILLER_380_1302 ();
 b15zdnd11an1n64x5 FILLER_380_1366 ();
 b15zdnd11an1n64x5 FILLER_380_1430 ();
 b15zdnd11an1n16x5 FILLER_380_1494 ();
 b15zdnd00an1n01x5 FILLER_380_1510 ();
 b15zdnd11an1n64x5 FILLER_380_1519 ();
 b15zdnd11an1n64x5 FILLER_380_1583 ();
 b15zdnd11an1n64x5 FILLER_380_1647 ();
 b15zdnd11an1n64x5 FILLER_380_1711 ();
 b15zdnd11an1n64x5 FILLER_380_1775 ();
 b15zdnd11an1n64x5 FILLER_380_1839 ();
 b15zdnd11an1n64x5 FILLER_380_1903 ();
 b15zdnd11an1n64x5 FILLER_380_1967 ();
 b15zdnd11an1n64x5 FILLER_380_2031 ();
 b15zdnd11an1n32x5 FILLER_380_2095 ();
 b15zdnd11an1n16x5 FILLER_380_2127 ();
 b15zdnd11an1n08x5 FILLER_380_2143 ();
 b15zdnd00an1n02x5 FILLER_380_2151 ();
 b15zdnd00an1n01x5 FILLER_380_2153 ();
 b15zdnd11an1n64x5 FILLER_380_2162 ();
 b15zdnd11an1n32x5 FILLER_380_2226 ();
 b15zdnd11an1n16x5 FILLER_380_2258 ();
 b15zdnd00an1n02x5 FILLER_380_2274 ();
 b15zdnd11an1n64x5 FILLER_381_0 ();
 b15zdnd11an1n64x5 FILLER_381_64 ();
 b15zdnd11an1n32x5 FILLER_381_128 ();
 b15zdnd11an1n16x5 FILLER_381_160 ();
 b15zdnd11an1n08x5 FILLER_381_176 ();
 b15zdnd11an1n04x5 FILLER_381_184 ();
 b15zdnd00an1n02x5 FILLER_381_188 ();
 b15zdnd11an1n16x5 FILLER_381_202 ();
 b15zdnd11an1n04x5 FILLER_381_218 ();
 b15zdnd00an1n02x5 FILLER_381_222 ();
 b15zdnd00an1n01x5 FILLER_381_224 ();
 b15zdnd11an1n64x5 FILLER_381_267 ();
 b15zdnd11an1n64x5 FILLER_381_331 ();
 b15zdnd11an1n64x5 FILLER_381_395 ();
 b15zdnd11an1n64x5 FILLER_381_459 ();
 b15zdnd11an1n64x5 FILLER_381_523 ();
 b15zdnd11an1n64x5 FILLER_381_587 ();
 b15zdnd11an1n64x5 FILLER_381_651 ();
 b15zdnd11an1n64x5 FILLER_381_715 ();
 b15zdnd11an1n64x5 FILLER_381_779 ();
 b15zdnd11an1n64x5 FILLER_381_843 ();
 b15zdnd11an1n64x5 FILLER_381_907 ();
 b15zdnd11an1n64x5 FILLER_381_971 ();
 b15zdnd11an1n64x5 FILLER_381_1035 ();
 b15zdnd11an1n64x5 FILLER_381_1099 ();
 b15zdnd11an1n64x5 FILLER_381_1163 ();
 b15zdnd11an1n64x5 FILLER_381_1227 ();
 b15zdnd11an1n64x5 FILLER_381_1291 ();
 b15zdnd11an1n64x5 FILLER_381_1355 ();
 b15zdnd11an1n64x5 FILLER_381_1419 ();
 b15zdnd11an1n64x5 FILLER_381_1483 ();
 b15zdnd11an1n64x5 FILLER_381_1547 ();
 b15zdnd11an1n64x5 FILLER_381_1611 ();
 b15zdnd11an1n64x5 FILLER_381_1675 ();
 b15zdnd11an1n64x5 FILLER_381_1739 ();
 b15zdnd11an1n64x5 FILLER_381_1803 ();
 b15zdnd11an1n64x5 FILLER_381_1867 ();
 b15zdnd11an1n64x5 FILLER_381_1931 ();
 b15zdnd11an1n64x5 FILLER_381_1995 ();
 b15zdnd11an1n64x5 FILLER_381_2059 ();
 b15zdnd11an1n64x5 FILLER_381_2123 ();
 b15zdnd11an1n64x5 FILLER_381_2187 ();
 b15zdnd11an1n32x5 FILLER_381_2251 ();
 b15zdnd00an1n01x5 FILLER_381_2283 ();
 b15zdnd11an1n64x5 FILLER_382_8 ();
 b15zdnd11an1n64x5 FILLER_382_72 ();
 b15zdnd11an1n32x5 FILLER_382_136 ();
 b15zdnd11an1n16x5 FILLER_382_168 ();
 b15zdnd11an1n04x5 FILLER_382_184 ();
 b15zdnd00an1n01x5 FILLER_382_188 ();
 b15zdnd11an1n16x5 FILLER_382_196 ();
 b15zdnd11an1n08x5 FILLER_382_212 ();
 b15zdnd00an1n02x5 FILLER_382_220 ();
 b15zdnd00an1n01x5 FILLER_382_222 ();
 b15zdnd11an1n64x5 FILLER_382_229 ();
 b15zdnd11an1n64x5 FILLER_382_293 ();
 b15zdnd11an1n64x5 FILLER_382_357 ();
 b15zdnd11an1n64x5 FILLER_382_421 ();
 b15zdnd11an1n64x5 FILLER_382_485 ();
 b15zdnd11an1n64x5 FILLER_382_549 ();
 b15zdnd11an1n64x5 FILLER_382_613 ();
 b15zdnd11an1n32x5 FILLER_382_677 ();
 b15zdnd11an1n08x5 FILLER_382_709 ();
 b15zdnd00an1n01x5 FILLER_382_717 ();
 b15zdnd11an1n64x5 FILLER_382_726 ();
 b15zdnd11an1n64x5 FILLER_382_790 ();
 b15zdnd11an1n64x5 FILLER_382_854 ();
 b15zdnd11an1n64x5 FILLER_382_918 ();
 b15zdnd11an1n64x5 FILLER_382_982 ();
 b15zdnd11an1n64x5 FILLER_382_1046 ();
 b15zdnd11an1n64x5 FILLER_382_1110 ();
 b15zdnd11an1n64x5 FILLER_382_1174 ();
 b15zdnd11an1n64x5 FILLER_382_1238 ();
 b15zdnd11an1n64x5 FILLER_382_1302 ();
 b15zdnd11an1n64x5 FILLER_382_1366 ();
 b15zdnd11an1n64x5 FILLER_382_1430 ();
 b15zdnd11an1n64x5 FILLER_382_1494 ();
 b15zdnd11an1n64x5 FILLER_382_1558 ();
 b15zdnd11an1n64x5 FILLER_382_1622 ();
 b15zdnd11an1n64x5 FILLER_382_1686 ();
 b15zdnd11an1n64x5 FILLER_382_1750 ();
 b15zdnd11an1n64x5 FILLER_382_1814 ();
 b15zdnd11an1n64x5 FILLER_382_1878 ();
 b15zdnd11an1n64x5 FILLER_382_1942 ();
 b15zdnd11an1n64x5 FILLER_382_2006 ();
 b15zdnd11an1n64x5 FILLER_382_2070 ();
 b15zdnd11an1n16x5 FILLER_382_2134 ();
 b15zdnd11an1n04x5 FILLER_382_2150 ();
 b15zdnd11an1n64x5 FILLER_382_2162 ();
 b15zdnd11an1n32x5 FILLER_382_2226 ();
 b15zdnd11an1n16x5 FILLER_382_2258 ();
 b15zdnd00an1n02x5 FILLER_382_2274 ();
 b15zdnd11an1n64x5 FILLER_383_0 ();
 b15zdnd11an1n64x5 FILLER_383_64 ();
 b15zdnd11an1n64x5 FILLER_383_128 ();
 b15zdnd11an1n64x5 FILLER_383_192 ();
 b15zdnd11an1n64x5 FILLER_383_256 ();
 b15zdnd11an1n64x5 FILLER_383_320 ();
 b15zdnd11an1n64x5 FILLER_383_384 ();
 b15zdnd11an1n64x5 FILLER_383_448 ();
 b15zdnd11an1n64x5 FILLER_383_512 ();
 b15zdnd11an1n64x5 FILLER_383_576 ();
 b15zdnd11an1n64x5 FILLER_383_640 ();
 b15zdnd11an1n64x5 FILLER_383_704 ();
 b15zdnd11an1n64x5 FILLER_383_768 ();
 b15zdnd11an1n64x5 FILLER_383_832 ();
 b15zdnd11an1n64x5 FILLER_383_896 ();
 b15zdnd11an1n64x5 FILLER_383_960 ();
 b15zdnd11an1n64x5 FILLER_383_1024 ();
 b15zdnd11an1n64x5 FILLER_383_1088 ();
 b15zdnd11an1n64x5 FILLER_383_1152 ();
 b15zdnd11an1n64x5 FILLER_383_1216 ();
 b15zdnd11an1n64x5 FILLER_383_1280 ();
 b15zdnd11an1n64x5 FILLER_383_1344 ();
 b15zdnd11an1n64x5 FILLER_383_1408 ();
 b15zdnd11an1n64x5 FILLER_383_1472 ();
 b15zdnd11an1n64x5 FILLER_383_1536 ();
 b15zdnd11an1n64x5 FILLER_383_1600 ();
 b15zdnd11an1n64x5 FILLER_383_1664 ();
 b15zdnd11an1n64x5 FILLER_383_1728 ();
 b15zdnd11an1n64x5 FILLER_383_1792 ();
 b15zdnd11an1n64x5 FILLER_383_1856 ();
 b15zdnd11an1n64x5 FILLER_383_1920 ();
 b15zdnd11an1n64x5 FILLER_383_1984 ();
 b15zdnd11an1n64x5 FILLER_383_2048 ();
 b15zdnd11an1n64x5 FILLER_383_2112 ();
 b15zdnd11an1n64x5 FILLER_383_2176 ();
 b15zdnd11an1n32x5 FILLER_383_2240 ();
 b15zdnd11an1n08x5 FILLER_383_2272 ();
 b15zdnd11an1n04x5 FILLER_383_2280 ();
 b15zdnd11an1n64x5 FILLER_384_8 ();
 b15zdnd11an1n64x5 FILLER_384_72 ();
 b15zdnd11an1n64x5 FILLER_384_136 ();
 b15zdnd11an1n64x5 FILLER_384_200 ();
 b15zdnd11an1n64x5 FILLER_384_264 ();
 b15zdnd11an1n64x5 FILLER_384_328 ();
 b15zdnd11an1n64x5 FILLER_384_392 ();
 b15zdnd11an1n64x5 FILLER_384_456 ();
 b15zdnd11an1n64x5 FILLER_384_520 ();
 b15zdnd11an1n64x5 FILLER_384_584 ();
 b15zdnd11an1n64x5 FILLER_384_648 ();
 b15zdnd11an1n04x5 FILLER_384_712 ();
 b15zdnd00an1n02x5 FILLER_384_716 ();
 b15zdnd11an1n64x5 FILLER_384_726 ();
 b15zdnd11an1n64x5 FILLER_384_790 ();
 b15zdnd11an1n64x5 FILLER_384_854 ();
 b15zdnd11an1n64x5 FILLER_384_918 ();
 b15zdnd11an1n64x5 FILLER_384_982 ();
 b15zdnd11an1n64x5 FILLER_384_1046 ();
 b15zdnd11an1n64x5 FILLER_384_1110 ();
 b15zdnd11an1n64x5 FILLER_384_1174 ();
 b15zdnd11an1n64x5 FILLER_384_1238 ();
 b15zdnd11an1n64x5 FILLER_384_1302 ();
 b15zdnd11an1n64x5 FILLER_384_1366 ();
 b15zdnd11an1n64x5 FILLER_384_1430 ();
 b15zdnd11an1n64x5 FILLER_384_1494 ();
 b15zdnd11an1n64x5 FILLER_384_1558 ();
 b15zdnd11an1n64x5 FILLER_384_1622 ();
 b15zdnd11an1n64x5 FILLER_384_1686 ();
 b15zdnd11an1n64x5 FILLER_384_1750 ();
 b15zdnd11an1n64x5 FILLER_384_1814 ();
 b15zdnd11an1n64x5 FILLER_384_1878 ();
 b15zdnd11an1n64x5 FILLER_384_1942 ();
 b15zdnd11an1n64x5 FILLER_384_2006 ();
 b15zdnd11an1n64x5 FILLER_384_2070 ();
 b15zdnd11an1n16x5 FILLER_384_2134 ();
 b15zdnd11an1n04x5 FILLER_384_2150 ();
 b15zdnd11an1n64x5 FILLER_384_2162 ();
 b15zdnd11an1n32x5 FILLER_384_2226 ();
 b15zdnd11an1n16x5 FILLER_384_2258 ();
 b15zdnd00an1n02x5 FILLER_384_2274 ();
 b15zdnd11an1n64x5 FILLER_385_0 ();
 b15zdnd11an1n64x5 FILLER_385_64 ();
 b15zdnd11an1n64x5 FILLER_385_128 ();
 b15zdnd11an1n64x5 FILLER_385_192 ();
 b15zdnd11an1n64x5 FILLER_385_256 ();
 b15zdnd11an1n64x5 FILLER_385_320 ();
 b15zdnd11an1n64x5 FILLER_385_384 ();
 b15zdnd11an1n64x5 FILLER_385_448 ();
 b15zdnd11an1n64x5 FILLER_385_512 ();
 b15zdnd11an1n64x5 FILLER_385_576 ();
 b15zdnd11an1n64x5 FILLER_385_640 ();
 b15zdnd11an1n64x5 FILLER_385_704 ();
 b15zdnd11an1n64x5 FILLER_385_768 ();
 b15zdnd11an1n64x5 FILLER_385_832 ();
 b15zdnd11an1n64x5 FILLER_385_896 ();
 b15zdnd11an1n64x5 FILLER_385_960 ();
 b15zdnd11an1n64x5 FILLER_385_1024 ();
 b15zdnd11an1n64x5 FILLER_385_1088 ();
 b15zdnd11an1n64x5 FILLER_385_1152 ();
 b15zdnd11an1n64x5 FILLER_385_1216 ();
 b15zdnd11an1n64x5 FILLER_385_1280 ();
 b15zdnd11an1n64x5 FILLER_385_1344 ();
 b15zdnd11an1n64x5 FILLER_385_1408 ();
 b15zdnd11an1n64x5 FILLER_385_1472 ();
 b15zdnd11an1n64x5 FILLER_385_1536 ();
 b15zdnd11an1n64x5 FILLER_385_1600 ();
 b15zdnd11an1n64x5 FILLER_385_1664 ();
 b15zdnd11an1n64x5 FILLER_385_1728 ();
 b15zdnd11an1n64x5 FILLER_385_1792 ();
 b15zdnd11an1n64x5 FILLER_385_1856 ();
 b15zdnd11an1n64x5 FILLER_385_1920 ();
 b15zdnd11an1n64x5 FILLER_385_1984 ();
 b15zdnd11an1n64x5 FILLER_385_2048 ();
 b15zdnd11an1n64x5 FILLER_385_2112 ();
 b15zdnd11an1n64x5 FILLER_385_2176 ();
 b15zdnd11an1n32x5 FILLER_385_2240 ();
 b15zdnd11an1n08x5 FILLER_385_2272 ();
 b15zdnd11an1n04x5 FILLER_385_2280 ();
 b15zdnd11an1n64x5 FILLER_386_8 ();
 b15zdnd11an1n64x5 FILLER_386_72 ();
 b15zdnd11an1n64x5 FILLER_386_136 ();
 b15zdnd11an1n64x5 FILLER_386_200 ();
 b15zdnd11an1n64x5 FILLER_386_264 ();
 b15zdnd11an1n64x5 FILLER_386_328 ();
 b15zdnd11an1n64x5 FILLER_386_392 ();
 b15zdnd11an1n64x5 FILLER_386_456 ();
 b15zdnd11an1n64x5 FILLER_386_520 ();
 b15zdnd11an1n64x5 FILLER_386_584 ();
 b15zdnd11an1n64x5 FILLER_386_648 ();
 b15zdnd11an1n04x5 FILLER_386_712 ();
 b15zdnd00an1n02x5 FILLER_386_716 ();
 b15zdnd11an1n32x5 FILLER_386_726 ();
 b15zdnd00an1n01x5 FILLER_386_758 ();
 b15zdnd11an1n64x5 FILLER_386_770 ();
 b15zdnd11an1n64x5 FILLER_386_834 ();
 b15zdnd11an1n64x5 FILLER_386_898 ();
 b15zdnd11an1n64x5 FILLER_386_962 ();
 b15zdnd11an1n64x5 FILLER_386_1026 ();
 b15zdnd11an1n64x5 FILLER_386_1090 ();
 b15zdnd11an1n64x5 FILLER_386_1154 ();
 b15zdnd11an1n64x5 FILLER_386_1218 ();
 b15zdnd11an1n64x5 FILLER_386_1282 ();
 b15zdnd11an1n64x5 FILLER_386_1346 ();
 b15zdnd11an1n64x5 FILLER_386_1410 ();
 b15zdnd11an1n64x5 FILLER_386_1474 ();
 b15zdnd11an1n64x5 FILLER_386_1538 ();
 b15zdnd11an1n64x5 FILLER_386_1602 ();
 b15zdnd11an1n64x5 FILLER_386_1666 ();
 b15zdnd11an1n64x5 FILLER_386_1730 ();
 b15zdnd11an1n64x5 FILLER_386_1794 ();
 b15zdnd11an1n64x5 FILLER_386_1858 ();
 b15zdnd11an1n64x5 FILLER_386_1922 ();
 b15zdnd11an1n64x5 FILLER_386_1986 ();
 b15zdnd11an1n64x5 FILLER_386_2050 ();
 b15zdnd11an1n32x5 FILLER_386_2114 ();
 b15zdnd11an1n08x5 FILLER_386_2146 ();
 b15zdnd11an1n64x5 FILLER_386_2162 ();
 b15zdnd11an1n32x5 FILLER_386_2226 ();
 b15zdnd11an1n16x5 FILLER_386_2258 ();
 b15zdnd00an1n02x5 FILLER_386_2274 ();
 b15zdnd11an1n64x5 FILLER_387_0 ();
 b15zdnd11an1n64x5 FILLER_387_64 ();
 b15zdnd11an1n64x5 FILLER_387_128 ();
 b15zdnd11an1n64x5 FILLER_387_192 ();
 b15zdnd11an1n64x5 FILLER_387_256 ();
 b15zdnd11an1n64x5 FILLER_387_320 ();
 b15zdnd11an1n64x5 FILLER_387_384 ();
 b15zdnd11an1n64x5 FILLER_387_448 ();
 b15zdnd11an1n64x5 FILLER_387_512 ();
 b15zdnd11an1n64x5 FILLER_387_576 ();
 b15zdnd11an1n64x5 FILLER_387_640 ();
 b15zdnd11an1n32x5 FILLER_387_704 ();
 b15zdnd11an1n08x5 FILLER_387_736 ();
 b15zdnd00an1n02x5 FILLER_387_744 ();
 b15zdnd11an1n64x5 FILLER_387_760 ();
 b15zdnd11an1n64x5 FILLER_387_824 ();
 b15zdnd11an1n64x5 FILLER_387_888 ();
 b15zdnd11an1n64x5 FILLER_387_952 ();
 b15zdnd11an1n64x5 FILLER_387_1016 ();
 b15zdnd11an1n64x5 FILLER_387_1080 ();
 b15zdnd11an1n64x5 FILLER_387_1144 ();
 b15zdnd11an1n64x5 FILLER_387_1208 ();
 b15zdnd11an1n64x5 FILLER_387_1272 ();
 b15zdnd11an1n64x5 FILLER_387_1336 ();
 b15zdnd11an1n64x5 FILLER_387_1400 ();
 b15zdnd11an1n64x5 FILLER_387_1464 ();
 b15zdnd11an1n64x5 FILLER_387_1528 ();
 b15zdnd11an1n64x5 FILLER_387_1592 ();
 b15zdnd11an1n64x5 FILLER_387_1656 ();
 b15zdnd11an1n64x5 FILLER_387_1720 ();
 b15zdnd11an1n64x5 FILLER_387_1784 ();
 b15zdnd11an1n16x5 FILLER_387_1848 ();
 b15zdnd00an1n02x5 FILLER_387_1864 ();
 b15zdnd00an1n01x5 FILLER_387_1866 ();
 b15zdnd11an1n64x5 FILLER_387_1881 ();
 b15zdnd11an1n64x5 FILLER_387_1945 ();
 b15zdnd11an1n64x5 FILLER_387_2009 ();
 b15zdnd11an1n64x5 FILLER_387_2073 ();
 b15zdnd11an1n64x5 FILLER_387_2137 ();
 b15zdnd11an1n64x5 FILLER_387_2201 ();
 b15zdnd11an1n16x5 FILLER_387_2265 ();
 b15zdnd00an1n02x5 FILLER_387_2281 ();
 b15zdnd00an1n01x5 FILLER_387_2283 ();
 b15zdnd11an1n64x5 FILLER_388_8 ();
 b15zdnd11an1n64x5 FILLER_388_72 ();
 b15zdnd11an1n64x5 FILLER_388_136 ();
 b15zdnd11an1n64x5 FILLER_388_200 ();
 b15zdnd11an1n64x5 FILLER_388_264 ();
 b15zdnd11an1n64x5 FILLER_388_328 ();
 b15zdnd11an1n64x5 FILLER_388_392 ();
 b15zdnd11an1n64x5 FILLER_388_456 ();
 b15zdnd11an1n64x5 FILLER_388_520 ();
 b15zdnd11an1n64x5 FILLER_388_584 ();
 b15zdnd11an1n64x5 FILLER_388_648 ();
 b15zdnd11an1n04x5 FILLER_388_712 ();
 b15zdnd00an1n02x5 FILLER_388_716 ();
 b15zdnd11an1n64x5 FILLER_388_726 ();
 b15zdnd11an1n64x5 FILLER_388_790 ();
 b15zdnd11an1n16x5 FILLER_388_854 ();
 b15zdnd11an1n08x5 FILLER_388_870 ();
 b15zdnd11an1n04x5 FILLER_388_878 ();
 b15zdnd00an1n02x5 FILLER_388_882 ();
 b15zdnd11an1n32x5 FILLER_388_898 ();
 b15zdnd11an1n04x5 FILLER_388_930 ();
 b15zdnd00an1n02x5 FILLER_388_934 ();
 b15zdnd00an1n01x5 FILLER_388_936 ();
 b15zdnd11an1n04x5 FILLER_388_948 ();
 b15zdnd11an1n64x5 FILLER_388_963 ();
 b15zdnd11an1n64x5 FILLER_388_1027 ();
 b15zdnd11an1n64x5 FILLER_388_1091 ();
 b15zdnd00an1n02x5 FILLER_388_1155 ();
 b15zdnd11an1n08x5 FILLER_388_1171 ();
 b15zdnd00an1n01x5 FILLER_388_1179 ();
 b15zdnd11an1n64x5 FILLER_388_1194 ();
 b15zdnd11an1n64x5 FILLER_388_1258 ();
 b15zdnd11an1n64x5 FILLER_388_1322 ();
 b15zdnd11an1n64x5 FILLER_388_1386 ();
 b15zdnd11an1n16x5 FILLER_388_1450 ();
 b15zdnd11an1n04x5 FILLER_388_1466 ();
 b15zdnd00an1n02x5 FILLER_388_1470 ();
 b15zdnd11an1n04x5 FILLER_388_1476 ();
 b15zdnd11an1n64x5 FILLER_388_1484 ();
 b15zdnd11an1n64x5 FILLER_388_1548 ();
 b15zdnd11an1n64x5 FILLER_388_1612 ();
 b15zdnd11an1n64x5 FILLER_388_1676 ();
 b15zdnd11an1n64x5 FILLER_388_1740 ();
 b15zdnd11an1n64x5 FILLER_388_1804 ();
 b15zdnd11an1n64x5 FILLER_388_1868 ();
 b15zdnd11an1n64x5 FILLER_388_1932 ();
 b15zdnd11an1n64x5 FILLER_388_1996 ();
 b15zdnd11an1n64x5 FILLER_388_2060 ();
 b15zdnd11an1n16x5 FILLER_388_2124 ();
 b15zdnd11an1n08x5 FILLER_388_2140 ();
 b15zdnd11an1n04x5 FILLER_388_2148 ();
 b15zdnd00an1n02x5 FILLER_388_2152 ();
 b15zdnd11an1n64x5 FILLER_388_2162 ();
 b15zdnd11an1n32x5 FILLER_388_2226 ();
 b15zdnd11an1n16x5 FILLER_388_2258 ();
 b15zdnd00an1n02x5 FILLER_388_2274 ();
 b15zdnd11an1n64x5 FILLER_389_0 ();
 b15zdnd11an1n64x5 FILLER_389_64 ();
 b15zdnd11an1n64x5 FILLER_389_128 ();
 b15zdnd11an1n64x5 FILLER_389_192 ();
 b15zdnd11an1n64x5 FILLER_389_256 ();
 b15zdnd11an1n64x5 FILLER_389_320 ();
 b15zdnd11an1n64x5 FILLER_389_384 ();
 b15zdnd11an1n64x5 FILLER_389_448 ();
 b15zdnd11an1n64x5 FILLER_389_512 ();
 b15zdnd11an1n64x5 FILLER_389_576 ();
 b15zdnd11an1n64x5 FILLER_389_640 ();
 b15zdnd11an1n32x5 FILLER_389_704 ();
 b15zdnd11an1n04x5 FILLER_389_736 ();
 b15zdnd00an1n01x5 FILLER_389_740 ();
 b15zdnd11an1n08x5 FILLER_389_752 ();
 b15zdnd00an1n02x5 FILLER_389_760 ();
 b15zdnd11an1n64x5 FILLER_389_776 ();
 b15zdnd11an1n32x5 FILLER_389_840 ();
 b15zdnd11an1n16x5 FILLER_389_872 ();
 b15zdnd11an1n04x5 FILLER_389_888 ();
 b15zdnd00an1n02x5 FILLER_389_892 ();
 b15zdnd11an1n32x5 FILLER_389_908 ();
 b15zdnd11an1n08x5 FILLER_389_940 ();
 b15zdnd11an1n04x5 FILLER_389_948 ();
 b15zdnd00an1n02x5 FILLER_389_952 ();
 b15zdnd00an1n01x5 FILLER_389_954 ();
 b15zdnd11an1n04x5 FILLER_389_969 ();
 b15zdnd00an1n01x5 FILLER_389_973 ();
 b15zdnd11an1n64x5 FILLER_389_988 ();
 b15zdnd11an1n64x5 FILLER_389_1052 ();
 b15zdnd11an1n16x5 FILLER_389_1116 ();
 b15zdnd11an1n08x5 FILLER_389_1132 ();
 b15zdnd11an1n16x5 FILLER_389_1154 ();
 b15zdnd11an1n64x5 FILLER_389_1184 ();
 b15zdnd11an1n64x5 FILLER_389_1248 ();
 b15zdnd00an1n01x5 FILLER_389_1312 ();
 b15zdnd11an1n08x5 FILLER_389_1327 ();
 b15zdnd11an1n04x5 FILLER_389_1335 ();
 b15zdnd11an1n64x5 FILLER_389_1353 ();
 b15zdnd11an1n32x5 FILLER_389_1417 ();
 b15zdnd11an1n16x5 FILLER_389_1449 ();
 b15zdnd00an1n02x5 FILLER_389_1465 ();
 b15zdnd11an1n64x5 FILLER_389_1509 ();
 b15zdnd11an1n16x5 FILLER_389_1573 ();
 b15zdnd11an1n04x5 FILLER_389_1589 ();
 b15zdnd00an1n01x5 FILLER_389_1593 ();
 b15zdnd11an1n04x5 FILLER_389_1608 ();
 b15zdnd11an1n16x5 FILLER_389_1626 ();
 b15zdnd11an1n04x5 FILLER_389_1653 ();
 b15zdnd11an1n16x5 FILLER_389_1668 ();
 b15zdnd11an1n08x5 FILLER_389_1684 ();
 b15zdnd11an1n04x5 FILLER_389_1692 ();
 b15zdnd11an1n04x5 FILLER_389_1710 ();
 b15zdnd11an1n64x5 FILLER_389_1728 ();
 b15zdnd11an1n32x5 FILLER_389_1792 ();
 b15zdnd11an1n16x5 FILLER_389_1824 ();
 b15zdnd00an1n01x5 FILLER_389_1840 ();
 b15zdnd11an1n04x5 FILLER_389_1855 ();
 b15zdnd11an1n04x5 FILLER_389_1873 ();
 b15zdnd11an1n32x5 FILLER_389_1891 ();
 b15zdnd11an1n08x5 FILLER_389_1923 ();
 b15zdnd11an1n04x5 FILLER_389_1931 ();
 b15zdnd00an1n02x5 FILLER_389_1935 ();
 b15zdnd11an1n64x5 FILLER_389_1948 ();
 b15zdnd11an1n64x5 FILLER_389_2012 ();
 b15zdnd11an1n08x5 FILLER_389_2076 ();
 b15zdnd00an1n02x5 FILLER_389_2084 ();
 b15zdnd11an1n08x5 FILLER_389_2100 ();
 b15zdnd11an1n64x5 FILLER_389_2122 ();
 b15zdnd11an1n64x5 FILLER_389_2186 ();
 b15zdnd11an1n32x5 FILLER_389_2250 ();
 b15zdnd00an1n02x5 FILLER_389_2282 ();
endmodule
