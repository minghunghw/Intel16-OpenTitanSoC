// ##############################################################################
// ## Intel Top Secret                                                         ##
// ##############################################################################
// ## Copyright © Intel Corporation.                                           ##
// ##                                                                          ##
// ## This is the property of Intel Corporation and may only be utilized       ##
// ## pursuant to a written Restricted Use Nondisclosure Agreement             ##
// ## with Intel Corporation.  It may not be used, reproduced, or              ##
// ## disclosed to others except in accordance with the terms and              ##
// ## conditions of such agreement.                                            ##
// ##                                                                          ##
// ## All products, processes, computer systems, dates, and figures            ##
// ## specified are preliminary based on current expectations, and are         ##
// ## subject to change without notice.                                        ##
// ##############################################################################
// ## Text_Tag % __Placeholder neutral1


`ifdef INTCNOPWR
      //do nothing
`else
      `define POWER_AWARE_MODE
`endif



// `timescale 1ps/1ps



primitive INTCseq_cdiar2ah_0( MGM_CLK0, clk `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
  output MGM_CLK0;
  input clk;
  `ifdef POWER_AWARE_MODE
  input vcc, vssx;
  `endif

  table
  `ifdef POWER_AWARE_MODE
  //clk vcc, vssx: MGM_CLK0
    1  1  0: 1;
    0  1  0: 0;
  `else
  //clk: MGM_CLK0
    1: 1;
    0: 0;
  `endif
  endtable

endprimitive


primitive INTCseq_cdiar2ah_1( MGM_C0, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
  output MGM_C0;
  input rb;
  `ifdef POWER_AWARE_MODE
  input vcc, vssx;
  `endif

  table
  `ifdef POWER_AWARE_MODE
  //rb vcc, vssx: MGM_C0
    0  1  0: 1;
    1  1  0: 0;
  `else
  //rb: MGM_C0
    0: 1;
    1: 0;
  `endif
  endtable

endprimitive


primitive INTCseq_cdiar2ah_N_IQ_FF_UDP( Q, C, P, CK, D `ifdef POWER_AWARE_MODE , vcc, vssx `endif , N );
   output Q;
   reg Q;
   input C, P, CK, D, N; 
   `ifdef POWER_AWARE_MODE
   input vcc, vssx;
   `endif
   table 
  `ifdef POWER_AWARE_MODE
   //C  P  CK D  PW GN N  :  Q  :  Q 
     0  0  n  ?  1  0  ?  :  ?  :  -;
     ?  0  n  ?  1  0  ?  :  0  :  0;
     0  ?  n  ?  1  0  ?  :  1  :  1;
     ?  0  r  0  1  0  ?  :  ?  :  0;
     1  0  ?  ?  1  0  ?  :  ?  :  0;
     0  ?  r  1  1  0  ?  :  ?  :  1;
     0  1  ?  ?  1  0  ?  :  ?  :  1;
     0  0  ?  *  1  0  ?  :  ?  :  -;
     0  ?  ?  *  1  0  ?  :  1  :  1;
     ?  0  ?  *  1  0  ?  :  0  :  0;
     0  *  ?  ?  1  0  ?  :  1  :  1;
     *  0  ?  ?  1  0  ?  :  0  :  0;
     ?  0  *  0  1  0  ?  :  0  :  0;
     0  ?  *  1  1  0  ?  :  1  :  1;
     ?  ?  ?  ?  1  0  *  :  ?  :  x;
  `else
   //C  P  CK D  N  :  Q  :  Q 
     0  0  n  ?  ?  :  ?  :  -;
     ?  0  n  ?  ?  :  0  :  0;
     0  ?  n  ?  ?  :  1  :  1;
     ?  0  r  0  ?  :  ?  :  0;
     1  0  ?  ?  ?  :  ?  :  0;
     0  ?  r  1  ?  :  ?  :  1;
     0  1  ?  ?  ?  :  ?  :  1;
     0  0  ?  *  ?  :  ?  :  -;
     0  ?  ?  *  ?  :  1  :  1;
     ?  0  ?  *  ?  :  0  :  0;
     0  *  ?  ?  ?  :  1  :  1;
     *  0  ?  ?  ?  :  0  :  0;
     ?  0  *  0  ?  :  0  :  0;
     0  ?  *  1  ?  :  1  :  1;
     ?  ?  ?  ?  *  :  ?  :  x;
  `endif

endtable
endprimitive



`celldefine
module INTCseq_cdiar2ah_func( clk, clkout, d, rb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, notifier;
   output clkout;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_D0, d, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( clkout, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_cdiar2ah_1( MGM_D0, d );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( clkout, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15cdiar2ah1n04x5( clk, clkout, d, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cdiar2ah_func b15cdiar2ah1n04x5_behav_inst(.clk(clk),.clkout(clkout),.d(d),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cdiar2ah_func b15cdiar2ah1n04x5_behav_inst(.clk(clk),.clkout(clkout),.d(d),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cdiar2ah_func b15cdiar2ah1n04x5_inst(.clk(clk_delay),.clkout(clkout),.d(d_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cdiar2ah_func b15cdiar2ah1n04x5_inst(.clk(clk_delay),.clkout(clkout),.d(d_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> clkout
      (posedge clk => (clkout : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> clkout
      (posedge clk => (clkout : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> clkout
      (negedge rb => (clkout +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> clkout
      (negedge rb => (clkout +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc rb --> clkout
      (negedge rb => (clkout +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> clkout
      (negedge rb => (clkout +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cdiar2ah1n08x5( clk, clkout, d, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cdiar2ah_func b15cdiar2ah1n08x5_behav_inst(.clk(clk),.clkout(clkout),.d(d),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cdiar2ah_func b15cdiar2ah1n08x5_behav_inst(.clk(clk),.clkout(clkout),.d(d),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cdiar2ah_func b15cdiar2ah1n08x5_inst(.clk(clk_delay),.clkout(clkout),.d(d_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cdiar2ah_func b15cdiar2ah1n08x5_inst(.clk(clk_delay),.clkout(clkout),.d(d_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> clkout
      (posedge clk => (clkout : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> clkout
      (posedge clk => (clkout : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> clkout
      (negedge rb => (clkout +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> clkout
      (negedge rb => (clkout +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc rb --> clkout
      (negedge rb => (clkout +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> clkout
      (negedge rb => (clkout +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_cdiyr2ah_func( clk, clkout, d, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, notifier;
   output clkout;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, d, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( clkout, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_0( MGM_D0, d );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( clkout, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15cdiyr2ah1n04x5( clk, clkout, d `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cdiyr2ah_func b15cdiyr2ah1n04x5_behav_inst(.clk(clk),.clkout(clkout),.d(d),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cdiyr2ah_func b15cdiyr2ah1n04x5_behav_inst(.clk(clk),.clkout(clkout),.d(d),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cdiyr2ah_func b15cdiyr2ah1n04x5_inst(.clk(clk_delay),.clkout(clkout),.d(d_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cdiyr2ah_func b15cdiyr2ah1n04x5_inst(.clk(clk_delay),.clkout(clkout),.d(d_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> clkout
      (posedge clk => (clkout : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> clkout
      (posedge clk => (clkout : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cdiyr2ah1n08x5( clk, clkout, d `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cdiyr2ah_func b15cdiyr2ah1n08x5_behav_inst(.clk(clk),.clkout(clkout),.d(d),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cdiyr2ah_func b15cdiyr2ah1n08x5_behav_inst(.clk(clk),.clkout(clkout),.d(d),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cdiyr2ah_func b15cdiyr2ah1n08x5_inst(.clk(clk_delay),.clkout(clkout),.d(d_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cdiyr2ah_func b15cdiyr2ah1n08x5_inst(.clk(clk_delay),.clkout(clkout),.d(d_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> clkout
      (posedge clk => (clkout : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> clkout
      (posedge clk => (clkout : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine


primitive INTCseq_cilao5ah_2( MGM_D0, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
  output MGM_D0;
  input en, te;
  `ifdef POWER_AWARE_MODE
  input vcc, vssx;
  `endif

  table
  `ifdef POWER_AWARE_MODE
  //en, te vcc, vssx: MGM_D0
    1  ?  1  0: 1;
    ?  1  1  0: 1;
    0  0  1  0: 0;
  `else
  //en, te: MGM_D0
    1  ?: 1;
    ?  1: 1;
    0  0: 0;
  `endif
  endtable

endprimitive


primitive INTCseq_cilao5ah_N_IQ_LATCH_UDP( Q, C, P, CK, D `ifdef POWER_AWARE_MODE , vcc, vssx `endif , N );
   output Q;
   reg Q;
   input C, P, CK, D, N; 
   `ifdef POWER_AWARE_MODE
   input vcc, vssx;
   `endif
   table 
  `ifdef POWER_AWARE_MODE
   //C  P  CK D  PW GN N  :  Q  :  Q 
     0  0  0  ?  1  0  ?  :  ?  :  -;
     ?  0  1  0  1  0  ?  :  ?  :  0;
     ?  0  ?  0  1  0  ?  :  0  :  0;
     ?  0  0  ?  1  0  ?  :  0  :  0;
     1  0  ?  ?  1  0  ?  :  ?  :  0;
     0  ?  1  1  1  0  ?  :  ?  :  1;
     0  ?  ?  1  1  0  ?  :  1  :  1;
     0  ?  0  ?  1  0  ?  :  1  :  1;
     0  1  ?  ?  1  0  ?  :  ?  :  1;
     ?  ?  ?  ?  1  0  *  :  ?  :  x;
  `else
   //C  P  CK D  N  :  Q  :  Q 
     0  0  0  ?  ?  :  ?  :  -;
     ?  0  1  0  ?  :  ?  :  0;
     ?  0  ?  0  ?  :  0  :  0;
     ?  0  0  ?  ?  :  0  :  0;
     1  0  ?  ?  ?  :  ?  :  0;
     0  ?  1  1  ?  :  ?  :  1;
     0  ?  ?  1  ?  :  1  :  1;
     0  ?  0  ?  ?  :  1  :  1;
     0  1  ?  ?  ?  :  ?  :  1;
     ?  ?  ?  ?  *  :  ?  :  x;
  `endif

endtable
endprimitive


primitive INTCseq_cilao5ah_3( clkout, IQ, clk `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
  output clkout;
  input IQ, clk;
  `ifdef POWER_AWARE_MODE
  input vcc, vssx;
  `endif

  table
  `ifdef POWER_AWARE_MODE
  //IQ, clk vcc, vssx: clkout
    1  1  1  0: 1;
    0  ?  1  0: 0;
    ?  0  1  0: 0;
  `else
  //IQ, clk: clkout
    1  1: 1;
    0  ?: 0;
    ?  0: 0;
  `endif
  endtable

endprimitive



`celldefine
module INTCseq_cilao5ah_func( clk, clkout, en, te, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te, notifier;
   output clkout;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_1( MGM_EN0, clk, vcc, vssx );
   INTCseq_cilao5ah_2( MGM_D0, en, te, vcc, vssx );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, 1'b0, 1'b0, MGM_EN0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cilao5ah_3( clkout, IQ, clk, vcc, vssx );
`else
   INTCseq_cdiar2ah_1( MGM_EN0, clk );
   INTCseq_cilao5ah_2( MGM_D0, en, te );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, 1'b0, 1'b0, MGM_EN0, MGM_D0, notifier );
   INTCseq_cilao5ah_3( clkout, IQ, clk );
`endif

endmodule
`endcelldefine



`celldefine
module b15cilao5ah1n02x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilao5ah_func b15cilao5ah1n02x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilao5ah_func b15cilao5ah1n02x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilao5ah_func b15cilao5ah1n02x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilao5ah_func b15cilao5ah1n02x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilao5ah1n04x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilao5ah_func b15cilao5ah1n04x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilao5ah_func b15cilao5ah1n04x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilao5ah_func b15cilao5ah1n04x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilao5ah_func b15cilao5ah1n04x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilao5ah1n06x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilao5ah_func b15cilao5ah1n06x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilao5ah_func b15cilao5ah1n06x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilao5ah_func b15cilao5ah1n06x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilao5ah_func b15cilao5ah1n06x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilao5ah1n08x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilao5ah_func b15cilao5ah1n08x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilao5ah_func b15cilao5ah1n08x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilao5ah_func b15cilao5ah1n08x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilao5ah_func b15cilao5ah1n08x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilao5ah1n12x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilao5ah_func b15cilao5ah1n12x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilao5ah_func b15cilao5ah1n12x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilao5ah_func b15cilao5ah1n12x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilao5ah_func b15cilao5ah1n12x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilao5ah1n16x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilao5ah_func b15cilao5ah1n16x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilao5ah_func b15cilao5ah1n16x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilao5ah_func b15cilao5ah1n16x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilao5ah_func b15cilao5ah1n16x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_cilb01ah_func( clk, clkout, en, te, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te, notifier;
   output clkout;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_1( MGM_EN0, clk, vcc, vssx );
   INTCseq_cilao5ah_2( MGM_D0, en, te, vcc, vssx );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, 1'b0, 1'b0, MGM_EN0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cilao5ah_3( clkout, IQ, clk, vcc, vssx );
`else
   INTCseq_cdiar2ah_1( MGM_EN0, clk );
   INTCseq_cilao5ah_2( MGM_D0, en, te );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, 1'b0, 1'b0, MGM_EN0, MGM_D0, notifier );
   INTCseq_cilao5ah_3( clkout, IQ, clk );
`endif

endmodule
`endcelldefine



`celldefine
module b15cilb01ah1n02x3( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n02x3_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n02x3_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n02x3_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n02x3_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb01ah1n02x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n02x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n02x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n02x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n02x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb01ah1n03x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n03x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n03x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n03x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n03x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb01ah1n04x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n04x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n04x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n04x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n04x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb01ah1n06x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n06x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n06x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n06x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n06x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb01ah1n08x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n08x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n08x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n08x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n08x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb01ah1n12x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n12x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n12x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n12x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n12x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb01ah1n16x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n16x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n16x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n16x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n16x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb01ah1n24x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n24x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n24x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n24x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n24x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb01ah1n32x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n32x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n32x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n32x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n32x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb01ah1n48x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n48x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n48x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n48x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n48x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb01ah1n64x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n64x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n64x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n64x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n64x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb01ah1n80x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n80x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n80x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb01ah_func b15cilb01ah1n80x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb01ah_func b15cilb01ah1n80x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_cilb05ah_func( clk, clkout, en, te, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te, notifier;
   output clkout;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_1( MGM_EN0, clk, vcc, vssx );
   INTCseq_cilao5ah_2( MGM_D0, en, te, vcc, vssx );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, 1'b0, 1'b0, MGM_EN0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cilao5ah_3( clkout, IQ, clk, vcc, vssx );
`else
   INTCseq_cdiar2ah_1( MGM_EN0, clk );
   INTCseq_cilao5ah_2( MGM_D0, en, te );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, 1'b0, 1'b0, MGM_EN0, MGM_D0, notifier );
   INTCseq_cilao5ah_3( clkout, IQ, clk );
`endif

endmodule
`endcelldefine



`celldefine
module b15cilb05ah1n02x3( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n02x3_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n02x3_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n02x3_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n02x3_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb05ah1n02x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n02x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n02x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n02x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n02x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb05ah1n03x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n03x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n03x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n03x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n03x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb05ah1n04x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n04x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n04x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n04x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n04x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb05ah1n06x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n06x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n06x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n06x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n06x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb05ah1n08x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n08x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n08x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n08x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n08x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb05ah1n12x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n12x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n12x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n12x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n12x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb05ah1n16x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n16x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n16x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n16x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n16x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb05ah1n24x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n24x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n24x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n24x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n24x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb05ah1n32x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n32x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n32x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n32x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n32x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb05ah1n48x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n48x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n48x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n48x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n48x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb05ah1n64x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n64x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n64x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n64x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n64x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb05ah1n80x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n80x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n80x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb05ah_func b15cilb05ah1n80x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb05ah_func b15cilb05ah1n80x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-LH
      $setuphold(posedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-LH
      $setuphold(posedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine


primitive INTCseq_cilb81ah_4( MGM_D0, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
  output MGM_D0;
  input en, te;
  `ifdef POWER_AWARE_MODE
  input vcc, vssx;
  `endif

  table
  `ifdef POWER_AWARE_MODE
  //en, te vcc, vssx: MGM_D0
    0  0  1  0: 1;
    1  ?  1  0: 0;
    ?  1  1  0: 0;
  `else
  //en, te: MGM_D0
    0  0: 1;
    1  ?: 0;
    ?  1: 0;
  `endif
  endtable

endprimitive



`celldefine
module INTCseq_cilb81ah_func( clk, clkout, en, te, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te, notifier;
   output clkout;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_EN0, clk, vcc, vssx );
   INTCseq_cilb81ah_4( MGM_D0, en, te, vcc, vssx );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, 1'b0, 1'b0, MGM_EN0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cilao5ah_2( clkout, IQ, clk, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_EN0, clk );
   INTCseq_cilb81ah_4( MGM_D0, en, te );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, 1'b0, 1'b0, MGM_EN0, MGM_D0, notifier );
   INTCseq_cilao5ah_2( clkout, IQ, clk );
`endif

endmodule
`endcelldefine



`celldefine
module b15cilb81ah1n02x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n02x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n02x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n02x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n02x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb81ah1n03x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n03x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n03x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n03x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n03x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb81ah1n04x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n04x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n04x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n04x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n04x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb81ah1n08x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n08x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n08x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n08x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n08x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb81ah1n12x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n12x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n12x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n12x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n12x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb81ah1n16x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n16x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n16x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n16x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n16x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb81ah1n24x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n24x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n24x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n24x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n24x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb81ah1n32x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n32x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n32x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n32x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n32x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15cilb81ah1n64x5( clk, clkout, en, te `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, en, te;
   output clkout;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n64x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n64x5_behav_inst(.clk(clk),.clkout(clkout),.en(en),.te(te),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire en_delay ;
   wire te_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_cilb81ah_func b15cilb81ah1n64x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_cilb81ah_func b15cilb81ah1n64x5_inst(.clk(clk_delay),.clkout(clkout),.en(en_delay),.te(te_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,en_delay);
   not MGM_G1(MGM_W1,te_delay);
   and MGM_G2(ENABLE_NOT_en_AND_NOT_te,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W2,en_delay);
   and MGM_G4(ENABLE_NOT_en_AND_te,te_delay,MGM_W2);
   not MGM_G5(MGM_W3,te_delay);
   and MGM_G6(ENABLE_en_AND_NOT_te,MGM_W3,en_delay);
   and MGM_G7(ENABLE_en_AND_te,te_delay,en_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(en==1'b0 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc negedge clk --> clkout
      (negedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b1 && te==1'b1)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      if(en==1'b0 && te==1'b0)
      // comb arc posedge clk --> clkout
      (posedge clk => (clkout:clk)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_NOT_te == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_en_AND_te == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,negedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold en- clk-HL
      $setuphold(negedge clk,posedge en,0.0,0.0,notifier,,,clk_delay,en_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,negedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      // setuphold te- clk-HL
      $setuphold(negedge clk,posedge te,0.0,0.0,notifier,,,clk_delay,te_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine


primitive INTCseq_fdw003ah_5( MGM_D0, d, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
  output MGM_D0;
  input d, si, ssb;
  `ifdef POWER_AWARE_MODE
  input vcc, vssx;
  `endif

  table
  `ifdef POWER_AWARE_MODE
  //d, si, ssb vcc, vssx: MGM_D0
    1  1  ?  1  0: 1;
    1  ?  1  1  0: 1;
    ?  1  0  1  0: 1;
    0  0  ?  1  0: 0;
    0  ?  1  1  0: 0;
    ?  0  0  1  0: 0;
  `else
  //d, si, ssb: MGM_D0
    1  1  ?: 1;
    1  ?  1: 1;
    ?  1  0: 1;
    0  0  ?: 0;
    0  ?  1: 0;
    ?  0  0: 0;
  `endif
  endtable

endprimitive



`celldefine
module INTCseq_fdw003ah_func( clk, d, o, rb, si, ssb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fdw003ah1n05x5( clk, d, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fdw003ah_func b15fdw003ah1n05x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fdw003ah_func b15fdw003ah1n05x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fdw003ah_func b15fdw003ah1n05x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fdw003ah_func b15fdw003ah1n05x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,rb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,rb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,rb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,rb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,rb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,rb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,rb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,rb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,rb_delay);
   and MGM_G38(ENABLE_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,rb_delay);
   and MGM_G40(ENABLE_rb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   and MGM_G42(MGM_W32,si_delay,MGM_W31);
   not MGM_G43(MGM_W33,ssb_delay);
   and MGM_G44(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W33,MGM_W32);
   not MGM_G45(MGM_W34,si_delay);
   and MGM_G46(MGM_W35,MGM_W34,d_delay);
   and MGM_G47(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G48(MGM_W36,si_delay,d_delay);
   not MGM_G49(MGM_W37,ssb_delay);
   and MGM_G50(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W37,MGM_W36);
   and MGM_G51(MGM_W38,si_delay,d_delay);
   and MGM_G52(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W38);
   not MGM_G53(MGM_W39,clk_delay);
   not MGM_G54(MGM_W40,d_delay);
   and MGM_G55(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G56(MGM_W42,si_delay);
   and MGM_G57(MGM_W43,MGM_W42,MGM_W41);
   not MGM_G58(MGM_W44,ssb_delay);
   and MGM_G59(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W45,clk_delay);
   not MGM_G61(MGM_W46,d_delay);
   and MGM_G62(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G63(MGM_W48,si_delay);
   and MGM_G64(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G65(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G66(MGM_W50,clk_delay);
   not MGM_G67(MGM_W51,d_delay);
   and MGM_G68(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G69(MGM_W53,si_delay,MGM_W52);
   not MGM_G70(MGM_W54,ssb_delay);
   and MGM_G71(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W54,MGM_W53);
   not MGM_G72(MGM_W55,clk_delay);
   not MGM_G73(MGM_W56,d_delay);
   and MGM_G74(MGM_W57,MGM_W56,MGM_W55);
   and MGM_G75(MGM_W58,si_delay,MGM_W57);
   and MGM_G76(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,clk_delay);
   and MGM_G78(MGM_W60,d_delay,MGM_W59);
   not MGM_G79(MGM_W61,si_delay);
   and MGM_G80(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G81(MGM_W63,ssb_delay);
   and MGM_G82(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G83(MGM_W64,clk_delay);
   and MGM_G84(MGM_W65,d_delay,MGM_W64);
   not MGM_G85(MGM_W66,si_delay);
   and MGM_G86(MGM_W67,MGM_W66,MGM_W65);
   and MGM_G87(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W67);
   not MGM_G88(MGM_W68,clk_delay);
   and MGM_G89(MGM_W69,d_delay,MGM_W68);
   and MGM_G90(MGM_W70,si_delay,MGM_W69);
   not MGM_G91(MGM_W71,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W71,MGM_W70);
   not MGM_G93(MGM_W72,clk_delay);
   and MGM_G94(MGM_W73,d_delay,MGM_W72);
   and MGM_G95(MGM_W74,si_delay,MGM_W73);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W74);
   not MGM_G97(MGM_W75,d_delay);
   and MGM_G98(MGM_W76,MGM_W75,clk_delay);
   not MGM_G99(MGM_W77,si_delay);
   and MGM_G100(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G101(MGM_W79,ssb_delay);
   and MGM_G102(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G103(MGM_W80,d_delay);
   and MGM_G104(MGM_W81,MGM_W80,clk_delay);
   not MGM_G105(MGM_W82,si_delay);
   and MGM_G106(MGM_W83,MGM_W82,MGM_W81);
   and MGM_G107(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W83);
   not MGM_G108(MGM_W84,d_delay);
   and MGM_G109(MGM_W85,MGM_W84,clk_delay);
   and MGM_G110(MGM_W86,si_delay,MGM_W85);
   not MGM_G111(MGM_W87,ssb_delay);
   and MGM_G112(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W87,MGM_W86);
   not MGM_G113(MGM_W88,d_delay);
   and MGM_G114(MGM_W89,MGM_W88,clk_delay);
   and MGM_G115(MGM_W90,si_delay,MGM_W89);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W90);
   and MGM_G117(MGM_W91,d_delay,clk_delay);
   not MGM_G118(MGM_W92,si_delay);
   and MGM_G119(MGM_W93,MGM_W92,MGM_W91);
   not MGM_G120(MGM_W94,ssb_delay);
   and MGM_G121(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W94,MGM_W93);
   and MGM_G122(MGM_W95,d_delay,clk_delay);
   not MGM_G123(MGM_W96,si_delay);
   and MGM_G124(MGM_W97,MGM_W96,MGM_W95);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W97);
   and MGM_G126(MGM_W98,d_delay,clk_delay);
   and MGM_G127(MGM_W99,si_delay,MGM_W98);
   not MGM_G128(MGM_W100,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W100,MGM_W99);
   and MGM_G130(MGM_W101,d_delay,clk_delay);
   and MGM_G131(MGM_W102,si_delay,MGM_W101);
   and MGM_G132(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W102);
   not MGM_G133(MGM_W103,d_delay);
   and MGM_G134(MGM_W104,rb_delay,MGM_W103);
   not MGM_G135(MGM_W105,ssb_delay);
   and MGM_G136(ENABLE_NOT_d_AND_rb_AND_NOT_ssb,MGM_W105,MGM_W104);
   and MGM_G137(MGM_W106,rb_delay,d_delay);
   not MGM_G138(MGM_W107,ssb_delay);
   and MGM_G139(ENABLE_d_AND_rb_AND_NOT_ssb,MGM_W107,MGM_W106);
   not MGM_G140(MGM_W108,d_delay);
   and MGM_G141(MGM_W109,rb_delay,MGM_W108);
   and MGM_G142(ENABLE_NOT_d_AND_rb_AND_si,si_delay,MGM_W109);
   and MGM_G143(MGM_W110,rb_delay,d_delay);
   not MGM_G144(MGM_W111,si_delay);
   and MGM_G145(ENABLE_d_AND_rb_AND_NOT_si,MGM_W111,MGM_W110);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fdw003ah1n10x5( clk, d, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fdw003ah_func b15fdw003ah1n10x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fdw003ah_func b15fdw003ah1n10x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fdw003ah_func b15fdw003ah1n10x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fdw003ah_func b15fdw003ah1n10x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,rb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,rb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,rb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,rb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,rb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,rb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,rb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,rb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,rb_delay);
   and MGM_G38(ENABLE_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,rb_delay);
   and MGM_G40(ENABLE_rb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   and MGM_G42(MGM_W32,si_delay,MGM_W31);
   not MGM_G43(MGM_W33,ssb_delay);
   and MGM_G44(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W33,MGM_W32);
   not MGM_G45(MGM_W34,si_delay);
   and MGM_G46(MGM_W35,MGM_W34,d_delay);
   and MGM_G47(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G48(MGM_W36,si_delay,d_delay);
   not MGM_G49(MGM_W37,ssb_delay);
   and MGM_G50(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W37,MGM_W36);
   and MGM_G51(MGM_W38,si_delay,d_delay);
   and MGM_G52(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W38);
   not MGM_G53(MGM_W39,clk_delay);
   not MGM_G54(MGM_W40,d_delay);
   and MGM_G55(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G56(MGM_W42,si_delay);
   and MGM_G57(MGM_W43,MGM_W42,MGM_W41);
   not MGM_G58(MGM_W44,ssb_delay);
   and MGM_G59(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W45,clk_delay);
   not MGM_G61(MGM_W46,d_delay);
   and MGM_G62(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G63(MGM_W48,si_delay);
   and MGM_G64(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G65(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G66(MGM_W50,clk_delay);
   not MGM_G67(MGM_W51,d_delay);
   and MGM_G68(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G69(MGM_W53,si_delay,MGM_W52);
   not MGM_G70(MGM_W54,ssb_delay);
   and MGM_G71(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W54,MGM_W53);
   not MGM_G72(MGM_W55,clk_delay);
   not MGM_G73(MGM_W56,d_delay);
   and MGM_G74(MGM_W57,MGM_W56,MGM_W55);
   and MGM_G75(MGM_W58,si_delay,MGM_W57);
   and MGM_G76(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,clk_delay);
   and MGM_G78(MGM_W60,d_delay,MGM_W59);
   not MGM_G79(MGM_W61,si_delay);
   and MGM_G80(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G81(MGM_W63,ssb_delay);
   and MGM_G82(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G83(MGM_W64,clk_delay);
   and MGM_G84(MGM_W65,d_delay,MGM_W64);
   not MGM_G85(MGM_W66,si_delay);
   and MGM_G86(MGM_W67,MGM_W66,MGM_W65);
   and MGM_G87(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W67);
   not MGM_G88(MGM_W68,clk_delay);
   and MGM_G89(MGM_W69,d_delay,MGM_W68);
   and MGM_G90(MGM_W70,si_delay,MGM_W69);
   not MGM_G91(MGM_W71,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W71,MGM_W70);
   not MGM_G93(MGM_W72,clk_delay);
   and MGM_G94(MGM_W73,d_delay,MGM_W72);
   and MGM_G95(MGM_W74,si_delay,MGM_W73);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W74);
   not MGM_G97(MGM_W75,d_delay);
   and MGM_G98(MGM_W76,MGM_W75,clk_delay);
   not MGM_G99(MGM_W77,si_delay);
   and MGM_G100(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G101(MGM_W79,ssb_delay);
   and MGM_G102(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G103(MGM_W80,d_delay);
   and MGM_G104(MGM_W81,MGM_W80,clk_delay);
   not MGM_G105(MGM_W82,si_delay);
   and MGM_G106(MGM_W83,MGM_W82,MGM_W81);
   and MGM_G107(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W83);
   not MGM_G108(MGM_W84,d_delay);
   and MGM_G109(MGM_W85,MGM_W84,clk_delay);
   and MGM_G110(MGM_W86,si_delay,MGM_W85);
   not MGM_G111(MGM_W87,ssb_delay);
   and MGM_G112(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W87,MGM_W86);
   not MGM_G113(MGM_W88,d_delay);
   and MGM_G114(MGM_W89,MGM_W88,clk_delay);
   and MGM_G115(MGM_W90,si_delay,MGM_W89);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W90);
   and MGM_G117(MGM_W91,d_delay,clk_delay);
   not MGM_G118(MGM_W92,si_delay);
   and MGM_G119(MGM_W93,MGM_W92,MGM_W91);
   not MGM_G120(MGM_W94,ssb_delay);
   and MGM_G121(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W94,MGM_W93);
   and MGM_G122(MGM_W95,d_delay,clk_delay);
   not MGM_G123(MGM_W96,si_delay);
   and MGM_G124(MGM_W97,MGM_W96,MGM_W95);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W97);
   and MGM_G126(MGM_W98,d_delay,clk_delay);
   and MGM_G127(MGM_W99,si_delay,MGM_W98);
   not MGM_G128(MGM_W100,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W100,MGM_W99);
   and MGM_G130(MGM_W101,d_delay,clk_delay);
   and MGM_G131(MGM_W102,si_delay,MGM_W101);
   and MGM_G132(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W102);
   not MGM_G133(MGM_W103,d_delay);
   and MGM_G134(MGM_W104,rb_delay,MGM_W103);
   not MGM_G135(MGM_W105,ssb_delay);
   and MGM_G136(ENABLE_NOT_d_AND_rb_AND_NOT_ssb,MGM_W105,MGM_W104);
   and MGM_G137(MGM_W106,rb_delay,d_delay);
   not MGM_G138(MGM_W107,ssb_delay);
   and MGM_G139(ENABLE_d_AND_rb_AND_NOT_ssb,MGM_W107,MGM_W106);
   not MGM_G140(MGM_W108,d_delay);
   and MGM_G141(MGM_W109,rb_delay,MGM_W108);
   and MGM_G142(ENABLE_NOT_d_AND_rb_AND_si,si_delay,MGM_W109);
   and MGM_G143(MGM_W110,rb_delay,d_delay);
   not MGM_G144(MGM_W111,si_delay);
   and MGM_G145(ENABLE_d_AND_rb_AND_NOT_si,MGM_W111,MGM_W110);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fdw003ah1n20x5( clk, d, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fdw003ah_func b15fdw003ah1n20x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fdw003ah_func b15fdw003ah1n20x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fdw003ah_func b15fdw003ah1n20x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fdw003ah_func b15fdw003ah1n20x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,rb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,rb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,rb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,rb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,rb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,rb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,rb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,rb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,rb_delay);
   and MGM_G38(ENABLE_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,rb_delay);
   and MGM_G40(ENABLE_rb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   and MGM_G42(MGM_W32,si_delay,MGM_W31);
   not MGM_G43(MGM_W33,ssb_delay);
   and MGM_G44(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W33,MGM_W32);
   not MGM_G45(MGM_W34,si_delay);
   and MGM_G46(MGM_W35,MGM_W34,d_delay);
   and MGM_G47(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G48(MGM_W36,si_delay,d_delay);
   not MGM_G49(MGM_W37,ssb_delay);
   and MGM_G50(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W37,MGM_W36);
   and MGM_G51(MGM_W38,si_delay,d_delay);
   and MGM_G52(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W38);
   not MGM_G53(MGM_W39,clk_delay);
   not MGM_G54(MGM_W40,d_delay);
   and MGM_G55(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G56(MGM_W42,si_delay);
   and MGM_G57(MGM_W43,MGM_W42,MGM_W41);
   not MGM_G58(MGM_W44,ssb_delay);
   and MGM_G59(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W45,clk_delay);
   not MGM_G61(MGM_W46,d_delay);
   and MGM_G62(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G63(MGM_W48,si_delay);
   and MGM_G64(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G65(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G66(MGM_W50,clk_delay);
   not MGM_G67(MGM_W51,d_delay);
   and MGM_G68(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G69(MGM_W53,si_delay,MGM_W52);
   not MGM_G70(MGM_W54,ssb_delay);
   and MGM_G71(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W54,MGM_W53);
   not MGM_G72(MGM_W55,clk_delay);
   not MGM_G73(MGM_W56,d_delay);
   and MGM_G74(MGM_W57,MGM_W56,MGM_W55);
   and MGM_G75(MGM_W58,si_delay,MGM_W57);
   and MGM_G76(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,clk_delay);
   and MGM_G78(MGM_W60,d_delay,MGM_W59);
   not MGM_G79(MGM_W61,si_delay);
   and MGM_G80(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G81(MGM_W63,ssb_delay);
   and MGM_G82(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G83(MGM_W64,clk_delay);
   and MGM_G84(MGM_W65,d_delay,MGM_W64);
   not MGM_G85(MGM_W66,si_delay);
   and MGM_G86(MGM_W67,MGM_W66,MGM_W65);
   and MGM_G87(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W67);
   not MGM_G88(MGM_W68,clk_delay);
   and MGM_G89(MGM_W69,d_delay,MGM_W68);
   and MGM_G90(MGM_W70,si_delay,MGM_W69);
   not MGM_G91(MGM_W71,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W71,MGM_W70);
   not MGM_G93(MGM_W72,clk_delay);
   and MGM_G94(MGM_W73,d_delay,MGM_W72);
   and MGM_G95(MGM_W74,si_delay,MGM_W73);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W74);
   not MGM_G97(MGM_W75,d_delay);
   and MGM_G98(MGM_W76,MGM_W75,clk_delay);
   not MGM_G99(MGM_W77,si_delay);
   and MGM_G100(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G101(MGM_W79,ssb_delay);
   and MGM_G102(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G103(MGM_W80,d_delay);
   and MGM_G104(MGM_W81,MGM_W80,clk_delay);
   not MGM_G105(MGM_W82,si_delay);
   and MGM_G106(MGM_W83,MGM_W82,MGM_W81);
   and MGM_G107(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W83);
   not MGM_G108(MGM_W84,d_delay);
   and MGM_G109(MGM_W85,MGM_W84,clk_delay);
   and MGM_G110(MGM_W86,si_delay,MGM_W85);
   not MGM_G111(MGM_W87,ssb_delay);
   and MGM_G112(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W87,MGM_W86);
   not MGM_G113(MGM_W88,d_delay);
   and MGM_G114(MGM_W89,MGM_W88,clk_delay);
   and MGM_G115(MGM_W90,si_delay,MGM_W89);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W90);
   and MGM_G117(MGM_W91,d_delay,clk_delay);
   not MGM_G118(MGM_W92,si_delay);
   and MGM_G119(MGM_W93,MGM_W92,MGM_W91);
   not MGM_G120(MGM_W94,ssb_delay);
   and MGM_G121(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W94,MGM_W93);
   and MGM_G122(MGM_W95,d_delay,clk_delay);
   not MGM_G123(MGM_W96,si_delay);
   and MGM_G124(MGM_W97,MGM_W96,MGM_W95);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W97);
   and MGM_G126(MGM_W98,d_delay,clk_delay);
   and MGM_G127(MGM_W99,si_delay,MGM_W98);
   not MGM_G128(MGM_W100,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W100,MGM_W99);
   and MGM_G130(MGM_W101,d_delay,clk_delay);
   and MGM_G131(MGM_W102,si_delay,MGM_W101);
   and MGM_G132(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W102);
   not MGM_G133(MGM_W103,d_delay);
   and MGM_G134(MGM_W104,rb_delay,MGM_W103);
   not MGM_G135(MGM_W105,ssb_delay);
   and MGM_G136(ENABLE_NOT_d_AND_rb_AND_NOT_ssb,MGM_W105,MGM_W104);
   and MGM_G137(MGM_W106,rb_delay,d_delay);
   not MGM_G138(MGM_W107,ssb_delay);
   and MGM_G139(ENABLE_d_AND_rb_AND_NOT_ssb,MGM_W107,MGM_W106);
   not MGM_G140(MGM_W108,d_delay);
   and MGM_G141(MGM_W109,rb_delay,MGM_W108);
   and MGM_G142(ENABLE_NOT_d_AND_rb_AND_si,si_delay,MGM_W109);
   and MGM_G143(MGM_W110,rb_delay,d_delay);
   not MGM_G144(MGM_W111,si_delay);
   and MGM_G145(ENABLE_d_AND_rb_AND_NOT_si,MGM_W111,MGM_W110);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fdw003ah1n30x5( clk, d, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fdw003ah_func b15fdw003ah1n30x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fdw003ah_func b15fdw003ah1n30x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fdw003ah_func b15fdw003ah1n30x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fdw003ah_func b15fdw003ah1n30x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,rb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,rb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,rb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,rb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,rb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,rb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,rb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,rb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,rb_delay);
   and MGM_G38(ENABLE_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,rb_delay);
   and MGM_G40(ENABLE_rb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   and MGM_G42(MGM_W32,si_delay,MGM_W31);
   not MGM_G43(MGM_W33,ssb_delay);
   and MGM_G44(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W33,MGM_W32);
   not MGM_G45(MGM_W34,si_delay);
   and MGM_G46(MGM_W35,MGM_W34,d_delay);
   and MGM_G47(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G48(MGM_W36,si_delay,d_delay);
   not MGM_G49(MGM_W37,ssb_delay);
   and MGM_G50(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W37,MGM_W36);
   and MGM_G51(MGM_W38,si_delay,d_delay);
   and MGM_G52(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W38);
   not MGM_G53(MGM_W39,clk_delay);
   not MGM_G54(MGM_W40,d_delay);
   and MGM_G55(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G56(MGM_W42,si_delay);
   and MGM_G57(MGM_W43,MGM_W42,MGM_W41);
   not MGM_G58(MGM_W44,ssb_delay);
   and MGM_G59(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W45,clk_delay);
   not MGM_G61(MGM_W46,d_delay);
   and MGM_G62(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G63(MGM_W48,si_delay);
   and MGM_G64(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G65(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G66(MGM_W50,clk_delay);
   not MGM_G67(MGM_W51,d_delay);
   and MGM_G68(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G69(MGM_W53,si_delay,MGM_W52);
   not MGM_G70(MGM_W54,ssb_delay);
   and MGM_G71(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W54,MGM_W53);
   not MGM_G72(MGM_W55,clk_delay);
   not MGM_G73(MGM_W56,d_delay);
   and MGM_G74(MGM_W57,MGM_W56,MGM_W55);
   and MGM_G75(MGM_W58,si_delay,MGM_W57);
   and MGM_G76(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,clk_delay);
   and MGM_G78(MGM_W60,d_delay,MGM_W59);
   not MGM_G79(MGM_W61,si_delay);
   and MGM_G80(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G81(MGM_W63,ssb_delay);
   and MGM_G82(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G83(MGM_W64,clk_delay);
   and MGM_G84(MGM_W65,d_delay,MGM_W64);
   not MGM_G85(MGM_W66,si_delay);
   and MGM_G86(MGM_W67,MGM_W66,MGM_W65);
   and MGM_G87(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W67);
   not MGM_G88(MGM_W68,clk_delay);
   and MGM_G89(MGM_W69,d_delay,MGM_W68);
   and MGM_G90(MGM_W70,si_delay,MGM_W69);
   not MGM_G91(MGM_W71,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W71,MGM_W70);
   not MGM_G93(MGM_W72,clk_delay);
   and MGM_G94(MGM_W73,d_delay,MGM_W72);
   and MGM_G95(MGM_W74,si_delay,MGM_W73);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W74);
   not MGM_G97(MGM_W75,d_delay);
   and MGM_G98(MGM_W76,MGM_W75,clk_delay);
   not MGM_G99(MGM_W77,si_delay);
   and MGM_G100(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G101(MGM_W79,ssb_delay);
   and MGM_G102(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G103(MGM_W80,d_delay);
   and MGM_G104(MGM_W81,MGM_W80,clk_delay);
   not MGM_G105(MGM_W82,si_delay);
   and MGM_G106(MGM_W83,MGM_W82,MGM_W81);
   and MGM_G107(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W83);
   not MGM_G108(MGM_W84,d_delay);
   and MGM_G109(MGM_W85,MGM_W84,clk_delay);
   and MGM_G110(MGM_W86,si_delay,MGM_W85);
   not MGM_G111(MGM_W87,ssb_delay);
   and MGM_G112(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W87,MGM_W86);
   not MGM_G113(MGM_W88,d_delay);
   and MGM_G114(MGM_W89,MGM_W88,clk_delay);
   and MGM_G115(MGM_W90,si_delay,MGM_W89);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W90);
   and MGM_G117(MGM_W91,d_delay,clk_delay);
   not MGM_G118(MGM_W92,si_delay);
   and MGM_G119(MGM_W93,MGM_W92,MGM_W91);
   not MGM_G120(MGM_W94,ssb_delay);
   and MGM_G121(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W94,MGM_W93);
   and MGM_G122(MGM_W95,d_delay,clk_delay);
   not MGM_G123(MGM_W96,si_delay);
   and MGM_G124(MGM_W97,MGM_W96,MGM_W95);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W97);
   and MGM_G126(MGM_W98,d_delay,clk_delay);
   and MGM_G127(MGM_W99,si_delay,MGM_W98);
   not MGM_G128(MGM_W100,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W100,MGM_W99);
   and MGM_G130(MGM_W101,d_delay,clk_delay);
   and MGM_G131(MGM_W102,si_delay,MGM_W101);
   and MGM_G132(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W102);
   not MGM_G133(MGM_W103,d_delay);
   and MGM_G134(MGM_W104,rb_delay,MGM_W103);
   not MGM_G135(MGM_W105,ssb_delay);
   and MGM_G136(ENABLE_NOT_d_AND_rb_AND_NOT_ssb,MGM_W105,MGM_W104);
   and MGM_G137(MGM_W106,rb_delay,d_delay);
   not MGM_G138(MGM_W107,ssb_delay);
   and MGM_G139(ENABLE_d_AND_rb_AND_NOT_ssb,MGM_W107,MGM_W106);
   not MGM_G140(MGM_W108,d_delay);
   and MGM_G141(MGM_W109,rb_delay,MGM_W108);
   and MGM_G142(ENABLE_NOT_d_AND_rb_AND_si,si_delay,MGM_W109);
   and MGM_G143(MGM_W110,rb_delay,d_delay);
   not MGM_G144(MGM_W111,si_delay);
   and MGM_G145(ENABLE_d_AND_rb_AND_NOT_si,MGM_W111,MGM_W110);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fhw000ah_func( clk, d, o, si, ssb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fhw000ah1n05x5( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fhw000ah_func b15fhw000ah1n05x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fhw000ah_func b15fhw000ah1n05x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fhw000ah_func b15fhw000ah1n05x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fhw000ah_func b15fhw000ah1n05x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fhw000ah1n10x5( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fhw000ah_func b15fhw000ah1n10x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fhw000ah_func b15fhw000ah1n10x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fhw000ah_func b15fhw000ah1n10x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fhw000ah_func b15fhw000ah1n10x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fhw000ah1n20x5( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fhw000ah_func b15fhw000ah1n20x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fhw000ah_func b15fhw000ah1n20x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fhw000ah_func b15fhw000ah1n20x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fhw000ah_func b15fhw000ah1n20x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fhw000ah1n30x5( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fhw000ah_func b15fhw000ah1n30x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fhw000ah_func b15fhw000ah1n30x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fhw000ah_func b15fhw000ah1n30x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fhw000ah_func b15fhw000ah1n30x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fmm200ah_func( clk, d, o, si, ssb, notifier, notifier0 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb, notifier, notifier0;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, 1'b0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier0 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D1, IQ1, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, 1'b0, 1'b0, MGM_CLK1, MGM_D1, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ2, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, 1'b0, 1'b0, MGM_CLK0, MGM_D0, notifier0 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk );
   INTCseq_cdiar2ah_0( MGM_D1, IQ1 );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, 1'b0, 1'b0, MGM_CLK1, MGM_D1, notifier );
   INTCseq_cdiar2ah_0( o, IQ2 );
`endif

endmodule
`endcelldefine



`celldefine
module b15fmm200ah1n04x5( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fmm200ah_func b15fmm200ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.notifier0(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fmm200ah_func b15fmm200ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.notifier0(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   reg notifier0;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fmm200ah_func b15fmm200ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.notifier0(notifier0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fmm200ah_func b15fmm200ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.notifier0(notifier0));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fmm203ah_func( clk, d, o, rb, si, ssb, notifier, notifier0 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb, notifier, notifier0;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier0 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C1, rb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D1, IQ1, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, MGM_C1, 1'b0, MGM_CLK1, MGM_D1, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ2, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, notifier0 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk );
   INTCseq_cdiar2ah_1( MGM_C1, rb );
   INTCseq_cdiar2ah_0( MGM_D1, IQ1 );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, MGM_C1, 1'b0, MGM_CLK1, MGM_D1, notifier );
   INTCseq_cdiar2ah_0( o, IQ2 );
`endif

endmodule
`endcelldefine



`celldefine
module b15fmm203ah1n04x5( clk, d, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fmm203ah_func b15fmm203ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.notifier0(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fmm203ah_func b15fmm203ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.notifier0(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   reg notifier0;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fmm203ah_func b15fmm203ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.notifier0(notifier0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fmm203ah_func b15fmm203ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.notifier0(notifier0));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,rb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,rb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,rb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,rb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,rb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,rb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,rb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,rb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,rb_delay);
   and MGM_G38(ENABLE_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,rb_delay);
   and MGM_G40(ENABLE_rb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   and MGM_G42(MGM_W32,si_delay,MGM_W31);
   not MGM_G43(MGM_W33,ssb_delay);
   and MGM_G44(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W33,MGM_W32);
   not MGM_G45(MGM_W34,si_delay);
   and MGM_G46(MGM_W35,MGM_W34,d_delay);
   and MGM_G47(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G48(MGM_W36,si_delay,d_delay);
   not MGM_G49(MGM_W37,ssb_delay);
   and MGM_G50(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W37,MGM_W36);
   and MGM_G51(MGM_W38,si_delay,d_delay);
   and MGM_G52(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W38);
   not MGM_G53(MGM_W39,clk_delay);
   not MGM_G54(MGM_W40,d_delay);
   and MGM_G55(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G56(MGM_W42,si_delay);
   and MGM_G57(MGM_W43,MGM_W42,MGM_W41);
   not MGM_G58(MGM_W44,ssb_delay);
   and MGM_G59(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W45,clk_delay);
   not MGM_G61(MGM_W46,d_delay);
   and MGM_G62(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G63(MGM_W48,si_delay);
   and MGM_G64(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G65(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G66(MGM_W50,clk_delay);
   not MGM_G67(MGM_W51,d_delay);
   and MGM_G68(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G69(MGM_W53,si_delay,MGM_W52);
   not MGM_G70(MGM_W54,ssb_delay);
   and MGM_G71(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W54,MGM_W53);
   not MGM_G72(MGM_W55,clk_delay);
   not MGM_G73(MGM_W56,d_delay);
   and MGM_G74(MGM_W57,MGM_W56,MGM_W55);
   and MGM_G75(MGM_W58,si_delay,MGM_W57);
   and MGM_G76(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,clk_delay);
   and MGM_G78(MGM_W60,d_delay,MGM_W59);
   not MGM_G79(MGM_W61,si_delay);
   and MGM_G80(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G81(MGM_W63,ssb_delay);
   and MGM_G82(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G83(MGM_W64,clk_delay);
   and MGM_G84(MGM_W65,d_delay,MGM_W64);
   not MGM_G85(MGM_W66,si_delay);
   and MGM_G86(MGM_W67,MGM_W66,MGM_W65);
   and MGM_G87(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W67);
   not MGM_G88(MGM_W68,clk_delay);
   and MGM_G89(MGM_W69,d_delay,MGM_W68);
   and MGM_G90(MGM_W70,si_delay,MGM_W69);
   not MGM_G91(MGM_W71,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W71,MGM_W70);
   not MGM_G93(MGM_W72,clk_delay);
   and MGM_G94(MGM_W73,d_delay,MGM_W72);
   and MGM_G95(MGM_W74,si_delay,MGM_W73);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W74);
   not MGM_G97(MGM_W75,d_delay);
   and MGM_G98(MGM_W76,MGM_W75,clk_delay);
   not MGM_G99(MGM_W77,si_delay);
   and MGM_G100(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G101(MGM_W79,ssb_delay);
   and MGM_G102(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G103(MGM_W80,d_delay);
   and MGM_G104(MGM_W81,MGM_W80,clk_delay);
   not MGM_G105(MGM_W82,si_delay);
   and MGM_G106(MGM_W83,MGM_W82,MGM_W81);
   and MGM_G107(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W83);
   not MGM_G108(MGM_W84,d_delay);
   and MGM_G109(MGM_W85,MGM_W84,clk_delay);
   and MGM_G110(MGM_W86,si_delay,MGM_W85);
   not MGM_G111(MGM_W87,ssb_delay);
   and MGM_G112(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W87,MGM_W86);
   not MGM_G113(MGM_W88,d_delay);
   and MGM_G114(MGM_W89,MGM_W88,clk_delay);
   and MGM_G115(MGM_W90,si_delay,MGM_W89);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W90);
   and MGM_G117(MGM_W91,d_delay,clk_delay);
   not MGM_G118(MGM_W92,si_delay);
   and MGM_G119(MGM_W93,MGM_W92,MGM_W91);
   not MGM_G120(MGM_W94,ssb_delay);
   and MGM_G121(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W94,MGM_W93);
   and MGM_G122(MGM_W95,d_delay,clk_delay);
   not MGM_G123(MGM_W96,si_delay);
   and MGM_G124(MGM_W97,MGM_W96,MGM_W95);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W97);
   and MGM_G126(MGM_W98,d_delay,clk_delay);
   and MGM_G127(MGM_W99,si_delay,MGM_W98);
   not MGM_G128(MGM_W100,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W100,MGM_W99);
   and MGM_G130(MGM_W101,d_delay,clk_delay);
   and MGM_G131(MGM_W102,si_delay,MGM_W101);
   and MGM_G132(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W102);
   not MGM_G133(MGM_W103,d_delay);
   and MGM_G134(MGM_W104,rb_delay,MGM_W103);
   not MGM_G135(MGM_W105,ssb_delay);
   and MGM_G136(ENABLE_NOT_d_AND_rb_AND_NOT_ssb,MGM_W105,MGM_W104);
   and MGM_G137(MGM_W106,rb_delay,d_delay);
   not MGM_G138(MGM_W107,ssb_delay);
   and MGM_G139(ENABLE_d_AND_rb_AND_NOT_ssb,MGM_W107,MGM_W106);
   not MGM_G140(MGM_W108,d_delay);
   and MGM_G141(MGM_W109,rb_delay,MGM_W108);
   and MGM_G142(ENABLE_NOT_d_AND_rb_AND_si,si_delay,MGM_W109);
   and MGM_G143(MGM_W110,rb_delay,d_delay);
   not MGM_G144(MGM_W111,si_delay);
   and MGM_G145(ENABLE_d_AND_rb_AND_NOT_si,MGM_W111,MGM_W110);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fmm20cah_func( clk, d, o, psb, si, ssb, notifier, notifier0 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, si, ssb, notifier, notifier0;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_P0, psb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, 1'b0, MGM_P0, MGM_CLK0, MGM_D0, vcc, vssx, notifier0 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_P1, psb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D1, IQ1, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, 1'b0, MGM_P1, MGM_CLK1, MGM_D1, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ2, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_P0, psb );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, 1'b0, MGM_P0, MGM_CLK0, MGM_D0, notifier0 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk );
   INTCseq_cdiar2ah_1( MGM_P1, psb );
   INTCseq_cdiar2ah_0( MGM_D1, IQ1 );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, 1'b0, MGM_P1, MGM_CLK1, MGM_D1, notifier );
   INTCseq_cdiar2ah_0( o, IQ2 );
`endif

endmodule
`endcelldefine



`celldefine
module b15fmm20cah1n04x5( clk, d, o, psb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fmm20cah_func b15fmm20cah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0),.notifier0(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fmm20cah_func b15fmm20cah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0),.notifier0(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   reg notifier0;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fmm20cah_func b15fmm20cah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.notifier0(notifier0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fmm20cah_func b15fmm20cah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.notifier0(notifier0));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,psb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,psb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,psb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,psb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,psb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,psb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,psb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,psb_delay);
   and MGM_G38(ENABLE_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,psb_delay);
   and MGM_G40(ENABLE_psb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   not MGM_G42(MGM_W32,si_delay);
   and MGM_G43(MGM_W33,MGM_W32,MGM_W31);
   not MGM_G44(MGM_W34,ssb_delay);
   and MGM_G45(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W34,MGM_W33);
   not MGM_G46(MGM_W35,d_delay);
   not MGM_G47(MGM_W36,si_delay);
   and MGM_G48(MGM_W37,MGM_W36,MGM_W35);
   and MGM_G49(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W37);
   not MGM_G50(MGM_W38,d_delay);
   and MGM_G51(MGM_W39,si_delay,MGM_W38);
   and MGM_G52(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W39);
   not MGM_G53(MGM_W40,si_delay);
   and MGM_G54(MGM_W41,MGM_W40,d_delay);
   not MGM_G55(MGM_W42,ssb_delay);
   and MGM_G56(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W42,MGM_W41);
   not MGM_G57(MGM_W43,clk_delay);
   not MGM_G58(MGM_W44,d_delay);
   and MGM_G59(MGM_W45,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W46,si_delay);
   and MGM_G61(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G62(MGM_W48,ssb_delay);
   and MGM_G63(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   not MGM_G64(MGM_W49,clk_delay);
   not MGM_G65(MGM_W50,d_delay);
   and MGM_G66(MGM_W51,MGM_W50,MGM_W49);
   not MGM_G67(MGM_W52,si_delay);
   and MGM_G68(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G69(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G70(MGM_W54,clk_delay);
   not MGM_G71(MGM_W55,d_delay);
   and MGM_G72(MGM_W56,MGM_W55,MGM_W54);
   and MGM_G73(MGM_W57,si_delay,MGM_W56);
   not MGM_G74(MGM_W58,ssb_delay);
   and MGM_G75(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W58,MGM_W57);
   not MGM_G76(MGM_W59,clk_delay);
   not MGM_G77(MGM_W60,d_delay);
   and MGM_G78(MGM_W61,MGM_W60,MGM_W59);
   and MGM_G79(MGM_W62,si_delay,MGM_W61);
   and MGM_G80(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W62);
   not MGM_G81(MGM_W63,clk_delay);
   and MGM_G82(MGM_W64,d_delay,MGM_W63);
   not MGM_G83(MGM_W65,si_delay);
   and MGM_G84(MGM_W66,MGM_W65,MGM_W64);
   not MGM_G85(MGM_W67,ssb_delay);
   and MGM_G86(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W67,MGM_W66);
   not MGM_G87(MGM_W68,clk_delay);
   and MGM_G88(MGM_W69,d_delay,MGM_W68);
   not MGM_G89(MGM_W70,si_delay);
   and MGM_G90(MGM_W71,MGM_W70,MGM_W69);
   and MGM_G91(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W71);
   not MGM_G92(MGM_W72,clk_delay);
   and MGM_G93(MGM_W73,d_delay,MGM_W72);
   and MGM_G94(MGM_W74,si_delay,MGM_W73);
   not MGM_G95(MGM_W75,ssb_delay);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G97(MGM_W76,clk_delay);
   and MGM_G98(MGM_W77,d_delay,MGM_W76);
   and MGM_G99(MGM_W78,si_delay,MGM_W77);
   and MGM_G100(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W78);
   not MGM_G101(MGM_W79,d_delay);
   and MGM_G102(MGM_W80,MGM_W79,clk_delay);
   not MGM_G103(MGM_W81,si_delay);
   and MGM_G104(MGM_W82,MGM_W81,MGM_W80);
   not MGM_G105(MGM_W83,ssb_delay);
   and MGM_G106(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W83,MGM_W82);
   not MGM_G107(MGM_W84,d_delay);
   and MGM_G108(MGM_W85,MGM_W84,clk_delay);
   not MGM_G109(MGM_W86,si_delay);
   and MGM_G110(MGM_W87,MGM_W86,MGM_W85);
   and MGM_G111(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W87);
   not MGM_G112(MGM_W88,d_delay);
   and MGM_G113(MGM_W89,MGM_W88,clk_delay);
   and MGM_G114(MGM_W90,si_delay,MGM_W89);
   not MGM_G115(MGM_W91,ssb_delay);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W91,MGM_W90);
   not MGM_G117(MGM_W92,d_delay);
   and MGM_G118(MGM_W93,MGM_W92,clk_delay);
   and MGM_G119(MGM_W94,si_delay,MGM_W93);
   and MGM_G120(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W94);
   and MGM_G121(MGM_W95,d_delay,clk_delay);
   not MGM_G122(MGM_W96,si_delay);
   and MGM_G123(MGM_W97,MGM_W96,MGM_W95);
   not MGM_G124(MGM_W98,ssb_delay);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W98,MGM_W97);
   and MGM_G126(MGM_W99,d_delay,clk_delay);
   not MGM_G127(MGM_W100,si_delay);
   and MGM_G128(MGM_W101,MGM_W100,MGM_W99);
   and MGM_G129(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W101);
   and MGM_G130(MGM_W102,d_delay,clk_delay);
   and MGM_G131(MGM_W103,si_delay,MGM_W102);
   not MGM_G132(MGM_W104,ssb_delay);
   and MGM_G133(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W104,MGM_W103);
   and MGM_G134(MGM_W105,d_delay,clk_delay);
   and MGM_G135(MGM_W106,si_delay,MGM_W105);
   and MGM_G136(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W106);
   not MGM_G137(MGM_W107,d_delay);
   and MGM_G138(MGM_W108,psb_delay,MGM_W107);
   not MGM_G139(MGM_W109,ssb_delay);
   and MGM_G140(ENABLE_NOT_d_AND_psb_AND_NOT_ssb,MGM_W109,MGM_W108);
   and MGM_G141(MGM_W110,psb_delay,d_delay);
   not MGM_G142(MGM_W111,ssb_delay);
   and MGM_G143(ENABLE_d_AND_psb_AND_NOT_ssb,MGM_W111,MGM_W110);
   not MGM_G144(MGM_W112,d_delay);
   and MGM_G145(MGM_W113,psb_delay,MGM_W112);
   and MGM_G146(ENABLE_NOT_d_AND_psb_AND_si,si_delay,MGM_W113);
   and MGM_G147(MGM_W114,psb_delay,d_delay);
   not MGM_G148(MGM_W115,si_delay);
   and MGM_G149(ENABLE_d_AND_psb_AND_NOT_si,MGM_W115,MGM_W114);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fmm300ah_func( clk, d, o, si, ssb, notifier, notifier0 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb, notifier, notifier0;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, 1'b0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier0 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D1, IQ1, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, 1'b0, 1'b0, MGM_CLK1, MGM_D1, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( MGM_CLK2, clk, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D2, IQ2, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ3, 1'b0, 1'b0, MGM_CLK2, MGM_D2, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ3, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, 1'b0, 1'b0, MGM_CLK0, MGM_D0, notifier0 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk );
   INTCseq_cdiar2ah_0( MGM_D1, IQ1 );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, 1'b0, 1'b0, MGM_CLK1, MGM_D1, notifier );
   INTCseq_cdiar2ah_0( MGM_CLK2, clk );
   INTCseq_cdiar2ah_0( MGM_D2, IQ2 );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ3, 1'b0, 1'b0, MGM_CLK2, MGM_D2, notifier );
   INTCseq_cdiar2ah_0( o, IQ3 );
`endif

endmodule
`endcelldefine



`celldefine
module b15fmm300ah1n04x5( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fmm300ah_func b15fmm300ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.notifier0(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fmm300ah_func b15fmm300ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.notifier0(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   reg notifier0;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fmm300ah_func b15fmm300ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.notifier0(notifier0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fmm300ah_func b15fmm300ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.notifier0(notifier0));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fmm303ah_func( clk, d, o, rb, si, ssb, notifier, notifier0 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb, notifier, notifier0;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier0 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C1, rb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D1, IQ1, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, MGM_C1, 1'b0, MGM_CLK1, MGM_D1, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( MGM_CLK2, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C2, rb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D2, IQ2, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ3, MGM_C2, 1'b0, MGM_CLK2, MGM_D2, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ3, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, notifier0 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk );
   INTCseq_cdiar2ah_1( MGM_C1, rb );
   INTCseq_cdiar2ah_0( MGM_D1, IQ1 );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, MGM_C1, 1'b0, MGM_CLK1, MGM_D1, notifier );
   INTCseq_cdiar2ah_0( MGM_CLK2, clk );
   INTCseq_cdiar2ah_1( MGM_C2, rb );
   INTCseq_cdiar2ah_0( MGM_D2, IQ2 );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ3, MGM_C2, 1'b0, MGM_CLK2, MGM_D2, notifier );
   INTCseq_cdiar2ah_0( o, IQ3 );
`endif

endmodule
`endcelldefine



`celldefine
module b15fmm303ah1n04x5( clk, d, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fmm303ah_func b15fmm303ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.notifier0(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fmm303ah_func b15fmm303ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.notifier0(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   reg notifier0;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fmm303ah_func b15fmm303ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.notifier0(notifier0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fmm303ah_func b15fmm303ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.notifier0(notifier0));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,rb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,rb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,rb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,rb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,rb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,rb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,rb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,rb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,rb_delay);
   and MGM_G38(ENABLE_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,rb_delay);
   and MGM_G40(ENABLE_rb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   and MGM_G42(MGM_W32,si_delay,MGM_W31);
   not MGM_G43(MGM_W33,ssb_delay);
   and MGM_G44(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W33,MGM_W32);
   not MGM_G45(MGM_W34,si_delay);
   and MGM_G46(MGM_W35,MGM_W34,d_delay);
   and MGM_G47(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G48(MGM_W36,si_delay,d_delay);
   not MGM_G49(MGM_W37,ssb_delay);
   and MGM_G50(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W37,MGM_W36);
   and MGM_G51(MGM_W38,si_delay,d_delay);
   and MGM_G52(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W38);
   not MGM_G53(MGM_W39,clk_delay);
   not MGM_G54(MGM_W40,d_delay);
   and MGM_G55(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G56(MGM_W42,si_delay);
   and MGM_G57(MGM_W43,MGM_W42,MGM_W41);
   not MGM_G58(MGM_W44,ssb_delay);
   and MGM_G59(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W45,clk_delay);
   not MGM_G61(MGM_W46,d_delay);
   and MGM_G62(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G63(MGM_W48,si_delay);
   and MGM_G64(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G65(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G66(MGM_W50,clk_delay);
   not MGM_G67(MGM_W51,d_delay);
   and MGM_G68(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G69(MGM_W53,si_delay,MGM_W52);
   not MGM_G70(MGM_W54,ssb_delay);
   and MGM_G71(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W54,MGM_W53);
   not MGM_G72(MGM_W55,clk_delay);
   not MGM_G73(MGM_W56,d_delay);
   and MGM_G74(MGM_W57,MGM_W56,MGM_W55);
   and MGM_G75(MGM_W58,si_delay,MGM_W57);
   and MGM_G76(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,clk_delay);
   and MGM_G78(MGM_W60,d_delay,MGM_W59);
   not MGM_G79(MGM_W61,si_delay);
   and MGM_G80(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G81(MGM_W63,ssb_delay);
   and MGM_G82(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G83(MGM_W64,clk_delay);
   and MGM_G84(MGM_W65,d_delay,MGM_W64);
   not MGM_G85(MGM_W66,si_delay);
   and MGM_G86(MGM_W67,MGM_W66,MGM_W65);
   and MGM_G87(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W67);
   not MGM_G88(MGM_W68,clk_delay);
   and MGM_G89(MGM_W69,d_delay,MGM_W68);
   and MGM_G90(MGM_W70,si_delay,MGM_W69);
   not MGM_G91(MGM_W71,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W71,MGM_W70);
   not MGM_G93(MGM_W72,clk_delay);
   and MGM_G94(MGM_W73,d_delay,MGM_W72);
   and MGM_G95(MGM_W74,si_delay,MGM_W73);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W74);
   not MGM_G97(MGM_W75,d_delay);
   and MGM_G98(MGM_W76,MGM_W75,clk_delay);
   not MGM_G99(MGM_W77,si_delay);
   and MGM_G100(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G101(MGM_W79,ssb_delay);
   and MGM_G102(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G103(MGM_W80,d_delay);
   and MGM_G104(MGM_W81,MGM_W80,clk_delay);
   not MGM_G105(MGM_W82,si_delay);
   and MGM_G106(MGM_W83,MGM_W82,MGM_W81);
   and MGM_G107(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W83);
   not MGM_G108(MGM_W84,d_delay);
   and MGM_G109(MGM_W85,MGM_W84,clk_delay);
   and MGM_G110(MGM_W86,si_delay,MGM_W85);
   not MGM_G111(MGM_W87,ssb_delay);
   and MGM_G112(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W87,MGM_W86);
   not MGM_G113(MGM_W88,d_delay);
   and MGM_G114(MGM_W89,MGM_W88,clk_delay);
   and MGM_G115(MGM_W90,si_delay,MGM_W89);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W90);
   and MGM_G117(MGM_W91,d_delay,clk_delay);
   not MGM_G118(MGM_W92,si_delay);
   and MGM_G119(MGM_W93,MGM_W92,MGM_W91);
   not MGM_G120(MGM_W94,ssb_delay);
   and MGM_G121(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W94,MGM_W93);
   and MGM_G122(MGM_W95,d_delay,clk_delay);
   not MGM_G123(MGM_W96,si_delay);
   and MGM_G124(MGM_W97,MGM_W96,MGM_W95);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W97);
   and MGM_G126(MGM_W98,d_delay,clk_delay);
   and MGM_G127(MGM_W99,si_delay,MGM_W98);
   not MGM_G128(MGM_W100,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W100,MGM_W99);
   and MGM_G130(MGM_W101,d_delay,clk_delay);
   and MGM_G131(MGM_W102,si_delay,MGM_W101);
   and MGM_G132(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W102);
   not MGM_G133(MGM_W103,d_delay);
   and MGM_G134(MGM_W104,rb_delay,MGM_W103);
   not MGM_G135(MGM_W105,ssb_delay);
   and MGM_G136(ENABLE_NOT_d_AND_rb_AND_NOT_ssb,MGM_W105,MGM_W104);
   and MGM_G137(MGM_W106,rb_delay,d_delay);
   not MGM_G138(MGM_W107,ssb_delay);
   and MGM_G139(ENABLE_d_AND_rb_AND_NOT_ssb,MGM_W107,MGM_W106);
   not MGM_G140(MGM_W108,d_delay);
   and MGM_G141(MGM_W109,rb_delay,MGM_W108);
   and MGM_G142(ENABLE_NOT_d_AND_rb_AND_si,si_delay,MGM_W109);
   and MGM_G143(MGM_W110,rb_delay,d_delay);
   not MGM_G144(MGM_W111,si_delay);
   and MGM_G145(ENABLE_d_AND_rb_AND_NOT_si,MGM_W111,MGM_W110);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fmm30cah_func( clk, d, o, psb, si, ssb, notifier, notifier0 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, si, ssb, notifier, notifier0;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_P0, psb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, 1'b0, MGM_P0, MGM_CLK0, MGM_D0, vcc, vssx, notifier0 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_P1, psb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D1, IQ1, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, 1'b0, MGM_P1, MGM_CLK1, MGM_D1, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( MGM_CLK2, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_P2, psb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D2, IQ2, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ3, 1'b0, MGM_P2, MGM_CLK2, MGM_D2, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ3, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_P0, psb );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, 1'b0, MGM_P0, MGM_CLK0, MGM_D0, notifier0 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk );
   INTCseq_cdiar2ah_1( MGM_P1, psb );
   INTCseq_cdiar2ah_0( MGM_D1, IQ1 );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, 1'b0, MGM_P1, MGM_CLK1, MGM_D1, notifier );
   INTCseq_cdiar2ah_0( MGM_CLK2, clk );
   INTCseq_cdiar2ah_1( MGM_P2, psb );
   INTCseq_cdiar2ah_0( MGM_D2, IQ2 );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ3, 1'b0, MGM_P2, MGM_CLK2, MGM_D2, notifier );
   INTCseq_cdiar2ah_0( o, IQ3 );
`endif

endmodule
`endcelldefine



`celldefine
module b15fmm30cah1n04x5( clk, d, o, psb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fmm30cah_func b15fmm30cah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0),.notifier0(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fmm30cah_func b15fmm30cah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0),.notifier0(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   reg notifier0;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fmm30cah_func b15fmm30cah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.notifier0(notifier0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fmm30cah_func b15fmm30cah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.notifier0(notifier0));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,psb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,psb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,psb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,psb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,psb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,psb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,psb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,psb_delay);
   and MGM_G38(ENABLE_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,psb_delay);
   and MGM_G40(ENABLE_psb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   not MGM_G42(MGM_W32,si_delay);
   and MGM_G43(MGM_W33,MGM_W32,MGM_W31);
   not MGM_G44(MGM_W34,ssb_delay);
   and MGM_G45(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W34,MGM_W33);
   not MGM_G46(MGM_W35,d_delay);
   not MGM_G47(MGM_W36,si_delay);
   and MGM_G48(MGM_W37,MGM_W36,MGM_W35);
   and MGM_G49(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W37);
   not MGM_G50(MGM_W38,d_delay);
   and MGM_G51(MGM_W39,si_delay,MGM_W38);
   and MGM_G52(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W39);
   not MGM_G53(MGM_W40,si_delay);
   and MGM_G54(MGM_W41,MGM_W40,d_delay);
   not MGM_G55(MGM_W42,ssb_delay);
   and MGM_G56(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W42,MGM_W41);
   not MGM_G57(MGM_W43,clk_delay);
   not MGM_G58(MGM_W44,d_delay);
   and MGM_G59(MGM_W45,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W46,si_delay);
   and MGM_G61(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G62(MGM_W48,ssb_delay);
   and MGM_G63(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   not MGM_G64(MGM_W49,clk_delay);
   not MGM_G65(MGM_W50,d_delay);
   and MGM_G66(MGM_W51,MGM_W50,MGM_W49);
   not MGM_G67(MGM_W52,si_delay);
   and MGM_G68(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G69(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G70(MGM_W54,clk_delay);
   not MGM_G71(MGM_W55,d_delay);
   and MGM_G72(MGM_W56,MGM_W55,MGM_W54);
   and MGM_G73(MGM_W57,si_delay,MGM_W56);
   not MGM_G74(MGM_W58,ssb_delay);
   and MGM_G75(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W58,MGM_W57);
   not MGM_G76(MGM_W59,clk_delay);
   not MGM_G77(MGM_W60,d_delay);
   and MGM_G78(MGM_W61,MGM_W60,MGM_W59);
   and MGM_G79(MGM_W62,si_delay,MGM_W61);
   and MGM_G80(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W62);
   not MGM_G81(MGM_W63,clk_delay);
   and MGM_G82(MGM_W64,d_delay,MGM_W63);
   not MGM_G83(MGM_W65,si_delay);
   and MGM_G84(MGM_W66,MGM_W65,MGM_W64);
   not MGM_G85(MGM_W67,ssb_delay);
   and MGM_G86(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W67,MGM_W66);
   not MGM_G87(MGM_W68,clk_delay);
   and MGM_G88(MGM_W69,d_delay,MGM_W68);
   not MGM_G89(MGM_W70,si_delay);
   and MGM_G90(MGM_W71,MGM_W70,MGM_W69);
   and MGM_G91(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W71);
   not MGM_G92(MGM_W72,clk_delay);
   and MGM_G93(MGM_W73,d_delay,MGM_W72);
   and MGM_G94(MGM_W74,si_delay,MGM_W73);
   not MGM_G95(MGM_W75,ssb_delay);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G97(MGM_W76,clk_delay);
   and MGM_G98(MGM_W77,d_delay,MGM_W76);
   and MGM_G99(MGM_W78,si_delay,MGM_W77);
   and MGM_G100(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W78);
   not MGM_G101(MGM_W79,d_delay);
   and MGM_G102(MGM_W80,MGM_W79,clk_delay);
   not MGM_G103(MGM_W81,si_delay);
   and MGM_G104(MGM_W82,MGM_W81,MGM_W80);
   not MGM_G105(MGM_W83,ssb_delay);
   and MGM_G106(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W83,MGM_W82);
   not MGM_G107(MGM_W84,d_delay);
   and MGM_G108(MGM_W85,MGM_W84,clk_delay);
   not MGM_G109(MGM_W86,si_delay);
   and MGM_G110(MGM_W87,MGM_W86,MGM_W85);
   and MGM_G111(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W87);
   not MGM_G112(MGM_W88,d_delay);
   and MGM_G113(MGM_W89,MGM_W88,clk_delay);
   and MGM_G114(MGM_W90,si_delay,MGM_W89);
   not MGM_G115(MGM_W91,ssb_delay);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W91,MGM_W90);
   not MGM_G117(MGM_W92,d_delay);
   and MGM_G118(MGM_W93,MGM_W92,clk_delay);
   and MGM_G119(MGM_W94,si_delay,MGM_W93);
   and MGM_G120(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W94);
   and MGM_G121(MGM_W95,d_delay,clk_delay);
   not MGM_G122(MGM_W96,si_delay);
   and MGM_G123(MGM_W97,MGM_W96,MGM_W95);
   not MGM_G124(MGM_W98,ssb_delay);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W98,MGM_W97);
   and MGM_G126(MGM_W99,d_delay,clk_delay);
   not MGM_G127(MGM_W100,si_delay);
   and MGM_G128(MGM_W101,MGM_W100,MGM_W99);
   and MGM_G129(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W101);
   and MGM_G130(MGM_W102,d_delay,clk_delay);
   and MGM_G131(MGM_W103,si_delay,MGM_W102);
   not MGM_G132(MGM_W104,ssb_delay);
   and MGM_G133(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W104,MGM_W103);
   and MGM_G134(MGM_W105,d_delay,clk_delay);
   and MGM_G135(MGM_W106,si_delay,MGM_W105);
   and MGM_G136(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W106);
   not MGM_G137(MGM_W107,d_delay);
   and MGM_G138(MGM_W108,psb_delay,MGM_W107);
   not MGM_G139(MGM_W109,ssb_delay);
   and MGM_G140(ENABLE_NOT_d_AND_psb_AND_NOT_ssb,MGM_W109,MGM_W108);
   and MGM_G141(MGM_W110,psb_delay,d_delay);
   not MGM_G142(MGM_W111,ssb_delay);
   and MGM_G143(ENABLE_d_AND_psb_AND_NOT_ssb,MGM_W111,MGM_W110);
   not MGM_G144(MGM_W112,d_delay);
   and MGM_G145(MGM_W113,psb_delay,MGM_W112);
   and MGM_G146(ENABLE_NOT_d_AND_psb_AND_si,si_delay,MGM_W113);
   and MGM_G147(MGM_W114,psb_delay,d_delay);
   not MGM_G148(MGM_W115,si_delay);
   and MGM_G149(ENABLE_d_AND_psb_AND_NOT_si,MGM_W115,MGM_W114);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b0))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fpn000ah_func( clk, d, o, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, d, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_0( MGM_D0, d );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fpn000ah1n02x5( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn000ah1n03x5( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn000ah1n04x5( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn000ah1n06x5( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn000ah1n08x5( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn000ah1n08x7( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n08x7_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n08x7_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n08x7_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n08x7_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn000ah1n12x5( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn000ah1n12x7( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n12x7_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n12x7_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n12x7_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n12x7_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn000ah1n16x5( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn000ah1n16x7( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n16x7_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n16x7_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn000ah_func b15fpn000ah1n16x7_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn000ah_func b15fpn000ah1n16x7_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine


primitive INTCseq_fpn010ah_N_IQN_FF_UDP( Q, C, P, CK, D `ifdef POWER_AWARE_MODE , vcc, vssx `endif , N );
   output Q;
   reg Q;
   input C, P, CK, D, N; 
   `ifdef POWER_AWARE_MODE
   input vcc, vssx;
   `endif
   table 
  `ifdef POWER_AWARE_MODE
   //C  P  CK D  PW GN N  :  Q  :  Q 
     0  0  n  ?  1  0  ?  :  ?  :  -;
     ?  0  n  ?  1  0  ?  :  1  :  1;
     0  ?  n  ?  1  0  ?  :  0  :  0;
     ?  0  r  0  1  0  ?  :  ?  :  1;
     1  0  ?  ?  1  0  ?  :  ?  :  1;
     0  ?  r  1  1  0  ?  :  ?  :  0;
     0  1  ?  ?  1  0  ?  :  ?  :  0;
     0  0  ?  *  1  0  ?  :  ?  :  -;
     0  ?  ?  *  1  0  ?  :  0  :  0;
     ?  0  ?  *  1  0  ?  :  1  :  1;
     0  *  ?  ?  1  0  ?  :  0  :  0;
     *  0  ?  ?  1  0  ?  :  1  :  1;
     ?  0  *  0  1  0  ?  :  1  :  1;
     0  ?  *  1  1  0  ?  :  0  :  0;
     ?  ?  ?  ?  1  0  *  :  ?  :  x;
  `else
   //C  P  CK D  N  :  Q  :  Q 
     0  0  n  ?  ?  :  ?  :  -;
     ?  0  n  ?  ?  :  1  :  1;
     0  ?  n  ?  ?  :  0  :  0;
     ?  0  r  0  ?  :  ?  :  1;
     1  0  ?  ?  ?  :  ?  :  1;
     0  ?  r  1  ?  :  ?  :  0;
     0  1  ?  ?  ?  :  ?  :  0;
     0  0  ?  *  ?  :  ?  :  -;
     0  ?  ?  *  ?  :  0  :  0;
     ?  0  ?  *  ?  :  1  :  1;
     0  *  ?  ?  ?  :  0  :  0;
     *  0  ?  ?  ?  :  1  :  1;
     ?  0  *  0  ?  :  1  :  1;
     0  ?  *  1  ?  :  0  :  0;
     ?  ?  ?  ?  *  :  ?  :  x;
  `endif

endtable
endprimitive



`celldefine
module INTCseq_fpn010ah_func( clk, d, o1, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, notifier;
   output o1;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, d, vcc, vssx );
   INTCseq_fpn010ah_N_IQN_FF_UDP( IQN, 1'b0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o1, IQN, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_0( MGM_D0, d );
   INTCseq_fpn010ah_N_IQN_FF_UDP( IQN, 1'b0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o1, IQN );
`endif

endmodule
`endcelldefine



`celldefine
module b15fpn010ah1n02x5( clk, d, o1 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o1;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn010ah_func b15fpn010ah1n02x5_behav_inst(.clk(clk),.d(d),.o1(o1),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn010ah_func b15fpn010ah1n02x5_behav_inst(.clk(clk),.d(d),.o1(o1),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn010ah_func b15fpn010ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn010ah_func b15fpn010ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn010ah1n03x5( clk, d, o1 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o1;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn010ah_func b15fpn010ah1n03x5_behav_inst(.clk(clk),.d(d),.o1(o1),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn010ah_func b15fpn010ah1n03x5_behav_inst(.clk(clk),.d(d),.o1(o1),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn010ah_func b15fpn010ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn010ah_func b15fpn010ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn010ah1n04x5( clk, d, o1 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o1;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn010ah_func b15fpn010ah1n04x5_behav_inst(.clk(clk),.d(d),.o1(o1),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn010ah_func b15fpn010ah1n04x5_behav_inst(.clk(clk),.d(d),.o1(o1),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn010ah_func b15fpn010ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn010ah_func b15fpn010ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn010ah1n06x5( clk, d, o1 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o1;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn010ah_func b15fpn010ah1n06x5_behav_inst(.clk(clk),.d(d),.o1(o1),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn010ah_func b15fpn010ah1n06x5_behav_inst(.clk(clk),.d(d),.o1(o1),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn010ah_func b15fpn010ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn010ah_func b15fpn010ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn010ah1n08x5( clk, d, o1 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o1;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn010ah_func b15fpn010ah1n08x5_behav_inst(.clk(clk),.d(d),.o1(o1),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn010ah_func b15fpn010ah1n08x5_behav_inst(.clk(clk),.d(d),.o1(o1),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn010ah_func b15fpn010ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn010ah_func b15fpn010ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn010ah1n12x5( clk, d, o1 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o1;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn010ah_func b15fpn010ah1n12x5_behav_inst(.clk(clk),.d(d),.o1(o1),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn010ah_func b15fpn010ah1n12x5_behav_inst(.clk(clk),.d(d),.o1(o1),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn010ah_func b15fpn010ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn010ah_func b15fpn010ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn010ah1n16x5( clk, d, o1 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o1;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn010ah_func b15fpn010ah1n16x5_behav_inst(.clk(clk),.d(d),.o1(o1),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn010ah_func b15fpn010ah1n16x5_behav_inst(.clk(clk),.d(d),.o1(o1),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn010ah_func b15fpn010ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn010ah_func b15fpn010ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine


primitive INTCseq_fpn040ah_6( int1, IQ, d, den `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
  output int1;
  input IQ, d, den;
  `ifdef POWER_AWARE_MODE
  input vcc, vssx;
  `endif

  table
  `ifdef POWER_AWARE_MODE
  //IQ, d, den vcc, vssx: int1
    1  1  ?  1  0: 1;
    1  ?  0  1  0: 1;
    ?  1  1  1  0: 1;
    0  0  ?  1  0: 0;
    0  ?  0  1  0: 0;
    ?  0  1  1  0: 0;
  `else
  //IQ, d, den: int1
    1  1  ?: 1;
    1  ?  0: 1;
    ?  1  1: 1;
    0  0  ?: 0;
    0  ?  0: 0;
    ?  0  1: 0;
  `endif
  endtable

endprimitive



`celldefine
module INTCseq_fpn040ah_func( clk, d, den, o, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, int1, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_fpn040ah_6( int1, IQ, d, den, vcc, vssx );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_0( MGM_D0, int1 );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_fpn040ah_6( int1, IQ, d, den );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fpn040ah1n02x5( clk, d, den, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn040ah_func b15fpn040ah1n02x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn040ah_func b15fpn040ah1n02x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn040ah_func b15fpn040ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn040ah_func b15fpn040ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_den,den_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_den,den_delay,d_delay);
   buf MGM_G3(ENABLE_den,den_delay);
   not MGM_G4(ENABLE_NOT_d,d_delay);
   buf MGM_G5(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den == 1'b1),
      negedge d &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den == 1'b1),
      posedge d &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d == 1'b1),
      negedge den &&& (ENABLE_NOT_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d == 1'b1),
      posedge den &&& (ENABLE_NOT_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d == 1'b1),
      negedge den &&& (ENABLE_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d == 1'b1),
      posedge den &&& (ENABLE_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn040ah1n03x5( clk, d, den, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn040ah_func b15fpn040ah1n03x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn040ah_func b15fpn040ah1n03x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn040ah_func b15fpn040ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn040ah_func b15fpn040ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_den,den_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_den,den_delay,d_delay);
   buf MGM_G3(ENABLE_den,den_delay);
   not MGM_G4(ENABLE_NOT_d,d_delay);
   buf MGM_G5(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den == 1'b1),
      negedge d &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den == 1'b1),
      posedge d &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d == 1'b1),
      negedge den &&& (ENABLE_NOT_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d == 1'b1),
      posedge den &&& (ENABLE_NOT_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d == 1'b1),
      negedge den &&& (ENABLE_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d == 1'b1),
      posedge den &&& (ENABLE_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn040ah1n04x5( clk, d, den, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn040ah_func b15fpn040ah1n04x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn040ah_func b15fpn040ah1n04x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn040ah_func b15fpn040ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn040ah_func b15fpn040ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_den,den_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_den,den_delay,d_delay);
   buf MGM_G3(ENABLE_den,den_delay);
   not MGM_G4(ENABLE_NOT_d,d_delay);
   buf MGM_G5(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den == 1'b1),
      negedge d &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den == 1'b1),
      posedge d &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d == 1'b1),
      negedge den &&& (ENABLE_NOT_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d == 1'b1),
      posedge den &&& (ENABLE_NOT_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d == 1'b1),
      negedge den &&& (ENABLE_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d == 1'b1),
      posedge den &&& (ENABLE_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn040ah1n06x5( clk, d, den, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn040ah_func b15fpn040ah1n06x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn040ah_func b15fpn040ah1n06x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn040ah_func b15fpn040ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn040ah_func b15fpn040ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_den,den_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_den,den_delay,d_delay);
   buf MGM_G3(ENABLE_den,den_delay);
   not MGM_G4(ENABLE_NOT_d,d_delay);
   buf MGM_G5(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den == 1'b1),
      negedge d &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den == 1'b1),
      posedge d &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d == 1'b1),
      negedge den &&& (ENABLE_NOT_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d == 1'b1),
      posedge den &&& (ENABLE_NOT_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d == 1'b1),
      negedge den &&& (ENABLE_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d == 1'b1),
      posedge den &&& (ENABLE_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn040ah1n08x5( clk, d, den, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn040ah_func b15fpn040ah1n08x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn040ah_func b15fpn040ah1n08x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn040ah_func b15fpn040ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn040ah_func b15fpn040ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_den,den_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_den,den_delay,d_delay);
   buf MGM_G3(ENABLE_den,den_delay);
   not MGM_G4(ENABLE_NOT_d,d_delay);
   buf MGM_G5(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den == 1'b1),
      negedge d &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den == 1'b1),
      posedge d &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d == 1'b1),
      negedge den &&& (ENABLE_NOT_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d == 1'b1),
      posedge den &&& (ENABLE_NOT_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d == 1'b1),
      negedge den &&& (ENABLE_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d == 1'b1),
      posedge den &&& (ENABLE_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn040ah1n12x5( clk, d, den, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn040ah_func b15fpn040ah1n12x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn040ah_func b15fpn040ah1n12x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn040ah_func b15fpn040ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn040ah_func b15fpn040ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_den,den_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_den,den_delay,d_delay);
   buf MGM_G3(ENABLE_den,den_delay);
   not MGM_G4(ENABLE_NOT_d,d_delay);
   buf MGM_G5(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den == 1'b1),
      negedge d &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den == 1'b1),
      posedge d &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d == 1'b1),
      negedge den &&& (ENABLE_NOT_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d == 1'b1),
      posedge den &&& (ENABLE_NOT_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d == 1'b1),
      negedge den &&& (ENABLE_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d == 1'b1),
      posedge den &&& (ENABLE_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn040ah1n16x5( clk, d, den, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn040ah_func b15fpn040ah1n16x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn040ah_func b15fpn040ah1n16x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn040ah_func b15fpn040ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn040ah_func b15fpn040ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_den,den_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_den,den_delay,d_delay);
   buf MGM_G3(ENABLE_den,den_delay);
   not MGM_G4(ENABLE_NOT_d,d_delay);
   buf MGM_G5(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den == 1'b1),
      negedge d &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den == 1'b1),
      posedge d &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d == 1'b1),
      negedge den &&& (ENABLE_NOT_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d == 1'b1),
      posedge den &&& (ENABLE_NOT_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d == 1'b1),
      negedge den &&& (ENABLE_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d == 1'b1),
      posedge den &&& (ENABLE_d == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fpn080ah_func( clkb, d, o, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_1( MGM_CLK0, clkb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, d, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_1( MGM_CLK0, clkb );
   INTCseq_cdiar2ah_0( MGM_D0, d );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fpn080ah1n02x5( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n02x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n02x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n02x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n02x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn080ah1n03x5( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n03x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n03x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n03x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n03x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn080ah1n04x5( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n04x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n04x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n04x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n04x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn080ah1n06x5( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n06x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n06x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n06x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n06x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn080ah1n08x5( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n08x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n08x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n08x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n08x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn080ah1n08x7( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n08x7_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n08x7_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n08x7_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n08x7_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn080ah1n12x5( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n12x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n12x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n12x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n12x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn080ah1n12x7( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n12x7_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n12x7_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n12x7_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n12x7_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn080ah1n16x5( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n16x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n16x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n16x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n16x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpn080ah1n16x7( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n16x7_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n16x7_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpn080ah_func b15fpn080ah1n16x7_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpn080ah_func b15fpn080ah1n16x7_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fpy000ah_func( clk, d, o, si, ssb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fpy000ah1n02x5( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy000ah1n03x5( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy000ah1n04x5( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy000ah1n06x5( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy000ah1n08x5( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy000ah1n08x7( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n08x7_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n08x7_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n08x7_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n08x7_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy000ah1n12x5( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy000ah1n12x7( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n12x7_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n12x7_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n12x7_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n12x7_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy000ah1n16x5( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy000ah1n16x7( clk, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n16x7_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n16x7_behav_inst(.clk(clk),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy000ah_func b15fpy000ah1n16x7_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy000ah_func b15fpy000ah1n16x7_inst(.clk(clk_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fpy010ah_func( clk, d, o1, si, ssb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb, notifier;
   output o1;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_fpn010ah_N_IQN_FF_UDP( IQN, 1'b0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o1, IQN, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_fpn010ah_N_IQN_FF_UDP( IQN, 1'b0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o1, IQN );
`endif

endmodule
`endcelldefine



`celldefine
module b15fpy010ah1n02x5( clk, d, o1, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o1;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy010ah_func b15fpy010ah1n02x5_behav_inst(.clk(clk),.d(d),.o1(o1),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy010ah_func b15fpy010ah1n02x5_behav_inst(.clk(clk),.d(d),.o1(o1),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy010ah_func b15fpy010ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy010ah_func b15fpy010ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy010ah1n03x5( clk, d, o1, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o1;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy010ah_func b15fpy010ah1n03x5_behav_inst(.clk(clk),.d(d),.o1(o1),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy010ah_func b15fpy010ah1n03x5_behav_inst(.clk(clk),.d(d),.o1(o1),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy010ah_func b15fpy010ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy010ah_func b15fpy010ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy010ah1n04x5( clk, d, o1, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o1;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy010ah_func b15fpy010ah1n04x5_behav_inst(.clk(clk),.d(d),.o1(o1),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy010ah_func b15fpy010ah1n04x5_behav_inst(.clk(clk),.d(d),.o1(o1),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy010ah_func b15fpy010ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy010ah_func b15fpy010ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy010ah1n06x5( clk, d, o1, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o1;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy010ah_func b15fpy010ah1n06x5_behav_inst(.clk(clk),.d(d),.o1(o1),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy010ah_func b15fpy010ah1n06x5_behav_inst(.clk(clk),.d(d),.o1(o1),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy010ah_func b15fpy010ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy010ah_func b15fpy010ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy010ah1n08x5( clk, d, o1, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o1;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy010ah_func b15fpy010ah1n08x5_behav_inst(.clk(clk),.d(d),.o1(o1),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy010ah_func b15fpy010ah1n08x5_behav_inst(.clk(clk),.d(d),.o1(o1),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy010ah_func b15fpy010ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy010ah_func b15fpy010ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy010ah1n12x5( clk, d, o1, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o1;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy010ah_func b15fpy010ah1n12x5_behav_inst(.clk(clk),.d(d),.o1(o1),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy010ah_func b15fpy010ah1n12x5_behav_inst(.clk(clk),.d(d),.o1(o1),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy010ah_func b15fpy010ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy010ah_func b15fpy010ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy010ah1n16x5( clk, d, o1, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, si, ssb;
   output o1;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy010ah_func b15fpy010ah1n16x5_behav_inst(.clk(clk),.d(d),.o1(o1),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy010ah_func b15fpy010ah1n16x5_behav_inst(.clk(clk),.d(d),.o1(o1),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy010ah_func b15fpy010ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy010ah_func b15fpy010ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o1(o1),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fpy040ah_func( clk, d, den, o, si, ssb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, si, ssb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, int2, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_fpn040ah_6( int1, IQ, d, den, vcc, vssx );
   INTCseq_fdw003ah_5( int2, int1, si, ssb, vcc, vssx );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_0( MGM_D0, int2 );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_fpn040ah_6( int1, IQ, d, den );
   INTCseq_fdw003ah_5( int2, int1, si, ssb );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fpy040ah1n02x5( clk, d, den, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy040ah_func b15fpy040ah1n02x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy040ah_func b15fpy040ah1n02x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy040ah_func b15fpy040ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy040ah_func b15fpy040ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,den_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   not MGM_G8(MGM_W7,den_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(MGM_W9,si_delay,MGM_W8);
   not MGM_G11(MGM_W10,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W10,MGM_W9);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,den_delay,MGM_W11);
   not MGM_G15(MGM_W13,si_delay);
   and MGM_G16(MGM_W14,MGM_W13,MGM_W12);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,den_delay,MGM_W16);
   not MGM_G21(MGM_W18,si_delay);
   and MGM_G22(MGM_W19,MGM_W18,MGM_W17);
   and MGM_G23(ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G24(MGM_W20,d_delay);
   and MGM_G25(MGM_W21,den_delay,MGM_W20);
   and MGM_G26(MGM_W22,si_delay,MGM_W21);
   not MGM_G27(MGM_W23,ssb_delay);
   and MGM_G28(ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W23,MGM_W22);
   not MGM_G29(MGM_W24,d_delay);
   and MGM_G30(MGM_W25,den_delay,MGM_W24);
   and MGM_G31(MGM_W26,si_delay,MGM_W25);
   and MGM_G32(ENABLE_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W26);
   not MGM_G33(MGM_W27,den_delay);
   and MGM_G34(MGM_W28,MGM_W27,d_delay);
   not MGM_G35(MGM_W29,si_delay);
   and MGM_G36(MGM_W30,MGM_W29,MGM_W28);
   not MGM_G37(MGM_W31,ssb_delay);
   and MGM_G38(ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W31,MGM_W30);
   not MGM_G39(MGM_W32,den_delay);
   and MGM_G40(MGM_W33,MGM_W32,d_delay);
   and MGM_G41(MGM_W34,si_delay,MGM_W33);
   not MGM_G42(MGM_W35,ssb_delay);
   and MGM_G43(ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W35,MGM_W34);
   and MGM_G44(MGM_W36,den_delay,d_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   not MGM_G47(MGM_W39,ssb_delay);
   and MGM_G48(ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W39,MGM_W38);
   and MGM_G49(MGM_W40,den_delay,d_delay);
   not MGM_G50(MGM_W41,si_delay);
   and MGM_G51(MGM_W42,MGM_W41,MGM_W40);
   and MGM_G52(ENABLE_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W42);
   and MGM_G53(MGM_W43,den_delay,d_delay);
   and MGM_G54(MGM_W44,si_delay,MGM_W43);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_d_AND_den_AND_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   and MGM_G57(MGM_W46,den_delay,d_delay);
   and MGM_G58(MGM_W47,si_delay,MGM_W46);
   and MGM_G59(ENABLE_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W47);
   not MGM_G60(MGM_W48,si_delay);
   and MGM_G61(MGM_W49,MGM_W48,den_delay);
   and MGM_G62(ENABLE_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   and MGM_G63(MGM_W50,si_delay,den_delay);
   and MGM_G64(ENABLE_den_AND_si_AND_ssb,ssb_delay,MGM_W50);
   not MGM_G65(MGM_W51,d_delay);
   not MGM_G66(MGM_W52,si_delay);
   and MGM_G67(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G68(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G69(MGM_W54,d_delay);
   and MGM_G70(MGM_W55,si_delay,MGM_W54);
   and MGM_G71(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W55);
   not MGM_G72(MGM_W56,si_delay);
   and MGM_G73(MGM_W57,MGM_W56,d_delay);
   and MGM_G74(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W57);
   and MGM_G75(MGM_W58,si_delay,d_delay);
   and MGM_G76(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,d_delay);
   not MGM_G78(MGM_W60,den_delay);
   and MGM_G79(MGM_W61,MGM_W60,MGM_W59);
   not MGM_G80(MGM_W62,ssb_delay);
   and MGM_G81(ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb,MGM_W62,MGM_W61);
   not MGM_G82(MGM_W63,d_delay);
   and MGM_G83(MGM_W64,den_delay,MGM_W63);
   not MGM_G84(MGM_W65,ssb_delay);
   and MGM_G85(ENABLE_NOT_d_AND_den_AND_NOT_ssb,MGM_W65,MGM_W64);
   not MGM_G86(MGM_W66,den_delay);
   and MGM_G87(MGM_W67,MGM_W66,d_delay);
   not MGM_G88(MGM_W68,ssb_delay);
   and MGM_G89(ENABLE_d_AND_NOT_den_AND_NOT_ssb,MGM_W68,MGM_W67);
   and MGM_G90(MGM_W69,den_delay,d_delay);
   not MGM_G91(MGM_W70,ssb_delay);
   and MGM_G92(ENABLE_d_AND_den_AND_NOT_ssb,MGM_W70,MGM_W69);
   not MGM_G93(MGM_W71,d_delay);
   not MGM_G94(MGM_W72,den_delay);
   and MGM_G95(MGM_W73,MGM_W72,MGM_W71);
   not MGM_G96(MGM_W74,si_delay);
   and MGM_G97(ENABLE_NOT_d_AND_NOT_den_AND_NOT_si,MGM_W74,MGM_W73);
   not MGM_G98(MGM_W75,d_delay);
   not MGM_G99(MGM_W76,den_delay);
   and MGM_G100(MGM_W77,MGM_W76,MGM_W75);
   and MGM_G101(ENABLE_NOT_d_AND_NOT_den_AND_si,si_delay,MGM_W77);
   not MGM_G102(MGM_W78,d_delay);
   and MGM_G103(MGM_W79,den_delay,MGM_W78);
   and MGM_G104(ENABLE_NOT_d_AND_den_AND_si,si_delay,MGM_W79);
   not MGM_G105(MGM_W80,den_delay);
   and MGM_G106(MGM_W81,MGM_W80,d_delay);
   not MGM_G107(MGM_W82,si_delay);
   and MGM_G108(ENABLE_d_AND_NOT_den_AND_NOT_si,MGM_W82,MGM_W81);
   not MGM_G109(MGM_W83,den_delay);
   and MGM_G110(MGM_W84,MGM_W83,d_delay);
   and MGM_G111(ENABLE_d_AND_NOT_den_AND_si,si_delay,MGM_W84);
   and MGM_G112(MGM_W85,den_delay,d_delay);
   not MGM_G113(MGM_W86,si_delay);
   and MGM_G114(ENABLE_d_AND_den_AND_NOT_si,MGM_W86,MGM_W85);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy040ah1n03x5( clk, d, den, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy040ah_func b15fpy040ah1n03x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy040ah_func b15fpy040ah1n03x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy040ah_func b15fpy040ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy040ah_func b15fpy040ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,den_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   not MGM_G8(MGM_W7,den_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(MGM_W9,si_delay,MGM_W8);
   not MGM_G11(MGM_W10,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W10,MGM_W9);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,den_delay,MGM_W11);
   not MGM_G15(MGM_W13,si_delay);
   and MGM_G16(MGM_W14,MGM_W13,MGM_W12);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,den_delay,MGM_W16);
   not MGM_G21(MGM_W18,si_delay);
   and MGM_G22(MGM_W19,MGM_W18,MGM_W17);
   and MGM_G23(ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G24(MGM_W20,d_delay);
   and MGM_G25(MGM_W21,den_delay,MGM_W20);
   and MGM_G26(MGM_W22,si_delay,MGM_W21);
   not MGM_G27(MGM_W23,ssb_delay);
   and MGM_G28(ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W23,MGM_W22);
   not MGM_G29(MGM_W24,d_delay);
   and MGM_G30(MGM_W25,den_delay,MGM_W24);
   and MGM_G31(MGM_W26,si_delay,MGM_W25);
   and MGM_G32(ENABLE_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W26);
   not MGM_G33(MGM_W27,den_delay);
   and MGM_G34(MGM_W28,MGM_W27,d_delay);
   not MGM_G35(MGM_W29,si_delay);
   and MGM_G36(MGM_W30,MGM_W29,MGM_W28);
   not MGM_G37(MGM_W31,ssb_delay);
   and MGM_G38(ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W31,MGM_W30);
   not MGM_G39(MGM_W32,den_delay);
   and MGM_G40(MGM_W33,MGM_W32,d_delay);
   and MGM_G41(MGM_W34,si_delay,MGM_W33);
   not MGM_G42(MGM_W35,ssb_delay);
   and MGM_G43(ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W35,MGM_W34);
   and MGM_G44(MGM_W36,den_delay,d_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   not MGM_G47(MGM_W39,ssb_delay);
   and MGM_G48(ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W39,MGM_W38);
   and MGM_G49(MGM_W40,den_delay,d_delay);
   not MGM_G50(MGM_W41,si_delay);
   and MGM_G51(MGM_W42,MGM_W41,MGM_W40);
   and MGM_G52(ENABLE_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W42);
   and MGM_G53(MGM_W43,den_delay,d_delay);
   and MGM_G54(MGM_W44,si_delay,MGM_W43);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_d_AND_den_AND_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   and MGM_G57(MGM_W46,den_delay,d_delay);
   and MGM_G58(MGM_W47,si_delay,MGM_W46);
   and MGM_G59(ENABLE_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W47);
   not MGM_G60(MGM_W48,si_delay);
   and MGM_G61(MGM_W49,MGM_W48,den_delay);
   and MGM_G62(ENABLE_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   and MGM_G63(MGM_W50,si_delay,den_delay);
   and MGM_G64(ENABLE_den_AND_si_AND_ssb,ssb_delay,MGM_W50);
   not MGM_G65(MGM_W51,d_delay);
   not MGM_G66(MGM_W52,si_delay);
   and MGM_G67(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G68(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G69(MGM_W54,d_delay);
   and MGM_G70(MGM_W55,si_delay,MGM_W54);
   and MGM_G71(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W55);
   not MGM_G72(MGM_W56,si_delay);
   and MGM_G73(MGM_W57,MGM_W56,d_delay);
   and MGM_G74(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W57);
   and MGM_G75(MGM_W58,si_delay,d_delay);
   and MGM_G76(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,d_delay);
   not MGM_G78(MGM_W60,den_delay);
   and MGM_G79(MGM_W61,MGM_W60,MGM_W59);
   not MGM_G80(MGM_W62,ssb_delay);
   and MGM_G81(ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb,MGM_W62,MGM_W61);
   not MGM_G82(MGM_W63,d_delay);
   and MGM_G83(MGM_W64,den_delay,MGM_W63);
   not MGM_G84(MGM_W65,ssb_delay);
   and MGM_G85(ENABLE_NOT_d_AND_den_AND_NOT_ssb,MGM_W65,MGM_W64);
   not MGM_G86(MGM_W66,den_delay);
   and MGM_G87(MGM_W67,MGM_W66,d_delay);
   not MGM_G88(MGM_W68,ssb_delay);
   and MGM_G89(ENABLE_d_AND_NOT_den_AND_NOT_ssb,MGM_W68,MGM_W67);
   and MGM_G90(MGM_W69,den_delay,d_delay);
   not MGM_G91(MGM_W70,ssb_delay);
   and MGM_G92(ENABLE_d_AND_den_AND_NOT_ssb,MGM_W70,MGM_W69);
   not MGM_G93(MGM_W71,d_delay);
   not MGM_G94(MGM_W72,den_delay);
   and MGM_G95(MGM_W73,MGM_W72,MGM_W71);
   not MGM_G96(MGM_W74,si_delay);
   and MGM_G97(ENABLE_NOT_d_AND_NOT_den_AND_NOT_si,MGM_W74,MGM_W73);
   not MGM_G98(MGM_W75,d_delay);
   not MGM_G99(MGM_W76,den_delay);
   and MGM_G100(MGM_W77,MGM_W76,MGM_W75);
   and MGM_G101(ENABLE_NOT_d_AND_NOT_den_AND_si,si_delay,MGM_W77);
   not MGM_G102(MGM_W78,d_delay);
   and MGM_G103(MGM_W79,den_delay,MGM_W78);
   and MGM_G104(ENABLE_NOT_d_AND_den_AND_si,si_delay,MGM_W79);
   not MGM_G105(MGM_W80,den_delay);
   and MGM_G106(MGM_W81,MGM_W80,d_delay);
   not MGM_G107(MGM_W82,si_delay);
   and MGM_G108(ENABLE_d_AND_NOT_den_AND_NOT_si,MGM_W82,MGM_W81);
   not MGM_G109(MGM_W83,den_delay);
   and MGM_G110(MGM_W84,MGM_W83,d_delay);
   and MGM_G111(ENABLE_d_AND_NOT_den_AND_si,si_delay,MGM_W84);
   and MGM_G112(MGM_W85,den_delay,d_delay);
   not MGM_G113(MGM_W86,si_delay);
   and MGM_G114(ENABLE_d_AND_den_AND_NOT_si,MGM_W86,MGM_W85);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy040ah1n04x5( clk, d, den, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy040ah_func b15fpy040ah1n04x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy040ah_func b15fpy040ah1n04x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy040ah_func b15fpy040ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy040ah_func b15fpy040ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,den_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   not MGM_G8(MGM_W7,den_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(MGM_W9,si_delay,MGM_W8);
   not MGM_G11(MGM_W10,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W10,MGM_W9);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,den_delay,MGM_W11);
   not MGM_G15(MGM_W13,si_delay);
   and MGM_G16(MGM_W14,MGM_W13,MGM_W12);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,den_delay,MGM_W16);
   not MGM_G21(MGM_W18,si_delay);
   and MGM_G22(MGM_W19,MGM_W18,MGM_W17);
   and MGM_G23(ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G24(MGM_W20,d_delay);
   and MGM_G25(MGM_W21,den_delay,MGM_W20);
   and MGM_G26(MGM_W22,si_delay,MGM_W21);
   not MGM_G27(MGM_W23,ssb_delay);
   and MGM_G28(ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W23,MGM_W22);
   not MGM_G29(MGM_W24,d_delay);
   and MGM_G30(MGM_W25,den_delay,MGM_W24);
   and MGM_G31(MGM_W26,si_delay,MGM_W25);
   and MGM_G32(ENABLE_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W26);
   not MGM_G33(MGM_W27,den_delay);
   and MGM_G34(MGM_W28,MGM_W27,d_delay);
   not MGM_G35(MGM_W29,si_delay);
   and MGM_G36(MGM_W30,MGM_W29,MGM_W28);
   not MGM_G37(MGM_W31,ssb_delay);
   and MGM_G38(ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W31,MGM_W30);
   not MGM_G39(MGM_W32,den_delay);
   and MGM_G40(MGM_W33,MGM_W32,d_delay);
   and MGM_G41(MGM_W34,si_delay,MGM_W33);
   not MGM_G42(MGM_W35,ssb_delay);
   and MGM_G43(ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W35,MGM_W34);
   and MGM_G44(MGM_W36,den_delay,d_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   not MGM_G47(MGM_W39,ssb_delay);
   and MGM_G48(ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W39,MGM_W38);
   and MGM_G49(MGM_W40,den_delay,d_delay);
   not MGM_G50(MGM_W41,si_delay);
   and MGM_G51(MGM_W42,MGM_W41,MGM_W40);
   and MGM_G52(ENABLE_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W42);
   and MGM_G53(MGM_W43,den_delay,d_delay);
   and MGM_G54(MGM_W44,si_delay,MGM_W43);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_d_AND_den_AND_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   and MGM_G57(MGM_W46,den_delay,d_delay);
   and MGM_G58(MGM_W47,si_delay,MGM_W46);
   and MGM_G59(ENABLE_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W47);
   not MGM_G60(MGM_W48,si_delay);
   and MGM_G61(MGM_W49,MGM_W48,den_delay);
   and MGM_G62(ENABLE_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   and MGM_G63(MGM_W50,si_delay,den_delay);
   and MGM_G64(ENABLE_den_AND_si_AND_ssb,ssb_delay,MGM_W50);
   not MGM_G65(MGM_W51,d_delay);
   not MGM_G66(MGM_W52,si_delay);
   and MGM_G67(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G68(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G69(MGM_W54,d_delay);
   and MGM_G70(MGM_W55,si_delay,MGM_W54);
   and MGM_G71(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W55);
   not MGM_G72(MGM_W56,si_delay);
   and MGM_G73(MGM_W57,MGM_W56,d_delay);
   and MGM_G74(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W57);
   and MGM_G75(MGM_W58,si_delay,d_delay);
   and MGM_G76(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,d_delay);
   not MGM_G78(MGM_W60,den_delay);
   and MGM_G79(MGM_W61,MGM_W60,MGM_W59);
   not MGM_G80(MGM_W62,ssb_delay);
   and MGM_G81(ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb,MGM_W62,MGM_W61);
   not MGM_G82(MGM_W63,d_delay);
   and MGM_G83(MGM_W64,den_delay,MGM_W63);
   not MGM_G84(MGM_W65,ssb_delay);
   and MGM_G85(ENABLE_NOT_d_AND_den_AND_NOT_ssb,MGM_W65,MGM_W64);
   not MGM_G86(MGM_W66,den_delay);
   and MGM_G87(MGM_W67,MGM_W66,d_delay);
   not MGM_G88(MGM_W68,ssb_delay);
   and MGM_G89(ENABLE_d_AND_NOT_den_AND_NOT_ssb,MGM_W68,MGM_W67);
   and MGM_G90(MGM_W69,den_delay,d_delay);
   not MGM_G91(MGM_W70,ssb_delay);
   and MGM_G92(ENABLE_d_AND_den_AND_NOT_ssb,MGM_W70,MGM_W69);
   not MGM_G93(MGM_W71,d_delay);
   not MGM_G94(MGM_W72,den_delay);
   and MGM_G95(MGM_W73,MGM_W72,MGM_W71);
   not MGM_G96(MGM_W74,si_delay);
   and MGM_G97(ENABLE_NOT_d_AND_NOT_den_AND_NOT_si,MGM_W74,MGM_W73);
   not MGM_G98(MGM_W75,d_delay);
   not MGM_G99(MGM_W76,den_delay);
   and MGM_G100(MGM_W77,MGM_W76,MGM_W75);
   and MGM_G101(ENABLE_NOT_d_AND_NOT_den_AND_si,si_delay,MGM_W77);
   not MGM_G102(MGM_W78,d_delay);
   and MGM_G103(MGM_W79,den_delay,MGM_W78);
   and MGM_G104(ENABLE_NOT_d_AND_den_AND_si,si_delay,MGM_W79);
   not MGM_G105(MGM_W80,den_delay);
   and MGM_G106(MGM_W81,MGM_W80,d_delay);
   not MGM_G107(MGM_W82,si_delay);
   and MGM_G108(ENABLE_d_AND_NOT_den_AND_NOT_si,MGM_W82,MGM_W81);
   not MGM_G109(MGM_W83,den_delay);
   and MGM_G110(MGM_W84,MGM_W83,d_delay);
   and MGM_G111(ENABLE_d_AND_NOT_den_AND_si,si_delay,MGM_W84);
   and MGM_G112(MGM_W85,den_delay,d_delay);
   not MGM_G113(MGM_W86,si_delay);
   and MGM_G114(ENABLE_d_AND_den_AND_NOT_si,MGM_W86,MGM_W85);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy040ah1n06x5( clk, d, den, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy040ah_func b15fpy040ah1n06x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy040ah_func b15fpy040ah1n06x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy040ah_func b15fpy040ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy040ah_func b15fpy040ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,den_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   not MGM_G8(MGM_W7,den_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(MGM_W9,si_delay,MGM_W8);
   not MGM_G11(MGM_W10,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W10,MGM_W9);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,den_delay,MGM_W11);
   not MGM_G15(MGM_W13,si_delay);
   and MGM_G16(MGM_W14,MGM_W13,MGM_W12);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,den_delay,MGM_W16);
   not MGM_G21(MGM_W18,si_delay);
   and MGM_G22(MGM_W19,MGM_W18,MGM_W17);
   and MGM_G23(ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G24(MGM_W20,d_delay);
   and MGM_G25(MGM_W21,den_delay,MGM_W20);
   and MGM_G26(MGM_W22,si_delay,MGM_W21);
   not MGM_G27(MGM_W23,ssb_delay);
   and MGM_G28(ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W23,MGM_W22);
   not MGM_G29(MGM_W24,d_delay);
   and MGM_G30(MGM_W25,den_delay,MGM_W24);
   and MGM_G31(MGM_W26,si_delay,MGM_W25);
   and MGM_G32(ENABLE_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W26);
   not MGM_G33(MGM_W27,den_delay);
   and MGM_G34(MGM_W28,MGM_W27,d_delay);
   not MGM_G35(MGM_W29,si_delay);
   and MGM_G36(MGM_W30,MGM_W29,MGM_W28);
   not MGM_G37(MGM_W31,ssb_delay);
   and MGM_G38(ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W31,MGM_W30);
   not MGM_G39(MGM_W32,den_delay);
   and MGM_G40(MGM_W33,MGM_W32,d_delay);
   and MGM_G41(MGM_W34,si_delay,MGM_W33);
   not MGM_G42(MGM_W35,ssb_delay);
   and MGM_G43(ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W35,MGM_W34);
   and MGM_G44(MGM_W36,den_delay,d_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   not MGM_G47(MGM_W39,ssb_delay);
   and MGM_G48(ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W39,MGM_W38);
   and MGM_G49(MGM_W40,den_delay,d_delay);
   not MGM_G50(MGM_W41,si_delay);
   and MGM_G51(MGM_W42,MGM_W41,MGM_W40);
   and MGM_G52(ENABLE_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W42);
   and MGM_G53(MGM_W43,den_delay,d_delay);
   and MGM_G54(MGM_W44,si_delay,MGM_W43);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_d_AND_den_AND_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   and MGM_G57(MGM_W46,den_delay,d_delay);
   and MGM_G58(MGM_W47,si_delay,MGM_W46);
   and MGM_G59(ENABLE_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W47);
   not MGM_G60(MGM_W48,si_delay);
   and MGM_G61(MGM_W49,MGM_W48,den_delay);
   and MGM_G62(ENABLE_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   and MGM_G63(MGM_W50,si_delay,den_delay);
   and MGM_G64(ENABLE_den_AND_si_AND_ssb,ssb_delay,MGM_W50);
   not MGM_G65(MGM_W51,d_delay);
   not MGM_G66(MGM_W52,si_delay);
   and MGM_G67(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G68(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G69(MGM_W54,d_delay);
   and MGM_G70(MGM_W55,si_delay,MGM_W54);
   and MGM_G71(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W55);
   not MGM_G72(MGM_W56,si_delay);
   and MGM_G73(MGM_W57,MGM_W56,d_delay);
   and MGM_G74(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W57);
   and MGM_G75(MGM_W58,si_delay,d_delay);
   and MGM_G76(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,d_delay);
   not MGM_G78(MGM_W60,den_delay);
   and MGM_G79(MGM_W61,MGM_W60,MGM_W59);
   not MGM_G80(MGM_W62,ssb_delay);
   and MGM_G81(ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb,MGM_W62,MGM_W61);
   not MGM_G82(MGM_W63,d_delay);
   and MGM_G83(MGM_W64,den_delay,MGM_W63);
   not MGM_G84(MGM_W65,ssb_delay);
   and MGM_G85(ENABLE_NOT_d_AND_den_AND_NOT_ssb,MGM_W65,MGM_W64);
   not MGM_G86(MGM_W66,den_delay);
   and MGM_G87(MGM_W67,MGM_W66,d_delay);
   not MGM_G88(MGM_W68,ssb_delay);
   and MGM_G89(ENABLE_d_AND_NOT_den_AND_NOT_ssb,MGM_W68,MGM_W67);
   and MGM_G90(MGM_W69,den_delay,d_delay);
   not MGM_G91(MGM_W70,ssb_delay);
   and MGM_G92(ENABLE_d_AND_den_AND_NOT_ssb,MGM_W70,MGM_W69);
   not MGM_G93(MGM_W71,d_delay);
   not MGM_G94(MGM_W72,den_delay);
   and MGM_G95(MGM_W73,MGM_W72,MGM_W71);
   not MGM_G96(MGM_W74,si_delay);
   and MGM_G97(ENABLE_NOT_d_AND_NOT_den_AND_NOT_si,MGM_W74,MGM_W73);
   not MGM_G98(MGM_W75,d_delay);
   not MGM_G99(MGM_W76,den_delay);
   and MGM_G100(MGM_W77,MGM_W76,MGM_W75);
   and MGM_G101(ENABLE_NOT_d_AND_NOT_den_AND_si,si_delay,MGM_W77);
   not MGM_G102(MGM_W78,d_delay);
   and MGM_G103(MGM_W79,den_delay,MGM_W78);
   and MGM_G104(ENABLE_NOT_d_AND_den_AND_si,si_delay,MGM_W79);
   not MGM_G105(MGM_W80,den_delay);
   and MGM_G106(MGM_W81,MGM_W80,d_delay);
   not MGM_G107(MGM_W82,si_delay);
   and MGM_G108(ENABLE_d_AND_NOT_den_AND_NOT_si,MGM_W82,MGM_W81);
   not MGM_G109(MGM_W83,den_delay);
   and MGM_G110(MGM_W84,MGM_W83,d_delay);
   and MGM_G111(ENABLE_d_AND_NOT_den_AND_si,si_delay,MGM_W84);
   and MGM_G112(MGM_W85,den_delay,d_delay);
   not MGM_G113(MGM_W86,si_delay);
   and MGM_G114(ENABLE_d_AND_den_AND_NOT_si,MGM_W86,MGM_W85);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy040ah1n08x5( clk, d, den, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy040ah_func b15fpy040ah1n08x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy040ah_func b15fpy040ah1n08x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy040ah_func b15fpy040ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy040ah_func b15fpy040ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,den_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   not MGM_G8(MGM_W7,den_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(MGM_W9,si_delay,MGM_W8);
   not MGM_G11(MGM_W10,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W10,MGM_W9);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,den_delay,MGM_W11);
   not MGM_G15(MGM_W13,si_delay);
   and MGM_G16(MGM_W14,MGM_W13,MGM_W12);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,den_delay,MGM_W16);
   not MGM_G21(MGM_W18,si_delay);
   and MGM_G22(MGM_W19,MGM_W18,MGM_W17);
   and MGM_G23(ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G24(MGM_W20,d_delay);
   and MGM_G25(MGM_W21,den_delay,MGM_W20);
   and MGM_G26(MGM_W22,si_delay,MGM_W21);
   not MGM_G27(MGM_W23,ssb_delay);
   and MGM_G28(ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W23,MGM_W22);
   not MGM_G29(MGM_W24,d_delay);
   and MGM_G30(MGM_W25,den_delay,MGM_W24);
   and MGM_G31(MGM_W26,si_delay,MGM_W25);
   and MGM_G32(ENABLE_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W26);
   not MGM_G33(MGM_W27,den_delay);
   and MGM_G34(MGM_W28,MGM_W27,d_delay);
   not MGM_G35(MGM_W29,si_delay);
   and MGM_G36(MGM_W30,MGM_W29,MGM_W28);
   not MGM_G37(MGM_W31,ssb_delay);
   and MGM_G38(ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W31,MGM_W30);
   not MGM_G39(MGM_W32,den_delay);
   and MGM_G40(MGM_W33,MGM_W32,d_delay);
   and MGM_G41(MGM_W34,si_delay,MGM_W33);
   not MGM_G42(MGM_W35,ssb_delay);
   and MGM_G43(ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W35,MGM_W34);
   and MGM_G44(MGM_W36,den_delay,d_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   not MGM_G47(MGM_W39,ssb_delay);
   and MGM_G48(ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W39,MGM_W38);
   and MGM_G49(MGM_W40,den_delay,d_delay);
   not MGM_G50(MGM_W41,si_delay);
   and MGM_G51(MGM_W42,MGM_W41,MGM_W40);
   and MGM_G52(ENABLE_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W42);
   and MGM_G53(MGM_W43,den_delay,d_delay);
   and MGM_G54(MGM_W44,si_delay,MGM_W43);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_d_AND_den_AND_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   and MGM_G57(MGM_W46,den_delay,d_delay);
   and MGM_G58(MGM_W47,si_delay,MGM_W46);
   and MGM_G59(ENABLE_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W47);
   not MGM_G60(MGM_W48,si_delay);
   and MGM_G61(MGM_W49,MGM_W48,den_delay);
   and MGM_G62(ENABLE_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   and MGM_G63(MGM_W50,si_delay,den_delay);
   and MGM_G64(ENABLE_den_AND_si_AND_ssb,ssb_delay,MGM_W50);
   not MGM_G65(MGM_W51,d_delay);
   not MGM_G66(MGM_W52,si_delay);
   and MGM_G67(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G68(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G69(MGM_W54,d_delay);
   and MGM_G70(MGM_W55,si_delay,MGM_W54);
   and MGM_G71(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W55);
   not MGM_G72(MGM_W56,si_delay);
   and MGM_G73(MGM_W57,MGM_W56,d_delay);
   and MGM_G74(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W57);
   and MGM_G75(MGM_W58,si_delay,d_delay);
   and MGM_G76(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,d_delay);
   not MGM_G78(MGM_W60,den_delay);
   and MGM_G79(MGM_W61,MGM_W60,MGM_W59);
   not MGM_G80(MGM_W62,ssb_delay);
   and MGM_G81(ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb,MGM_W62,MGM_W61);
   not MGM_G82(MGM_W63,d_delay);
   and MGM_G83(MGM_W64,den_delay,MGM_W63);
   not MGM_G84(MGM_W65,ssb_delay);
   and MGM_G85(ENABLE_NOT_d_AND_den_AND_NOT_ssb,MGM_W65,MGM_W64);
   not MGM_G86(MGM_W66,den_delay);
   and MGM_G87(MGM_W67,MGM_W66,d_delay);
   not MGM_G88(MGM_W68,ssb_delay);
   and MGM_G89(ENABLE_d_AND_NOT_den_AND_NOT_ssb,MGM_W68,MGM_W67);
   and MGM_G90(MGM_W69,den_delay,d_delay);
   not MGM_G91(MGM_W70,ssb_delay);
   and MGM_G92(ENABLE_d_AND_den_AND_NOT_ssb,MGM_W70,MGM_W69);
   not MGM_G93(MGM_W71,d_delay);
   not MGM_G94(MGM_W72,den_delay);
   and MGM_G95(MGM_W73,MGM_W72,MGM_W71);
   not MGM_G96(MGM_W74,si_delay);
   and MGM_G97(ENABLE_NOT_d_AND_NOT_den_AND_NOT_si,MGM_W74,MGM_W73);
   not MGM_G98(MGM_W75,d_delay);
   not MGM_G99(MGM_W76,den_delay);
   and MGM_G100(MGM_W77,MGM_W76,MGM_W75);
   and MGM_G101(ENABLE_NOT_d_AND_NOT_den_AND_si,si_delay,MGM_W77);
   not MGM_G102(MGM_W78,d_delay);
   and MGM_G103(MGM_W79,den_delay,MGM_W78);
   and MGM_G104(ENABLE_NOT_d_AND_den_AND_si,si_delay,MGM_W79);
   not MGM_G105(MGM_W80,den_delay);
   and MGM_G106(MGM_W81,MGM_W80,d_delay);
   not MGM_G107(MGM_W82,si_delay);
   and MGM_G108(ENABLE_d_AND_NOT_den_AND_NOT_si,MGM_W82,MGM_W81);
   not MGM_G109(MGM_W83,den_delay);
   and MGM_G110(MGM_W84,MGM_W83,d_delay);
   and MGM_G111(ENABLE_d_AND_NOT_den_AND_si,si_delay,MGM_W84);
   and MGM_G112(MGM_W85,den_delay,d_delay);
   not MGM_G113(MGM_W86,si_delay);
   and MGM_G114(ENABLE_d_AND_den_AND_NOT_si,MGM_W86,MGM_W85);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy040ah1n12x5( clk, d, den, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy040ah_func b15fpy040ah1n12x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy040ah_func b15fpy040ah1n12x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy040ah_func b15fpy040ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy040ah_func b15fpy040ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,den_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   not MGM_G8(MGM_W7,den_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(MGM_W9,si_delay,MGM_W8);
   not MGM_G11(MGM_W10,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W10,MGM_W9);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,den_delay,MGM_W11);
   not MGM_G15(MGM_W13,si_delay);
   and MGM_G16(MGM_W14,MGM_W13,MGM_W12);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,den_delay,MGM_W16);
   not MGM_G21(MGM_W18,si_delay);
   and MGM_G22(MGM_W19,MGM_W18,MGM_W17);
   and MGM_G23(ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G24(MGM_W20,d_delay);
   and MGM_G25(MGM_W21,den_delay,MGM_W20);
   and MGM_G26(MGM_W22,si_delay,MGM_W21);
   not MGM_G27(MGM_W23,ssb_delay);
   and MGM_G28(ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W23,MGM_W22);
   not MGM_G29(MGM_W24,d_delay);
   and MGM_G30(MGM_W25,den_delay,MGM_W24);
   and MGM_G31(MGM_W26,si_delay,MGM_W25);
   and MGM_G32(ENABLE_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W26);
   not MGM_G33(MGM_W27,den_delay);
   and MGM_G34(MGM_W28,MGM_W27,d_delay);
   not MGM_G35(MGM_W29,si_delay);
   and MGM_G36(MGM_W30,MGM_W29,MGM_W28);
   not MGM_G37(MGM_W31,ssb_delay);
   and MGM_G38(ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W31,MGM_W30);
   not MGM_G39(MGM_W32,den_delay);
   and MGM_G40(MGM_W33,MGM_W32,d_delay);
   and MGM_G41(MGM_W34,si_delay,MGM_W33);
   not MGM_G42(MGM_W35,ssb_delay);
   and MGM_G43(ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W35,MGM_W34);
   and MGM_G44(MGM_W36,den_delay,d_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   not MGM_G47(MGM_W39,ssb_delay);
   and MGM_G48(ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W39,MGM_W38);
   and MGM_G49(MGM_W40,den_delay,d_delay);
   not MGM_G50(MGM_W41,si_delay);
   and MGM_G51(MGM_W42,MGM_W41,MGM_W40);
   and MGM_G52(ENABLE_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W42);
   and MGM_G53(MGM_W43,den_delay,d_delay);
   and MGM_G54(MGM_W44,si_delay,MGM_W43);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_d_AND_den_AND_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   and MGM_G57(MGM_W46,den_delay,d_delay);
   and MGM_G58(MGM_W47,si_delay,MGM_W46);
   and MGM_G59(ENABLE_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W47);
   not MGM_G60(MGM_W48,si_delay);
   and MGM_G61(MGM_W49,MGM_W48,den_delay);
   and MGM_G62(ENABLE_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   and MGM_G63(MGM_W50,si_delay,den_delay);
   and MGM_G64(ENABLE_den_AND_si_AND_ssb,ssb_delay,MGM_W50);
   not MGM_G65(MGM_W51,d_delay);
   not MGM_G66(MGM_W52,si_delay);
   and MGM_G67(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G68(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G69(MGM_W54,d_delay);
   and MGM_G70(MGM_W55,si_delay,MGM_W54);
   and MGM_G71(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W55);
   not MGM_G72(MGM_W56,si_delay);
   and MGM_G73(MGM_W57,MGM_W56,d_delay);
   and MGM_G74(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W57);
   and MGM_G75(MGM_W58,si_delay,d_delay);
   and MGM_G76(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,d_delay);
   not MGM_G78(MGM_W60,den_delay);
   and MGM_G79(MGM_W61,MGM_W60,MGM_W59);
   not MGM_G80(MGM_W62,ssb_delay);
   and MGM_G81(ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb,MGM_W62,MGM_W61);
   not MGM_G82(MGM_W63,d_delay);
   and MGM_G83(MGM_W64,den_delay,MGM_W63);
   not MGM_G84(MGM_W65,ssb_delay);
   and MGM_G85(ENABLE_NOT_d_AND_den_AND_NOT_ssb,MGM_W65,MGM_W64);
   not MGM_G86(MGM_W66,den_delay);
   and MGM_G87(MGM_W67,MGM_W66,d_delay);
   not MGM_G88(MGM_W68,ssb_delay);
   and MGM_G89(ENABLE_d_AND_NOT_den_AND_NOT_ssb,MGM_W68,MGM_W67);
   and MGM_G90(MGM_W69,den_delay,d_delay);
   not MGM_G91(MGM_W70,ssb_delay);
   and MGM_G92(ENABLE_d_AND_den_AND_NOT_ssb,MGM_W70,MGM_W69);
   not MGM_G93(MGM_W71,d_delay);
   not MGM_G94(MGM_W72,den_delay);
   and MGM_G95(MGM_W73,MGM_W72,MGM_W71);
   not MGM_G96(MGM_W74,si_delay);
   and MGM_G97(ENABLE_NOT_d_AND_NOT_den_AND_NOT_si,MGM_W74,MGM_W73);
   not MGM_G98(MGM_W75,d_delay);
   not MGM_G99(MGM_W76,den_delay);
   and MGM_G100(MGM_W77,MGM_W76,MGM_W75);
   and MGM_G101(ENABLE_NOT_d_AND_NOT_den_AND_si,si_delay,MGM_W77);
   not MGM_G102(MGM_W78,d_delay);
   and MGM_G103(MGM_W79,den_delay,MGM_W78);
   and MGM_G104(ENABLE_NOT_d_AND_den_AND_si,si_delay,MGM_W79);
   not MGM_G105(MGM_W80,den_delay);
   and MGM_G106(MGM_W81,MGM_W80,d_delay);
   not MGM_G107(MGM_W82,si_delay);
   and MGM_G108(ENABLE_d_AND_NOT_den_AND_NOT_si,MGM_W82,MGM_W81);
   not MGM_G109(MGM_W83,den_delay);
   and MGM_G110(MGM_W84,MGM_W83,d_delay);
   and MGM_G111(ENABLE_d_AND_NOT_den_AND_si,si_delay,MGM_W84);
   and MGM_G112(MGM_W85,den_delay,d_delay);
   not MGM_G113(MGM_W86,si_delay);
   and MGM_G114(ENABLE_d_AND_den_AND_NOT_si,MGM_W86,MGM_W85);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy040ah1n16x5( clk, d, den, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy040ah_func b15fpy040ah1n16x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy040ah_func b15fpy040ah1n16x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy040ah_func b15fpy040ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy040ah_func b15fpy040ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,den_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   not MGM_G8(MGM_W7,den_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(MGM_W9,si_delay,MGM_W8);
   not MGM_G11(MGM_W10,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W10,MGM_W9);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,den_delay,MGM_W11);
   not MGM_G15(MGM_W13,si_delay);
   and MGM_G16(MGM_W14,MGM_W13,MGM_W12);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,den_delay,MGM_W16);
   not MGM_G21(MGM_W18,si_delay);
   and MGM_G22(MGM_W19,MGM_W18,MGM_W17);
   and MGM_G23(ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G24(MGM_W20,d_delay);
   and MGM_G25(MGM_W21,den_delay,MGM_W20);
   and MGM_G26(MGM_W22,si_delay,MGM_W21);
   not MGM_G27(MGM_W23,ssb_delay);
   and MGM_G28(ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W23,MGM_W22);
   not MGM_G29(MGM_W24,d_delay);
   and MGM_G30(MGM_W25,den_delay,MGM_W24);
   and MGM_G31(MGM_W26,si_delay,MGM_W25);
   and MGM_G32(ENABLE_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W26);
   not MGM_G33(MGM_W27,den_delay);
   and MGM_G34(MGM_W28,MGM_W27,d_delay);
   not MGM_G35(MGM_W29,si_delay);
   and MGM_G36(MGM_W30,MGM_W29,MGM_W28);
   not MGM_G37(MGM_W31,ssb_delay);
   and MGM_G38(ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W31,MGM_W30);
   not MGM_G39(MGM_W32,den_delay);
   and MGM_G40(MGM_W33,MGM_W32,d_delay);
   and MGM_G41(MGM_W34,si_delay,MGM_W33);
   not MGM_G42(MGM_W35,ssb_delay);
   and MGM_G43(ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W35,MGM_W34);
   and MGM_G44(MGM_W36,den_delay,d_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   not MGM_G47(MGM_W39,ssb_delay);
   and MGM_G48(ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W39,MGM_W38);
   and MGM_G49(MGM_W40,den_delay,d_delay);
   not MGM_G50(MGM_W41,si_delay);
   and MGM_G51(MGM_W42,MGM_W41,MGM_W40);
   and MGM_G52(ENABLE_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W42);
   and MGM_G53(MGM_W43,den_delay,d_delay);
   and MGM_G54(MGM_W44,si_delay,MGM_W43);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_d_AND_den_AND_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   and MGM_G57(MGM_W46,den_delay,d_delay);
   and MGM_G58(MGM_W47,si_delay,MGM_W46);
   and MGM_G59(ENABLE_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W47);
   not MGM_G60(MGM_W48,si_delay);
   and MGM_G61(MGM_W49,MGM_W48,den_delay);
   and MGM_G62(ENABLE_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   and MGM_G63(MGM_W50,si_delay,den_delay);
   and MGM_G64(ENABLE_den_AND_si_AND_ssb,ssb_delay,MGM_W50);
   not MGM_G65(MGM_W51,d_delay);
   not MGM_G66(MGM_W52,si_delay);
   and MGM_G67(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G68(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G69(MGM_W54,d_delay);
   and MGM_G70(MGM_W55,si_delay,MGM_W54);
   and MGM_G71(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W55);
   not MGM_G72(MGM_W56,si_delay);
   and MGM_G73(MGM_W57,MGM_W56,d_delay);
   and MGM_G74(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W57);
   and MGM_G75(MGM_W58,si_delay,d_delay);
   and MGM_G76(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,d_delay);
   not MGM_G78(MGM_W60,den_delay);
   and MGM_G79(MGM_W61,MGM_W60,MGM_W59);
   not MGM_G80(MGM_W62,ssb_delay);
   and MGM_G81(ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb,MGM_W62,MGM_W61);
   not MGM_G82(MGM_W63,d_delay);
   and MGM_G83(MGM_W64,den_delay,MGM_W63);
   not MGM_G84(MGM_W65,ssb_delay);
   and MGM_G85(ENABLE_NOT_d_AND_den_AND_NOT_ssb,MGM_W65,MGM_W64);
   not MGM_G86(MGM_W66,den_delay);
   and MGM_G87(MGM_W67,MGM_W66,d_delay);
   not MGM_G88(MGM_W68,ssb_delay);
   and MGM_G89(ENABLE_d_AND_NOT_den_AND_NOT_ssb,MGM_W68,MGM_W67);
   and MGM_G90(MGM_W69,den_delay,d_delay);
   not MGM_G91(MGM_W70,ssb_delay);
   and MGM_G92(ENABLE_d_AND_den_AND_NOT_ssb,MGM_W70,MGM_W69);
   not MGM_G93(MGM_W71,d_delay);
   not MGM_G94(MGM_W72,den_delay);
   and MGM_G95(MGM_W73,MGM_W72,MGM_W71);
   not MGM_G96(MGM_W74,si_delay);
   and MGM_G97(ENABLE_NOT_d_AND_NOT_den_AND_NOT_si,MGM_W74,MGM_W73);
   not MGM_G98(MGM_W75,d_delay);
   not MGM_G99(MGM_W76,den_delay);
   and MGM_G100(MGM_W77,MGM_W76,MGM_W75);
   and MGM_G101(ENABLE_NOT_d_AND_NOT_den_AND_si,si_delay,MGM_W77);
   not MGM_G102(MGM_W78,d_delay);
   and MGM_G103(MGM_W79,den_delay,MGM_W78);
   and MGM_G104(ENABLE_NOT_d_AND_den_AND_si,si_delay,MGM_W79);
   not MGM_G105(MGM_W80,den_delay);
   and MGM_G106(MGM_W81,MGM_W80,d_delay);
   not MGM_G107(MGM_W82,si_delay);
   and MGM_G108(ENABLE_d_AND_NOT_den_AND_NOT_si,MGM_W82,MGM_W81);
   not MGM_G109(MGM_W83,den_delay);
   and MGM_G110(MGM_W84,MGM_W83,d_delay);
   and MGM_G111(ENABLE_d_AND_NOT_den_AND_si,si_delay,MGM_W84);
   and MGM_G112(MGM_W85,den_delay,d_delay);
   not MGM_G113(MGM_W86,si_delay);
   and MGM_G114(ENABLE_d_AND_den_AND_NOT_si,MGM_W86,MGM_W85);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_den_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_den_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fpy080ah_func( clkb, d, o, si, ssb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, si, ssb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_1( MGM_CLK0, clkb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_1( MGM_CLK0, clkb );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fpy080ah1n02x5( clkb, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n02x5_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n02x5_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n02x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n02x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy080ah1n03x5( clkb, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n03x5_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n03x5_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n03x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n03x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy080ah1n04x5( clkb, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n04x5_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n04x5_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n04x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n04x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy080ah1n06x5( clkb, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n06x5_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n06x5_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n06x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n06x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy080ah1n08x5( clkb, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n08x5_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n08x5_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n08x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n08x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy080ah1n08x7( clkb, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n08x7_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n08x7_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n08x7_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n08x7_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy080ah1n12x5( clkb, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n12x5_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n12x5_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n12x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n12x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy080ah1n12x7( clkb, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n12x7_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n12x7_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n12x7_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n12x7_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy080ah1n16x5( clkb, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n16x5_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n16x5_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n16x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n16x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy080ah1n16x7( clkb, d, o, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n16x7_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n16x7_behav_inst(.clkb(clkb),.d(d),.o(o),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy080ah_func b15fpy080ah1n16x7_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy080ah_func b15fpy080ah1n16x7_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,si_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,ssb_delay);
   and MGM_G4(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W4,d_delay);
   not MGM_G6(MGM_W5,si_delay);
   and MGM_G7(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G8(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d_delay);
   and MGM_G10(MGM_W8,si_delay,MGM_W7);
   not MGM_G11(MGM_W9,ssb_delay);
   and MGM_G12(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W9,MGM_W8);
   not MGM_G13(MGM_W10,d_delay);
   and MGM_G14(MGM_W11,si_delay,MGM_W10);
   and MGM_G15(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W11);
   not MGM_G16(MGM_W12,si_delay);
   and MGM_G17(MGM_W13,MGM_W12,d_delay);
   not MGM_G18(MGM_W14,ssb_delay);
   and MGM_G19(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W14,MGM_W13);
   not MGM_G20(MGM_W15,si_delay);
   and MGM_G21(MGM_W16,MGM_W15,d_delay);
   and MGM_G22(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W16);
   and MGM_G23(MGM_W17,si_delay,d_delay);
   not MGM_G24(MGM_W18,ssb_delay);
   and MGM_G25(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   and MGM_G26(MGM_W19,si_delay,d_delay);
   and MGM_G27(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W19);
   not MGM_G28(MGM_W20,si_delay);
   and MGM_G29(ENABLE_NOT_si_AND_ssb,ssb_delay,MGM_W20);
   and MGM_G30(ENABLE_si_AND_ssb,ssb_delay,si_delay);
   not MGM_G31(MGM_W21,d_delay);
   not MGM_G32(MGM_W22,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_NOT_ssb,MGM_W22,MGM_W21);
   not MGM_G34(MGM_W23,ssb_delay);
   and MGM_G35(ENABLE_d_AND_NOT_ssb,MGM_W23,d_delay);
   not MGM_G36(MGM_W24,d_delay);
   and MGM_G37(ENABLE_NOT_d_AND_si,si_delay,MGM_W24);
   not MGM_G38(MGM_W25,si_delay);
   and MGM_G39(ENABLE_d_AND_NOT_si,MGM_W25,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fpy200ah_func( clk, d1, d2, o1, o2, si1, si2, ssb, notifier0, notifier1 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, si1, si2, ssb, notifier0, notifier1;
   output o1, o2;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d2, si2, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, 1'b0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier1 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D1, d1, si1, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, 1'b0, 1'b0, MGM_CLK1, MGM_D1, vcc, vssx, notifier0 );
   INTCseq_cdiar2ah_0( o1, IQ1, vcc, vssx );
   INTCseq_cdiar2ah_0( o2, IQ2, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_fdw003ah_5( MGM_D0, d2, si2, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, 1'b0, 1'b0, MGM_CLK0, MGM_D0, notifier1 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk );
   INTCseq_fdw003ah_5( MGM_D1, d1, si1, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, 1'b0, 1'b0, MGM_CLK1, MGM_D1, notifier0 );
   INTCseq_cdiar2ah_0( o1, IQ1 );
   INTCseq_cdiar2ah_0( o2, IQ2 );
`endif

endmodule
`endcelldefine



`celldefine
module b15fpy200ah1n02x5( clk, d1, d2, o1, o2, si1, si2, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, si1, si2, ssb;
   output o1, o2;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy200ah_func b15fpy200ah1n02x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.d1(d1),.d2(d2),.si1(si1),.si2(si2),.notifier0(1'b0),.notifier1(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy200ah_func b15fpy200ah1n02x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.d1(d1),.d2(d2),.si1(si1),.si2(si2),.notifier0(1'b0),.notifier1(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire ssb_delay ;
   wire d1_delay ;
   wire d2_delay ;
   wire si1_delay ;
   wire si2_delay ;
   reg notifier;
   reg notifier0;
   reg notifier1;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
     notifier1 = (notifier1 !== notifier) ? notifier : ~notifier1;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy200ah_func b15fpy200ah1n02x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.d1(d1_delay),.d2(d2_delay),.si1(si1_delay),.si2(si2_delay),.notifier0(notifier0),.notifier1(notifier1),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy200ah_func b15fpy200ah1n02x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.d1(d1_delay),.d2(d2_delay),.si1(si1_delay),.si2(si2_delay),.notifier0(notifier0),.notifier1(notifier1));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d1_delay);
   not MGM_G1(MGM_W1,d2_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,si1_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,si2_delay);
   and MGM_G6(MGM_W6,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W7,ssb_delay);
   and MGM_G8(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W7,MGM_W6);
   not MGM_G9(MGM_W8,d1_delay);
   not MGM_G10(MGM_W9,d2_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   not MGM_G12(MGM_W11,si1_delay);
   and MGM_G13(MGM_W12,MGM_W11,MGM_W10);
   not MGM_G14(MGM_W13,si2_delay);
   and MGM_G15(MGM_W14,MGM_W13,MGM_W12);
   and MGM_G16(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W14);
   not MGM_G17(MGM_W15,d1_delay);
   not MGM_G18(MGM_W16,d2_delay);
   and MGM_G19(MGM_W17,MGM_W16,MGM_W15);
   not MGM_G20(MGM_W18,si1_delay);
   and MGM_G21(MGM_W19,MGM_W18,MGM_W17);
   and MGM_G22(MGM_W20,si2_delay,MGM_W19);
   not MGM_G23(MGM_W21,ssb_delay);
   and MGM_G24(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W21,MGM_W20);
   not MGM_G25(MGM_W22,d1_delay);
   not MGM_G26(MGM_W23,d2_delay);
   and MGM_G27(MGM_W24,MGM_W23,MGM_W22);
   not MGM_G28(MGM_W25,si1_delay);
   and MGM_G29(MGM_W26,MGM_W25,MGM_W24);
   and MGM_G30(MGM_W27,si2_delay,MGM_W26);
   and MGM_G31(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G32(MGM_W28,d1_delay);
   not MGM_G33(MGM_W29,d2_delay);
   and MGM_G34(MGM_W30,MGM_W29,MGM_W28);
   and MGM_G35(MGM_W31,si1_delay,MGM_W30);
   not MGM_G36(MGM_W32,si2_delay);
   and MGM_G37(MGM_W33,MGM_W32,MGM_W31);
   not MGM_G38(MGM_W34,ssb_delay);
   and MGM_G39(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W34,MGM_W33);
   not MGM_G40(MGM_W35,d1_delay);
   not MGM_G41(MGM_W36,d2_delay);
   and MGM_G42(MGM_W37,MGM_W36,MGM_W35);
   and MGM_G43(MGM_W38,si1_delay,MGM_W37);
   not MGM_G44(MGM_W39,si2_delay);
   and MGM_G45(MGM_W40,MGM_W39,MGM_W38);
   and MGM_G46(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G47(MGM_W41,d1_delay);
   not MGM_G48(MGM_W42,d2_delay);
   and MGM_G49(MGM_W43,MGM_W42,MGM_W41);
   and MGM_G50(MGM_W44,si1_delay,MGM_W43);
   and MGM_G51(MGM_W45,si2_delay,MGM_W44);
   not MGM_G52(MGM_W46,ssb_delay);
   and MGM_G53(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W46,MGM_W45);
   not MGM_G54(MGM_W47,d1_delay);
   not MGM_G55(MGM_W48,d2_delay);
   and MGM_G56(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G57(MGM_W50,si1_delay,MGM_W49);
   and MGM_G58(MGM_W51,si2_delay,MGM_W50);
   and MGM_G59(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W51);
   not MGM_G60(MGM_W52,d1_delay);
   and MGM_G61(MGM_W53,d2_delay,MGM_W52);
   not MGM_G62(MGM_W54,si1_delay);
   and MGM_G63(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G64(MGM_W56,si2_delay);
   and MGM_G65(MGM_W57,MGM_W56,MGM_W55);
   not MGM_G66(MGM_W58,ssb_delay);
   and MGM_G67(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W58,MGM_W57);
   not MGM_G68(MGM_W59,d1_delay);
   and MGM_G69(MGM_W60,d2_delay,MGM_W59);
   not MGM_G70(MGM_W61,si1_delay);
   and MGM_G71(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G72(MGM_W63,si2_delay);
   and MGM_G73(MGM_W64,MGM_W63,MGM_W62);
   and MGM_G74(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W64);
   not MGM_G75(MGM_W65,d1_delay);
   and MGM_G76(MGM_W66,d2_delay,MGM_W65);
   not MGM_G77(MGM_W67,si1_delay);
   and MGM_G78(MGM_W68,MGM_W67,MGM_W66);
   and MGM_G79(MGM_W69,si2_delay,MGM_W68);
   not MGM_G80(MGM_W70,ssb_delay);
   and MGM_G81(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W70,MGM_W69);
   not MGM_G82(MGM_W71,d1_delay);
   and MGM_G83(MGM_W72,d2_delay,MGM_W71);
   not MGM_G84(MGM_W73,si1_delay);
   and MGM_G85(MGM_W74,MGM_W73,MGM_W72);
   and MGM_G86(MGM_W75,si2_delay,MGM_W74);
   and MGM_G87(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W75);
   not MGM_G88(MGM_W76,d1_delay);
   and MGM_G89(MGM_W77,d2_delay,MGM_W76);
   and MGM_G90(MGM_W78,si1_delay,MGM_W77);
   not MGM_G91(MGM_W79,si2_delay);
   and MGM_G92(MGM_W80,MGM_W79,MGM_W78);
   not MGM_G93(MGM_W81,ssb_delay);
   and MGM_G94(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W81,MGM_W80);
   not MGM_G95(MGM_W82,d1_delay);
   and MGM_G96(MGM_W83,d2_delay,MGM_W82);
   and MGM_G97(MGM_W84,si1_delay,MGM_W83);
   not MGM_G98(MGM_W85,si2_delay);
   and MGM_G99(MGM_W86,MGM_W85,MGM_W84);
   and MGM_G100(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W86);
   not MGM_G101(MGM_W87,d1_delay);
   and MGM_G102(MGM_W88,d2_delay,MGM_W87);
   and MGM_G103(MGM_W89,si1_delay,MGM_W88);
   and MGM_G104(MGM_W90,si2_delay,MGM_W89);
   not MGM_G105(MGM_W91,ssb_delay);
   and MGM_G106(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W91,MGM_W90);
   not MGM_G107(MGM_W92,d1_delay);
   and MGM_G108(MGM_W93,d2_delay,MGM_W92);
   and MGM_G109(MGM_W94,si1_delay,MGM_W93);
   and MGM_G110(MGM_W95,si2_delay,MGM_W94);
   and MGM_G111(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W95);
   not MGM_G112(MGM_W96,d2_delay);
   and MGM_G113(MGM_W97,MGM_W96,d1_delay);
   not MGM_G114(MGM_W98,si1_delay);
   and MGM_G115(MGM_W99,MGM_W98,MGM_W97);
   not MGM_G116(MGM_W100,si2_delay);
   and MGM_G117(MGM_W101,MGM_W100,MGM_W99);
   not MGM_G118(MGM_W102,ssb_delay);
   and MGM_G119(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W102,MGM_W101);
   not MGM_G120(MGM_W103,d2_delay);
   and MGM_G121(MGM_W104,MGM_W103,d1_delay);
   not MGM_G122(MGM_W105,si1_delay);
   and MGM_G123(MGM_W106,MGM_W105,MGM_W104);
   not MGM_G124(MGM_W107,si2_delay);
   and MGM_G125(MGM_W108,MGM_W107,MGM_W106);
   and MGM_G126(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W108);
   not MGM_G127(MGM_W109,d2_delay);
   and MGM_G128(MGM_W110,MGM_W109,d1_delay);
   not MGM_G129(MGM_W111,si1_delay);
   and MGM_G130(MGM_W112,MGM_W111,MGM_W110);
   and MGM_G131(MGM_W113,si2_delay,MGM_W112);
   not MGM_G132(MGM_W114,ssb_delay);
   and MGM_G133(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W114,MGM_W113);
   not MGM_G134(MGM_W115,d2_delay);
   and MGM_G135(MGM_W116,MGM_W115,d1_delay);
   not MGM_G136(MGM_W117,si1_delay);
   and MGM_G137(MGM_W118,MGM_W117,MGM_W116);
   and MGM_G138(MGM_W119,si2_delay,MGM_W118);
   and MGM_G139(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W119);
   not MGM_G140(MGM_W120,d2_delay);
   and MGM_G141(MGM_W121,MGM_W120,d1_delay);
   and MGM_G142(MGM_W122,si1_delay,MGM_W121);
   not MGM_G143(MGM_W123,si2_delay);
   and MGM_G144(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G145(MGM_W125,ssb_delay);
   and MGM_G146(ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W125,MGM_W124);
   not MGM_G147(MGM_W126,d2_delay);
   and MGM_G148(MGM_W127,MGM_W126,d1_delay);
   and MGM_G149(MGM_W128,si1_delay,MGM_W127);
   not MGM_G150(MGM_W129,si2_delay);
   and MGM_G151(MGM_W130,MGM_W129,MGM_W128);
   and MGM_G152(ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W130);
   not MGM_G153(MGM_W131,d2_delay);
   and MGM_G154(MGM_W132,MGM_W131,d1_delay);
   and MGM_G155(MGM_W133,si1_delay,MGM_W132);
   and MGM_G156(MGM_W134,si2_delay,MGM_W133);
   not MGM_G157(MGM_W135,ssb_delay);
   and MGM_G158(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W135,MGM_W134);
   not MGM_G159(MGM_W136,d2_delay);
   and MGM_G160(MGM_W137,MGM_W136,d1_delay);
   and MGM_G161(MGM_W138,si1_delay,MGM_W137);
   and MGM_G162(MGM_W139,si2_delay,MGM_W138);
   and MGM_G163(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W139);
   and MGM_G164(MGM_W140,d2_delay,d1_delay);
   not MGM_G165(MGM_W141,si1_delay);
   and MGM_G166(MGM_W142,MGM_W141,MGM_W140);
   not MGM_G167(MGM_W143,si2_delay);
   and MGM_G168(MGM_W144,MGM_W143,MGM_W142);
   not MGM_G169(MGM_W145,ssb_delay);
   and MGM_G170(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W145,MGM_W144);
   and MGM_G171(MGM_W146,d2_delay,d1_delay);
   not MGM_G172(MGM_W147,si1_delay);
   and MGM_G173(MGM_W148,MGM_W147,MGM_W146);
   not MGM_G174(MGM_W149,si2_delay);
   and MGM_G175(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G176(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W150);
   and MGM_G177(MGM_W151,d2_delay,d1_delay);
   not MGM_G178(MGM_W152,si1_delay);
   and MGM_G179(MGM_W153,MGM_W152,MGM_W151);
   and MGM_G180(MGM_W154,si2_delay,MGM_W153);
   not MGM_G181(MGM_W155,ssb_delay);
   and MGM_G182(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W155,MGM_W154);
   and MGM_G183(MGM_W156,d2_delay,d1_delay);
   not MGM_G184(MGM_W157,si1_delay);
   and MGM_G185(MGM_W158,MGM_W157,MGM_W156);
   and MGM_G186(MGM_W159,si2_delay,MGM_W158);
   and MGM_G187(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W159);
   and MGM_G188(MGM_W160,d2_delay,d1_delay);
   and MGM_G189(MGM_W161,si1_delay,MGM_W160);
   not MGM_G190(MGM_W162,si2_delay);
   and MGM_G191(MGM_W163,MGM_W162,MGM_W161);
   not MGM_G192(MGM_W164,ssb_delay);
   and MGM_G193(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W164,MGM_W163);
   and MGM_G194(MGM_W165,d2_delay,d1_delay);
   and MGM_G195(MGM_W166,si1_delay,MGM_W165);
   not MGM_G196(MGM_W167,si2_delay);
   and MGM_G197(MGM_W168,MGM_W167,MGM_W166);
   and MGM_G198(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W168);
   and MGM_G199(MGM_W169,d2_delay,d1_delay);
   and MGM_G200(MGM_W170,si1_delay,MGM_W169);
   and MGM_G201(MGM_W171,si2_delay,MGM_W170);
   not MGM_G202(MGM_W172,ssb_delay);
   and MGM_G203(ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W172,MGM_W171);
   and MGM_G204(MGM_W173,d2_delay,d1_delay);
   and MGM_G205(MGM_W174,si1_delay,MGM_W173);
   and MGM_G206(MGM_W175,si2_delay,MGM_W174);
   and MGM_G207(ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W175);
   not MGM_G208(MGM_W176,d1_delay);
   not MGM_G209(MGM_W177,d2_delay);
   and MGM_G210(MGM_W178,MGM_W177,MGM_W176);
   not MGM_G211(MGM_W179,si1_delay);
   and MGM_G212(MGM_W180,MGM_W179,MGM_W178);
   and MGM_G213(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2,si2_delay,MGM_W180);
   not MGM_G214(MGM_W181,d1_delay);
   not MGM_G215(MGM_W182,d2_delay);
   and MGM_G216(MGM_W183,MGM_W182,MGM_W181);
   and MGM_G217(MGM_W184,si1_delay,MGM_W183);
   not MGM_G218(MGM_W185,si2_delay);
   and MGM_G219(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2,MGM_W185,MGM_W184);
   not MGM_G220(MGM_W186,d1_delay);
   not MGM_G221(MGM_W187,d2_delay);
   and MGM_G222(MGM_W188,MGM_W187,MGM_W186);
   and MGM_G223(MGM_W189,si1_delay,MGM_W188);
   and MGM_G224(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2,si2_delay,MGM_W189);
   not MGM_G225(MGM_W190,d1_delay);
   and MGM_G226(MGM_W191,d2_delay,MGM_W190);
   not MGM_G227(MGM_W192,si1_delay);
   and MGM_G228(MGM_W193,MGM_W192,MGM_W191);
   not MGM_G229(MGM_W194,si2_delay);
   and MGM_G230(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2,MGM_W194,MGM_W193);
   not MGM_G231(MGM_W195,d1_delay);
   and MGM_G232(MGM_W196,d2_delay,MGM_W195);
   and MGM_G233(MGM_W197,si1_delay,MGM_W196);
   not MGM_G234(MGM_W198,si2_delay);
   and MGM_G235(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2,MGM_W198,MGM_W197);
   not MGM_G236(MGM_W199,d1_delay);
   and MGM_G237(MGM_W200,d2_delay,MGM_W199);
   and MGM_G238(MGM_W201,si1_delay,MGM_W200);
   and MGM_G239(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2,si2_delay,MGM_W201);
   not MGM_G240(MGM_W202,d2_delay);
   and MGM_G241(MGM_W203,MGM_W202,d1_delay);
   not MGM_G242(MGM_W204,si1_delay);
   and MGM_G243(MGM_W205,MGM_W204,MGM_W203);
   not MGM_G244(MGM_W206,si2_delay);
   and MGM_G245(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2,MGM_W206,MGM_W205);
   not MGM_G246(MGM_W207,d2_delay);
   and MGM_G247(MGM_W208,MGM_W207,d1_delay);
   not MGM_G248(MGM_W209,si1_delay);
   and MGM_G249(MGM_W210,MGM_W209,MGM_W208);
   and MGM_G250(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2,si2_delay,MGM_W210);
   not MGM_G251(MGM_W211,d2_delay);
   and MGM_G252(MGM_W212,MGM_W211,d1_delay);
   and MGM_G253(MGM_W213,si1_delay,MGM_W212);
   and MGM_G254(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2,si2_delay,MGM_W213);
   and MGM_G255(MGM_W214,d2_delay,d1_delay);
   not MGM_G256(MGM_W215,si1_delay);
   and MGM_G257(MGM_W216,MGM_W215,MGM_W214);
   not MGM_G258(MGM_W217,si2_delay);
   and MGM_G259(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2,MGM_W217,MGM_W216);
   and MGM_G260(MGM_W218,d2_delay,d1_delay);
   not MGM_G261(MGM_W219,si1_delay);
   and MGM_G262(MGM_W220,MGM_W219,MGM_W218);
   and MGM_G263(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2,si2_delay,MGM_W220);
   and MGM_G264(MGM_W221,d2_delay,d1_delay);
   and MGM_G265(MGM_W222,si1_delay,MGM_W221);
   not MGM_G266(MGM_W223,si2_delay);
   and MGM_G267(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2,MGM_W223,MGM_W222);
   buf MGM_G268(ENABLE_ssb,ssb_delay);
   not MGM_G269(ENABLE_NOT_ssb,ssb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk,0.0,0,notifier);
      
      $width(posedge clk,0.0,0,notifier);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,negedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,posedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy200ah1n03x5( clk, d1, d2, o1, o2, si1, si2, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, si1, si2, ssb;
   output o1, o2;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy200ah_func b15fpy200ah1n03x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.d1(d1),.d2(d2),.si1(si1),.si2(si2),.notifier0(1'b0),.notifier1(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy200ah_func b15fpy200ah1n03x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.d1(d1),.d2(d2),.si1(si1),.si2(si2),.notifier0(1'b0),.notifier1(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire ssb_delay ;
   wire d1_delay ;
   wire d2_delay ;
   wire si1_delay ;
   wire si2_delay ;
   reg notifier;
   reg notifier0;
   reg notifier1;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
     notifier1 = (notifier1 !== notifier) ? notifier : ~notifier1;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy200ah_func b15fpy200ah1n03x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.d1(d1_delay),.d2(d2_delay),.si1(si1_delay),.si2(si2_delay),.notifier0(notifier0),.notifier1(notifier1),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy200ah_func b15fpy200ah1n03x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.d1(d1_delay),.d2(d2_delay),.si1(si1_delay),.si2(si2_delay),.notifier0(notifier0),.notifier1(notifier1));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d1_delay);
   not MGM_G1(MGM_W1,d2_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,si1_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,si2_delay);
   and MGM_G6(MGM_W6,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W7,ssb_delay);
   and MGM_G8(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W7,MGM_W6);
   not MGM_G9(MGM_W8,d1_delay);
   not MGM_G10(MGM_W9,d2_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   not MGM_G12(MGM_W11,si1_delay);
   and MGM_G13(MGM_W12,MGM_W11,MGM_W10);
   not MGM_G14(MGM_W13,si2_delay);
   and MGM_G15(MGM_W14,MGM_W13,MGM_W12);
   and MGM_G16(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W14);
   not MGM_G17(MGM_W15,d1_delay);
   not MGM_G18(MGM_W16,d2_delay);
   and MGM_G19(MGM_W17,MGM_W16,MGM_W15);
   not MGM_G20(MGM_W18,si1_delay);
   and MGM_G21(MGM_W19,MGM_W18,MGM_W17);
   and MGM_G22(MGM_W20,si2_delay,MGM_W19);
   not MGM_G23(MGM_W21,ssb_delay);
   and MGM_G24(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W21,MGM_W20);
   not MGM_G25(MGM_W22,d1_delay);
   not MGM_G26(MGM_W23,d2_delay);
   and MGM_G27(MGM_W24,MGM_W23,MGM_W22);
   not MGM_G28(MGM_W25,si1_delay);
   and MGM_G29(MGM_W26,MGM_W25,MGM_W24);
   and MGM_G30(MGM_W27,si2_delay,MGM_W26);
   and MGM_G31(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G32(MGM_W28,d1_delay);
   not MGM_G33(MGM_W29,d2_delay);
   and MGM_G34(MGM_W30,MGM_W29,MGM_W28);
   and MGM_G35(MGM_W31,si1_delay,MGM_W30);
   not MGM_G36(MGM_W32,si2_delay);
   and MGM_G37(MGM_W33,MGM_W32,MGM_W31);
   not MGM_G38(MGM_W34,ssb_delay);
   and MGM_G39(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W34,MGM_W33);
   not MGM_G40(MGM_W35,d1_delay);
   not MGM_G41(MGM_W36,d2_delay);
   and MGM_G42(MGM_W37,MGM_W36,MGM_W35);
   and MGM_G43(MGM_W38,si1_delay,MGM_W37);
   not MGM_G44(MGM_W39,si2_delay);
   and MGM_G45(MGM_W40,MGM_W39,MGM_W38);
   and MGM_G46(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G47(MGM_W41,d1_delay);
   not MGM_G48(MGM_W42,d2_delay);
   and MGM_G49(MGM_W43,MGM_W42,MGM_W41);
   and MGM_G50(MGM_W44,si1_delay,MGM_W43);
   and MGM_G51(MGM_W45,si2_delay,MGM_W44);
   not MGM_G52(MGM_W46,ssb_delay);
   and MGM_G53(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W46,MGM_W45);
   not MGM_G54(MGM_W47,d1_delay);
   not MGM_G55(MGM_W48,d2_delay);
   and MGM_G56(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G57(MGM_W50,si1_delay,MGM_W49);
   and MGM_G58(MGM_W51,si2_delay,MGM_W50);
   and MGM_G59(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W51);
   not MGM_G60(MGM_W52,d1_delay);
   and MGM_G61(MGM_W53,d2_delay,MGM_W52);
   not MGM_G62(MGM_W54,si1_delay);
   and MGM_G63(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G64(MGM_W56,si2_delay);
   and MGM_G65(MGM_W57,MGM_W56,MGM_W55);
   not MGM_G66(MGM_W58,ssb_delay);
   and MGM_G67(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W58,MGM_W57);
   not MGM_G68(MGM_W59,d1_delay);
   and MGM_G69(MGM_W60,d2_delay,MGM_W59);
   not MGM_G70(MGM_W61,si1_delay);
   and MGM_G71(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G72(MGM_W63,si2_delay);
   and MGM_G73(MGM_W64,MGM_W63,MGM_W62);
   and MGM_G74(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W64);
   not MGM_G75(MGM_W65,d1_delay);
   and MGM_G76(MGM_W66,d2_delay,MGM_W65);
   not MGM_G77(MGM_W67,si1_delay);
   and MGM_G78(MGM_W68,MGM_W67,MGM_W66);
   and MGM_G79(MGM_W69,si2_delay,MGM_W68);
   not MGM_G80(MGM_W70,ssb_delay);
   and MGM_G81(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W70,MGM_W69);
   not MGM_G82(MGM_W71,d1_delay);
   and MGM_G83(MGM_W72,d2_delay,MGM_W71);
   not MGM_G84(MGM_W73,si1_delay);
   and MGM_G85(MGM_W74,MGM_W73,MGM_W72);
   and MGM_G86(MGM_W75,si2_delay,MGM_W74);
   and MGM_G87(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W75);
   not MGM_G88(MGM_W76,d1_delay);
   and MGM_G89(MGM_W77,d2_delay,MGM_W76);
   and MGM_G90(MGM_W78,si1_delay,MGM_W77);
   not MGM_G91(MGM_W79,si2_delay);
   and MGM_G92(MGM_W80,MGM_W79,MGM_W78);
   not MGM_G93(MGM_W81,ssb_delay);
   and MGM_G94(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W81,MGM_W80);
   not MGM_G95(MGM_W82,d1_delay);
   and MGM_G96(MGM_W83,d2_delay,MGM_W82);
   and MGM_G97(MGM_W84,si1_delay,MGM_W83);
   not MGM_G98(MGM_W85,si2_delay);
   and MGM_G99(MGM_W86,MGM_W85,MGM_W84);
   and MGM_G100(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W86);
   not MGM_G101(MGM_W87,d1_delay);
   and MGM_G102(MGM_W88,d2_delay,MGM_W87);
   and MGM_G103(MGM_W89,si1_delay,MGM_W88);
   and MGM_G104(MGM_W90,si2_delay,MGM_W89);
   not MGM_G105(MGM_W91,ssb_delay);
   and MGM_G106(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W91,MGM_W90);
   not MGM_G107(MGM_W92,d1_delay);
   and MGM_G108(MGM_W93,d2_delay,MGM_W92);
   and MGM_G109(MGM_W94,si1_delay,MGM_W93);
   and MGM_G110(MGM_W95,si2_delay,MGM_W94);
   and MGM_G111(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W95);
   not MGM_G112(MGM_W96,d2_delay);
   and MGM_G113(MGM_W97,MGM_W96,d1_delay);
   not MGM_G114(MGM_W98,si1_delay);
   and MGM_G115(MGM_W99,MGM_W98,MGM_W97);
   not MGM_G116(MGM_W100,si2_delay);
   and MGM_G117(MGM_W101,MGM_W100,MGM_W99);
   not MGM_G118(MGM_W102,ssb_delay);
   and MGM_G119(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W102,MGM_W101);
   not MGM_G120(MGM_W103,d2_delay);
   and MGM_G121(MGM_W104,MGM_W103,d1_delay);
   not MGM_G122(MGM_W105,si1_delay);
   and MGM_G123(MGM_W106,MGM_W105,MGM_W104);
   not MGM_G124(MGM_W107,si2_delay);
   and MGM_G125(MGM_W108,MGM_W107,MGM_W106);
   and MGM_G126(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W108);
   not MGM_G127(MGM_W109,d2_delay);
   and MGM_G128(MGM_W110,MGM_W109,d1_delay);
   not MGM_G129(MGM_W111,si1_delay);
   and MGM_G130(MGM_W112,MGM_W111,MGM_W110);
   and MGM_G131(MGM_W113,si2_delay,MGM_W112);
   not MGM_G132(MGM_W114,ssb_delay);
   and MGM_G133(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W114,MGM_W113);
   not MGM_G134(MGM_W115,d2_delay);
   and MGM_G135(MGM_W116,MGM_W115,d1_delay);
   not MGM_G136(MGM_W117,si1_delay);
   and MGM_G137(MGM_W118,MGM_W117,MGM_W116);
   and MGM_G138(MGM_W119,si2_delay,MGM_W118);
   and MGM_G139(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W119);
   not MGM_G140(MGM_W120,d2_delay);
   and MGM_G141(MGM_W121,MGM_W120,d1_delay);
   and MGM_G142(MGM_W122,si1_delay,MGM_W121);
   not MGM_G143(MGM_W123,si2_delay);
   and MGM_G144(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G145(MGM_W125,ssb_delay);
   and MGM_G146(ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W125,MGM_W124);
   not MGM_G147(MGM_W126,d2_delay);
   and MGM_G148(MGM_W127,MGM_W126,d1_delay);
   and MGM_G149(MGM_W128,si1_delay,MGM_W127);
   not MGM_G150(MGM_W129,si2_delay);
   and MGM_G151(MGM_W130,MGM_W129,MGM_W128);
   and MGM_G152(ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W130);
   not MGM_G153(MGM_W131,d2_delay);
   and MGM_G154(MGM_W132,MGM_W131,d1_delay);
   and MGM_G155(MGM_W133,si1_delay,MGM_W132);
   and MGM_G156(MGM_W134,si2_delay,MGM_W133);
   not MGM_G157(MGM_W135,ssb_delay);
   and MGM_G158(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W135,MGM_W134);
   not MGM_G159(MGM_W136,d2_delay);
   and MGM_G160(MGM_W137,MGM_W136,d1_delay);
   and MGM_G161(MGM_W138,si1_delay,MGM_W137);
   and MGM_G162(MGM_W139,si2_delay,MGM_W138);
   and MGM_G163(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W139);
   and MGM_G164(MGM_W140,d2_delay,d1_delay);
   not MGM_G165(MGM_W141,si1_delay);
   and MGM_G166(MGM_W142,MGM_W141,MGM_W140);
   not MGM_G167(MGM_W143,si2_delay);
   and MGM_G168(MGM_W144,MGM_W143,MGM_W142);
   not MGM_G169(MGM_W145,ssb_delay);
   and MGM_G170(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W145,MGM_W144);
   and MGM_G171(MGM_W146,d2_delay,d1_delay);
   not MGM_G172(MGM_W147,si1_delay);
   and MGM_G173(MGM_W148,MGM_W147,MGM_W146);
   not MGM_G174(MGM_W149,si2_delay);
   and MGM_G175(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G176(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W150);
   and MGM_G177(MGM_W151,d2_delay,d1_delay);
   not MGM_G178(MGM_W152,si1_delay);
   and MGM_G179(MGM_W153,MGM_W152,MGM_W151);
   and MGM_G180(MGM_W154,si2_delay,MGM_W153);
   not MGM_G181(MGM_W155,ssb_delay);
   and MGM_G182(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W155,MGM_W154);
   and MGM_G183(MGM_W156,d2_delay,d1_delay);
   not MGM_G184(MGM_W157,si1_delay);
   and MGM_G185(MGM_W158,MGM_W157,MGM_W156);
   and MGM_G186(MGM_W159,si2_delay,MGM_W158);
   and MGM_G187(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W159);
   and MGM_G188(MGM_W160,d2_delay,d1_delay);
   and MGM_G189(MGM_W161,si1_delay,MGM_W160);
   not MGM_G190(MGM_W162,si2_delay);
   and MGM_G191(MGM_W163,MGM_W162,MGM_W161);
   not MGM_G192(MGM_W164,ssb_delay);
   and MGM_G193(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W164,MGM_W163);
   and MGM_G194(MGM_W165,d2_delay,d1_delay);
   and MGM_G195(MGM_W166,si1_delay,MGM_W165);
   not MGM_G196(MGM_W167,si2_delay);
   and MGM_G197(MGM_W168,MGM_W167,MGM_W166);
   and MGM_G198(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W168);
   and MGM_G199(MGM_W169,d2_delay,d1_delay);
   and MGM_G200(MGM_W170,si1_delay,MGM_W169);
   and MGM_G201(MGM_W171,si2_delay,MGM_W170);
   not MGM_G202(MGM_W172,ssb_delay);
   and MGM_G203(ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W172,MGM_W171);
   and MGM_G204(MGM_W173,d2_delay,d1_delay);
   and MGM_G205(MGM_W174,si1_delay,MGM_W173);
   and MGM_G206(MGM_W175,si2_delay,MGM_W174);
   and MGM_G207(ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W175);
   not MGM_G208(MGM_W176,d1_delay);
   not MGM_G209(MGM_W177,d2_delay);
   and MGM_G210(MGM_W178,MGM_W177,MGM_W176);
   not MGM_G211(MGM_W179,si1_delay);
   and MGM_G212(MGM_W180,MGM_W179,MGM_W178);
   and MGM_G213(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2,si2_delay,MGM_W180);
   not MGM_G214(MGM_W181,d1_delay);
   not MGM_G215(MGM_W182,d2_delay);
   and MGM_G216(MGM_W183,MGM_W182,MGM_W181);
   and MGM_G217(MGM_W184,si1_delay,MGM_W183);
   not MGM_G218(MGM_W185,si2_delay);
   and MGM_G219(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2,MGM_W185,MGM_W184);
   not MGM_G220(MGM_W186,d1_delay);
   not MGM_G221(MGM_W187,d2_delay);
   and MGM_G222(MGM_W188,MGM_W187,MGM_W186);
   and MGM_G223(MGM_W189,si1_delay,MGM_W188);
   and MGM_G224(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2,si2_delay,MGM_W189);
   not MGM_G225(MGM_W190,d1_delay);
   and MGM_G226(MGM_W191,d2_delay,MGM_W190);
   not MGM_G227(MGM_W192,si1_delay);
   and MGM_G228(MGM_W193,MGM_W192,MGM_W191);
   not MGM_G229(MGM_W194,si2_delay);
   and MGM_G230(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2,MGM_W194,MGM_W193);
   not MGM_G231(MGM_W195,d1_delay);
   and MGM_G232(MGM_W196,d2_delay,MGM_W195);
   and MGM_G233(MGM_W197,si1_delay,MGM_W196);
   not MGM_G234(MGM_W198,si2_delay);
   and MGM_G235(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2,MGM_W198,MGM_W197);
   not MGM_G236(MGM_W199,d1_delay);
   and MGM_G237(MGM_W200,d2_delay,MGM_W199);
   and MGM_G238(MGM_W201,si1_delay,MGM_W200);
   and MGM_G239(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2,si2_delay,MGM_W201);
   not MGM_G240(MGM_W202,d2_delay);
   and MGM_G241(MGM_W203,MGM_W202,d1_delay);
   not MGM_G242(MGM_W204,si1_delay);
   and MGM_G243(MGM_W205,MGM_W204,MGM_W203);
   not MGM_G244(MGM_W206,si2_delay);
   and MGM_G245(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2,MGM_W206,MGM_W205);
   not MGM_G246(MGM_W207,d2_delay);
   and MGM_G247(MGM_W208,MGM_W207,d1_delay);
   not MGM_G248(MGM_W209,si1_delay);
   and MGM_G249(MGM_W210,MGM_W209,MGM_W208);
   and MGM_G250(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2,si2_delay,MGM_W210);
   not MGM_G251(MGM_W211,d2_delay);
   and MGM_G252(MGM_W212,MGM_W211,d1_delay);
   and MGM_G253(MGM_W213,si1_delay,MGM_W212);
   and MGM_G254(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2,si2_delay,MGM_W213);
   and MGM_G255(MGM_W214,d2_delay,d1_delay);
   not MGM_G256(MGM_W215,si1_delay);
   and MGM_G257(MGM_W216,MGM_W215,MGM_W214);
   not MGM_G258(MGM_W217,si2_delay);
   and MGM_G259(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2,MGM_W217,MGM_W216);
   and MGM_G260(MGM_W218,d2_delay,d1_delay);
   not MGM_G261(MGM_W219,si1_delay);
   and MGM_G262(MGM_W220,MGM_W219,MGM_W218);
   and MGM_G263(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2,si2_delay,MGM_W220);
   and MGM_G264(MGM_W221,d2_delay,d1_delay);
   and MGM_G265(MGM_W222,si1_delay,MGM_W221);
   not MGM_G266(MGM_W223,si2_delay);
   and MGM_G267(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2,MGM_W223,MGM_W222);
   buf MGM_G268(ENABLE_ssb,ssb_delay);
   not MGM_G269(ENABLE_NOT_ssb,ssb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk,0.0,0,notifier);
      
      $width(posedge clk,0.0,0,notifier);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,negedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,posedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy200ah1n04x5( clk, d1, d2, o1, o2, si1, si2, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, si1, si2, ssb;
   output o1, o2;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy200ah_func b15fpy200ah1n04x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.d1(d1),.d2(d2),.si1(si1),.si2(si2),.notifier0(1'b0),.notifier1(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy200ah_func b15fpy200ah1n04x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.d1(d1),.d2(d2),.si1(si1),.si2(si2),.notifier0(1'b0),.notifier1(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire ssb_delay ;
   wire d1_delay ;
   wire d2_delay ;
   wire si1_delay ;
   wire si2_delay ;
   reg notifier;
   reg notifier0;
   reg notifier1;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
     notifier1 = (notifier1 !== notifier) ? notifier : ~notifier1;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy200ah_func b15fpy200ah1n04x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.d1(d1_delay),.d2(d2_delay),.si1(si1_delay),.si2(si2_delay),.notifier0(notifier0),.notifier1(notifier1),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy200ah_func b15fpy200ah1n04x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.d1(d1_delay),.d2(d2_delay),.si1(si1_delay),.si2(si2_delay),.notifier0(notifier0),.notifier1(notifier1));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d1_delay);
   not MGM_G1(MGM_W1,d2_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,si1_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,si2_delay);
   and MGM_G6(MGM_W6,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W7,ssb_delay);
   and MGM_G8(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W7,MGM_W6);
   not MGM_G9(MGM_W8,d1_delay);
   not MGM_G10(MGM_W9,d2_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   not MGM_G12(MGM_W11,si1_delay);
   and MGM_G13(MGM_W12,MGM_W11,MGM_W10);
   not MGM_G14(MGM_W13,si2_delay);
   and MGM_G15(MGM_W14,MGM_W13,MGM_W12);
   and MGM_G16(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W14);
   not MGM_G17(MGM_W15,d1_delay);
   not MGM_G18(MGM_W16,d2_delay);
   and MGM_G19(MGM_W17,MGM_W16,MGM_W15);
   not MGM_G20(MGM_W18,si1_delay);
   and MGM_G21(MGM_W19,MGM_W18,MGM_W17);
   and MGM_G22(MGM_W20,si2_delay,MGM_W19);
   not MGM_G23(MGM_W21,ssb_delay);
   and MGM_G24(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W21,MGM_W20);
   not MGM_G25(MGM_W22,d1_delay);
   not MGM_G26(MGM_W23,d2_delay);
   and MGM_G27(MGM_W24,MGM_W23,MGM_W22);
   not MGM_G28(MGM_W25,si1_delay);
   and MGM_G29(MGM_W26,MGM_W25,MGM_W24);
   and MGM_G30(MGM_W27,si2_delay,MGM_W26);
   and MGM_G31(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G32(MGM_W28,d1_delay);
   not MGM_G33(MGM_W29,d2_delay);
   and MGM_G34(MGM_W30,MGM_W29,MGM_W28);
   and MGM_G35(MGM_W31,si1_delay,MGM_W30);
   not MGM_G36(MGM_W32,si2_delay);
   and MGM_G37(MGM_W33,MGM_W32,MGM_W31);
   not MGM_G38(MGM_W34,ssb_delay);
   and MGM_G39(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W34,MGM_W33);
   not MGM_G40(MGM_W35,d1_delay);
   not MGM_G41(MGM_W36,d2_delay);
   and MGM_G42(MGM_W37,MGM_W36,MGM_W35);
   and MGM_G43(MGM_W38,si1_delay,MGM_W37);
   not MGM_G44(MGM_W39,si2_delay);
   and MGM_G45(MGM_W40,MGM_W39,MGM_W38);
   and MGM_G46(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G47(MGM_W41,d1_delay);
   not MGM_G48(MGM_W42,d2_delay);
   and MGM_G49(MGM_W43,MGM_W42,MGM_W41);
   and MGM_G50(MGM_W44,si1_delay,MGM_W43);
   and MGM_G51(MGM_W45,si2_delay,MGM_W44);
   not MGM_G52(MGM_W46,ssb_delay);
   and MGM_G53(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W46,MGM_W45);
   not MGM_G54(MGM_W47,d1_delay);
   not MGM_G55(MGM_W48,d2_delay);
   and MGM_G56(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G57(MGM_W50,si1_delay,MGM_W49);
   and MGM_G58(MGM_W51,si2_delay,MGM_W50);
   and MGM_G59(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W51);
   not MGM_G60(MGM_W52,d1_delay);
   and MGM_G61(MGM_W53,d2_delay,MGM_W52);
   not MGM_G62(MGM_W54,si1_delay);
   and MGM_G63(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G64(MGM_W56,si2_delay);
   and MGM_G65(MGM_W57,MGM_W56,MGM_W55);
   not MGM_G66(MGM_W58,ssb_delay);
   and MGM_G67(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W58,MGM_W57);
   not MGM_G68(MGM_W59,d1_delay);
   and MGM_G69(MGM_W60,d2_delay,MGM_W59);
   not MGM_G70(MGM_W61,si1_delay);
   and MGM_G71(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G72(MGM_W63,si2_delay);
   and MGM_G73(MGM_W64,MGM_W63,MGM_W62);
   and MGM_G74(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W64);
   not MGM_G75(MGM_W65,d1_delay);
   and MGM_G76(MGM_W66,d2_delay,MGM_W65);
   not MGM_G77(MGM_W67,si1_delay);
   and MGM_G78(MGM_W68,MGM_W67,MGM_W66);
   and MGM_G79(MGM_W69,si2_delay,MGM_W68);
   not MGM_G80(MGM_W70,ssb_delay);
   and MGM_G81(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W70,MGM_W69);
   not MGM_G82(MGM_W71,d1_delay);
   and MGM_G83(MGM_W72,d2_delay,MGM_W71);
   not MGM_G84(MGM_W73,si1_delay);
   and MGM_G85(MGM_W74,MGM_W73,MGM_W72);
   and MGM_G86(MGM_W75,si2_delay,MGM_W74);
   and MGM_G87(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W75);
   not MGM_G88(MGM_W76,d1_delay);
   and MGM_G89(MGM_W77,d2_delay,MGM_W76);
   and MGM_G90(MGM_W78,si1_delay,MGM_W77);
   not MGM_G91(MGM_W79,si2_delay);
   and MGM_G92(MGM_W80,MGM_W79,MGM_W78);
   not MGM_G93(MGM_W81,ssb_delay);
   and MGM_G94(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W81,MGM_W80);
   not MGM_G95(MGM_W82,d1_delay);
   and MGM_G96(MGM_W83,d2_delay,MGM_W82);
   and MGM_G97(MGM_W84,si1_delay,MGM_W83);
   not MGM_G98(MGM_W85,si2_delay);
   and MGM_G99(MGM_W86,MGM_W85,MGM_W84);
   and MGM_G100(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W86);
   not MGM_G101(MGM_W87,d1_delay);
   and MGM_G102(MGM_W88,d2_delay,MGM_W87);
   and MGM_G103(MGM_W89,si1_delay,MGM_W88);
   and MGM_G104(MGM_W90,si2_delay,MGM_W89);
   not MGM_G105(MGM_W91,ssb_delay);
   and MGM_G106(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W91,MGM_W90);
   not MGM_G107(MGM_W92,d1_delay);
   and MGM_G108(MGM_W93,d2_delay,MGM_W92);
   and MGM_G109(MGM_W94,si1_delay,MGM_W93);
   and MGM_G110(MGM_W95,si2_delay,MGM_W94);
   and MGM_G111(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W95);
   not MGM_G112(MGM_W96,d2_delay);
   and MGM_G113(MGM_W97,MGM_W96,d1_delay);
   not MGM_G114(MGM_W98,si1_delay);
   and MGM_G115(MGM_W99,MGM_W98,MGM_W97);
   not MGM_G116(MGM_W100,si2_delay);
   and MGM_G117(MGM_W101,MGM_W100,MGM_W99);
   not MGM_G118(MGM_W102,ssb_delay);
   and MGM_G119(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W102,MGM_W101);
   not MGM_G120(MGM_W103,d2_delay);
   and MGM_G121(MGM_W104,MGM_W103,d1_delay);
   not MGM_G122(MGM_W105,si1_delay);
   and MGM_G123(MGM_W106,MGM_W105,MGM_W104);
   not MGM_G124(MGM_W107,si2_delay);
   and MGM_G125(MGM_W108,MGM_W107,MGM_W106);
   and MGM_G126(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W108);
   not MGM_G127(MGM_W109,d2_delay);
   and MGM_G128(MGM_W110,MGM_W109,d1_delay);
   not MGM_G129(MGM_W111,si1_delay);
   and MGM_G130(MGM_W112,MGM_W111,MGM_W110);
   and MGM_G131(MGM_W113,si2_delay,MGM_W112);
   not MGM_G132(MGM_W114,ssb_delay);
   and MGM_G133(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W114,MGM_W113);
   not MGM_G134(MGM_W115,d2_delay);
   and MGM_G135(MGM_W116,MGM_W115,d1_delay);
   not MGM_G136(MGM_W117,si1_delay);
   and MGM_G137(MGM_W118,MGM_W117,MGM_W116);
   and MGM_G138(MGM_W119,si2_delay,MGM_W118);
   and MGM_G139(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W119);
   not MGM_G140(MGM_W120,d2_delay);
   and MGM_G141(MGM_W121,MGM_W120,d1_delay);
   and MGM_G142(MGM_W122,si1_delay,MGM_W121);
   not MGM_G143(MGM_W123,si2_delay);
   and MGM_G144(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G145(MGM_W125,ssb_delay);
   and MGM_G146(ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W125,MGM_W124);
   not MGM_G147(MGM_W126,d2_delay);
   and MGM_G148(MGM_W127,MGM_W126,d1_delay);
   and MGM_G149(MGM_W128,si1_delay,MGM_W127);
   not MGM_G150(MGM_W129,si2_delay);
   and MGM_G151(MGM_W130,MGM_W129,MGM_W128);
   and MGM_G152(ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W130);
   not MGM_G153(MGM_W131,d2_delay);
   and MGM_G154(MGM_W132,MGM_W131,d1_delay);
   and MGM_G155(MGM_W133,si1_delay,MGM_W132);
   and MGM_G156(MGM_W134,si2_delay,MGM_W133);
   not MGM_G157(MGM_W135,ssb_delay);
   and MGM_G158(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W135,MGM_W134);
   not MGM_G159(MGM_W136,d2_delay);
   and MGM_G160(MGM_W137,MGM_W136,d1_delay);
   and MGM_G161(MGM_W138,si1_delay,MGM_W137);
   and MGM_G162(MGM_W139,si2_delay,MGM_W138);
   and MGM_G163(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W139);
   and MGM_G164(MGM_W140,d2_delay,d1_delay);
   not MGM_G165(MGM_W141,si1_delay);
   and MGM_G166(MGM_W142,MGM_W141,MGM_W140);
   not MGM_G167(MGM_W143,si2_delay);
   and MGM_G168(MGM_W144,MGM_W143,MGM_W142);
   not MGM_G169(MGM_W145,ssb_delay);
   and MGM_G170(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W145,MGM_W144);
   and MGM_G171(MGM_W146,d2_delay,d1_delay);
   not MGM_G172(MGM_W147,si1_delay);
   and MGM_G173(MGM_W148,MGM_W147,MGM_W146);
   not MGM_G174(MGM_W149,si2_delay);
   and MGM_G175(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G176(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W150);
   and MGM_G177(MGM_W151,d2_delay,d1_delay);
   not MGM_G178(MGM_W152,si1_delay);
   and MGM_G179(MGM_W153,MGM_W152,MGM_W151);
   and MGM_G180(MGM_W154,si2_delay,MGM_W153);
   not MGM_G181(MGM_W155,ssb_delay);
   and MGM_G182(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W155,MGM_W154);
   and MGM_G183(MGM_W156,d2_delay,d1_delay);
   not MGM_G184(MGM_W157,si1_delay);
   and MGM_G185(MGM_W158,MGM_W157,MGM_W156);
   and MGM_G186(MGM_W159,si2_delay,MGM_W158);
   and MGM_G187(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W159);
   and MGM_G188(MGM_W160,d2_delay,d1_delay);
   and MGM_G189(MGM_W161,si1_delay,MGM_W160);
   not MGM_G190(MGM_W162,si2_delay);
   and MGM_G191(MGM_W163,MGM_W162,MGM_W161);
   not MGM_G192(MGM_W164,ssb_delay);
   and MGM_G193(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W164,MGM_W163);
   and MGM_G194(MGM_W165,d2_delay,d1_delay);
   and MGM_G195(MGM_W166,si1_delay,MGM_W165);
   not MGM_G196(MGM_W167,si2_delay);
   and MGM_G197(MGM_W168,MGM_W167,MGM_W166);
   and MGM_G198(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W168);
   and MGM_G199(MGM_W169,d2_delay,d1_delay);
   and MGM_G200(MGM_W170,si1_delay,MGM_W169);
   and MGM_G201(MGM_W171,si2_delay,MGM_W170);
   not MGM_G202(MGM_W172,ssb_delay);
   and MGM_G203(ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W172,MGM_W171);
   and MGM_G204(MGM_W173,d2_delay,d1_delay);
   and MGM_G205(MGM_W174,si1_delay,MGM_W173);
   and MGM_G206(MGM_W175,si2_delay,MGM_W174);
   and MGM_G207(ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W175);
   not MGM_G208(MGM_W176,d1_delay);
   not MGM_G209(MGM_W177,d2_delay);
   and MGM_G210(MGM_W178,MGM_W177,MGM_W176);
   not MGM_G211(MGM_W179,si1_delay);
   and MGM_G212(MGM_W180,MGM_W179,MGM_W178);
   and MGM_G213(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2,si2_delay,MGM_W180);
   not MGM_G214(MGM_W181,d1_delay);
   not MGM_G215(MGM_W182,d2_delay);
   and MGM_G216(MGM_W183,MGM_W182,MGM_W181);
   and MGM_G217(MGM_W184,si1_delay,MGM_W183);
   not MGM_G218(MGM_W185,si2_delay);
   and MGM_G219(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2,MGM_W185,MGM_W184);
   not MGM_G220(MGM_W186,d1_delay);
   not MGM_G221(MGM_W187,d2_delay);
   and MGM_G222(MGM_W188,MGM_W187,MGM_W186);
   and MGM_G223(MGM_W189,si1_delay,MGM_W188);
   and MGM_G224(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2,si2_delay,MGM_W189);
   not MGM_G225(MGM_W190,d1_delay);
   and MGM_G226(MGM_W191,d2_delay,MGM_W190);
   not MGM_G227(MGM_W192,si1_delay);
   and MGM_G228(MGM_W193,MGM_W192,MGM_W191);
   not MGM_G229(MGM_W194,si2_delay);
   and MGM_G230(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2,MGM_W194,MGM_W193);
   not MGM_G231(MGM_W195,d1_delay);
   and MGM_G232(MGM_W196,d2_delay,MGM_W195);
   and MGM_G233(MGM_W197,si1_delay,MGM_W196);
   not MGM_G234(MGM_W198,si2_delay);
   and MGM_G235(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2,MGM_W198,MGM_W197);
   not MGM_G236(MGM_W199,d1_delay);
   and MGM_G237(MGM_W200,d2_delay,MGM_W199);
   and MGM_G238(MGM_W201,si1_delay,MGM_W200);
   and MGM_G239(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2,si2_delay,MGM_W201);
   not MGM_G240(MGM_W202,d2_delay);
   and MGM_G241(MGM_W203,MGM_W202,d1_delay);
   not MGM_G242(MGM_W204,si1_delay);
   and MGM_G243(MGM_W205,MGM_W204,MGM_W203);
   not MGM_G244(MGM_W206,si2_delay);
   and MGM_G245(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2,MGM_W206,MGM_W205);
   not MGM_G246(MGM_W207,d2_delay);
   and MGM_G247(MGM_W208,MGM_W207,d1_delay);
   not MGM_G248(MGM_W209,si1_delay);
   and MGM_G249(MGM_W210,MGM_W209,MGM_W208);
   and MGM_G250(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2,si2_delay,MGM_W210);
   not MGM_G251(MGM_W211,d2_delay);
   and MGM_G252(MGM_W212,MGM_W211,d1_delay);
   and MGM_G253(MGM_W213,si1_delay,MGM_W212);
   and MGM_G254(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2,si2_delay,MGM_W213);
   and MGM_G255(MGM_W214,d2_delay,d1_delay);
   not MGM_G256(MGM_W215,si1_delay);
   and MGM_G257(MGM_W216,MGM_W215,MGM_W214);
   not MGM_G258(MGM_W217,si2_delay);
   and MGM_G259(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2,MGM_W217,MGM_W216);
   and MGM_G260(MGM_W218,d2_delay,d1_delay);
   not MGM_G261(MGM_W219,si1_delay);
   and MGM_G262(MGM_W220,MGM_W219,MGM_W218);
   and MGM_G263(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2,si2_delay,MGM_W220);
   and MGM_G264(MGM_W221,d2_delay,d1_delay);
   and MGM_G265(MGM_W222,si1_delay,MGM_W221);
   not MGM_G266(MGM_W223,si2_delay);
   and MGM_G267(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2,MGM_W223,MGM_W222);
   buf MGM_G268(ENABLE_ssb,ssb_delay);
   not MGM_G269(ENABLE_NOT_ssb,ssb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk,0.0,0,notifier);
      
      $width(posedge clk,0.0,0,notifier);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,negedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,posedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy200ah1n08x5( clk, d1, d2, o1, o2, si1, si2, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, si1, si2, ssb;
   output o1, o2;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy200ah_func b15fpy200ah1n08x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.d1(d1),.d2(d2),.si1(si1),.si2(si2),.notifier0(1'b0),.notifier1(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy200ah_func b15fpy200ah1n08x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.d1(d1),.d2(d2),.si1(si1),.si2(si2),.notifier0(1'b0),.notifier1(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire ssb_delay ;
   wire d1_delay ;
   wire d2_delay ;
   wire si1_delay ;
   wire si2_delay ;
   reg notifier;
   reg notifier0;
   reg notifier1;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
     notifier1 = (notifier1 !== notifier) ? notifier : ~notifier1;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy200ah_func b15fpy200ah1n08x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.d1(d1_delay),.d2(d2_delay),.si1(si1_delay),.si2(si2_delay),.notifier0(notifier0),.notifier1(notifier1),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy200ah_func b15fpy200ah1n08x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.d1(d1_delay),.d2(d2_delay),.si1(si1_delay),.si2(si2_delay),.notifier0(notifier0),.notifier1(notifier1));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d1_delay);
   not MGM_G1(MGM_W1,d2_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,si1_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,si2_delay);
   and MGM_G6(MGM_W6,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W7,ssb_delay);
   and MGM_G8(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W7,MGM_W6);
   not MGM_G9(MGM_W8,d1_delay);
   not MGM_G10(MGM_W9,d2_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   not MGM_G12(MGM_W11,si1_delay);
   and MGM_G13(MGM_W12,MGM_W11,MGM_W10);
   not MGM_G14(MGM_W13,si2_delay);
   and MGM_G15(MGM_W14,MGM_W13,MGM_W12);
   and MGM_G16(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W14);
   not MGM_G17(MGM_W15,d1_delay);
   not MGM_G18(MGM_W16,d2_delay);
   and MGM_G19(MGM_W17,MGM_W16,MGM_W15);
   not MGM_G20(MGM_W18,si1_delay);
   and MGM_G21(MGM_W19,MGM_W18,MGM_W17);
   and MGM_G22(MGM_W20,si2_delay,MGM_W19);
   not MGM_G23(MGM_W21,ssb_delay);
   and MGM_G24(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W21,MGM_W20);
   not MGM_G25(MGM_W22,d1_delay);
   not MGM_G26(MGM_W23,d2_delay);
   and MGM_G27(MGM_W24,MGM_W23,MGM_W22);
   not MGM_G28(MGM_W25,si1_delay);
   and MGM_G29(MGM_W26,MGM_W25,MGM_W24);
   and MGM_G30(MGM_W27,si2_delay,MGM_W26);
   and MGM_G31(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G32(MGM_W28,d1_delay);
   not MGM_G33(MGM_W29,d2_delay);
   and MGM_G34(MGM_W30,MGM_W29,MGM_W28);
   and MGM_G35(MGM_W31,si1_delay,MGM_W30);
   not MGM_G36(MGM_W32,si2_delay);
   and MGM_G37(MGM_W33,MGM_W32,MGM_W31);
   not MGM_G38(MGM_W34,ssb_delay);
   and MGM_G39(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W34,MGM_W33);
   not MGM_G40(MGM_W35,d1_delay);
   not MGM_G41(MGM_W36,d2_delay);
   and MGM_G42(MGM_W37,MGM_W36,MGM_W35);
   and MGM_G43(MGM_W38,si1_delay,MGM_W37);
   not MGM_G44(MGM_W39,si2_delay);
   and MGM_G45(MGM_W40,MGM_W39,MGM_W38);
   and MGM_G46(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G47(MGM_W41,d1_delay);
   not MGM_G48(MGM_W42,d2_delay);
   and MGM_G49(MGM_W43,MGM_W42,MGM_W41);
   and MGM_G50(MGM_W44,si1_delay,MGM_W43);
   and MGM_G51(MGM_W45,si2_delay,MGM_W44);
   not MGM_G52(MGM_W46,ssb_delay);
   and MGM_G53(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W46,MGM_W45);
   not MGM_G54(MGM_W47,d1_delay);
   not MGM_G55(MGM_W48,d2_delay);
   and MGM_G56(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G57(MGM_W50,si1_delay,MGM_W49);
   and MGM_G58(MGM_W51,si2_delay,MGM_W50);
   and MGM_G59(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W51);
   not MGM_G60(MGM_W52,d1_delay);
   and MGM_G61(MGM_W53,d2_delay,MGM_W52);
   not MGM_G62(MGM_W54,si1_delay);
   and MGM_G63(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G64(MGM_W56,si2_delay);
   and MGM_G65(MGM_W57,MGM_W56,MGM_W55);
   not MGM_G66(MGM_W58,ssb_delay);
   and MGM_G67(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W58,MGM_W57);
   not MGM_G68(MGM_W59,d1_delay);
   and MGM_G69(MGM_W60,d2_delay,MGM_W59);
   not MGM_G70(MGM_W61,si1_delay);
   and MGM_G71(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G72(MGM_W63,si2_delay);
   and MGM_G73(MGM_W64,MGM_W63,MGM_W62);
   and MGM_G74(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W64);
   not MGM_G75(MGM_W65,d1_delay);
   and MGM_G76(MGM_W66,d2_delay,MGM_W65);
   not MGM_G77(MGM_W67,si1_delay);
   and MGM_G78(MGM_W68,MGM_W67,MGM_W66);
   and MGM_G79(MGM_W69,si2_delay,MGM_W68);
   not MGM_G80(MGM_W70,ssb_delay);
   and MGM_G81(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W70,MGM_W69);
   not MGM_G82(MGM_W71,d1_delay);
   and MGM_G83(MGM_W72,d2_delay,MGM_W71);
   not MGM_G84(MGM_W73,si1_delay);
   and MGM_G85(MGM_W74,MGM_W73,MGM_W72);
   and MGM_G86(MGM_W75,si2_delay,MGM_W74);
   and MGM_G87(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W75);
   not MGM_G88(MGM_W76,d1_delay);
   and MGM_G89(MGM_W77,d2_delay,MGM_W76);
   and MGM_G90(MGM_W78,si1_delay,MGM_W77);
   not MGM_G91(MGM_W79,si2_delay);
   and MGM_G92(MGM_W80,MGM_W79,MGM_W78);
   not MGM_G93(MGM_W81,ssb_delay);
   and MGM_G94(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W81,MGM_W80);
   not MGM_G95(MGM_W82,d1_delay);
   and MGM_G96(MGM_W83,d2_delay,MGM_W82);
   and MGM_G97(MGM_W84,si1_delay,MGM_W83);
   not MGM_G98(MGM_W85,si2_delay);
   and MGM_G99(MGM_W86,MGM_W85,MGM_W84);
   and MGM_G100(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W86);
   not MGM_G101(MGM_W87,d1_delay);
   and MGM_G102(MGM_W88,d2_delay,MGM_W87);
   and MGM_G103(MGM_W89,si1_delay,MGM_W88);
   and MGM_G104(MGM_W90,si2_delay,MGM_W89);
   not MGM_G105(MGM_W91,ssb_delay);
   and MGM_G106(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W91,MGM_W90);
   not MGM_G107(MGM_W92,d1_delay);
   and MGM_G108(MGM_W93,d2_delay,MGM_W92);
   and MGM_G109(MGM_W94,si1_delay,MGM_W93);
   and MGM_G110(MGM_W95,si2_delay,MGM_W94);
   and MGM_G111(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W95);
   not MGM_G112(MGM_W96,d2_delay);
   and MGM_G113(MGM_W97,MGM_W96,d1_delay);
   not MGM_G114(MGM_W98,si1_delay);
   and MGM_G115(MGM_W99,MGM_W98,MGM_W97);
   not MGM_G116(MGM_W100,si2_delay);
   and MGM_G117(MGM_W101,MGM_W100,MGM_W99);
   not MGM_G118(MGM_W102,ssb_delay);
   and MGM_G119(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W102,MGM_W101);
   not MGM_G120(MGM_W103,d2_delay);
   and MGM_G121(MGM_W104,MGM_W103,d1_delay);
   not MGM_G122(MGM_W105,si1_delay);
   and MGM_G123(MGM_W106,MGM_W105,MGM_W104);
   not MGM_G124(MGM_W107,si2_delay);
   and MGM_G125(MGM_W108,MGM_W107,MGM_W106);
   and MGM_G126(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W108);
   not MGM_G127(MGM_W109,d2_delay);
   and MGM_G128(MGM_W110,MGM_W109,d1_delay);
   not MGM_G129(MGM_W111,si1_delay);
   and MGM_G130(MGM_W112,MGM_W111,MGM_W110);
   and MGM_G131(MGM_W113,si2_delay,MGM_W112);
   not MGM_G132(MGM_W114,ssb_delay);
   and MGM_G133(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W114,MGM_W113);
   not MGM_G134(MGM_W115,d2_delay);
   and MGM_G135(MGM_W116,MGM_W115,d1_delay);
   not MGM_G136(MGM_W117,si1_delay);
   and MGM_G137(MGM_W118,MGM_W117,MGM_W116);
   and MGM_G138(MGM_W119,si2_delay,MGM_W118);
   and MGM_G139(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W119);
   not MGM_G140(MGM_W120,d2_delay);
   and MGM_G141(MGM_W121,MGM_W120,d1_delay);
   and MGM_G142(MGM_W122,si1_delay,MGM_W121);
   not MGM_G143(MGM_W123,si2_delay);
   and MGM_G144(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G145(MGM_W125,ssb_delay);
   and MGM_G146(ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W125,MGM_W124);
   not MGM_G147(MGM_W126,d2_delay);
   and MGM_G148(MGM_W127,MGM_W126,d1_delay);
   and MGM_G149(MGM_W128,si1_delay,MGM_W127);
   not MGM_G150(MGM_W129,si2_delay);
   and MGM_G151(MGM_W130,MGM_W129,MGM_W128);
   and MGM_G152(ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W130);
   not MGM_G153(MGM_W131,d2_delay);
   and MGM_G154(MGM_W132,MGM_W131,d1_delay);
   and MGM_G155(MGM_W133,si1_delay,MGM_W132);
   and MGM_G156(MGM_W134,si2_delay,MGM_W133);
   not MGM_G157(MGM_W135,ssb_delay);
   and MGM_G158(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W135,MGM_W134);
   not MGM_G159(MGM_W136,d2_delay);
   and MGM_G160(MGM_W137,MGM_W136,d1_delay);
   and MGM_G161(MGM_W138,si1_delay,MGM_W137);
   and MGM_G162(MGM_W139,si2_delay,MGM_W138);
   and MGM_G163(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W139);
   and MGM_G164(MGM_W140,d2_delay,d1_delay);
   not MGM_G165(MGM_W141,si1_delay);
   and MGM_G166(MGM_W142,MGM_W141,MGM_W140);
   not MGM_G167(MGM_W143,si2_delay);
   and MGM_G168(MGM_W144,MGM_W143,MGM_W142);
   not MGM_G169(MGM_W145,ssb_delay);
   and MGM_G170(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W145,MGM_W144);
   and MGM_G171(MGM_W146,d2_delay,d1_delay);
   not MGM_G172(MGM_W147,si1_delay);
   and MGM_G173(MGM_W148,MGM_W147,MGM_W146);
   not MGM_G174(MGM_W149,si2_delay);
   and MGM_G175(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G176(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W150);
   and MGM_G177(MGM_W151,d2_delay,d1_delay);
   not MGM_G178(MGM_W152,si1_delay);
   and MGM_G179(MGM_W153,MGM_W152,MGM_W151);
   and MGM_G180(MGM_W154,si2_delay,MGM_W153);
   not MGM_G181(MGM_W155,ssb_delay);
   and MGM_G182(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W155,MGM_W154);
   and MGM_G183(MGM_W156,d2_delay,d1_delay);
   not MGM_G184(MGM_W157,si1_delay);
   and MGM_G185(MGM_W158,MGM_W157,MGM_W156);
   and MGM_G186(MGM_W159,si2_delay,MGM_W158);
   and MGM_G187(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W159);
   and MGM_G188(MGM_W160,d2_delay,d1_delay);
   and MGM_G189(MGM_W161,si1_delay,MGM_W160);
   not MGM_G190(MGM_W162,si2_delay);
   and MGM_G191(MGM_W163,MGM_W162,MGM_W161);
   not MGM_G192(MGM_W164,ssb_delay);
   and MGM_G193(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W164,MGM_W163);
   and MGM_G194(MGM_W165,d2_delay,d1_delay);
   and MGM_G195(MGM_W166,si1_delay,MGM_W165);
   not MGM_G196(MGM_W167,si2_delay);
   and MGM_G197(MGM_W168,MGM_W167,MGM_W166);
   and MGM_G198(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W168);
   and MGM_G199(MGM_W169,d2_delay,d1_delay);
   and MGM_G200(MGM_W170,si1_delay,MGM_W169);
   and MGM_G201(MGM_W171,si2_delay,MGM_W170);
   not MGM_G202(MGM_W172,ssb_delay);
   and MGM_G203(ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W172,MGM_W171);
   and MGM_G204(MGM_W173,d2_delay,d1_delay);
   and MGM_G205(MGM_W174,si1_delay,MGM_W173);
   and MGM_G206(MGM_W175,si2_delay,MGM_W174);
   and MGM_G207(ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W175);
   not MGM_G208(MGM_W176,d1_delay);
   not MGM_G209(MGM_W177,d2_delay);
   and MGM_G210(MGM_W178,MGM_W177,MGM_W176);
   not MGM_G211(MGM_W179,si1_delay);
   and MGM_G212(MGM_W180,MGM_W179,MGM_W178);
   and MGM_G213(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2,si2_delay,MGM_W180);
   not MGM_G214(MGM_W181,d1_delay);
   not MGM_G215(MGM_W182,d2_delay);
   and MGM_G216(MGM_W183,MGM_W182,MGM_W181);
   and MGM_G217(MGM_W184,si1_delay,MGM_W183);
   not MGM_G218(MGM_W185,si2_delay);
   and MGM_G219(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2,MGM_W185,MGM_W184);
   not MGM_G220(MGM_W186,d1_delay);
   not MGM_G221(MGM_W187,d2_delay);
   and MGM_G222(MGM_W188,MGM_W187,MGM_W186);
   and MGM_G223(MGM_W189,si1_delay,MGM_W188);
   and MGM_G224(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2,si2_delay,MGM_W189);
   not MGM_G225(MGM_W190,d1_delay);
   and MGM_G226(MGM_W191,d2_delay,MGM_W190);
   not MGM_G227(MGM_W192,si1_delay);
   and MGM_G228(MGM_W193,MGM_W192,MGM_W191);
   not MGM_G229(MGM_W194,si2_delay);
   and MGM_G230(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2,MGM_W194,MGM_W193);
   not MGM_G231(MGM_W195,d1_delay);
   and MGM_G232(MGM_W196,d2_delay,MGM_W195);
   and MGM_G233(MGM_W197,si1_delay,MGM_W196);
   not MGM_G234(MGM_W198,si2_delay);
   and MGM_G235(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2,MGM_W198,MGM_W197);
   not MGM_G236(MGM_W199,d1_delay);
   and MGM_G237(MGM_W200,d2_delay,MGM_W199);
   and MGM_G238(MGM_W201,si1_delay,MGM_W200);
   and MGM_G239(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2,si2_delay,MGM_W201);
   not MGM_G240(MGM_W202,d2_delay);
   and MGM_G241(MGM_W203,MGM_W202,d1_delay);
   not MGM_G242(MGM_W204,si1_delay);
   and MGM_G243(MGM_W205,MGM_W204,MGM_W203);
   not MGM_G244(MGM_W206,si2_delay);
   and MGM_G245(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2,MGM_W206,MGM_W205);
   not MGM_G246(MGM_W207,d2_delay);
   and MGM_G247(MGM_W208,MGM_W207,d1_delay);
   not MGM_G248(MGM_W209,si1_delay);
   and MGM_G249(MGM_W210,MGM_W209,MGM_W208);
   and MGM_G250(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2,si2_delay,MGM_W210);
   not MGM_G251(MGM_W211,d2_delay);
   and MGM_G252(MGM_W212,MGM_W211,d1_delay);
   and MGM_G253(MGM_W213,si1_delay,MGM_W212);
   and MGM_G254(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2,si2_delay,MGM_W213);
   and MGM_G255(MGM_W214,d2_delay,d1_delay);
   not MGM_G256(MGM_W215,si1_delay);
   and MGM_G257(MGM_W216,MGM_W215,MGM_W214);
   not MGM_G258(MGM_W217,si2_delay);
   and MGM_G259(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2,MGM_W217,MGM_W216);
   and MGM_G260(MGM_W218,d2_delay,d1_delay);
   not MGM_G261(MGM_W219,si1_delay);
   and MGM_G262(MGM_W220,MGM_W219,MGM_W218);
   and MGM_G263(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2,si2_delay,MGM_W220);
   and MGM_G264(MGM_W221,d2_delay,d1_delay);
   and MGM_G265(MGM_W222,si1_delay,MGM_W221);
   not MGM_G266(MGM_W223,si2_delay);
   and MGM_G267(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2,MGM_W223,MGM_W222);
   buf MGM_G268(ENABLE_ssb,ssb_delay);
   not MGM_G269(ENABLE_NOT_ssb,ssb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk,0.0,0,notifier);
      
      $width(posedge clk,0.0,0,notifier);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,negedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,posedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fpy400ah_func( clk, d1, d2, d3, d4, o1, o2, o3, o4, si1, si2, si3, si4, ssb, notifier0, notifier1, notifier2, notifier3 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, d3, d4, si1, si2, si3, si4, ssb, notifier0, notifier1, notifier2, notifier3;
   output o1, o2, o3, o4;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d4, si4, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ4, 1'b0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier3 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D1, d3, si3, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ3, 1'b0, 1'b0, MGM_CLK1, MGM_D1, vcc, vssx, notifier2 );
   INTCseq_cdiar2ah_0( MGM_CLK2, clk, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D2, d2, si2, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, 1'b0, 1'b0, MGM_CLK2, MGM_D2, vcc, vssx, notifier1 );
   INTCseq_cdiar2ah_0( MGM_CLK3, clk, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D3, d1, si1, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, 1'b0, 1'b0, MGM_CLK3, MGM_D3, vcc, vssx, notifier0 );
   INTCseq_cdiar2ah_0( o1, IQ1, vcc, vssx );
   INTCseq_cdiar2ah_0( o2, IQ2, vcc, vssx );
   INTCseq_cdiar2ah_0( o3, IQ3, vcc, vssx );
   INTCseq_cdiar2ah_0( o4, IQ4, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_fdw003ah_5( MGM_D0, d4, si4, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ4, 1'b0, 1'b0, MGM_CLK0, MGM_D0, notifier3 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk );
   INTCseq_fdw003ah_5( MGM_D1, d3, si3, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ3, 1'b0, 1'b0, MGM_CLK1, MGM_D1, notifier2 );
   INTCseq_cdiar2ah_0( MGM_CLK2, clk );
   INTCseq_fdw003ah_5( MGM_D2, d2, si2, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, 1'b0, 1'b0, MGM_CLK2, MGM_D2, notifier1 );
   INTCseq_cdiar2ah_0( MGM_CLK3, clk );
   INTCseq_fdw003ah_5( MGM_D3, d1, si1, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, 1'b0, 1'b0, MGM_CLK3, MGM_D3, notifier0 );
   INTCseq_cdiar2ah_0( o1, IQ1 );
   INTCseq_cdiar2ah_0( o2, IQ2 );
   INTCseq_cdiar2ah_0( o3, IQ3 );
   INTCseq_cdiar2ah_0( o4, IQ4 );
`endif

endmodule
`endcelldefine



`celldefine
module b15fpy400ah1d02x5( clk, d1, d2, d3, d4, o1, o2, o3, o4, si1, si2, si3, si4, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, d3, d4, si1, si2, si3, si4, ssb;
   output o1, o2, o3, o4;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy400ah_func b15fpy400ah1d02x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.si1(si1),.si2(si2),.si3(si3),.si4(si4),.notifier0(1'b0),.notifier1(1'b0),.notifier2(1'b0),.notifier3(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy400ah_func b15fpy400ah1d02x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.si1(si1),.si2(si2),.si3(si3),.si4(si4),.notifier0(1'b0),.notifier1(1'b0),.notifier2(1'b0),.notifier3(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire ssb_delay ;
   wire d1_delay ;
   wire d2_delay ;
   wire d3_delay ;
   wire d4_delay ;
   wire si1_delay ;
   wire si2_delay ;
   wire si3_delay ;
   wire si4_delay ;
   reg notifier;
   reg notifier0;
   reg notifier1;
   reg notifier2;
   reg notifier3;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
     notifier1 = (notifier1 !== notifier) ? notifier : ~notifier1;
     notifier2 = (notifier2 !== notifier) ? notifier : ~notifier2;
     notifier3 = (notifier3 !== notifier) ? notifier : ~notifier3;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy400ah_func b15fpy400ah1d02x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1_delay),.d2(d2_delay),.d3(d3_delay),.d4(d4_delay),.si1(si1_delay),.si2(si2_delay),.si3(si3_delay),.si4(si4_delay),.notifier0(notifier0),.notifier1(notifier1),.notifier2(notifier2),.notifier3(notifier3),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy400ah_func b15fpy400ah1d02x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1_delay),.d2(d2_delay),.d3(d3_delay),.d4(d4_delay),.si1(si1_delay),.si2(si2_delay),.si3(si3_delay),.si4(si4_delay),.notifier0(notifier0),.notifier1(notifier1),.notifier2(notifier2),.notifier3(notifier3));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d1_delay);
   not MGM_G1(MGM_W1,d2_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,d3_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,d4_delay);
   and MGM_G6(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G7(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G8(MGM_W7,si1_delay);
   not MGM_G9(MGM_W8,si2_delay);
   and MGM_G10(MGM_W9,MGM_W8,MGM_W7);
   not MGM_G11(MGM_W10,si3_delay);
   and MGM_G12(MGM_W11,MGM_W10,MGM_W9);
   not MGM_G13(MGM_W12,si4_delay);
   and MGM_G14(MGM_W13,MGM_W12,MGM_W11);
   not MGM_G15(MGM_W14,ssb_delay);
   and MGM_G16(ENABLE_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4_AND_NOT_ssb,MGM_W14,MGM_W13);
   and MGM_G17(MGM_W15,d2_delay,d1_delay);
   and MGM_G18(MGM_W16,d3_delay,MGM_W15);
   and MGM_G19(MGM_W17,d4_delay,MGM_W16);
   and MGM_G20(ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_ssb,ssb_delay,MGM_W17);
   and MGM_G21(MGM_W18,si2_delay,si1_delay);
   and MGM_G22(MGM_W19,si3_delay,MGM_W18);
   and MGM_G23(MGM_W20,si4_delay,MGM_W19);
   not MGM_G24(MGM_W21,ssb_delay);
   and MGM_G25(ENABLE_si1_AND_si2_AND_si3_AND_si4_AND_NOT_ssb,MGM_W21,MGM_W20);
   not MGM_G26(MGM_W22,d1_delay);
   not MGM_G27(MGM_W23,d2_delay);
   and MGM_G28(MGM_W24,MGM_W23,MGM_W22);
   not MGM_G29(MGM_W25,d3_delay);
   and MGM_G30(MGM_W26,MGM_W25,MGM_W24);
   not MGM_G31(MGM_W27,d4_delay);
   and MGM_G32(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G33(MGM_W29,si1_delay,MGM_W28);
   and MGM_G34(MGM_W30,si2_delay,MGM_W29);
   and MGM_G35(MGM_W31,si3_delay,MGM_W30);
   and MGM_G36(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4,si4_delay,MGM_W31);
   and MGM_G37(MGM_W32,d2_delay,d1_delay);
   and MGM_G38(MGM_W33,d3_delay,MGM_W32);
   and MGM_G39(MGM_W34,d4_delay,MGM_W33);
   not MGM_G40(MGM_W35,si1_delay);
   and MGM_G41(MGM_W36,MGM_W35,MGM_W34);
   not MGM_G42(MGM_W37,si2_delay);
   and MGM_G43(MGM_W38,MGM_W37,MGM_W36);
   not MGM_G44(MGM_W39,si3_delay);
   and MGM_G45(MGM_W40,MGM_W39,MGM_W38);
   not MGM_G46(MGM_W41,si4_delay);
   and MGM_G47(ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4,MGM_W41,MGM_W40);
   buf MGM_G48(ENABLE_ssb,ssb_delay);
   not MGM_G49(ENABLE_NOT_ssb,ssb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b0 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b0 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b1 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b1 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b0 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b0 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b1 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b1 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_si1_AND_si2_AND_si3_AND_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_si1_AND_si2_AND_si3_AND_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk,0.0,0,notifier);
      
      $width(posedge clk,0.0,0,notifier);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,negedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,posedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d3 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,d3_delay);
      
      // setuphold d3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d3 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,d3_delay);
      
      // setuphold d4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d4 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,d4_delay);
      
      // setuphold d4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d4 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,d4_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si3 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,si3_delay);
      
      // setuphold si3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si3 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,si3_delay);
      
      // setuphold si4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si4 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,si4_delay);
      
      // setuphold si4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si4 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,si4_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy400ah1d03x5( clk, d1, d2, d3, d4, o1, o2, o3, o4, si1, si2, si3, si4, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, d3, d4, si1, si2, si3, si4, ssb;
   output o1, o2, o3, o4;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy400ah_func b15fpy400ah1d03x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.si1(si1),.si2(si2),.si3(si3),.si4(si4),.notifier0(1'b0),.notifier1(1'b0),.notifier2(1'b0),.notifier3(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy400ah_func b15fpy400ah1d03x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.si1(si1),.si2(si2),.si3(si3),.si4(si4),.notifier0(1'b0),.notifier1(1'b0),.notifier2(1'b0),.notifier3(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire ssb_delay ;
   wire d1_delay ;
   wire d2_delay ;
   wire d3_delay ;
   wire d4_delay ;
   wire si1_delay ;
   wire si2_delay ;
   wire si3_delay ;
   wire si4_delay ;
   reg notifier;
   reg notifier0;
   reg notifier1;
   reg notifier2;
   reg notifier3;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
     notifier1 = (notifier1 !== notifier) ? notifier : ~notifier1;
     notifier2 = (notifier2 !== notifier) ? notifier : ~notifier2;
     notifier3 = (notifier3 !== notifier) ? notifier : ~notifier3;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy400ah_func b15fpy400ah1d03x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1_delay),.d2(d2_delay),.d3(d3_delay),.d4(d4_delay),.si1(si1_delay),.si2(si2_delay),.si3(si3_delay),.si4(si4_delay),.notifier0(notifier0),.notifier1(notifier1),.notifier2(notifier2),.notifier3(notifier3),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy400ah_func b15fpy400ah1d03x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1_delay),.d2(d2_delay),.d3(d3_delay),.d4(d4_delay),.si1(si1_delay),.si2(si2_delay),.si3(si3_delay),.si4(si4_delay),.notifier0(notifier0),.notifier1(notifier1),.notifier2(notifier2),.notifier3(notifier3));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d1_delay);
   not MGM_G1(MGM_W1,d2_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,d3_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,d4_delay);
   and MGM_G6(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G7(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G8(MGM_W7,si1_delay);
   not MGM_G9(MGM_W8,si2_delay);
   and MGM_G10(MGM_W9,MGM_W8,MGM_W7);
   not MGM_G11(MGM_W10,si3_delay);
   and MGM_G12(MGM_W11,MGM_W10,MGM_W9);
   not MGM_G13(MGM_W12,si4_delay);
   and MGM_G14(MGM_W13,MGM_W12,MGM_W11);
   not MGM_G15(MGM_W14,ssb_delay);
   and MGM_G16(ENABLE_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4_AND_NOT_ssb,MGM_W14,MGM_W13);
   and MGM_G17(MGM_W15,d2_delay,d1_delay);
   and MGM_G18(MGM_W16,d3_delay,MGM_W15);
   and MGM_G19(MGM_W17,d4_delay,MGM_W16);
   and MGM_G20(ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_ssb,ssb_delay,MGM_W17);
   and MGM_G21(MGM_W18,si2_delay,si1_delay);
   and MGM_G22(MGM_W19,si3_delay,MGM_W18);
   and MGM_G23(MGM_W20,si4_delay,MGM_W19);
   not MGM_G24(MGM_W21,ssb_delay);
   and MGM_G25(ENABLE_si1_AND_si2_AND_si3_AND_si4_AND_NOT_ssb,MGM_W21,MGM_W20);
   not MGM_G26(MGM_W22,d1_delay);
   not MGM_G27(MGM_W23,d2_delay);
   and MGM_G28(MGM_W24,MGM_W23,MGM_W22);
   not MGM_G29(MGM_W25,d3_delay);
   and MGM_G30(MGM_W26,MGM_W25,MGM_W24);
   not MGM_G31(MGM_W27,d4_delay);
   and MGM_G32(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G33(MGM_W29,si1_delay,MGM_W28);
   and MGM_G34(MGM_W30,si2_delay,MGM_W29);
   and MGM_G35(MGM_W31,si3_delay,MGM_W30);
   and MGM_G36(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4,si4_delay,MGM_W31);
   and MGM_G37(MGM_W32,d2_delay,d1_delay);
   and MGM_G38(MGM_W33,d3_delay,MGM_W32);
   and MGM_G39(MGM_W34,d4_delay,MGM_W33);
   not MGM_G40(MGM_W35,si1_delay);
   and MGM_G41(MGM_W36,MGM_W35,MGM_W34);
   not MGM_G42(MGM_W37,si2_delay);
   and MGM_G43(MGM_W38,MGM_W37,MGM_W36);
   not MGM_G44(MGM_W39,si3_delay);
   and MGM_G45(MGM_W40,MGM_W39,MGM_W38);
   not MGM_G46(MGM_W41,si4_delay);
   and MGM_G47(ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4,MGM_W41,MGM_W40);
   buf MGM_G48(ENABLE_ssb,ssb_delay);
   not MGM_G49(ENABLE_NOT_ssb,ssb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b0 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b0 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b1 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b1 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b0 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b0 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b1 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b1 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_si1_AND_si2_AND_si3_AND_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_si1_AND_si2_AND_si3_AND_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk,0.0,0,notifier);
      
      $width(posedge clk,0.0,0,notifier);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,negedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,posedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d3 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,d3_delay);
      
      // setuphold d3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d3 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,d3_delay);
      
      // setuphold d4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d4 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,d4_delay);
      
      // setuphold d4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d4 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,d4_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si3 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,si3_delay);
      
      // setuphold si3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si3 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,si3_delay);
      
      // setuphold si4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si4 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,si4_delay);
      
      // setuphold si4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si4 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,si4_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy400ah1d04x5( clk, d1, d2, d3, d4, o1, o2, o3, o4, si1, si2, si3, si4, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, d3, d4, si1, si2, si3, si4, ssb;
   output o1, o2, o3, o4;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy400ah_func b15fpy400ah1d04x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.si1(si1),.si2(si2),.si3(si3),.si4(si4),.notifier0(1'b0),.notifier1(1'b0),.notifier2(1'b0),.notifier3(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy400ah_func b15fpy400ah1d04x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.si1(si1),.si2(si2),.si3(si3),.si4(si4),.notifier0(1'b0),.notifier1(1'b0),.notifier2(1'b0),.notifier3(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire ssb_delay ;
   wire d1_delay ;
   wire d2_delay ;
   wire d3_delay ;
   wire d4_delay ;
   wire si1_delay ;
   wire si2_delay ;
   wire si3_delay ;
   wire si4_delay ;
   reg notifier;
   reg notifier0;
   reg notifier1;
   reg notifier2;
   reg notifier3;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
     notifier1 = (notifier1 !== notifier) ? notifier : ~notifier1;
     notifier2 = (notifier2 !== notifier) ? notifier : ~notifier2;
     notifier3 = (notifier3 !== notifier) ? notifier : ~notifier3;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy400ah_func b15fpy400ah1d04x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1_delay),.d2(d2_delay),.d3(d3_delay),.d4(d4_delay),.si1(si1_delay),.si2(si2_delay),.si3(si3_delay),.si4(si4_delay),.notifier0(notifier0),.notifier1(notifier1),.notifier2(notifier2),.notifier3(notifier3),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy400ah_func b15fpy400ah1d04x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1_delay),.d2(d2_delay),.d3(d3_delay),.d4(d4_delay),.si1(si1_delay),.si2(si2_delay),.si3(si3_delay),.si4(si4_delay),.notifier0(notifier0),.notifier1(notifier1),.notifier2(notifier2),.notifier3(notifier3));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d1_delay);
   not MGM_G1(MGM_W1,d2_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,d3_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,d4_delay);
   and MGM_G6(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G7(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G8(MGM_W7,si1_delay);
   not MGM_G9(MGM_W8,si2_delay);
   and MGM_G10(MGM_W9,MGM_W8,MGM_W7);
   not MGM_G11(MGM_W10,si3_delay);
   and MGM_G12(MGM_W11,MGM_W10,MGM_W9);
   not MGM_G13(MGM_W12,si4_delay);
   and MGM_G14(MGM_W13,MGM_W12,MGM_W11);
   not MGM_G15(MGM_W14,ssb_delay);
   and MGM_G16(ENABLE_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4_AND_NOT_ssb,MGM_W14,MGM_W13);
   and MGM_G17(MGM_W15,d2_delay,d1_delay);
   and MGM_G18(MGM_W16,d3_delay,MGM_W15);
   and MGM_G19(MGM_W17,d4_delay,MGM_W16);
   and MGM_G20(ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_ssb,ssb_delay,MGM_W17);
   and MGM_G21(MGM_W18,si2_delay,si1_delay);
   and MGM_G22(MGM_W19,si3_delay,MGM_W18);
   and MGM_G23(MGM_W20,si4_delay,MGM_W19);
   not MGM_G24(MGM_W21,ssb_delay);
   and MGM_G25(ENABLE_si1_AND_si2_AND_si3_AND_si4_AND_NOT_ssb,MGM_W21,MGM_W20);
   not MGM_G26(MGM_W22,d1_delay);
   not MGM_G27(MGM_W23,d2_delay);
   and MGM_G28(MGM_W24,MGM_W23,MGM_W22);
   not MGM_G29(MGM_W25,d3_delay);
   and MGM_G30(MGM_W26,MGM_W25,MGM_W24);
   not MGM_G31(MGM_W27,d4_delay);
   and MGM_G32(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G33(MGM_W29,si1_delay,MGM_W28);
   and MGM_G34(MGM_W30,si2_delay,MGM_W29);
   and MGM_G35(MGM_W31,si3_delay,MGM_W30);
   and MGM_G36(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4,si4_delay,MGM_W31);
   and MGM_G37(MGM_W32,d2_delay,d1_delay);
   and MGM_G38(MGM_W33,d3_delay,MGM_W32);
   and MGM_G39(MGM_W34,d4_delay,MGM_W33);
   not MGM_G40(MGM_W35,si1_delay);
   and MGM_G41(MGM_W36,MGM_W35,MGM_W34);
   not MGM_G42(MGM_W37,si2_delay);
   and MGM_G43(MGM_W38,MGM_W37,MGM_W36);
   not MGM_G44(MGM_W39,si3_delay);
   and MGM_G45(MGM_W40,MGM_W39,MGM_W38);
   not MGM_G46(MGM_W41,si4_delay);
   and MGM_G47(ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4,MGM_W41,MGM_W40);
   buf MGM_G48(ENABLE_ssb,ssb_delay);
   not MGM_G49(ENABLE_NOT_ssb,ssb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b0 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b0 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b1 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b1 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b0 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b0 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b1 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b1 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_si1_AND_si2_AND_si3_AND_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_si1_AND_si2_AND_si3_AND_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk,0.0,0,notifier);
      
      $width(posedge clk,0.0,0,notifier);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,negedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,posedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d3 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,d3_delay);
      
      // setuphold d3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d3 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,d3_delay);
      
      // setuphold d4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d4 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,d4_delay);
      
      // setuphold d4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d4 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,d4_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si3 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,si3_delay);
      
      // setuphold si3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si3 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,si3_delay);
      
      // setuphold si4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si4 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,si4_delay);
      
      // setuphold si4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si4 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,si4_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fpy400ah1d08x5( clk, d1, d2, d3, d4, o1, o2, o3, o4, si1, si2, si3, si4, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, d3, d4, si1, si2, si3, si4, ssb;
   output o1, o2, o3, o4;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy400ah_func b15fpy400ah1d08x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.si1(si1),.si2(si2),.si3(si3),.si4(si4),.notifier0(1'b0),.notifier1(1'b0),.notifier2(1'b0),.notifier3(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy400ah_func b15fpy400ah1d08x5_behav_inst(.clk(clk),.ssb(ssb),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.si1(si1),.si2(si2),.si3(si3),.si4(si4),.notifier0(1'b0),.notifier1(1'b0),.notifier2(1'b0),.notifier3(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire ssb_delay ;
   wire d1_delay ;
   wire d2_delay ;
   wire d3_delay ;
   wire d4_delay ;
   wire si1_delay ;
   wire si2_delay ;
   wire si3_delay ;
   wire si4_delay ;
   reg notifier;
   reg notifier0;
   reg notifier1;
   reg notifier2;
   reg notifier3;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
     notifier1 = (notifier1 !== notifier) ? notifier : ~notifier1;
     notifier2 = (notifier2 !== notifier) ? notifier : ~notifier2;
     notifier3 = (notifier3 !== notifier) ? notifier : ~notifier3;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fpy400ah_func b15fpy400ah1d08x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1_delay),.d2(d2_delay),.d3(d3_delay),.d4(d4_delay),.si1(si1_delay),.si2(si2_delay),.si3(si3_delay),.si4(si4_delay),.notifier0(notifier0),.notifier1(notifier1),.notifier2(notifier2),.notifier3(notifier3),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fpy400ah_func b15fpy400ah1d08x5_inst(.clk(clk_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1_delay),.d2(d2_delay),.d3(d3_delay),.d4(d4_delay),.si1(si1_delay),.si2(si2_delay),.si3(si3_delay),.si4(si4_delay),.notifier0(notifier0),.notifier1(notifier1),.notifier2(notifier2),.notifier3(notifier3));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d1_delay);
   not MGM_G1(MGM_W1,d2_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G3(MGM_W3,d3_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,d4_delay);
   and MGM_G6(MGM_W6,MGM_W5,MGM_W4);
   and MGM_G7(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G8(MGM_W7,si1_delay);
   not MGM_G9(MGM_W8,si2_delay);
   and MGM_G10(MGM_W9,MGM_W8,MGM_W7);
   not MGM_G11(MGM_W10,si3_delay);
   and MGM_G12(MGM_W11,MGM_W10,MGM_W9);
   not MGM_G13(MGM_W12,si4_delay);
   and MGM_G14(MGM_W13,MGM_W12,MGM_W11);
   not MGM_G15(MGM_W14,ssb_delay);
   and MGM_G16(ENABLE_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4_AND_NOT_ssb,MGM_W14,MGM_W13);
   and MGM_G17(MGM_W15,d2_delay,d1_delay);
   and MGM_G18(MGM_W16,d3_delay,MGM_W15);
   and MGM_G19(MGM_W17,d4_delay,MGM_W16);
   and MGM_G20(ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_ssb,ssb_delay,MGM_W17);
   and MGM_G21(MGM_W18,si2_delay,si1_delay);
   and MGM_G22(MGM_W19,si3_delay,MGM_W18);
   and MGM_G23(MGM_W20,si4_delay,MGM_W19);
   not MGM_G24(MGM_W21,ssb_delay);
   and MGM_G25(ENABLE_si1_AND_si2_AND_si3_AND_si4_AND_NOT_ssb,MGM_W21,MGM_W20);
   not MGM_G26(MGM_W22,d1_delay);
   not MGM_G27(MGM_W23,d2_delay);
   and MGM_G28(MGM_W24,MGM_W23,MGM_W22);
   not MGM_G29(MGM_W25,d3_delay);
   and MGM_G30(MGM_W26,MGM_W25,MGM_W24);
   not MGM_G31(MGM_W27,d4_delay);
   and MGM_G32(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G33(MGM_W29,si1_delay,MGM_W28);
   and MGM_G34(MGM_W30,si2_delay,MGM_W29);
   and MGM_G35(MGM_W31,si3_delay,MGM_W30);
   and MGM_G36(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4,si4_delay,MGM_W31);
   and MGM_G37(MGM_W32,d2_delay,d1_delay);
   and MGM_G38(MGM_W33,d3_delay,MGM_W32);
   and MGM_G39(MGM_W34,d4_delay,MGM_W33);
   not MGM_G40(MGM_W35,si1_delay);
   and MGM_G41(MGM_W36,MGM_W35,MGM_W34);
   not MGM_G42(MGM_W37,si2_delay);
   and MGM_G43(MGM_W38,MGM_W37,MGM_W36);
   not MGM_G44(MGM_W39,si3_delay);
   and MGM_G45(MGM_W40,MGM_W39,MGM_W38);
   not MGM_G46(MGM_W41,si4_delay);
   and MGM_G47(ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4,MGM_W41,MGM_W40);
   buf MGM_G48(ENABLE_ssb,ssb_delay);
   not MGM_G49(ENABLE_NOT_ssb,ssb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b0 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b0 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b1 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && si3==1'b1 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b0 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b0 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b1 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && si4==1'b1 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_si1_AND_si2_AND_si3_AND_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_si1_AND_si2_AND_si3_AND_si4_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk,0.0,0,notifier);
      
      $width(posedge clk,0.0,0,notifier);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,negedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,posedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d1 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d2 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d3 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,d3_delay);
      
      // setuphold d3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d3 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,d3_delay);
      
      // setuphold d4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      negedge d4 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,d4_delay);
      
      // setuphold d4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb == 1'b1),
      posedge d4 &&& (ENABLE_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,d4_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si1 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si2 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si3 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,si3_delay);
      
      // setuphold si3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si3 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,si3_delay);
      
      // setuphold si4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      negedge si4 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,si4_delay);
      
      // setuphold si4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb == 1'b1),
      posedge si4 &&& (ENABLE_NOT_ssb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,si4_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fqn003ah_func( clk, d, o, rb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, d, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_cdiar2ah_0( MGM_D0, d );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fqn003ah1n02x5( clk, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn003ah_func b15fqn003ah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn003ah_func b15fqn003ah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn003ah_func b15fqn003ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn003ah_func b15fqn003ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn003ah1n03x5( clk, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn003ah_func b15fqn003ah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn003ah_func b15fqn003ah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn003ah_func b15fqn003ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn003ah_func b15fqn003ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn003ah1n04x5( clk, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn003ah_func b15fqn003ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn003ah_func b15fqn003ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn003ah_func b15fqn003ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn003ah_func b15fqn003ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn003ah1n06x5( clk, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn003ah_func b15fqn003ah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn003ah_func b15fqn003ah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn003ah_func b15fqn003ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn003ah_func b15fqn003ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn003ah1n08x5( clk, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn003ah_func b15fqn003ah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn003ah_func b15fqn003ah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn003ah_func b15fqn003ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn003ah_func b15fqn003ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn003ah1n12x5( clk, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn003ah_func b15fqn003ah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn003ah_func b15fqn003ah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn003ah_func b15fqn003ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn003ah_func b15fqn003ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn003ah1n16x5( clk, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn003ah_func b15fqn003ah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn003ah_func b15fqn003ah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn003ah_func b15fqn003ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn003ah_func b15fqn003ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fqn00cah_func( clk, d, o, psb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_P0, psb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, d, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, MGM_P0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_P0, psb );
   INTCseq_cdiar2ah_0( MGM_D0, d );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, MGM_P0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fqn00cah1n02x5( clk, d, o, psb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00cah_func b15fqn00cah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00cah_func b15fqn00cah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00cah_func b15fqn00cah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00cah_func b15fqn00cah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_psb,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_psb,psb_delay,d_delay);
   buf MGM_G3(ENABLE_psb,psb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb == 1'b1),
      negedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb == 1'b1),
      posedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb,posedge clk,0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn00cah1n03x5( clk, d, o, psb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00cah_func b15fqn00cah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00cah_func b15fqn00cah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00cah_func b15fqn00cah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00cah_func b15fqn00cah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_psb,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_psb,psb_delay,d_delay);
   buf MGM_G3(ENABLE_psb,psb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb == 1'b1),
      negedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb == 1'b1),
      posedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb,posedge clk,0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn00cah1n04x5( clk, d, o, psb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00cah_func b15fqn00cah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00cah_func b15fqn00cah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00cah_func b15fqn00cah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00cah_func b15fqn00cah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_psb,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_psb,psb_delay,d_delay);
   buf MGM_G3(ENABLE_psb,psb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb == 1'b1),
      negedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb == 1'b1),
      posedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb,posedge clk,0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn00cah1n06x5( clk, d, o, psb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00cah_func b15fqn00cah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00cah_func b15fqn00cah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00cah_func b15fqn00cah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00cah_func b15fqn00cah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_psb,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_psb,psb_delay,d_delay);
   buf MGM_G3(ENABLE_psb,psb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb == 1'b1),
      negedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb == 1'b1),
      posedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb,posedge clk,0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn00cah1n08x5( clk, d, o, psb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00cah_func b15fqn00cah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00cah_func b15fqn00cah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00cah_func b15fqn00cah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00cah_func b15fqn00cah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_psb,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_psb,psb_delay,d_delay);
   buf MGM_G3(ENABLE_psb,psb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb == 1'b1),
      negedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb == 1'b1),
      posedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb,posedge clk,0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn00cah1n12x5( clk, d, o, psb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00cah_func b15fqn00cah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00cah_func b15fqn00cah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00cah_func b15fqn00cah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00cah_func b15fqn00cah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_psb,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_psb,psb_delay,d_delay);
   buf MGM_G3(ENABLE_psb,psb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb == 1'b1),
      negedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb == 1'b1),
      posedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb,posedge clk,0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn00cah1n16x5( clk, d, o, psb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00cah_func b15fqn00cah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00cah_func b15fqn00cah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00cah_func b15fqn00cah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00cah_func b15fqn00cah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_psb,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_psb,psb_delay,d_delay);
   buf MGM_G3(ENABLE_psb,psb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   not MGM_G9(MGM_W4,d_delay);
   and MGM_G10(ENABLE_clk_AND_NOT_d,MGM_W4,clk_delay);
   and MGM_G11(ENABLE_clk_AND_d,d_delay,clk_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb == 1'b1),
      negedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb == 1'b1),
      posedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb,posedge clk,0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine


primitive INTCseq_fqn00fah_LN_IQ_FF_UDP( Q, C, P, CK, D `ifdef POWER_AWARE_MODE , vcc, vssx `endif , N );
   output Q;
   reg Q;
   input C, P, CK, D, N; 
   `ifdef POWER_AWARE_MODE
   input vcc, vssx;
   `endif
   table 
  `ifdef POWER_AWARE_MODE
   //C  P  CK D  PW GN N  :  Q  :  Q 
     0  0  n  ?  1  0  ?  :  ?  :  -;
     ?  0  n  ?  1  0  ?  :  0  :  0;
     0  ?  n  ?  1  0  ?  :  1  :  1;
     ?  0  r  0  1  0  ?  :  ?  :  0;
     1  ?  ?  ?  1  0  ?  :  ?  :  0;
     0  ?  r  1  1  0  ?  :  ?  :  1;
     0  1  ?  ?  1  0  ?  :  ?  :  1;
     0  0  ?  *  1  0  ?  :  ?  :  -;
     0  ?  ?  *  1  0  ?  :  1  :  1;
     ?  0  ?  *  1  0  ?  :  0  :  0;
     0  *  ?  ?  1  0  ?  :  1  :  1;
     *  0  ?  ?  1  0  ?  :  0  :  0;
     ?  0  *  0  1  0  ?  :  0  :  0;
     0  ?  *  1  1  0  ?  :  1  :  1;
     ?  ?  ?  ?  1  0  *  :  ?  :  x;
  `else
   //C  P  CK D  N  :  Q  :  Q 
     0  0  n  ?  ?  :  ?  :  -;
     ?  0  n  ?  ?  :  0  :  0;
     0  ?  n  ?  ?  :  1  :  1;
     ?  0  r  0  ?  :  ?  :  0;
     1  ?  ?  ?  ?  :  ?  :  0;
     0  ?  r  1  ?  :  ?  :  1;
     0  1  ?  ?  ?  :  ?  :  1;
     0  0  ?  *  ?  :  ?  :  -;
     0  ?  ?  *  ?  :  1  :  1;
     ?  0  ?  *  ?  :  0  :  0;
     0  *  ?  ?  ?  :  1  :  1;
     *  0  ?  ?  ?  :  0  :  0;
     ?  0  *  0  ?  :  0  :  0;
     0  ?  *  1  ?  :  1  :  1;
     ?  ?  ?  ?  *  :  ?  :  x;
  `endif

endtable
endprimitive



`celldefine
module INTCseq_fqn00fah_func( clk, d, o, psb, rb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_P0, psb, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, d, vcc, vssx );
   INTCseq_fqn00fah_LN_IQ_FF_UDP( IQ, MGM_C0, MGM_P0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_P0, psb );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_cdiar2ah_0( MGM_D0, d );
   INTCseq_fqn00fah_LN_IQ_FF_UDP( IQ, MGM_C0, MGM_P0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fqn00fah1n02x5( clk, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00fah_func b15fqn00fah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00fah_func b15fqn00fah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00fah_func b15fqn00fah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00fah_func b15fqn00fah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clk_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clk_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clk_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,d_delay);
   and MGM_G15(MGM_W9,MGM_W8,clk_delay);
   and MGM_G16(ENABLE_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W9);
   and MGM_G17(MGM_W10,d_delay,clk_delay);
   and MGM_G18(ENABLE_clk_AND_d_AND_rb,rb_delay,MGM_W10);
   not MGM_G19(MGM_W11,clk_delay);
   not MGM_G20(MGM_W12,d_delay);
   and MGM_G21(ENABLE_NOT_clk_AND_NOT_d,MGM_W12,MGM_W11);
   not MGM_G22(MGM_W13,clk_delay);
   and MGM_G23(ENABLE_NOT_clk_AND_d,d_delay,MGM_W13);
   not MGM_G24(MGM_W14,d_delay);
   and MGM_G25(ENABLE_clk_AND_NOT_d,MGM_W14,clk_delay);
   and MGM_G26(ENABLE_clk_AND_d,d_delay,clk_delay);
   buf MGM_G27(ENABLE_psb,psb_delay);
   not MGM_G28(MGM_W15,clk_delay);
   not MGM_G29(MGM_W16,d_delay);
   and MGM_G30(MGM_W17,MGM_W16,MGM_W15);
   and MGM_G31(ENABLE_NOT_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W17);
   not MGM_G32(MGM_W18,clk_delay);
   and MGM_G33(MGM_W19,d_delay,MGM_W18);
   and MGM_G34(ENABLE_NOT_clk_AND_d_AND_psb,psb_delay,MGM_W19);
   not MGM_G35(MGM_W20,d_delay);
   and MGM_G36(MGM_W21,MGM_W20,clk_delay);
   and MGM_G37(ENABLE_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W21);
   and MGM_G38(MGM_W22,d_delay,clk_delay);
   and MGM_G39(ENABLE_clk_AND_d_AND_psb,psb_delay,MGM_W22);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      posedge clk &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      posedge clk &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn00fah1n03x5( clk, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00fah_func b15fqn00fah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00fah_func b15fqn00fah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00fah_func b15fqn00fah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00fah_func b15fqn00fah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clk_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clk_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clk_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,d_delay);
   and MGM_G15(MGM_W9,MGM_W8,clk_delay);
   and MGM_G16(ENABLE_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W9);
   and MGM_G17(MGM_W10,d_delay,clk_delay);
   and MGM_G18(ENABLE_clk_AND_d_AND_rb,rb_delay,MGM_W10);
   not MGM_G19(MGM_W11,clk_delay);
   not MGM_G20(MGM_W12,d_delay);
   and MGM_G21(ENABLE_NOT_clk_AND_NOT_d,MGM_W12,MGM_W11);
   not MGM_G22(MGM_W13,clk_delay);
   and MGM_G23(ENABLE_NOT_clk_AND_d,d_delay,MGM_W13);
   not MGM_G24(MGM_W14,d_delay);
   and MGM_G25(ENABLE_clk_AND_NOT_d,MGM_W14,clk_delay);
   and MGM_G26(ENABLE_clk_AND_d,d_delay,clk_delay);
   buf MGM_G27(ENABLE_psb,psb_delay);
   not MGM_G28(MGM_W15,clk_delay);
   not MGM_G29(MGM_W16,d_delay);
   and MGM_G30(MGM_W17,MGM_W16,MGM_W15);
   and MGM_G31(ENABLE_NOT_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W17);
   not MGM_G32(MGM_W18,clk_delay);
   and MGM_G33(MGM_W19,d_delay,MGM_W18);
   and MGM_G34(ENABLE_NOT_clk_AND_d_AND_psb,psb_delay,MGM_W19);
   not MGM_G35(MGM_W20,d_delay);
   and MGM_G36(MGM_W21,MGM_W20,clk_delay);
   and MGM_G37(ENABLE_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W21);
   and MGM_G38(MGM_W22,d_delay,clk_delay);
   and MGM_G39(ENABLE_clk_AND_d_AND_psb,psb_delay,MGM_W22);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      posedge clk &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      posedge clk &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn00fah1n04x5( clk, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00fah_func b15fqn00fah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00fah_func b15fqn00fah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00fah_func b15fqn00fah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00fah_func b15fqn00fah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clk_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clk_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clk_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,d_delay);
   and MGM_G15(MGM_W9,MGM_W8,clk_delay);
   and MGM_G16(ENABLE_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W9);
   and MGM_G17(MGM_W10,d_delay,clk_delay);
   and MGM_G18(ENABLE_clk_AND_d_AND_rb,rb_delay,MGM_W10);
   not MGM_G19(MGM_W11,clk_delay);
   not MGM_G20(MGM_W12,d_delay);
   and MGM_G21(ENABLE_NOT_clk_AND_NOT_d,MGM_W12,MGM_W11);
   not MGM_G22(MGM_W13,clk_delay);
   and MGM_G23(ENABLE_NOT_clk_AND_d,d_delay,MGM_W13);
   not MGM_G24(MGM_W14,d_delay);
   and MGM_G25(ENABLE_clk_AND_NOT_d,MGM_W14,clk_delay);
   and MGM_G26(ENABLE_clk_AND_d,d_delay,clk_delay);
   buf MGM_G27(ENABLE_psb,psb_delay);
   not MGM_G28(MGM_W15,clk_delay);
   not MGM_G29(MGM_W16,d_delay);
   and MGM_G30(MGM_W17,MGM_W16,MGM_W15);
   and MGM_G31(ENABLE_NOT_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W17);
   not MGM_G32(MGM_W18,clk_delay);
   and MGM_G33(MGM_W19,d_delay,MGM_W18);
   and MGM_G34(ENABLE_NOT_clk_AND_d_AND_psb,psb_delay,MGM_W19);
   not MGM_G35(MGM_W20,d_delay);
   and MGM_G36(MGM_W21,MGM_W20,clk_delay);
   and MGM_G37(ENABLE_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W21);
   and MGM_G38(MGM_W22,d_delay,clk_delay);
   and MGM_G39(ENABLE_clk_AND_d_AND_psb,psb_delay,MGM_W22);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      posedge clk &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      posedge clk &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn00fah1n06x5( clk, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00fah_func b15fqn00fah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00fah_func b15fqn00fah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00fah_func b15fqn00fah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00fah_func b15fqn00fah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clk_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clk_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clk_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,d_delay);
   and MGM_G15(MGM_W9,MGM_W8,clk_delay);
   and MGM_G16(ENABLE_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W9);
   and MGM_G17(MGM_W10,d_delay,clk_delay);
   and MGM_G18(ENABLE_clk_AND_d_AND_rb,rb_delay,MGM_W10);
   not MGM_G19(MGM_W11,clk_delay);
   not MGM_G20(MGM_W12,d_delay);
   and MGM_G21(ENABLE_NOT_clk_AND_NOT_d,MGM_W12,MGM_W11);
   not MGM_G22(MGM_W13,clk_delay);
   and MGM_G23(ENABLE_NOT_clk_AND_d,d_delay,MGM_W13);
   not MGM_G24(MGM_W14,d_delay);
   and MGM_G25(ENABLE_clk_AND_NOT_d,MGM_W14,clk_delay);
   and MGM_G26(ENABLE_clk_AND_d,d_delay,clk_delay);
   buf MGM_G27(ENABLE_psb,psb_delay);
   not MGM_G28(MGM_W15,clk_delay);
   not MGM_G29(MGM_W16,d_delay);
   and MGM_G30(MGM_W17,MGM_W16,MGM_W15);
   and MGM_G31(ENABLE_NOT_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W17);
   not MGM_G32(MGM_W18,clk_delay);
   and MGM_G33(MGM_W19,d_delay,MGM_W18);
   and MGM_G34(ENABLE_NOT_clk_AND_d_AND_psb,psb_delay,MGM_W19);
   not MGM_G35(MGM_W20,d_delay);
   and MGM_G36(MGM_W21,MGM_W20,clk_delay);
   and MGM_G37(ENABLE_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W21);
   and MGM_G38(MGM_W22,d_delay,clk_delay);
   and MGM_G39(ENABLE_clk_AND_d_AND_psb,psb_delay,MGM_W22);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      posedge clk &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      posedge clk &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn00fah1n08x5( clk, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00fah_func b15fqn00fah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00fah_func b15fqn00fah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00fah_func b15fqn00fah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00fah_func b15fqn00fah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clk_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clk_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clk_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,d_delay);
   and MGM_G15(MGM_W9,MGM_W8,clk_delay);
   and MGM_G16(ENABLE_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W9);
   and MGM_G17(MGM_W10,d_delay,clk_delay);
   and MGM_G18(ENABLE_clk_AND_d_AND_rb,rb_delay,MGM_W10);
   not MGM_G19(MGM_W11,clk_delay);
   not MGM_G20(MGM_W12,d_delay);
   and MGM_G21(ENABLE_NOT_clk_AND_NOT_d,MGM_W12,MGM_W11);
   not MGM_G22(MGM_W13,clk_delay);
   and MGM_G23(ENABLE_NOT_clk_AND_d,d_delay,MGM_W13);
   not MGM_G24(MGM_W14,d_delay);
   and MGM_G25(ENABLE_clk_AND_NOT_d,MGM_W14,clk_delay);
   and MGM_G26(ENABLE_clk_AND_d,d_delay,clk_delay);
   buf MGM_G27(ENABLE_psb,psb_delay);
   not MGM_G28(MGM_W15,clk_delay);
   not MGM_G29(MGM_W16,d_delay);
   and MGM_G30(MGM_W17,MGM_W16,MGM_W15);
   and MGM_G31(ENABLE_NOT_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W17);
   not MGM_G32(MGM_W18,clk_delay);
   and MGM_G33(MGM_W19,d_delay,MGM_W18);
   and MGM_G34(ENABLE_NOT_clk_AND_d_AND_psb,psb_delay,MGM_W19);
   not MGM_G35(MGM_W20,d_delay);
   and MGM_G36(MGM_W21,MGM_W20,clk_delay);
   and MGM_G37(ENABLE_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W21);
   and MGM_G38(MGM_W22,d_delay,clk_delay);
   and MGM_G39(ENABLE_clk_AND_d_AND_psb,psb_delay,MGM_W22);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      posedge clk &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      posedge clk &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn00fah1n12x5( clk, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00fah_func b15fqn00fah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00fah_func b15fqn00fah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00fah_func b15fqn00fah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00fah_func b15fqn00fah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clk_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clk_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clk_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,d_delay);
   and MGM_G15(MGM_W9,MGM_W8,clk_delay);
   and MGM_G16(ENABLE_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W9);
   and MGM_G17(MGM_W10,d_delay,clk_delay);
   and MGM_G18(ENABLE_clk_AND_d_AND_rb,rb_delay,MGM_W10);
   not MGM_G19(MGM_W11,clk_delay);
   not MGM_G20(MGM_W12,d_delay);
   and MGM_G21(ENABLE_NOT_clk_AND_NOT_d,MGM_W12,MGM_W11);
   not MGM_G22(MGM_W13,clk_delay);
   and MGM_G23(ENABLE_NOT_clk_AND_d,d_delay,MGM_W13);
   not MGM_G24(MGM_W14,d_delay);
   and MGM_G25(ENABLE_clk_AND_NOT_d,MGM_W14,clk_delay);
   and MGM_G26(ENABLE_clk_AND_d,d_delay,clk_delay);
   buf MGM_G27(ENABLE_psb,psb_delay);
   not MGM_G28(MGM_W15,clk_delay);
   not MGM_G29(MGM_W16,d_delay);
   and MGM_G30(MGM_W17,MGM_W16,MGM_W15);
   and MGM_G31(ENABLE_NOT_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W17);
   not MGM_G32(MGM_W18,clk_delay);
   and MGM_G33(MGM_W19,d_delay,MGM_W18);
   and MGM_G34(ENABLE_NOT_clk_AND_d_AND_psb,psb_delay,MGM_W19);
   not MGM_G35(MGM_W20,d_delay);
   and MGM_G36(MGM_W21,MGM_W20,clk_delay);
   and MGM_G37(ENABLE_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W21);
   and MGM_G38(MGM_W22,d_delay,clk_delay);
   and MGM_G39(ENABLE_clk_AND_d_AND_psb,psb_delay,MGM_W22);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      posedge clk &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      posedge clk &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn00fah1n16x5( clk, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00fah_func b15fqn00fah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00fah_func b15fqn00fah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn00fah_func b15fqn00fah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn00fah_func b15fqn00fah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clk_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clk_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clk_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,d_delay);
   and MGM_G15(MGM_W9,MGM_W8,clk_delay);
   and MGM_G16(ENABLE_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W9);
   and MGM_G17(MGM_W10,d_delay,clk_delay);
   and MGM_G18(ENABLE_clk_AND_d_AND_rb,rb_delay,MGM_W10);
   not MGM_G19(MGM_W11,clk_delay);
   not MGM_G20(MGM_W12,d_delay);
   and MGM_G21(ENABLE_NOT_clk_AND_NOT_d,MGM_W12,MGM_W11);
   not MGM_G22(MGM_W13,clk_delay);
   and MGM_G23(ENABLE_NOT_clk_AND_d,d_delay,MGM_W13);
   not MGM_G24(MGM_W14,d_delay);
   and MGM_G25(ENABLE_clk_AND_NOT_d,MGM_W14,clk_delay);
   and MGM_G26(ENABLE_clk_AND_d,d_delay,clk_delay);
   buf MGM_G27(ENABLE_psb,psb_delay);
   not MGM_G28(MGM_W15,clk_delay);
   not MGM_G29(MGM_W16,d_delay);
   and MGM_G30(MGM_W17,MGM_W16,MGM_W15);
   and MGM_G31(ENABLE_NOT_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W17);
   not MGM_G32(MGM_W18,clk_delay);
   and MGM_G33(MGM_W19,d_delay,MGM_W18);
   and MGM_G34(ENABLE_NOT_clk_AND_d_AND_psb,psb_delay,MGM_W19);
   not MGM_G35(MGM_W20,d_delay);
   and MGM_G36(MGM_W21,MGM_W20,clk_delay);
   and MGM_G37(ENABLE_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W21);
   and MGM_G38(MGM_W22,d_delay,clk_delay);
   and MGM_G39(ENABLE_clk_AND_d_AND_psb,psb_delay,MGM_W22);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      posedge clk &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      posedge clk &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fqn043ah_func( clk, d, den, o, rb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, int1, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_fpn040ah_6( int1, IQ, d, den, vcc, vssx );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_cdiar2ah_0( MGM_D0, int1 );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_fpn040ah_6( int1, IQ, d, den );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fqn043ah1n02x5( clk, d, den, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn043ah_func b15fqn043ah1n02x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn043ah_func b15fqn043ah1n02x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn043ah_func b15fqn043ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn043ah_func b15fqn043ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,den_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_den_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,den_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_den_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_den_AND_rb,rb_delay,den_delay);
   not MGM_G6(MGM_W3,d_delay);
   and MGM_G7(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W3);
   and MGM_G8(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G9(ENABLE_den,den_delay);
   not MGM_G10(MGM_W4,clk_delay);
   not MGM_G11(MGM_W5,d_delay);
   and MGM_G12(MGM_W6,MGM_W5,MGM_W4);
   not MGM_G13(MGM_W7,den_delay);
   and MGM_G14(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den,MGM_W7,MGM_W6);
   not MGM_G15(MGM_W8,clk_delay);
   not MGM_G16(MGM_W9,d_delay);
   and MGM_G17(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G18(ENABLE_NOT_clk_AND_NOT_d_AND_den,den_delay,MGM_W10);
   not MGM_G19(MGM_W11,clk_delay);
   and MGM_G20(MGM_W12,d_delay,MGM_W11);
   not MGM_G21(MGM_W13,den_delay);
   and MGM_G22(ENABLE_NOT_clk_AND_d_AND_NOT_den,MGM_W13,MGM_W12);
   not MGM_G23(MGM_W14,clk_delay);
   and MGM_G24(MGM_W15,d_delay,MGM_W14);
   and MGM_G25(ENABLE_NOT_clk_AND_d_AND_den,den_delay,MGM_W15);
   not MGM_G26(MGM_W16,d_delay);
   and MGM_G27(MGM_W17,MGM_W16,clk_delay);
   not MGM_G28(MGM_W18,den_delay);
   and MGM_G29(ENABLE_clk_AND_NOT_d_AND_NOT_den,MGM_W18,MGM_W17);
   not MGM_G30(MGM_W19,d_delay);
   and MGM_G31(MGM_W20,MGM_W19,clk_delay);
   and MGM_G32(ENABLE_clk_AND_NOT_d_AND_den,den_delay,MGM_W20);
   and MGM_G33(MGM_W21,d_delay,clk_delay);
   not MGM_G34(MGM_W22,den_delay);
   and MGM_G35(ENABLE_clk_AND_d_AND_NOT_den,MGM_W22,MGM_W21);
   and MGM_G36(MGM_W23,d_delay,clk_delay);
   and MGM_G37(ENABLE_clk_AND_d_AND_den,den_delay,MGM_W23);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_den == 1'b1),
      posedge clk &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn043ah1n03x5( clk, d, den, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn043ah_func b15fqn043ah1n03x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn043ah_func b15fqn043ah1n03x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn043ah_func b15fqn043ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn043ah_func b15fqn043ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,den_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_den_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,den_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_den_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_den_AND_rb,rb_delay,den_delay);
   not MGM_G6(MGM_W3,d_delay);
   and MGM_G7(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W3);
   and MGM_G8(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G9(ENABLE_den,den_delay);
   not MGM_G10(MGM_W4,clk_delay);
   not MGM_G11(MGM_W5,d_delay);
   and MGM_G12(MGM_W6,MGM_W5,MGM_W4);
   not MGM_G13(MGM_W7,den_delay);
   and MGM_G14(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den,MGM_W7,MGM_W6);
   not MGM_G15(MGM_W8,clk_delay);
   not MGM_G16(MGM_W9,d_delay);
   and MGM_G17(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G18(ENABLE_NOT_clk_AND_NOT_d_AND_den,den_delay,MGM_W10);
   not MGM_G19(MGM_W11,clk_delay);
   and MGM_G20(MGM_W12,d_delay,MGM_W11);
   not MGM_G21(MGM_W13,den_delay);
   and MGM_G22(ENABLE_NOT_clk_AND_d_AND_NOT_den,MGM_W13,MGM_W12);
   not MGM_G23(MGM_W14,clk_delay);
   and MGM_G24(MGM_W15,d_delay,MGM_W14);
   and MGM_G25(ENABLE_NOT_clk_AND_d_AND_den,den_delay,MGM_W15);
   not MGM_G26(MGM_W16,d_delay);
   and MGM_G27(MGM_W17,MGM_W16,clk_delay);
   not MGM_G28(MGM_W18,den_delay);
   and MGM_G29(ENABLE_clk_AND_NOT_d_AND_NOT_den,MGM_W18,MGM_W17);
   not MGM_G30(MGM_W19,d_delay);
   and MGM_G31(MGM_W20,MGM_W19,clk_delay);
   and MGM_G32(ENABLE_clk_AND_NOT_d_AND_den,den_delay,MGM_W20);
   and MGM_G33(MGM_W21,d_delay,clk_delay);
   not MGM_G34(MGM_W22,den_delay);
   and MGM_G35(ENABLE_clk_AND_d_AND_NOT_den,MGM_W22,MGM_W21);
   and MGM_G36(MGM_W23,d_delay,clk_delay);
   and MGM_G37(ENABLE_clk_AND_d_AND_den,den_delay,MGM_W23);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_den == 1'b1),
      posedge clk &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn043ah1n04x5( clk, d, den, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn043ah_func b15fqn043ah1n04x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn043ah_func b15fqn043ah1n04x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn043ah_func b15fqn043ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn043ah_func b15fqn043ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,den_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_den_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,den_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_den_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_den_AND_rb,rb_delay,den_delay);
   not MGM_G6(MGM_W3,d_delay);
   and MGM_G7(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W3);
   and MGM_G8(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G9(ENABLE_den,den_delay);
   not MGM_G10(MGM_W4,clk_delay);
   not MGM_G11(MGM_W5,d_delay);
   and MGM_G12(MGM_W6,MGM_W5,MGM_W4);
   not MGM_G13(MGM_W7,den_delay);
   and MGM_G14(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den,MGM_W7,MGM_W6);
   not MGM_G15(MGM_W8,clk_delay);
   not MGM_G16(MGM_W9,d_delay);
   and MGM_G17(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G18(ENABLE_NOT_clk_AND_NOT_d_AND_den,den_delay,MGM_W10);
   not MGM_G19(MGM_W11,clk_delay);
   and MGM_G20(MGM_W12,d_delay,MGM_W11);
   not MGM_G21(MGM_W13,den_delay);
   and MGM_G22(ENABLE_NOT_clk_AND_d_AND_NOT_den,MGM_W13,MGM_W12);
   not MGM_G23(MGM_W14,clk_delay);
   and MGM_G24(MGM_W15,d_delay,MGM_W14);
   and MGM_G25(ENABLE_NOT_clk_AND_d_AND_den,den_delay,MGM_W15);
   not MGM_G26(MGM_W16,d_delay);
   and MGM_G27(MGM_W17,MGM_W16,clk_delay);
   not MGM_G28(MGM_W18,den_delay);
   and MGM_G29(ENABLE_clk_AND_NOT_d_AND_NOT_den,MGM_W18,MGM_W17);
   not MGM_G30(MGM_W19,d_delay);
   and MGM_G31(MGM_W20,MGM_W19,clk_delay);
   and MGM_G32(ENABLE_clk_AND_NOT_d_AND_den,den_delay,MGM_W20);
   and MGM_G33(MGM_W21,d_delay,clk_delay);
   not MGM_G34(MGM_W22,den_delay);
   and MGM_G35(ENABLE_clk_AND_d_AND_NOT_den,MGM_W22,MGM_W21);
   and MGM_G36(MGM_W23,d_delay,clk_delay);
   and MGM_G37(ENABLE_clk_AND_d_AND_den,den_delay,MGM_W23);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_den == 1'b1),
      posedge clk &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn043ah1n06x5( clk, d, den, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn043ah_func b15fqn043ah1n06x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn043ah_func b15fqn043ah1n06x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn043ah_func b15fqn043ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn043ah_func b15fqn043ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,den_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_den_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,den_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_den_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_den_AND_rb,rb_delay,den_delay);
   not MGM_G6(MGM_W3,d_delay);
   and MGM_G7(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W3);
   and MGM_G8(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G9(ENABLE_den,den_delay);
   not MGM_G10(MGM_W4,clk_delay);
   not MGM_G11(MGM_W5,d_delay);
   and MGM_G12(MGM_W6,MGM_W5,MGM_W4);
   not MGM_G13(MGM_W7,den_delay);
   and MGM_G14(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den,MGM_W7,MGM_W6);
   not MGM_G15(MGM_W8,clk_delay);
   not MGM_G16(MGM_W9,d_delay);
   and MGM_G17(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G18(ENABLE_NOT_clk_AND_NOT_d_AND_den,den_delay,MGM_W10);
   not MGM_G19(MGM_W11,clk_delay);
   and MGM_G20(MGM_W12,d_delay,MGM_W11);
   not MGM_G21(MGM_W13,den_delay);
   and MGM_G22(ENABLE_NOT_clk_AND_d_AND_NOT_den,MGM_W13,MGM_W12);
   not MGM_G23(MGM_W14,clk_delay);
   and MGM_G24(MGM_W15,d_delay,MGM_W14);
   and MGM_G25(ENABLE_NOT_clk_AND_d_AND_den,den_delay,MGM_W15);
   not MGM_G26(MGM_W16,d_delay);
   and MGM_G27(MGM_W17,MGM_W16,clk_delay);
   not MGM_G28(MGM_W18,den_delay);
   and MGM_G29(ENABLE_clk_AND_NOT_d_AND_NOT_den,MGM_W18,MGM_W17);
   not MGM_G30(MGM_W19,d_delay);
   and MGM_G31(MGM_W20,MGM_W19,clk_delay);
   and MGM_G32(ENABLE_clk_AND_NOT_d_AND_den,den_delay,MGM_W20);
   and MGM_G33(MGM_W21,d_delay,clk_delay);
   not MGM_G34(MGM_W22,den_delay);
   and MGM_G35(ENABLE_clk_AND_d_AND_NOT_den,MGM_W22,MGM_W21);
   and MGM_G36(MGM_W23,d_delay,clk_delay);
   and MGM_G37(ENABLE_clk_AND_d_AND_den,den_delay,MGM_W23);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_den == 1'b1),
      posedge clk &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn043ah1n08x5( clk, d, den, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn043ah_func b15fqn043ah1n08x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn043ah_func b15fqn043ah1n08x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn043ah_func b15fqn043ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn043ah_func b15fqn043ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,den_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_den_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,den_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_den_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_den_AND_rb,rb_delay,den_delay);
   not MGM_G6(MGM_W3,d_delay);
   and MGM_G7(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W3);
   and MGM_G8(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G9(ENABLE_den,den_delay);
   not MGM_G10(MGM_W4,clk_delay);
   not MGM_G11(MGM_W5,d_delay);
   and MGM_G12(MGM_W6,MGM_W5,MGM_W4);
   not MGM_G13(MGM_W7,den_delay);
   and MGM_G14(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den,MGM_W7,MGM_W6);
   not MGM_G15(MGM_W8,clk_delay);
   not MGM_G16(MGM_W9,d_delay);
   and MGM_G17(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G18(ENABLE_NOT_clk_AND_NOT_d_AND_den,den_delay,MGM_W10);
   not MGM_G19(MGM_W11,clk_delay);
   and MGM_G20(MGM_W12,d_delay,MGM_W11);
   not MGM_G21(MGM_W13,den_delay);
   and MGM_G22(ENABLE_NOT_clk_AND_d_AND_NOT_den,MGM_W13,MGM_W12);
   not MGM_G23(MGM_W14,clk_delay);
   and MGM_G24(MGM_W15,d_delay,MGM_W14);
   and MGM_G25(ENABLE_NOT_clk_AND_d_AND_den,den_delay,MGM_W15);
   not MGM_G26(MGM_W16,d_delay);
   and MGM_G27(MGM_W17,MGM_W16,clk_delay);
   not MGM_G28(MGM_W18,den_delay);
   and MGM_G29(ENABLE_clk_AND_NOT_d_AND_NOT_den,MGM_W18,MGM_W17);
   not MGM_G30(MGM_W19,d_delay);
   and MGM_G31(MGM_W20,MGM_W19,clk_delay);
   and MGM_G32(ENABLE_clk_AND_NOT_d_AND_den,den_delay,MGM_W20);
   and MGM_G33(MGM_W21,d_delay,clk_delay);
   not MGM_G34(MGM_W22,den_delay);
   and MGM_G35(ENABLE_clk_AND_d_AND_NOT_den,MGM_W22,MGM_W21);
   and MGM_G36(MGM_W23,d_delay,clk_delay);
   and MGM_G37(ENABLE_clk_AND_d_AND_den,den_delay,MGM_W23);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_den == 1'b1),
      posedge clk &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn043ah1n12x5( clk, d, den, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn043ah_func b15fqn043ah1n12x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn043ah_func b15fqn043ah1n12x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn043ah_func b15fqn043ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn043ah_func b15fqn043ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,den_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_den_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,den_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_den_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_den_AND_rb,rb_delay,den_delay);
   not MGM_G6(MGM_W3,d_delay);
   and MGM_G7(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W3);
   and MGM_G8(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G9(ENABLE_den,den_delay);
   not MGM_G10(MGM_W4,clk_delay);
   not MGM_G11(MGM_W5,d_delay);
   and MGM_G12(MGM_W6,MGM_W5,MGM_W4);
   not MGM_G13(MGM_W7,den_delay);
   and MGM_G14(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den,MGM_W7,MGM_W6);
   not MGM_G15(MGM_W8,clk_delay);
   not MGM_G16(MGM_W9,d_delay);
   and MGM_G17(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G18(ENABLE_NOT_clk_AND_NOT_d_AND_den,den_delay,MGM_W10);
   not MGM_G19(MGM_W11,clk_delay);
   and MGM_G20(MGM_W12,d_delay,MGM_W11);
   not MGM_G21(MGM_W13,den_delay);
   and MGM_G22(ENABLE_NOT_clk_AND_d_AND_NOT_den,MGM_W13,MGM_W12);
   not MGM_G23(MGM_W14,clk_delay);
   and MGM_G24(MGM_W15,d_delay,MGM_W14);
   and MGM_G25(ENABLE_NOT_clk_AND_d_AND_den,den_delay,MGM_W15);
   not MGM_G26(MGM_W16,d_delay);
   and MGM_G27(MGM_W17,MGM_W16,clk_delay);
   not MGM_G28(MGM_W18,den_delay);
   and MGM_G29(ENABLE_clk_AND_NOT_d_AND_NOT_den,MGM_W18,MGM_W17);
   not MGM_G30(MGM_W19,d_delay);
   and MGM_G31(MGM_W20,MGM_W19,clk_delay);
   and MGM_G32(ENABLE_clk_AND_NOT_d_AND_den,den_delay,MGM_W20);
   and MGM_G33(MGM_W21,d_delay,clk_delay);
   not MGM_G34(MGM_W22,den_delay);
   and MGM_G35(ENABLE_clk_AND_d_AND_NOT_den,MGM_W22,MGM_W21);
   and MGM_G36(MGM_W23,d_delay,clk_delay);
   and MGM_G37(ENABLE_clk_AND_d_AND_den,den_delay,MGM_W23);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_den == 1'b1),
      posedge clk &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn043ah1n16x5( clk, d, den, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn043ah_func b15fqn043ah1n16x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn043ah_func b15fqn043ah1n16x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn043ah_func b15fqn043ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn043ah_func b15fqn043ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,den_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_den_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,den_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_den_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_den_AND_rb,rb_delay,den_delay);
   not MGM_G6(MGM_W3,d_delay);
   and MGM_G7(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W3);
   and MGM_G8(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G9(ENABLE_den,den_delay);
   not MGM_G10(MGM_W4,clk_delay);
   not MGM_G11(MGM_W5,d_delay);
   and MGM_G12(MGM_W6,MGM_W5,MGM_W4);
   not MGM_G13(MGM_W7,den_delay);
   and MGM_G14(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den,MGM_W7,MGM_W6);
   not MGM_G15(MGM_W8,clk_delay);
   not MGM_G16(MGM_W9,d_delay);
   and MGM_G17(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G18(ENABLE_NOT_clk_AND_NOT_d_AND_den,den_delay,MGM_W10);
   not MGM_G19(MGM_W11,clk_delay);
   and MGM_G20(MGM_W12,d_delay,MGM_W11);
   not MGM_G21(MGM_W13,den_delay);
   and MGM_G22(ENABLE_NOT_clk_AND_d_AND_NOT_den,MGM_W13,MGM_W12);
   not MGM_G23(MGM_W14,clk_delay);
   and MGM_G24(MGM_W15,d_delay,MGM_W14);
   and MGM_G25(ENABLE_NOT_clk_AND_d_AND_den,den_delay,MGM_W15);
   not MGM_G26(MGM_W16,d_delay);
   and MGM_G27(MGM_W17,MGM_W16,clk_delay);
   not MGM_G28(MGM_W18,den_delay);
   and MGM_G29(ENABLE_clk_AND_NOT_d_AND_NOT_den,MGM_W18,MGM_W17);
   not MGM_G30(MGM_W19,d_delay);
   and MGM_G31(MGM_W20,MGM_W19,clk_delay);
   and MGM_G32(ENABLE_clk_AND_NOT_d_AND_den,den_delay,MGM_W20);
   and MGM_G33(MGM_W21,d_delay,clk_delay);
   not MGM_G34(MGM_W22,den_delay);
   and MGM_G35(ENABLE_clk_AND_d_AND_NOT_den,MGM_W22,MGM_W21);
   and MGM_G36(MGM_W23,d_delay,clk_delay);
   and MGM_G37(ENABLE_clk_AND_d_AND_den,den_delay,MGM_W23);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_den == 1'b1),
      posedge clk &&& (ENABLE_den == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fqn08fah_func( clkb, d, o, psb, rb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, psb, rb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_1( MGM_CLK0, clkb, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_P0, psb, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, d, vcc, vssx );
   INTCseq_fqn00fah_LN_IQ_FF_UDP( IQ, MGM_C0, MGM_P0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_1( MGM_CLK0, clkb );
   INTCseq_cdiar2ah_1( MGM_P0, psb );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_cdiar2ah_0( MGM_D0, d );
   INTCseq_fqn00fah_LN_IQ_FF_UDP( IQ, MGM_C0, MGM_P0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fqn08fah1n02x5( clkb, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn08fah_func b15fqn08fah1n02x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn08fah_func b15fqn08fah1n02x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn08fah_func b15fqn08fah1n02x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn08fah_func b15fqn08fah1n02x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clkb_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clkb_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clkb_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clkb_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,d_delay);
   and MGM_G15(MGM_W9,MGM_W8,clkb_delay);
   and MGM_G16(ENABLE_clkb_AND_NOT_d_AND_rb,rb_delay,MGM_W9);
   and MGM_G17(MGM_W10,d_delay,clkb_delay);
   and MGM_G18(ENABLE_clkb_AND_d_AND_rb,rb_delay,MGM_W10);
   not MGM_G19(MGM_W11,clkb_delay);
   not MGM_G20(MGM_W12,d_delay);
   and MGM_G21(ENABLE_NOT_clkb_AND_NOT_d,MGM_W12,MGM_W11);
   not MGM_G22(MGM_W13,clkb_delay);
   and MGM_G23(ENABLE_NOT_clkb_AND_d,d_delay,MGM_W13);
   not MGM_G24(MGM_W14,d_delay);
   and MGM_G25(ENABLE_clkb_AND_NOT_d,MGM_W14,clkb_delay);
   and MGM_G26(ENABLE_clkb_AND_d,d_delay,clkb_delay);
   buf MGM_G27(ENABLE_psb,psb_delay);
   not MGM_G28(MGM_W15,clkb_delay);
   not MGM_G29(MGM_W16,d_delay);
   and MGM_G30(MGM_W17,MGM_W16,MGM_W15);
   and MGM_G31(ENABLE_NOT_clkb_AND_NOT_d_AND_psb,psb_delay,MGM_W17);
   not MGM_G32(MGM_W18,clkb_delay);
   and MGM_G33(MGM_W19,d_delay,MGM_W18);
   and MGM_G34(ENABLE_NOT_clkb_AND_d_AND_psb,psb_delay,MGM_W19);
   not MGM_G35(MGM_W20,d_delay);
   and MGM_G36(MGM_W21,MGM_W20,clkb_delay);
   and MGM_G37(ENABLE_clkb_AND_NOT_d_AND_psb,psb_delay,MGM_W21);
   and MGM_G38(MGM_W22,d_delay,clkb_delay);
   and MGM_G39(ENABLE_clkb_AND_d_AND_psb,psb_delay,MGM_W22);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      negedge clkb &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      negedge clkb &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn08fah1n04x5( clkb, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn08fah_func b15fqn08fah1n04x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn08fah_func b15fqn08fah1n04x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn08fah_func b15fqn08fah1n04x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn08fah_func b15fqn08fah1n04x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clkb_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clkb_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clkb_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clkb_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,d_delay);
   and MGM_G15(MGM_W9,MGM_W8,clkb_delay);
   and MGM_G16(ENABLE_clkb_AND_NOT_d_AND_rb,rb_delay,MGM_W9);
   and MGM_G17(MGM_W10,d_delay,clkb_delay);
   and MGM_G18(ENABLE_clkb_AND_d_AND_rb,rb_delay,MGM_W10);
   not MGM_G19(MGM_W11,clkb_delay);
   not MGM_G20(MGM_W12,d_delay);
   and MGM_G21(ENABLE_NOT_clkb_AND_NOT_d,MGM_W12,MGM_W11);
   not MGM_G22(MGM_W13,clkb_delay);
   and MGM_G23(ENABLE_NOT_clkb_AND_d,d_delay,MGM_W13);
   not MGM_G24(MGM_W14,d_delay);
   and MGM_G25(ENABLE_clkb_AND_NOT_d,MGM_W14,clkb_delay);
   and MGM_G26(ENABLE_clkb_AND_d,d_delay,clkb_delay);
   buf MGM_G27(ENABLE_psb,psb_delay);
   not MGM_G28(MGM_W15,clkb_delay);
   not MGM_G29(MGM_W16,d_delay);
   and MGM_G30(MGM_W17,MGM_W16,MGM_W15);
   and MGM_G31(ENABLE_NOT_clkb_AND_NOT_d_AND_psb,psb_delay,MGM_W17);
   not MGM_G32(MGM_W18,clkb_delay);
   and MGM_G33(MGM_W19,d_delay,MGM_W18);
   and MGM_G34(ENABLE_NOT_clkb_AND_d_AND_psb,psb_delay,MGM_W19);
   not MGM_G35(MGM_W20,d_delay);
   and MGM_G36(MGM_W21,MGM_W20,clkb_delay);
   and MGM_G37(ENABLE_clkb_AND_NOT_d_AND_psb,psb_delay,MGM_W21);
   and MGM_G38(MGM_W22,d_delay,clkb_delay);
   and MGM_G39(ENABLE_clkb_AND_d_AND_psb,psb_delay,MGM_W22);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      negedge clkb &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      negedge clkb &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn08fah1n08x5( clkb, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn08fah_func b15fqn08fah1n08x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn08fah_func b15fqn08fah1n08x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn08fah_func b15fqn08fah1n08x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn08fah_func b15fqn08fah1n08x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clkb_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clkb_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clkb_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clkb_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,d_delay);
   and MGM_G15(MGM_W9,MGM_W8,clkb_delay);
   and MGM_G16(ENABLE_clkb_AND_NOT_d_AND_rb,rb_delay,MGM_W9);
   and MGM_G17(MGM_W10,d_delay,clkb_delay);
   and MGM_G18(ENABLE_clkb_AND_d_AND_rb,rb_delay,MGM_W10);
   not MGM_G19(MGM_W11,clkb_delay);
   not MGM_G20(MGM_W12,d_delay);
   and MGM_G21(ENABLE_NOT_clkb_AND_NOT_d,MGM_W12,MGM_W11);
   not MGM_G22(MGM_W13,clkb_delay);
   and MGM_G23(ENABLE_NOT_clkb_AND_d,d_delay,MGM_W13);
   not MGM_G24(MGM_W14,d_delay);
   and MGM_G25(ENABLE_clkb_AND_NOT_d,MGM_W14,clkb_delay);
   and MGM_G26(ENABLE_clkb_AND_d,d_delay,clkb_delay);
   buf MGM_G27(ENABLE_psb,psb_delay);
   not MGM_G28(MGM_W15,clkb_delay);
   not MGM_G29(MGM_W16,d_delay);
   and MGM_G30(MGM_W17,MGM_W16,MGM_W15);
   and MGM_G31(ENABLE_NOT_clkb_AND_NOT_d_AND_psb,psb_delay,MGM_W17);
   not MGM_G32(MGM_W18,clkb_delay);
   and MGM_G33(MGM_W19,d_delay,MGM_W18);
   and MGM_G34(ENABLE_NOT_clkb_AND_d_AND_psb,psb_delay,MGM_W19);
   not MGM_G35(MGM_W20,d_delay);
   and MGM_G36(MGM_W21,MGM_W20,clkb_delay);
   and MGM_G37(ENABLE_clkb_AND_NOT_d_AND_psb,psb_delay,MGM_W21);
   and MGM_G38(MGM_W22,d_delay,clkb_delay);
   and MGM_G39(ENABLE_clkb_AND_d_AND_psb,psb_delay,MGM_W22);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      negedge clkb &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      negedge clkb &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqn08fah1n16x5( clkb, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn08fah_func b15fqn08fah1n16x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn08fah_func b15fqn08fah1n16x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqn08fah_func b15fqn08fah1n16x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqn08fah_func b15fqn08fah1n16x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clkb_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clkb_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clkb_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clkb_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,d_delay);
   and MGM_G15(MGM_W9,MGM_W8,clkb_delay);
   and MGM_G16(ENABLE_clkb_AND_NOT_d_AND_rb,rb_delay,MGM_W9);
   and MGM_G17(MGM_W10,d_delay,clkb_delay);
   and MGM_G18(ENABLE_clkb_AND_d_AND_rb,rb_delay,MGM_W10);
   not MGM_G19(MGM_W11,clkb_delay);
   not MGM_G20(MGM_W12,d_delay);
   and MGM_G21(ENABLE_NOT_clkb_AND_NOT_d,MGM_W12,MGM_W11);
   not MGM_G22(MGM_W13,clkb_delay);
   and MGM_G23(ENABLE_NOT_clkb_AND_d,d_delay,MGM_W13);
   not MGM_G24(MGM_W14,d_delay);
   and MGM_G25(ENABLE_clkb_AND_NOT_d,MGM_W14,clkb_delay);
   and MGM_G26(ENABLE_clkb_AND_d,d_delay,clkb_delay);
   buf MGM_G27(ENABLE_psb,psb_delay);
   not MGM_G28(MGM_W15,clkb_delay);
   not MGM_G29(MGM_W16,d_delay);
   and MGM_G30(MGM_W17,MGM_W16,MGM_W15);
   and MGM_G31(ENABLE_NOT_clkb_AND_NOT_d_AND_psb,psb_delay,MGM_W17);
   not MGM_G32(MGM_W18,clkb_delay);
   and MGM_G33(MGM_W19,d_delay,MGM_W18);
   and MGM_G34(ENABLE_NOT_clkb_AND_d_AND_psb,psb_delay,MGM_W19);
   not MGM_G35(MGM_W20,d_delay);
   and MGM_G36(MGM_W21,MGM_W20,clkb_delay);
   and MGM_G37(ENABLE_clkb_AND_NOT_d_AND_psb,psb_delay,MGM_W21);
   and MGM_G38(MGM_W22,d_delay,clkb_delay);
   and MGM_G39(ENABLE_clkb_AND_d_AND_psb,psb_delay,MGM_W22);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      negedge clkb &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      negedge clkb &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fqy003ah_func( clk, d, o, rb, si, ssb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fqy003ah1n02x5( clk, d, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy003ah_func b15fqy003ah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy003ah_func b15fqy003ah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy003ah_func b15fqy003ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy003ah_func b15fqy003ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,rb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,rb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,rb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,rb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,rb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,rb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,rb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,rb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,rb_delay);
   and MGM_G38(ENABLE_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,rb_delay);
   and MGM_G40(ENABLE_rb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   and MGM_G42(MGM_W32,si_delay,MGM_W31);
   not MGM_G43(MGM_W33,ssb_delay);
   and MGM_G44(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W33,MGM_W32);
   not MGM_G45(MGM_W34,si_delay);
   and MGM_G46(MGM_W35,MGM_W34,d_delay);
   and MGM_G47(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G48(MGM_W36,si_delay,d_delay);
   not MGM_G49(MGM_W37,ssb_delay);
   and MGM_G50(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W37,MGM_W36);
   and MGM_G51(MGM_W38,si_delay,d_delay);
   and MGM_G52(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W38);
   not MGM_G53(MGM_W39,clk_delay);
   not MGM_G54(MGM_W40,d_delay);
   and MGM_G55(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G56(MGM_W42,si_delay);
   and MGM_G57(MGM_W43,MGM_W42,MGM_W41);
   not MGM_G58(MGM_W44,ssb_delay);
   and MGM_G59(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W45,clk_delay);
   not MGM_G61(MGM_W46,d_delay);
   and MGM_G62(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G63(MGM_W48,si_delay);
   and MGM_G64(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G65(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G66(MGM_W50,clk_delay);
   not MGM_G67(MGM_W51,d_delay);
   and MGM_G68(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G69(MGM_W53,si_delay,MGM_W52);
   not MGM_G70(MGM_W54,ssb_delay);
   and MGM_G71(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W54,MGM_W53);
   not MGM_G72(MGM_W55,clk_delay);
   not MGM_G73(MGM_W56,d_delay);
   and MGM_G74(MGM_W57,MGM_W56,MGM_W55);
   and MGM_G75(MGM_W58,si_delay,MGM_W57);
   and MGM_G76(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,clk_delay);
   and MGM_G78(MGM_W60,d_delay,MGM_W59);
   not MGM_G79(MGM_W61,si_delay);
   and MGM_G80(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G81(MGM_W63,ssb_delay);
   and MGM_G82(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G83(MGM_W64,clk_delay);
   and MGM_G84(MGM_W65,d_delay,MGM_W64);
   not MGM_G85(MGM_W66,si_delay);
   and MGM_G86(MGM_W67,MGM_W66,MGM_W65);
   and MGM_G87(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W67);
   not MGM_G88(MGM_W68,clk_delay);
   and MGM_G89(MGM_W69,d_delay,MGM_W68);
   and MGM_G90(MGM_W70,si_delay,MGM_W69);
   not MGM_G91(MGM_W71,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W71,MGM_W70);
   not MGM_G93(MGM_W72,clk_delay);
   and MGM_G94(MGM_W73,d_delay,MGM_W72);
   and MGM_G95(MGM_W74,si_delay,MGM_W73);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W74);
   not MGM_G97(MGM_W75,d_delay);
   and MGM_G98(MGM_W76,MGM_W75,clk_delay);
   not MGM_G99(MGM_W77,si_delay);
   and MGM_G100(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G101(MGM_W79,ssb_delay);
   and MGM_G102(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G103(MGM_W80,d_delay);
   and MGM_G104(MGM_W81,MGM_W80,clk_delay);
   not MGM_G105(MGM_W82,si_delay);
   and MGM_G106(MGM_W83,MGM_W82,MGM_W81);
   and MGM_G107(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W83);
   not MGM_G108(MGM_W84,d_delay);
   and MGM_G109(MGM_W85,MGM_W84,clk_delay);
   and MGM_G110(MGM_W86,si_delay,MGM_W85);
   not MGM_G111(MGM_W87,ssb_delay);
   and MGM_G112(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W87,MGM_W86);
   not MGM_G113(MGM_W88,d_delay);
   and MGM_G114(MGM_W89,MGM_W88,clk_delay);
   and MGM_G115(MGM_W90,si_delay,MGM_W89);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W90);
   and MGM_G117(MGM_W91,d_delay,clk_delay);
   not MGM_G118(MGM_W92,si_delay);
   and MGM_G119(MGM_W93,MGM_W92,MGM_W91);
   not MGM_G120(MGM_W94,ssb_delay);
   and MGM_G121(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W94,MGM_W93);
   and MGM_G122(MGM_W95,d_delay,clk_delay);
   not MGM_G123(MGM_W96,si_delay);
   and MGM_G124(MGM_W97,MGM_W96,MGM_W95);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W97);
   and MGM_G126(MGM_W98,d_delay,clk_delay);
   and MGM_G127(MGM_W99,si_delay,MGM_W98);
   not MGM_G128(MGM_W100,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W100,MGM_W99);
   and MGM_G130(MGM_W101,d_delay,clk_delay);
   and MGM_G131(MGM_W102,si_delay,MGM_W101);
   and MGM_G132(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W102);
   not MGM_G133(MGM_W103,d_delay);
   and MGM_G134(MGM_W104,rb_delay,MGM_W103);
   not MGM_G135(MGM_W105,ssb_delay);
   and MGM_G136(ENABLE_NOT_d_AND_rb_AND_NOT_ssb,MGM_W105,MGM_W104);
   and MGM_G137(MGM_W106,rb_delay,d_delay);
   not MGM_G138(MGM_W107,ssb_delay);
   and MGM_G139(ENABLE_d_AND_rb_AND_NOT_ssb,MGM_W107,MGM_W106);
   not MGM_G140(MGM_W108,d_delay);
   and MGM_G141(MGM_W109,rb_delay,MGM_W108);
   and MGM_G142(ENABLE_NOT_d_AND_rb_AND_si,si_delay,MGM_W109);
   and MGM_G143(MGM_W110,rb_delay,d_delay);
   not MGM_G144(MGM_W111,si_delay);
   and MGM_G145(ENABLE_d_AND_rb_AND_NOT_si,MGM_W111,MGM_W110);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy003ah1n03x5( clk, d, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy003ah_func b15fqy003ah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy003ah_func b15fqy003ah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy003ah_func b15fqy003ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy003ah_func b15fqy003ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,rb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,rb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,rb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,rb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,rb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,rb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,rb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,rb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,rb_delay);
   and MGM_G38(ENABLE_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,rb_delay);
   and MGM_G40(ENABLE_rb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   and MGM_G42(MGM_W32,si_delay,MGM_W31);
   not MGM_G43(MGM_W33,ssb_delay);
   and MGM_G44(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W33,MGM_W32);
   not MGM_G45(MGM_W34,si_delay);
   and MGM_G46(MGM_W35,MGM_W34,d_delay);
   and MGM_G47(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G48(MGM_W36,si_delay,d_delay);
   not MGM_G49(MGM_W37,ssb_delay);
   and MGM_G50(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W37,MGM_W36);
   and MGM_G51(MGM_W38,si_delay,d_delay);
   and MGM_G52(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W38);
   not MGM_G53(MGM_W39,clk_delay);
   not MGM_G54(MGM_W40,d_delay);
   and MGM_G55(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G56(MGM_W42,si_delay);
   and MGM_G57(MGM_W43,MGM_W42,MGM_W41);
   not MGM_G58(MGM_W44,ssb_delay);
   and MGM_G59(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W45,clk_delay);
   not MGM_G61(MGM_W46,d_delay);
   and MGM_G62(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G63(MGM_W48,si_delay);
   and MGM_G64(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G65(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G66(MGM_W50,clk_delay);
   not MGM_G67(MGM_W51,d_delay);
   and MGM_G68(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G69(MGM_W53,si_delay,MGM_W52);
   not MGM_G70(MGM_W54,ssb_delay);
   and MGM_G71(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W54,MGM_W53);
   not MGM_G72(MGM_W55,clk_delay);
   not MGM_G73(MGM_W56,d_delay);
   and MGM_G74(MGM_W57,MGM_W56,MGM_W55);
   and MGM_G75(MGM_W58,si_delay,MGM_W57);
   and MGM_G76(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,clk_delay);
   and MGM_G78(MGM_W60,d_delay,MGM_W59);
   not MGM_G79(MGM_W61,si_delay);
   and MGM_G80(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G81(MGM_W63,ssb_delay);
   and MGM_G82(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G83(MGM_W64,clk_delay);
   and MGM_G84(MGM_W65,d_delay,MGM_W64);
   not MGM_G85(MGM_W66,si_delay);
   and MGM_G86(MGM_W67,MGM_W66,MGM_W65);
   and MGM_G87(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W67);
   not MGM_G88(MGM_W68,clk_delay);
   and MGM_G89(MGM_W69,d_delay,MGM_W68);
   and MGM_G90(MGM_W70,si_delay,MGM_W69);
   not MGM_G91(MGM_W71,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W71,MGM_W70);
   not MGM_G93(MGM_W72,clk_delay);
   and MGM_G94(MGM_W73,d_delay,MGM_W72);
   and MGM_G95(MGM_W74,si_delay,MGM_W73);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W74);
   not MGM_G97(MGM_W75,d_delay);
   and MGM_G98(MGM_W76,MGM_W75,clk_delay);
   not MGM_G99(MGM_W77,si_delay);
   and MGM_G100(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G101(MGM_W79,ssb_delay);
   and MGM_G102(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G103(MGM_W80,d_delay);
   and MGM_G104(MGM_W81,MGM_W80,clk_delay);
   not MGM_G105(MGM_W82,si_delay);
   and MGM_G106(MGM_W83,MGM_W82,MGM_W81);
   and MGM_G107(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W83);
   not MGM_G108(MGM_W84,d_delay);
   and MGM_G109(MGM_W85,MGM_W84,clk_delay);
   and MGM_G110(MGM_W86,si_delay,MGM_W85);
   not MGM_G111(MGM_W87,ssb_delay);
   and MGM_G112(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W87,MGM_W86);
   not MGM_G113(MGM_W88,d_delay);
   and MGM_G114(MGM_W89,MGM_W88,clk_delay);
   and MGM_G115(MGM_W90,si_delay,MGM_W89);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W90);
   and MGM_G117(MGM_W91,d_delay,clk_delay);
   not MGM_G118(MGM_W92,si_delay);
   and MGM_G119(MGM_W93,MGM_W92,MGM_W91);
   not MGM_G120(MGM_W94,ssb_delay);
   and MGM_G121(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W94,MGM_W93);
   and MGM_G122(MGM_W95,d_delay,clk_delay);
   not MGM_G123(MGM_W96,si_delay);
   and MGM_G124(MGM_W97,MGM_W96,MGM_W95);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W97);
   and MGM_G126(MGM_W98,d_delay,clk_delay);
   and MGM_G127(MGM_W99,si_delay,MGM_W98);
   not MGM_G128(MGM_W100,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W100,MGM_W99);
   and MGM_G130(MGM_W101,d_delay,clk_delay);
   and MGM_G131(MGM_W102,si_delay,MGM_W101);
   and MGM_G132(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W102);
   not MGM_G133(MGM_W103,d_delay);
   and MGM_G134(MGM_W104,rb_delay,MGM_W103);
   not MGM_G135(MGM_W105,ssb_delay);
   and MGM_G136(ENABLE_NOT_d_AND_rb_AND_NOT_ssb,MGM_W105,MGM_W104);
   and MGM_G137(MGM_W106,rb_delay,d_delay);
   not MGM_G138(MGM_W107,ssb_delay);
   and MGM_G139(ENABLE_d_AND_rb_AND_NOT_ssb,MGM_W107,MGM_W106);
   not MGM_G140(MGM_W108,d_delay);
   and MGM_G141(MGM_W109,rb_delay,MGM_W108);
   and MGM_G142(ENABLE_NOT_d_AND_rb_AND_si,si_delay,MGM_W109);
   and MGM_G143(MGM_W110,rb_delay,d_delay);
   not MGM_G144(MGM_W111,si_delay);
   and MGM_G145(ENABLE_d_AND_rb_AND_NOT_si,MGM_W111,MGM_W110);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy003ah1n04x5( clk, d, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy003ah_func b15fqy003ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy003ah_func b15fqy003ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy003ah_func b15fqy003ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy003ah_func b15fqy003ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,rb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,rb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,rb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,rb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,rb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,rb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,rb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,rb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,rb_delay);
   and MGM_G38(ENABLE_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,rb_delay);
   and MGM_G40(ENABLE_rb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   and MGM_G42(MGM_W32,si_delay,MGM_W31);
   not MGM_G43(MGM_W33,ssb_delay);
   and MGM_G44(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W33,MGM_W32);
   not MGM_G45(MGM_W34,si_delay);
   and MGM_G46(MGM_W35,MGM_W34,d_delay);
   and MGM_G47(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G48(MGM_W36,si_delay,d_delay);
   not MGM_G49(MGM_W37,ssb_delay);
   and MGM_G50(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W37,MGM_W36);
   and MGM_G51(MGM_W38,si_delay,d_delay);
   and MGM_G52(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W38);
   not MGM_G53(MGM_W39,clk_delay);
   not MGM_G54(MGM_W40,d_delay);
   and MGM_G55(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G56(MGM_W42,si_delay);
   and MGM_G57(MGM_W43,MGM_W42,MGM_W41);
   not MGM_G58(MGM_W44,ssb_delay);
   and MGM_G59(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W45,clk_delay);
   not MGM_G61(MGM_W46,d_delay);
   and MGM_G62(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G63(MGM_W48,si_delay);
   and MGM_G64(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G65(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G66(MGM_W50,clk_delay);
   not MGM_G67(MGM_W51,d_delay);
   and MGM_G68(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G69(MGM_W53,si_delay,MGM_W52);
   not MGM_G70(MGM_W54,ssb_delay);
   and MGM_G71(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W54,MGM_W53);
   not MGM_G72(MGM_W55,clk_delay);
   not MGM_G73(MGM_W56,d_delay);
   and MGM_G74(MGM_W57,MGM_W56,MGM_W55);
   and MGM_G75(MGM_W58,si_delay,MGM_W57);
   and MGM_G76(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,clk_delay);
   and MGM_G78(MGM_W60,d_delay,MGM_W59);
   not MGM_G79(MGM_W61,si_delay);
   and MGM_G80(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G81(MGM_W63,ssb_delay);
   and MGM_G82(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G83(MGM_W64,clk_delay);
   and MGM_G84(MGM_W65,d_delay,MGM_W64);
   not MGM_G85(MGM_W66,si_delay);
   and MGM_G86(MGM_W67,MGM_W66,MGM_W65);
   and MGM_G87(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W67);
   not MGM_G88(MGM_W68,clk_delay);
   and MGM_G89(MGM_W69,d_delay,MGM_W68);
   and MGM_G90(MGM_W70,si_delay,MGM_W69);
   not MGM_G91(MGM_W71,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W71,MGM_W70);
   not MGM_G93(MGM_W72,clk_delay);
   and MGM_G94(MGM_W73,d_delay,MGM_W72);
   and MGM_G95(MGM_W74,si_delay,MGM_W73);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W74);
   not MGM_G97(MGM_W75,d_delay);
   and MGM_G98(MGM_W76,MGM_W75,clk_delay);
   not MGM_G99(MGM_W77,si_delay);
   and MGM_G100(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G101(MGM_W79,ssb_delay);
   and MGM_G102(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G103(MGM_W80,d_delay);
   and MGM_G104(MGM_W81,MGM_W80,clk_delay);
   not MGM_G105(MGM_W82,si_delay);
   and MGM_G106(MGM_W83,MGM_W82,MGM_W81);
   and MGM_G107(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W83);
   not MGM_G108(MGM_W84,d_delay);
   and MGM_G109(MGM_W85,MGM_W84,clk_delay);
   and MGM_G110(MGM_W86,si_delay,MGM_W85);
   not MGM_G111(MGM_W87,ssb_delay);
   and MGM_G112(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W87,MGM_W86);
   not MGM_G113(MGM_W88,d_delay);
   and MGM_G114(MGM_W89,MGM_W88,clk_delay);
   and MGM_G115(MGM_W90,si_delay,MGM_W89);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W90);
   and MGM_G117(MGM_W91,d_delay,clk_delay);
   not MGM_G118(MGM_W92,si_delay);
   and MGM_G119(MGM_W93,MGM_W92,MGM_W91);
   not MGM_G120(MGM_W94,ssb_delay);
   and MGM_G121(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W94,MGM_W93);
   and MGM_G122(MGM_W95,d_delay,clk_delay);
   not MGM_G123(MGM_W96,si_delay);
   and MGM_G124(MGM_W97,MGM_W96,MGM_W95);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W97);
   and MGM_G126(MGM_W98,d_delay,clk_delay);
   and MGM_G127(MGM_W99,si_delay,MGM_W98);
   not MGM_G128(MGM_W100,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W100,MGM_W99);
   and MGM_G130(MGM_W101,d_delay,clk_delay);
   and MGM_G131(MGM_W102,si_delay,MGM_W101);
   and MGM_G132(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W102);
   not MGM_G133(MGM_W103,d_delay);
   and MGM_G134(MGM_W104,rb_delay,MGM_W103);
   not MGM_G135(MGM_W105,ssb_delay);
   and MGM_G136(ENABLE_NOT_d_AND_rb_AND_NOT_ssb,MGM_W105,MGM_W104);
   and MGM_G137(MGM_W106,rb_delay,d_delay);
   not MGM_G138(MGM_W107,ssb_delay);
   and MGM_G139(ENABLE_d_AND_rb_AND_NOT_ssb,MGM_W107,MGM_W106);
   not MGM_G140(MGM_W108,d_delay);
   and MGM_G141(MGM_W109,rb_delay,MGM_W108);
   and MGM_G142(ENABLE_NOT_d_AND_rb_AND_si,si_delay,MGM_W109);
   and MGM_G143(MGM_W110,rb_delay,d_delay);
   not MGM_G144(MGM_W111,si_delay);
   and MGM_G145(ENABLE_d_AND_rb_AND_NOT_si,MGM_W111,MGM_W110);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy003ah1n06x5( clk, d, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy003ah_func b15fqy003ah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy003ah_func b15fqy003ah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy003ah_func b15fqy003ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy003ah_func b15fqy003ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,rb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,rb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,rb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,rb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,rb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,rb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,rb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,rb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,rb_delay);
   and MGM_G38(ENABLE_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,rb_delay);
   and MGM_G40(ENABLE_rb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   and MGM_G42(MGM_W32,si_delay,MGM_W31);
   not MGM_G43(MGM_W33,ssb_delay);
   and MGM_G44(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W33,MGM_W32);
   not MGM_G45(MGM_W34,si_delay);
   and MGM_G46(MGM_W35,MGM_W34,d_delay);
   and MGM_G47(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G48(MGM_W36,si_delay,d_delay);
   not MGM_G49(MGM_W37,ssb_delay);
   and MGM_G50(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W37,MGM_W36);
   and MGM_G51(MGM_W38,si_delay,d_delay);
   and MGM_G52(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W38);
   not MGM_G53(MGM_W39,clk_delay);
   not MGM_G54(MGM_W40,d_delay);
   and MGM_G55(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G56(MGM_W42,si_delay);
   and MGM_G57(MGM_W43,MGM_W42,MGM_W41);
   not MGM_G58(MGM_W44,ssb_delay);
   and MGM_G59(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W45,clk_delay);
   not MGM_G61(MGM_W46,d_delay);
   and MGM_G62(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G63(MGM_W48,si_delay);
   and MGM_G64(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G65(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G66(MGM_W50,clk_delay);
   not MGM_G67(MGM_W51,d_delay);
   and MGM_G68(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G69(MGM_W53,si_delay,MGM_W52);
   not MGM_G70(MGM_W54,ssb_delay);
   and MGM_G71(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W54,MGM_W53);
   not MGM_G72(MGM_W55,clk_delay);
   not MGM_G73(MGM_W56,d_delay);
   and MGM_G74(MGM_W57,MGM_W56,MGM_W55);
   and MGM_G75(MGM_W58,si_delay,MGM_W57);
   and MGM_G76(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,clk_delay);
   and MGM_G78(MGM_W60,d_delay,MGM_W59);
   not MGM_G79(MGM_W61,si_delay);
   and MGM_G80(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G81(MGM_W63,ssb_delay);
   and MGM_G82(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G83(MGM_W64,clk_delay);
   and MGM_G84(MGM_W65,d_delay,MGM_W64);
   not MGM_G85(MGM_W66,si_delay);
   and MGM_G86(MGM_W67,MGM_W66,MGM_W65);
   and MGM_G87(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W67);
   not MGM_G88(MGM_W68,clk_delay);
   and MGM_G89(MGM_W69,d_delay,MGM_W68);
   and MGM_G90(MGM_W70,si_delay,MGM_W69);
   not MGM_G91(MGM_W71,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W71,MGM_W70);
   not MGM_G93(MGM_W72,clk_delay);
   and MGM_G94(MGM_W73,d_delay,MGM_W72);
   and MGM_G95(MGM_W74,si_delay,MGM_W73);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W74);
   not MGM_G97(MGM_W75,d_delay);
   and MGM_G98(MGM_W76,MGM_W75,clk_delay);
   not MGM_G99(MGM_W77,si_delay);
   and MGM_G100(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G101(MGM_W79,ssb_delay);
   and MGM_G102(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G103(MGM_W80,d_delay);
   and MGM_G104(MGM_W81,MGM_W80,clk_delay);
   not MGM_G105(MGM_W82,si_delay);
   and MGM_G106(MGM_W83,MGM_W82,MGM_W81);
   and MGM_G107(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W83);
   not MGM_G108(MGM_W84,d_delay);
   and MGM_G109(MGM_W85,MGM_W84,clk_delay);
   and MGM_G110(MGM_W86,si_delay,MGM_W85);
   not MGM_G111(MGM_W87,ssb_delay);
   and MGM_G112(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W87,MGM_W86);
   not MGM_G113(MGM_W88,d_delay);
   and MGM_G114(MGM_W89,MGM_W88,clk_delay);
   and MGM_G115(MGM_W90,si_delay,MGM_W89);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W90);
   and MGM_G117(MGM_W91,d_delay,clk_delay);
   not MGM_G118(MGM_W92,si_delay);
   and MGM_G119(MGM_W93,MGM_W92,MGM_W91);
   not MGM_G120(MGM_W94,ssb_delay);
   and MGM_G121(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W94,MGM_W93);
   and MGM_G122(MGM_W95,d_delay,clk_delay);
   not MGM_G123(MGM_W96,si_delay);
   and MGM_G124(MGM_W97,MGM_W96,MGM_W95);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W97);
   and MGM_G126(MGM_W98,d_delay,clk_delay);
   and MGM_G127(MGM_W99,si_delay,MGM_W98);
   not MGM_G128(MGM_W100,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W100,MGM_W99);
   and MGM_G130(MGM_W101,d_delay,clk_delay);
   and MGM_G131(MGM_W102,si_delay,MGM_W101);
   and MGM_G132(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W102);
   not MGM_G133(MGM_W103,d_delay);
   and MGM_G134(MGM_W104,rb_delay,MGM_W103);
   not MGM_G135(MGM_W105,ssb_delay);
   and MGM_G136(ENABLE_NOT_d_AND_rb_AND_NOT_ssb,MGM_W105,MGM_W104);
   and MGM_G137(MGM_W106,rb_delay,d_delay);
   not MGM_G138(MGM_W107,ssb_delay);
   and MGM_G139(ENABLE_d_AND_rb_AND_NOT_ssb,MGM_W107,MGM_W106);
   not MGM_G140(MGM_W108,d_delay);
   and MGM_G141(MGM_W109,rb_delay,MGM_W108);
   and MGM_G142(ENABLE_NOT_d_AND_rb_AND_si,si_delay,MGM_W109);
   and MGM_G143(MGM_W110,rb_delay,d_delay);
   not MGM_G144(MGM_W111,si_delay);
   and MGM_G145(ENABLE_d_AND_rb_AND_NOT_si,MGM_W111,MGM_W110);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy003ah1n08x5( clk, d, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy003ah_func b15fqy003ah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy003ah_func b15fqy003ah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy003ah_func b15fqy003ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy003ah_func b15fqy003ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,rb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,rb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,rb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,rb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,rb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,rb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,rb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,rb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,rb_delay);
   and MGM_G38(ENABLE_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,rb_delay);
   and MGM_G40(ENABLE_rb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   and MGM_G42(MGM_W32,si_delay,MGM_W31);
   not MGM_G43(MGM_W33,ssb_delay);
   and MGM_G44(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W33,MGM_W32);
   not MGM_G45(MGM_W34,si_delay);
   and MGM_G46(MGM_W35,MGM_W34,d_delay);
   and MGM_G47(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G48(MGM_W36,si_delay,d_delay);
   not MGM_G49(MGM_W37,ssb_delay);
   and MGM_G50(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W37,MGM_W36);
   and MGM_G51(MGM_W38,si_delay,d_delay);
   and MGM_G52(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W38);
   not MGM_G53(MGM_W39,clk_delay);
   not MGM_G54(MGM_W40,d_delay);
   and MGM_G55(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G56(MGM_W42,si_delay);
   and MGM_G57(MGM_W43,MGM_W42,MGM_W41);
   not MGM_G58(MGM_W44,ssb_delay);
   and MGM_G59(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W45,clk_delay);
   not MGM_G61(MGM_W46,d_delay);
   and MGM_G62(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G63(MGM_W48,si_delay);
   and MGM_G64(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G65(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G66(MGM_W50,clk_delay);
   not MGM_G67(MGM_W51,d_delay);
   and MGM_G68(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G69(MGM_W53,si_delay,MGM_W52);
   not MGM_G70(MGM_W54,ssb_delay);
   and MGM_G71(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W54,MGM_W53);
   not MGM_G72(MGM_W55,clk_delay);
   not MGM_G73(MGM_W56,d_delay);
   and MGM_G74(MGM_W57,MGM_W56,MGM_W55);
   and MGM_G75(MGM_W58,si_delay,MGM_W57);
   and MGM_G76(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,clk_delay);
   and MGM_G78(MGM_W60,d_delay,MGM_W59);
   not MGM_G79(MGM_W61,si_delay);
   and MGM_G80(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G81(MGM_W63,ssb_delay);
   and MGM_G82(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G83(MGM_W64,clk_delay);
   and MGM_G84(MGM_W65,d_delay,MGM_W64);
   not MGM_G85(MGM_W66,si_delay);
   and MGM_G86(MGM_W67,MGM_W66,MGM_W65);
   and MGM_G87(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W67);
   not MGM_G88(MGM_W68,clk_delay);
   and MGM_G89(MGM_W69,d_delay,MGM_W68);
   and MGM_G90(MGM_W70,si_delay,MGM_W69);
   not MGM_G91(MGM_W71,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W71,MGM_W70);
   not MGM_G93(MGM_W72,clk_delay);
   and MGM_G94(MGM_W73,d_delay,MGM_W72);
   and MGM_G95(MGM_W74,si_delay,MGM_W73);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W74);
   not MGM_G97(MGM_W75,d_delay);
   and MGM_G98(MGM_W76,MGM_W75,clk_delay);
   not MGM_G99(MGM_W77,si_delay);
   and MGM_G100(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G101(MGM_W79,ssb_delay);
   and MGM_G102(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G103(MGM_W80,d_delay);
   and MGM_G104(MGM_W81,MGM_W80,clk_delay);
   not MGM_G105(MGM_W82,si_delay);
   and MGM_G106(MGM_W83,MGM_W82,MGM_W81);
   and MGM_G107(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W83);
   not MGM_G108(MGM_W84,d_delay);
   and MGM_G109(MGM_W85,MGM_W84,clk_delay);
   and MGM_G110(MGM_W86,si_delay,MGM_W85);
   not MGM_G111(MGM_W87,ssb_delay);
   and MGM_G112(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W87,MGM_W86);
   not MGM_G113(MGM_W88,d_delay);
   and MGM_G114(MGM_W89,MGM_W88,clk_delay);
   and MGM_G115(MGM_W90,si_delay,MGM_W89);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W90);
   and MGM_G117(MGM_W91,d_delay,clk_delay);
   not MGM_G118(MGM_W92,si_delay);
   and MGM_G119(MGM_W93,MGM_W92,MGM_W91);
   not MGM_G120(MGM_W94,ssb_delay);
   and MGM_G121(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W94,MGM_W93);
   and MGM_G122(MGM_W95,d_delay,clk_delay);
   not MGM_G123(MGM_W96,si_delay);
   and MGM_G124(MGM_W97,MGM_W96,MGM_W95);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W97);
   and MGM_G126(MGM_W98,d_delay,clk_delay);
   and MGM_G127(MGM_W99,si_delay,MGM_W98);
   not MGM_G128(MGM_W100,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W100,MGM_W99);
   and MGM_G130(MGM_W101,d_delay,clk_delay);
   and MGM_G131(MGM_W102,si_delay,MGM_W101);
   and MGM_G132(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W102);
   not MGM_G133(MGM_W103,d_delay);
   and MGM_G134(MGM_W104,rb_delay,MGM_W103);
   not MGM_G135(MGM_W105,ssb_delay);
   and MGM_G136(ENABLE_NOT_d_AND_rb_AND_NOT_ssb,MGM_W105,MGM_W104);
   and MGM_G137(MGM_W106,rb_delay,d_delay);
   not MGM_G138(MGM_W107,ssb_delay);
   and MGM_G139(ENABLE_d_AND_rb_AND_NOT_ssb,MGM_W107,MGM_W106);
   not MGM_G140(MGM_W108,d_delay);
   and MGM_G141(MGM_W109,rb_delay,MGM_W108);
   and MGM_G142(ENABLE_NOT_d_AND_rb_AND_si,si_delay,MGM_W109);
   and MGM_G143(MGM_W110,rb_delay,d_delay);
   not MGM_G144(MGM_W111,si_delay);
   and MGM_G145(ENABLE_d_AND_rb_AND_NOT_si,MGM_W111,MGM_W110);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy003ah1n12x5( clk, d, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy003ah_func b15fqy003ah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy003ah_func b15fqy003ah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy003ah_func b15fqy003ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy003ah_func b15fqy003ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,rb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,rb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,rb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,rb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,rb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,rb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,rb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,rb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,rb_delay);
   and MGM_G38(ENABLE_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,rb_delay);
   and MGM_G40(ENABLE_rb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   and MGM_G42(MGM_W32,si_delay,MGM_W31);
   not MGM_G43(MGM_W33,ssb_delay);
   and MGM_G44(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W33,MGM_W32);
   not MGM_G45(MGM_W34,si_delay);
   and MGM_G46(MGM_W35,MGM_W34,d_delay);
   and MGM_G47(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G48(MGM_W36,si_delay,d_delay);
   not MGM_G49(MGM_W37,ssb_delay);
   and MGM_G50(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W37,MGM_W36);
   and MGM_G51(MGM_W38,si_delay,d_delay);
   and MGM_G52(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W38);
   not MGM_G53(MGM_W39,clk_delay);
   not MGM_G54(MGM_W40,d_delay);
   and MGM_G55(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G56(MGM_W42,si_delay);
   and MGM_G57(MGM_W43,MGM_W42,MGM_W41);
   not MGM_G58(MGM_W44,ssb_delay);
   and MGM_G59(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W45,clk_delay);
   not MGM_G61(MGM_W46,d_delay);
   and MGM_G62(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G63(MGM_W48,si_delay);
   and MGM_G64(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G65(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G66(MGM_W50,clk_delay);
   not MGM_G67(MGM_W51,d_delay);
   and MGM_G68(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G69(MGM_W53,si_delay,MGM_W52);
   not MGM_G70(MGM_W54,ssb_delay);
   and MGM_G71(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W54,MGM_W53);
   not MGM_G72(MGM_W55,clk_delay);
   not MGM_G73(MGM_W56,d_delay);
   and MGM_G74(MGM_W57,MGM_W56,MGM_W55);
   and MGM_G75(MGM_W58,si_delay,MGM_W57);
   and MGM_G76(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,clk_delay);
   and MGM_G78(MGM_W60,d_delay,MGM_W59);
   not MGM_G79(MGM_W61,si_delay);
   and MGM_G80(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G81(MGM_W63,ssb_delay);
   and MGM_G82(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G83(MGM_W64,clk_delay);
   and MGM_G84(MGM_W65,d_delay,MGM_W64);
   not MGM_G85(MGM_W66,si_delay);
   and MGM_G86(MGM_W67,MGM_W66,MGM_W65);
   and MGM_G87(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W67);
   not MGM_G88(MGM_W68,clk_delay);
   and MGM_G89(MGM_W69,d_delay,MGM_W68);
   and MGM_G90(MGM_W70,si_delay,MGM_W69);
   not MGM_G91(MGM_W71,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W71,MGM_W70);
   not MGM_G93(MGM_W72,clk_delay);
   and MGM_G94(MGM_W73,d_delay,MGM_W72);
   and MGM_G95(MGM_W74,si_delay,MGM_W73);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W74);
   not MGM_G97(MGM_W75,d_delay);
   and MGM_G98(MGM_W76,MGM_W75,clk_delay);
   not MGM_G99(MGM_W77,si_delay);
   and MGM_G100(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G101(MGM_W79,ssb_delay);
   and MGM_G102(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G103(MGM_W80,d_delay);
   and MGM_G104(MGM_W81,MGM_W80,clk_delay);
   not MGM_G105(MGM_W82,si_delay);
   and MGM_G106(MGM_W83,MGM_W82,MGM_W81);
   and MGM_G107(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W83);
   not MGM_G108(MGM_W84,d_delay);
   and MGM_G109(MGM_W85,MGM_W84,clk_delay);
   and MGM_G110(MGM_W86,si_delay,MGM_W85);
   not MGM_G111(MGM_W87,ssb_delay);
   and MGM_G112(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W87,MGM_W86);
   not MGM_G113(MGM_W88,d_delay);
   and MGM_G114(MGM_W89,MGM_W88,clk_delay);
   and MGM_G115(MGM_W90,si_delay,MGM_W89);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W90);
   and MGM_G117(MGM_W91,d_delay,clk_delay);
   not MGM_G118(MGM_W92,si_delay);
   and MGM_G119(MGM_W93,MGM_W92,MGM_W91);
   not MGM_G120(MGM_W94,ssb_delay);
   and MGM_G121(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W94,MGM_W93);
   and MGM_G122(MGM_W95,d_delay,clk_delay);
   not MGM_G123(MGM_W96,si_delay);
   and MGM_G124(MGM_W97,MGM_W96,MGM_W95);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W97);
   and MGM_G126(MGM_W98,d_delay,clk_delay);
   and MGM_G127(MGM_W99,si_delay,MGM_W98);
   not MGM_G128(MGM_W100,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W100,MGM_W99);
   and MGM_G130(MGM_W101,d_delay,clk_delay);
   and MGM_G131(MGM_W102,si_delay,MGM_W101);
   and MGM_G132(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W102);
   not MGM_G133(MGM_W103,d_delay);
   and MGM_G134(MGM_W104,rb_delay,MGM_W103);
   not MGM_G135(MGM_W105,ssb_delay);
   and MGM_G136(ENABLE_NOT_d_AND_rb_AND_NOT_ssb,MGM_W105,MGM_W104);
   and MGM_G137(MGM_W106,rb_delay,d_delay);
   not MGM_G138(MGM_W107,ssb_delay);
   and MGM_G139(ENABLE_d_AND_rb_AND_NOT_ssb,MGM_W107,MGM_W106);
   not MGM_G140(MGM_W108,d_delay);
   and MGM_G141(MGM_W109,rb_delay,MGM_W108);
   and MGM_G142(ENABLE_NOT_d_AND_rb_AND_si,si_delay,MGM_W109);
   and MGM_G143(MGM_W110,rb_delay,d_delay);
   not MGM_G144(MGM_W111,si_delay);
   and MGM_G145(ENABLE_d_AND_rb_AND_NOT_si,MGM_W111,MGM_W110);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy003ah1n16x5( clk, d, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy003ah_func b15fqy003ah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy003ah_func b15fqy003ah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy003ah_func b15fqy003ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy003ah_func b15fqy003ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,rb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,rb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,rb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,rb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,rb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,rb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,rb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,rb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,rb_delay);
   and MGM_G38(ENABLE_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,rb_delay);
   and MGM_G40(ENABLE_rb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   and MGM_G42(MGM_W32,si_delay,MGM_W31);
   not MGM_G43(MGM_W33,ssb_delay);
   and MGM_G44(ENABLE_NOT_d_AND_si_AND_NOT_ssb,MGM_W33,MGM_W32);
   not MGM_G45(MGM_W34,si_delay);
   and MGM_G46(MGM_W35,MGM_W34,d_delay);
   and MGM_G47(ENABLE_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G48(MGM_W36,si_delay,d_delay);
   not MGM_G49(MGM_W37,ssb_delay);
   and MGM_G50(ENABLE_d_AND_si_AND_NOT_ssb,MGM_W37,MGM_W36);
   and MGM_G51(MGM_W38,si_delay,d_delay);
   and MGM_G52(ENABLE_d_AND_si_AND_ssb,ssb_delay,MGM_W38);
   not MGM_G53(MGM_W39,clk_delay);
   not MGM_G54(MGM_W40,d_delay);
   and MGM_G55(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G56(MGM_W42,si_delay);
   and MGM_G57(MGM_W43,MGM_W42,MGM_W41);
   not MGM_G58(MGM_W44,ssb_delay);
   and MGM_G59(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W45,clk_delay);
   not MGM_G61(MGM_W46,d_delay);
   and MGM_G62(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G63(MGM_W48,si_delay);
   and MGM_G64(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G65(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G66(MGM_W50,clk_delay);
   not MGM_G67(MGM_W51,d_delay);
   and MGM_G68(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G69(MGM_W53,si_delay,MGM_W52);
   not MGM_G70(MGM_W54,ssb_delay);
   and MGM_G71(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W54,MGM_W53);
   not MGM_G72(MGM_W55,clk_delay);
   not MGM_G73(MGM_W56,d_delay);
   and MGM_G74(MGM_W57,MGM_W56,MGM_W55);
   and MGM_G75(MGM_W58,si_delay,MGM_W57);
   and MGM_G76(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W58);
   not MGM_G77(MGM_W59,clk_delay);
   and MGM_G78(MGM_W60,d_delay,MGM_W59);
   not MGM_G79(MGM_W61,si_delay);
   and MGM_G80(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G81(MGM_W63,ssb_delay);
   and MGM_G82(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G83(MGM_W64,clk_delay);
   and MGM_G84(MGM_W65,d_delay,MGM_W64);
   not MGM_G85(MGM_W66,si_delay);
   and MGM_G86(MGM_W67,MGM_W66,MGM_W65);
   and MGM_G87(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W67);
   not MGM_G88(MGM_W68,clk_delay);
   and MGM_G89(MGM_W69,d_delay,MGM_W68);
   and MGM_G90(MGM_W70,si_delay,MGM_W69);
   not MGM_G91(MGM_W71,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W71,MGM_W70);
   not MGM_G93(MGM_W72,clk_delay);
   and MGM_G94(MGM_W73,d_delay,MGM_W72);
   and MGM_G95(MGM_W74,si_delay,MGM_W73);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W74);
   not MGM_G97(MGM_W75,d_delay);
   and MGM_G98(MGM_W76,MGM_W75,clk_delay);
   not MGM_G99(MGM_W77,si_delay);
   and MGM_G100(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G101(MGM_W79,ssb_delay);
   and MGM_G102(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G103(MGM_W80,d_delay);
   and MGM_G104(MGM_W81,MGM_W80,clk_delay);
   not MGM_G105(MGM_W82,si_delay);
   and MGM_G106(MGM_W83,MGM_W82,MGM_W81);
   and MGM_G107(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W83);
   not MGM_G108(MGM_W84,d_delay);
   and MGM_G109(MGM_W85,MGM_W84,clk_delay);
   and MGM_G110(MGM_W86,si_delay,MGM_W85);
   not MGM_G111(MGM_W87,ssb_delay);
   and MGM_G112(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W87,MGM_W86);
   not MGM_G113(MGM_W88,d_delay);
   and MGM_G114(MGM_W89,MGM_W88,clk_delay);
   and MGM_G115(MGM_W90,si_delay,MGM_W89);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W90);
   and MGM_G117(MGM_W91,d_delay,clk_delay);
   not MGM_G118(MGM_W92,si_delay);
   and MGM_G119(MGM_W93,MGM_W92,MGM_W91);
   not MGM_G120(MGM_W94,ssb_delay);
   and MGM_G121(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W94,MGM_W93);
   and MGM_G122(MGM_W95,d_delay,clk_delay);
   not MGM_G123(MGM_W96,si_delay);
   and MGM_G124(MGM_W97,MGM_W96,MGM_W95);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W97);
   and MGM_G126(MGM_W98,d_delay,clk_delay);
   and MGM_G127(MGM_W99,si_delay,MGM_W98);
   not MGM_G128(MGM_W100,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W100,MGM_W99);
   and MGM_G130(MGM_W101,d_delay,clk_delay);
   and MGM_G131(MGM_W102,si_delay,MGM_W101);
   and MGM_G132(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W102);
   not MGM_G133(MGM_W103,d_delay);
   and MGM_G134(MGM_W104,rb_delay,MGM_W103);
   not MGM_G135(MGM_W105,ssb_delay);
   and MGM_G136(ENABLE_NOT_d_AND_rb_AND_NOT_ssb,MGM_W105,MGM_W104);
   and MGM_G137(MGM_W106,rb_delay,d_delay);
   not MGM_G138(MGM_W107,ssb_delay);
   and MGM_G139(ENABLE_d_AND_rb_AND_NOT_ssb,MGM_W107,MGM_W106);
   not MGM_G140(MGM_W108,d_delay);
   and MGM_G141(MGM_W109,rb_delay,MGM_W108);
   and MGM_G142(ENABLE_NOT_d_AND_rb_AND_si,si_delay,MGM_W109);
   and MGM_G143(MGM_W110,rb_delay,d_delay);
   not MGM_G144(MGM_W111,si_delay);
   and MGM_G145(ENABLE_d_AND_rb_AND_NOT_si,MGM_W111,MGM_W110);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fqy00cah_func( clk, d, o, psb, si, ssb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, si, ssb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_P0, psb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, MGM_P0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_P0, psb );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, 1'b0, MGM_P0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fqy00cah1n02x5( clk, d, o, psb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00cah_func b15fqy00cah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00cah_func b15fqy00cah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00cah_func b15fqy00cah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00cah_func b15fqy00cah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,psb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,psb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,psb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,psb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,psb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,psb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,psb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,psb_delay);
   and MGM_G38(ENABLE_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,psb_delay);
   and MGM_G40(ENABLE_psb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   not MGM_G42(MGM_W32,si_delay);
   and MGM_G43(MGM_W33,MGM_W32,MGM_W31);
   not MGM_G44(MGM_W34,ssb_delay);
   and MGM_G45(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W34,MGM_W33);
   not MGM_G46(MGM_W35,d_delay);
   not MGM_G47(MGM_W36,si_delay);
   and MGM_G48(MGM_W37,MGM_W36,MGM_W35);
   and MGM_G49(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W37);
   not MGM_G50(MGM_W38,d_delay);
   and MGM_G51(MGM_W39,si_delay,MGM_W38);
   and MGM_G52(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W39);
   not MGM_G53(MGM_W40,si_delay);
   and MGM_G54(MGM_W41,MGM_W40,d_delay);
   not MGM_G55(MGM_W42,ssb_delay);
   and MGM_G56(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W42,MGM_W41);
   not MGM_G57(MGM_W43,clk_delay);
   not MGM_G58(MGM_W44,d_delay);
   and MGM_G59(MGM_W45,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W46,si_delay);
   and MGM_G61(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G62(MGM_W48,ssb_delay);
   and MGM_G63(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   not MGM_G64(MGM_W49,clk_delay);
   not MGM_G65(MGM_W50,d_delay);
   and MGM_G66(MGM_W51,MGM_W50,MGM_W49);
   not MGM_G67(MGM_W52,si_delay);
   and MGM_G68(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G69(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G70(MGM_W54,clk_delay);
   not MGM_G71(MGM_W55,d_delay);
   and MGM_G72(MGM_W56,MGM_W55,MGM_W54);
   and MGM_G73(MGM_W57,si_delay,MGM_W56);
   not MGM_G74(MGM_W58,ssb_delay);
   and MGM_G75(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W58,MGM_W57);
   not MGM_G76(MGM_W59,clk_delay);
   not MGM_G77(MGM_W60,d_delay);
   and MGM_G78(MGM_W61,MGM_W60,MGM_W59);
   and MGM_G79(MGM_W62,si_delay,MGM_W61);
   and MGM_G80(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W62);
   not MGM_G81(MGM_W63,clk_delay);
   and MGM_G82(MGM_W64,d_delay,MGM_W63);
   not MGM_G83(MGM_W65,si_delay);
   and MGM_G84(MGM_W66,MGM_W65,MGM_W64);
   not MGM_G85(MGM_W67,ssb_delay);
   and MGM_G86(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W67,MGM_W66);
   not MGM_G87(MGM_W68,clk_delay);
   and MGM_G88(MGM_W69,d_delay,MGM_W68);
   not MGM_G89(MGM_W70,si_delay);
   and MGM_G90(MGM_W71,MGM_W70,MGM_W69);
   and MGM_G91(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W71);
   not MGM_G92(MGM_W72,clk_delay);
   and MGM_G93(MGM_W73,d_delay,MGM_W72);
   and MGM_G94(MGM_W74,si_delay,MGM_W73);
   not MGM_G95(MGM_W75,ssb_delay);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G97(MGM_W76,clk_delay);
   and MGM_G98(MGM_W77,d_delay,MGM_W76);
   and MGM_G99(MGM_W78,si_delay,MGM_W77);
   and MGM_G100(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W78);
   not MGM_G101(MGM_W79,d_delay);
   and MGM_G102(MGM_W80,MGM_W79,clk_delay);
   not MGM_G103(MGM_W81,si_delay);
   and MGM_G104(MGM_W82,MGM_W81,MGM_W80);
   not MGM_G105(MGM_W83,ssb_delay);
   and MGM_G106(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W83,MGM_W82);
   not MGM_G107(MGM_W84,d_delay);
   and MGM_G108(MGM_W85,MGM_W84,clk_delay);
   not MGM_G109(MGM_W86,si_delay);
   and MGM_G110(MGM_W87,MGM_W86,MGM_W85);
   and MGM_G111(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W87);
   not MGM_G112(MGM_W88,d_delay);
   and MGM_G113(MGM_W89,MGM_W88,clk_delay);
   and MGM_G114(MGM_W90,si_delay,MGM_W89);
   not MGM_G115(MGM_W91,ssb_delay);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W91,MGM_W90);
   not MGM_G117(MGM_W92,d_delay);
   and MGM_G118(MGM_W93,MGM_W92,clk_delay);
   and MGM_G119(MGM_W94,si_delay,MGM_W93);
   and MGM_G120(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W94);
   and MGM_G121(MGM_W95,d_delay,clk_delay);
   not MGM_G122(MGM_W96,si_delay);
   and MGM_G123(MGM_W97,MGM_W96,MGM_W95);
   not MGM_G124(MGM_W98,ssb_delay);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W98,MGM_W97);
   and MGM_G126(MGM_W99,d_delay,clk_delay);
   not MGM_G127(MGM_W100,si_delay);
   and MGM_G128(MGM_W101,MGM_W100,MGM_W99);
   and MGM_G129(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W101);
   and MGM_G130(MGM_W102,d_delay,clk_delay);
   and MGM_G131(MGM_W103,si_delay,MGM_W102);
   not MGM_G132(MGM_W104,ssb_delay);
   and MGM_G133(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W104,MGM_W103);
   and MGM_G134(MGM_W105,d_delay,clk_delay);
   and MGM_G135(MGM_W106,si_delay,MGM_W105);
   and MGM_G136(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W106);
   not MGM_G137(MGM_W107,d_delay);
   and MGM_G138(MGM_W108,psb_delay,MGM_W107);
   not MGM_G139(MGM_W109,ssb_delay);
   and MGM_G140(ENABLE_NOT_d_AND_psb_AND_NOT_ssb,MGM_W109,MGM_W108);
   and MGM_G141(MGM_W110,psb_delay,d_delay);
   not MGM_G142(MGM_W111,ssb_delay);
   and MGM_G143(ENABLE_d_AND_psb_AND_NOT_ssb,MGM_W111,MGM_W110);
   not MGM_G144(MGM_W112,d_delay);
   and MGM_G145(MGM_W113,psb_delay,MGM_W112);
   and MGM_G146(ENABLE_NOT_d_AND_psb_AND_si,si_delay,MGM_W113);
   and MGM_G147(MGM_W114,psb_delay,d_delay);
   not MGM_G148(MGM_W115,si_delay);
   and MGM_G149(ENABLE_d_AND_psb_AND_NOT_si,MGM_W115,MGM_W114);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy00cah1n03x5( clk, d, o, psb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00cah_func b15fqy00cah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00cah_func b15fqy00cah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00cah_func b15fqy00cah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00cah_func b15fqy00cah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,psb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,psb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,psb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,psb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,psb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,psb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,psb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,psb_delay);
   and MGM_G38(ENABLE_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,psb_delay);
   and MGM_G40(ENABLE_psb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   not MGM_G42(MGM_W32,si_delay);
   and MGM_G43(MGM_W33,MGM_W32,MGM_W31);
   not MGM_G44(MGM_W34,ssb_delay);
   and MGM_G45(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W34,MGM_W33);
   not MGM_G46(MGM_W35,d_delay);
   not MGM_G47(MGM_W36,si_delay);
   and MGM_G48(MGM_W37,MGM_W36,MGM_W35);
   and MGM_G49(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W37);
   not MGM_G50(MGM_W38,d_delay);
   and MGM_G51(MGM_W39,si_delay,MGM_W38);
   and MGM_G52(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W39);
   not MGM_G53(MGM_W40,si_delay);
   and MGM_G54(MGM_W41,MGM_W40,d_delay);
   not MGM_G55(MGM_W42,ssb_delay);
   and MGM_G56(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W42,MGM_W41);
   not MGM_G57(MGM_W43,clk_delay);
   not MGM_G58(MGM_W44,d_delay);
   and MGM_G59(MGM_W45,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W46,si_delay);
   and MGM_G61(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G62(MGM_W48,ssb_delay);
   and MGM_G63(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   not MGM_G64(MGM_W49,clk_delay);
   not MGM_G65(MGM_W50,d_delay);
   and MGM_G66(MGM_W51,MGM_W50,MGM_W49);
   not MGM_G67(MGM_W52,si_delay);
   and MGM_G68(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G69(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G70(MGM_W54,clk_delay);
   not MGM_G71(MGM_W55,d_delay);
   and MGM_G72(MGM_W56,MGM_W55,MGM_W54);
   and MGM_G73(MGM_W57,si_delay,MGM_W56);
   not MGM_G74(MGM_W58,ssb_delay);
   and MGM_G75(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W58,MGM_W57);
   not MGM_G76(MGM_W59,clk_delay);
   not MGM_G77(MGM_W60,d_delay);
   and MGM_G78(MGM_W61,MGM_W60,MGM_W59);
   and MGM_G79(MGM_W62,si_delay,MGM_W61);
   and MGM_G80(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W62);
   not MGM_G81(MGM_W63,clk_delay);
   and MGM_G82(MGM_W64,d_delay,MGM_W63);
   not MGM_G83(MGM_W65,si_delay);
   and MGM_G84(MGM_W66,MGM_W65,MGM_W64);
   not MGM_G85(MGM_W67,ssb_delay);
   and MGM_G86(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W67,MGM_W66);
   not MGM_G87(MGM_W68,clk_delay);
   and MGM_G88(MGM_W69,d_delay,MGM_W68);
   not MGM_G89(MGM_W70,si_delay);
   and MGM_G90(MGM_W71,MGM_W70,MGM_W69);
   and MGM_G91(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W71);
   not MGM_G92(MGM_W72,clk_delay);
   and MGM_G93(MGM_W73,d_delay,MGM_W72);
   and MGM_G94(MGM_W74,si_delay,MGM_W73);
   not MGM_G95(MGM_W75,ssb_delay);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G97(MGM_W76,clk_delay);
   and MGM_G98(MGM_W77,d_delay,MGM_W76);
   and MGM_G99(MGM_W78,si_delay,MGM_W77);
   and MGM_G100(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W78);
   not MGM_G101(MGM_W79,d_delay);
   and MGM_G102(MGM_W80,MGM_W79,clk_delay);
   not MGM_G103(MGM_W81,si_delay);
   and MGM_G104(MGM_W82,MGM_W81,MGM_W80);
   not MGM_G105(MGM_W83,ssb_delay);
   and MGM_G106(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W83,MGM_W82);
   not MGM_G107(MGM_W84,d_delay);
   and MGM_G108(MGM_W85,MGM_W84,clk_delay);
   not MGM_G109(MGM_W86,si_delay);
   and MGM_G110(MGM_W87,MGM_W86,MGM_W85);
   and MGM_G111(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W87);
   not MGM_G112(MGM_W88,d_delay);
   and MGM_G113(MGM_W89,MGM_W88,clk_delay);
   and MGM_G114(MGM_W90,si_delay,MGM_W89);
   not MGM_G115(MGM_W91,ssb_delay);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W91,MGM_W90);
   not MGM_G117(MGM_W92,d_delay);
   and MGM_G118(MGM_W93,MGM_W92,clk_delay);
   and MGM_G119(MGM_W94,si_delay,MGM_W93);
   and MGM_G120(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W94);
   and MGM_G121(MGM_W95,d_delay,clk_delay);
   not MGM_G122(MGM_W96,si_delay);
   and MGM_G123(MGM_W97,MGM_W96,MGM_W95);
   not MGM_G124(MGM_W98,ssb_delay);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W98,MGM_W97);
   and MGM_G126(MGM_W99,d_delay,clk_delay);
   not MGM_G127(MGM_W100,si_delay);
   and MGM_G128(MGM_W101,MGM_W100,MGM_W99);
   and MGM_G129(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W101);
   and MGM_G130(MGM_W102,d_delay,clk_delay);
   and MGM_G131(MGM_W103,si_delay,MGM_W102);
   not MGM_G132(MGM_W104,ssb_delay);
   and MGM_G133(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W104,MGM_W103);
   and MGM_G134(MGM_W105,d_delay,clk_delay);
   and MGM_G135(MGM_W106,si_delay,MGM_W105);
   and MGM_G136(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W106);
   not MGM_G137(MGM_W107,d_delay);
   and MGM_G138(MGM_W108,psb_delay,MGM_W107);
   not MGM_G139(MGM_W109,ssb_delay);
   and MGM_G140(ENABLE_NOT_d_AND_psb_AND_NOT_ssb,MGM_W109,MGM_W108);
   and MGM_G141(MGM_W110,psb_delay,d_delay);
   not MGM_G142(MGM_W111,ssb_delay);
   and MGM_G143(ENABLE_d_AND_psb_AND_NOT_ssb,MGM_W111,MGM_W110);
   not MGM_G144(MGM_W112,d_delay);
   and MGM_G145(MGM_W113,psb_delay,MGM_W112);
   and MGM_G146(ENABLE_NOT_d_AND_psb_AND_si,si_delay,MGM_W113);
   and MGM_G147(MGM_W114,psb_delay,d_delay);
   not MGM_G148(MGM_W115,si_delay);
   and MGM_G149(ENABLE_d_AND_psb_AND_NOT_si,MGM_W115,MGM_W114);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy00cah1n04x5( clk, d, o, psb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00cah_func b15fqy00cah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00cah_func b15fqy00cah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00cah_func b15fqy00cah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00cah_func b15fqy00cah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,psb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,psb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,psb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,psb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,psb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,psb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,psb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,psb_delay);
   and MGM_G38(ENABLE_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,psb_delay);
   and MGM_G40(ENABLE_psb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   not MGM_G42(MGM_W32,si_delay);
   and MGM_G43(MGM_W33,MGM_W32,MGM_W31);
   not MGM_G44(MGM_W34,ssb_delay);
   and MGM_G45(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W34,MGM_W33);
   not MGM_G46(MGM_W35,d_delay);
   not MGM_G47(MGM_W36,si_delay);
   and MGM_G48(MGM_W37,MGM_W36,MGM_W35);
   and MGM_G49(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W37);
   not MGM_G50(MGM_W38,d_delay);
   and MGM_G51(MGM_W39,si_delay,MGM_W38);
   and MGM_G52(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W39);
   not MGM_G53(MGM_W40,si_delay);
   and MGM_G54(MGM_W41,MGM_W40,d_delay);
   not MGM_G55(MGM_W42,ssb_delay);
   and MGM_G56(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W42,MGM_W41);
   not MGM_G57(MGM_W43,clk_delay);
   not MGM_G58(MGM_W44,d_delay);
   and MGM_G59(MGM_W45,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W46,si_delay);
   and MGM_G61(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G62(MGM_W48,ssb_delay);
   and MGM_G63(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   not MGM_G64(MGM_W49,clk_delay);
   not MGM_G65(MGM_W50,d_delay);
   and MGM_G66(MGM_W51,MGM_W50,MGM_W49);
   not MGM_G67(MGM_W52,si_delay);
   and MGM_G68(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G69(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G70(MGM_W54,clk_delay);
   not MGM_G71(MGM_W55,d_delay);
   and MGM_G72(MGM_W56,MGM_W55,MGM_W54);
   and MGM_G73(MGM_W57,si_delay,MGM_W56);
   not MGM_G74(MGM_W58,ssb_delay);
   and MGM_G75(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W58,MGM_W57);
   not MGM_G76(MGM_W59,clk_delay);
   not MGM_G77(MGM_W60,d_delay);
   and MGM_G78(MGM_W61,MGM_W60,MGM_W59);
   and MGM_G79(MGM_W62,si_delay,MGM_W61);
   and MGM_G80(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W62);
   not MGM_G81(MGM_W63,clk_delay);
   and MGM_G82(MGM_W64,d_delay,MGM_W63);
   not MGM_G83(MGM_W65,si_delay);
   and MGM_G84(MGM_W66,MGM_W65,MGM_W64);
   not MGM_G85(MGM_W67,ssb_delay);
   and MGM_G86(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W67,MGM_W66);
   not MGM_G87(MGM_W68,clk_delay);
   and MGM_G88(MGM_W69,d_delay,MGM_W68);
   not MGM_G89(MGM_W70,si_delay);
   and MGM_G90(MGM_W71,MGM_W70,MGM_W69);
   and MGM_G91(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W71);
   not MGM_G92(MGM_W72,clk_delay);
   and MGM_G93(MGM_W73,d_delay,MGM_W72);
   and MGM_G94(MGM_W74,si_delay,MGM_W73);
   not MGM_G95(MGM_W75,ssb_delay);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G97(MGM_W76,clk_delay);
   and MGM_G98(MGM_W77,d_delay,MGM_W76);
   and MGM_G99(MGM_W78,si_delay,MGM_W77);
   and MGM_G100(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W78);
   not MGM_G101(MGM_W79,d_delay);
   and MGM_G102(MGM_W80,MGM_W79,clk_delay);
   not MGM_G103(MGM_W81,si_delay);
   and MGM_G104(MGM_W82,MGM_W81,MGM_W80);
   not MGM_G105(MGM_W83,ssb_delay);
   and MGM_G106(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W83,MGM_W82);
   not MGM_G107(MGM_W84,d_delay);
   and MGM_G108(MGM_W85,MGM_W84,clk_delay);
   not MGM_G109(MGM_W86,si_delay);
   and MGM_G110(MGM_W87,MGM_W86,MGM_W85);
   and MGM_G111(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W87);
   not MGM_G112(MGM_W88,d_delay);
   and MGM_G113(MGM_W89,MGM_W88,clk_delay);
   and MGM_G114(MGM_W90,si_delay,MGM_W89);
   not MGM_G115(MGM_W91,ssb_delay);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W91,MGM_W90);
   not MGM_G117(MGM_W92,d_delay);
   and MGM_G118(MGM_W93,MGM_W92,clk_delay);
   and MGM_G119(MGM_W94,si_delay,MGM_W93);
   and MGM_G120(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W94);
   and MGM_G121(MGM_W95,d_delay,clk_delay);
   not MGM_G122(MGM_W96,si_delay);
   and MGM_G123(MGM_W97,MGM_W96,MGM_W95);
   not MGM_G124(MGM_W98,ssb_delay);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W98,MGM_W97);
   and MGM_G126(MGM_W99,d_delay,clk_delay);
   not MGM_G127(MGM_W100,si_delay);
   and MGM_G128(MGM_W101,MGM_W100,MGM_W99);
   and MGM_G129(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W101);
   and MGM_G130(MGM_W102,d_delay,clk_delay);
   and MGM_G131(MGM_W103,si_delay,MGM_W102);
   not MGM_G132(MGM_W104,ssb_delay);
   and MGM_G133(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W104,MGM_W103);
   and MGM_G134(MGM_W105,d_delay,clk_delay);
   and MGM_G135(MGM_W106,si_delay,MGM_W105);
   and MGM_G136(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W106);
   not MGM_G137(MGM_W107,d_delay);
   and MGM_G138(MGM_W108,psb_delay,MGM_W107);
   not MGM_G139(MGM_W109,ssb_delay);
   and MGM_G140(ENABLE_NOT_d_AND_psb_AND_NOT_ssb,MGM_W109,MGM_W108);
   and MGM_G141(MGM_W110,psb_delay,d_delay);
   not MGM_G142(MGM_W111,ssb_delay);
   and MGM_G143(ENABLE_d_AND_psb_AND_NOT_ssb,MGM_W111,MGM_W110);
   not MGM_G144(MGM_W112,d_delay);
   and MGM_G145(MGM_W113,psb_delay,MGM_W112);
   and MGM_G146(ENABLE_NOT_d_AND_psb_AND_si,si_delay,MGM_W113);
   and MGM_G147(MGM_W114,psb_delay,d_delay);
   not MGM_G148(MGM_W115,si_delay);
   and MGM_G149(ENABLE_d_AND_psb_AND_NOT_si,MGM_W115,MGM_W114);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy00cah1n06x5( clk, d, o, psb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00cah_func b15fqy00cah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00cah_func b15fqy00cah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00cah_func b15fqy00cah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00cah_func b15fqy00cah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,psb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,psb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,psb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,psb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,psb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,psb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,psb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,psb_delay);
   and MGM_G38(ENABLE_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,psb_delay);
   and MGM_G40(ENABLE_psb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   not MGM_G42(MGM_W32,si_delay);
   and MGM_G43(MGM_W33,MGM_W32,MGM_W31);
   not MGM_G44(MGM_W34,ssb_delay);
   and MGM_G45(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W34,MGM_W33);
   not MGM_G46(MGM_W35,d_delay);
   not MGM_G47(MGM_W36,si_delay);
   and MGM_G48(MGM_W37,MGM_W36,MGM_W35);
   and MGM_G49(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W37);
   not MGM_G50(MGM_W38,d_delay);
   and MGM_G51(MGM_W39,si_delay,MGM_W38);
   and MGM_G52(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W39);
   not MGM_G53(MGM_W40,si_delay);
   and MGM_G54(MGM_W41,MGM_W40,d_delay);
   not MGM_G55(MGM_W42,ssb_delay);
   and MGM_G56(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W42,MGM_W41);
   not MGM_G57(MGM_W43,clk_delay);
   not MGM_G58(MGM_W44,d_delay);
   and MGM_G59(MGM_W45,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W46,si_delay);
   and MGM_G61(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G62(MGM_W48,ssb_delay);
   and MGM_G63(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   not MGM_G64(MGM_W49,clk_delay);
   not MGM_G65(MGM_W50,d_delay);
   and MGM_G66(MGM_W51,MGM_W50,MGM_W49);
   not MGM_G67(MGM_W52,si_delay);
   and MGM_G68(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G69(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G70(MGM_W54,clk_delay);
   not MGM_G71(MGM_W55,d_delay);
   and MGM_G72(MGM_W56,MGM_W55,MGM_W54);
   and MGM_G73(MGM_W57,si_delay,MGM_W56);
   not MGM_G74(MGM_W58,ssb_delay);
   and MGM_G75(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W58,MGM_W57);
   not MGM_G76(MGM_W59,clk_delay);
   not MGM_G77(MGM_W60,d_delay);
   and MGM_G78(MGM_W61,MGM_W60,MGM_W59);
   and MGM_G79(MGM_W62,si_delay,MGM_W61);
   and MGM_G80(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W62);
   not MGM_G81(MGM_W63,clk_delay);
   and MGM_G82(MGM_W64,d_delay,MGM_W63);
   not MGM_G83(MGM_W65,si_delay);
   and MGM_G84(MGM_W66,MGM_W65,MGM_W64);
   not MGM_G85(MGM_W67,ssb_delay);
   and MGM_G86(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W67,MGM_W66);
   not MGM_G87(MGM_W68,clk_delay);
   and MGM_G88(MGM_W69,d_delay,MGM_W68);
   not MGM_G89(MGM_W70,si_delay);
   and MGM_G90(MGM_W71,MGM_W70,MGM_W69);
   and MGM_G91(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W71);
   not MGM_G92(MGM_W72,clk_delay);
   and MGM_G93(MGM_W73,d_delay,MGM_W72);
   and MGM_G94(MGM_W74,si_delay,MGM_W73);
   not MGM_G95(MGM_W75,ssb_delay);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G97(MGM_W76,clk_delay);
   and MGM_G98(MGM_W77,d_delay,MGM_W76);
   and MGM_G99(MGM_W78,si_delay,MGM_W77);
   and MGM_G100(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W78);
   not MGM_G101(MGM_W79,d_delay);
   and MGM_G102(MGM_W80,MGM_W79,clk_delay);
   not MGM_G103(MGM_W81,si_delay);
   and MGM_G104(MGM_W82,MGM_W81,MGM_W80);
   not MGM_G105(MGM_W83,ssb_delay);
   and MGM_G106(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W83,MGM_W82);
   not MGM_G107(MGM_W84,d_delay);
   and MGM_G108(MGM_W85,MGM_W84,clk_delay);
   not MGM_G109(MGM_W86,si_delay);
   and MGM_G110(MGM_W87,MGM_W86,MGM_W85);
   and MGM_G111(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W87);
   not MGM_G112(MGM_W88,d_delay);
   and MGM_G113(MGM_W89,MGM_W88,clk_delay);
   and MGM_G114(MGM_W90,si_delay,MGM_W89);
   not MGM_G115(MGM_W91,ssb_delay);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W91,MGM_W90);
   not MGM_G117(MGM_W92,d_delay);
   and MGM_G118(MGM_W93,MGM_W92,clk_delay);
   and MGM_G119(MGM_W94,si_delay,MGM_W93);
   and MGM_G120(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W94);
   and MGM_G121(MGM_W95,d_delay,clk_delay);
   not MGM_G122(MGM_W96,si_delay);
   and MGM_G123(MGM_W97,MGM_W96,MGM_W95);
   not MGM_G124(MGM_W98,ssb_delay);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W98,MGM_W97);
   and MGM_G126(MGM_W99,d_delay,clk_delay);
   not MGM_G127(MGM_W100,si_delay);
   and MGM_G128(MGM_W101,MGM_W100,MGM_W99);
   and MGM_G129(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W101);
   and MGM_G130(MGM_W102,d_delay,clk_delay);
   and MGM_G131(MGM_W103,si_delay,MGM_W102);
   not MGM_G132(MGM_W104,ssb_delay);
   and MGM_G133(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W104,MGM_W103);
   and MGM_G134(MGM_W105,d_delay,clk_delay);
   and MGM_G135(MGM_W106,si_delay,MGM_W105);
   and MGM_G136(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W106);
   not MGM_G137(MGM_W107,d_delay);
   and MGM_G138(MGM_W108,psb_delay,MGM_W107);
   not MGM_G139(MGM_W109,ssb_delay);
   and MGM_G140(ENABLE_NOT_d_AND_psb_AND_NOT_ssb,MGM_W109,MGM_W108);
   and MGM_G141(MGM_W110,psb_delay,d_delay);
   not MGM_G142(MGM_W111,ssb_delay);
   and MGM_G143(ENABLE_d_AND_psb_AND_NOT_ssb,MGM_W111,MGM_W110);
   not MGM_G144(MGM_W112,d_delay);
   and MGM_G145(MGM_W113,psb_delay,MGM_W112);
   and MGM_G146(ENABLE_NOT_d_AND_psb_AND_si,si_delay,MGM_W113);
   and MGM_G147(MGM_W114,psb_delay,d_delay);
   not MGM_G148(MGM_W115,si_delay);
   and MGM_G149(ENABLE_d_AND_psb_AND_NOT_si,MGM_W115,MGM_W114);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy00cah1n08x5( clk, d, o, psb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00cah_func b15fqy00cah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00cah_func b15fqy00cah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00cah_func b15fqy00cah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00cah_func b15fqy00cah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,psb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,psb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,psb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,psb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,psb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,psb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,psb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,psb_delay);
   and MGM_G38(ENABLE_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,psb_delay);
   and MGM_G40(ENABLE_psb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   not MGM_G42(MGM_W32,si_delay);
   and MGM_G43(MGM_W33,MGM_W32,MGM_W31);
   not MGM_G44(MGM_W34,ssb_delay);
   and MGM_G45(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W34,MGM_W33);
   not MGM_G46(MGM_W35,d_delay);
   not MGM_G47(MGM_W36,si_delay);
   and MGM_G48(MGM_W37,MGM_W36,MGM_W35);
   and MGM_G49(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W37);
   not MGM_G50(MGM_W38,d_delay);
   and MGM_G51(MGM_W39,si_delay,MGM_W38);
   and MGM_G52(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W39);
   not MGM_G53(MGM_W40,si_delay);
   and MGM_G54(MGM_W41,MGM_W40,d_delay);
   not MGM_G55(MGM_W42,ssb_delay);
   and MGM_G56(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W42,MGM_W41);
   not MGM_G57(MGM_W43,clk_delay);
   not MGM_G58(MGM_W44,d_delay);
   and MGM_G59(MGM_W45,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W46,si_delay);
   and MGM_G61(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G62(MGM_W48,ssb_delay);
   and MGM_G63(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   not MGM_G64(MGM_W49,clk_delay);
   not MGM_G65(MGM_W50,d_delay);
   and MGM_G66(MGM_W51,MGM_W50,MGM_W49);
   not MGM_G67(MGM_W52,si_delay);
   and MGM_G68(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G69(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G70(MGM_W54,clk_delay);
   not MGM_G71(MGM_W55,d_delay);
   and MGM_G72(MGM_W56,MGM_W55,MGM_W54);
   and MGM_G73(MGM_W57,si_delay,MGM_W56);
   not MGM_G74(MGM_W58,ssb_delay);
   and MGM_G75(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W58,MGM_W57);
   not MGM_G76(MGM_W59,clk_delay);
   not MGM_G77(MGM_W60,d_delay);
   and MGM_G78(MGM_W61,MGM_W60,MGM_W59);
   and MGM_G79(MGM_W62,si_delay,MGM_W61);
   and MGM_G80(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W62);
   not MGM_G81(MGM_W63,clk_delay);
   and MGM_G82(MGM_W64,d_delay,MGM_W63);
   not MGM_G83(MGM_W65,si_delay);
   and MGM_G84(MGM_W66,MGM_W65,MGM_W64);
   not MGM_G85(MGM_W67,ssb_delay);
   and MGM_G86(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W67,MGM_W66);
   not MGM_G87(MGM_W68,clk_delay);
   and MGM_G88(MGM_W69,d_delay,MGM_W68);
   not MGM_G89(MGM_W70,si_delay);
   and MGM_G90(MGM_W71,MGM_W70,MGM_W69);
   and MGM_G91(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W71);
   not MGM_G92(MGM_W72,clk_delay);
   and MGM_G93(MGM_W73,d_delay,MGM_W72);
   and MGM_G94(MGM_W74,si_delay,MGM_W73);
   not MGM_G95(MGM_W75,ssb_delay);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G97(MGM_W76,clk_delay);
   and MGM_G98(MGM_W77,d_delay,MGM_W76);
   and MGM_G99(MGM_W78,si_delay,MGM_W77);
   and MGM_G100(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W78);
   not MGM_G101(MGM_W79,d_delay);
   and MGM_G102(MGM_W80,MGM_W79,clk_delay);
   not MGM_G103(MGM_W81,si_delay);
   and MGM_G104(MGM_W82,MGM_W81,MGM_W80);
   not MGM_G105(MGM_W83,ssb_delay);
   and MGM_G106(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W83,MGM_W82);
   not MGM_G107(MGM_W84,d_delay);
   and MGM_G108(MGM_W85,MGM_W84,clk_delay);
   not MGM_G109(MGM_W86,si_delay);
   and MGM_G110(MGM_W87,MGM_W86,MGM_W85);
   and MGM_G111(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W87);
   not MGM_G112(MGM_W88,d_delay);
   and MGM_G113(MGM_W89,MGM_W88,clk_delay);
   and MGM_G114(MGM_W90,si_delay,MGM_W89);
   not MGM_G115(MGM_W91,ssb_delay);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W91,MGM_W90);
   not MGM_G117(MGM_W92,d_delay);
   and MGM_G118(MGM_W93,MGM_W92,clk_delay);
   and MGM_G119(MGM_W94,si_delay,MGM_W93);
   and MGM_G120(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W94);
   and MGM_G121(MGM_W95,d_delay,clk_delay);
   not MGM_G122(MGM_W96,si_delay);
   and MGM_G123(MGM_W97,MGM_W96,MGM_W95);
   not MGM_G124(MGM_W98,ssb_delay);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W98,MGM_W97);
   and MGM_G126(MGM_W99,d_delay,clk_delay);
   not MGM_G127(MGM_W100,si_delay);
   and MGM_G128(MGM_W101,MGM_W100,MGM_W99);
   and MGM_G129(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W101);
   and MGM_G130(MGM_W102,d_delay,clk_delay);
   and MGM_G131(MGM_W103,si_delay,MGM_W102);
   not MGM_G132(MGM_W104,ssb_delay);
   and MGM_G133(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W104,MGM_W103);
   and MGM_G134(MGM_W105,d_delay,clk_delay);
   and MGM_G135(MGM_W106,si_delay,MGM_W105);
   and MGM_G136(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W106);
   not MGM_G137(MGM_W107,d_delay);
   and MGM_G138(MGM_W108,psb_delay,MGM_W107);
   not MGM_G139(MGM_W109,ssb_delay);
   and MGM_G140(ENABLE_NOT_d_AND_psb_AND_NOT_ssb,MGM_W109,MGM_W108);
   and MGM_G141(MGM_W110,psb_delay,d_delay);
   not MGM_G142(MGM_W111,ssb_delay);
   and MGM_G143(ENABLE_d_AND_psb_AND_NOT_ssb,MGM_W111,MGM_W110);
   not MGM_G144(MGM_W112,d_delay);
   and MGM_G145(MGM_W113,psb_delay,MGM_W112);
   and MGM_G146(ENABLE_NOT_d_AND_psb_AND_si,si_delay,MGM_W113);
   and MGM_G147(MGM_W114,psb_delay,d_delay);
   not MGM_G148(MGM_W115,si_delay);
   and MGM_G149(ENABLE_d_AND_psb_AND_NOT_si,MGM_W115,MGM_W114);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy00cah1n12x5( clk, d, o, psb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00cah_func b15fqy00cah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00cah_func b15fqy00cah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00cah_func b15fqy00cah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00cah_func b15fqy00cah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,psb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,psb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,psb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,psb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,psb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,psb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,psb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,psb_delay);
   and MGM_G38(ENABLE_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,psb_delay);
   and MGM_G40(ENABLE_psb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   not MGM_G42(MGM_W32,si_delay);
   and MGM_G43(MGM_W33,MGM_W32,MGM_W31);
   not MGM_G44(MGM_W34,ssb_delay);
   and MGM_G45(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W34,MGM_W33);
   not MGM_G46(MGM_W35,d_delay);
   not MGM_G47(MGM_W36,si_delay);
   and MGM_G48(MGM_W37,MGM_W36,MGM_W35);
   and MGM_G49(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W37);
   not MGM_G50(MGM_W38,d_delay);
   and MGM_G51(MGM_W39,si_delay,MGM_W38);
   and MGM_G52(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W39);
   not MGM_G53(MGM_W40,si_delay);
   and MGM_G54(MGM_W41,MGM_W40,d_delay);
   not MGM_G55(MGM_W42,ssb_delay);
   and MGM_G56(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W42,MGM_W41);
   not MGM_G57(MGM_W43,clk_delay);
   not MGM_G58(MGM_W44,d_delay);
   and MGM_G59(MGM_W45,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W46,si_delay);
   and MGM_G61(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G62(MGM_W48,ssb_delay);
   and MGM_G63(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   not MGM_G64(MGM_W49,clk_delay);
   not MGM_G65(MGM_W50,d_delay);
   and MGM_G66(MGM_W51,MGM_W50,MGM_W49);
   not MGM_G67(MGM_W52,si_delay);
   and MGM_G68(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G69(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G70(MGM_W54,clk_delay);
   not MGM_G71(MGM_W55,d_delay);
   and MGM_G72(MGM_W56,MGM_W55,MGM_W54);
   and MGM_G73(MGM_W57,si_delay,MGM_W56);
   not MGM_G74(MGM_W58,ssb_delay);
   and MGM_G75(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W58,MGM_W57);
   not MGM_G76(MGM_W59,clk_delay);
   not MGM_G77(MGM_W60,d_delay);
   and MGM_G78(MGM_W61,MGM_W60,MGM_W59);
   and MGM_G79(MGM_W62,si_delay,MGM_W61);
   and MGM_G80(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W62);
   not MGM_G81(MGM_W63,clk_delay);
   and MGM_G82(MGM_W64,d_delay,MGM_W63);
   not MGM_G83(MGM_W65,si_delay);
   and MGM_G84(MGM_W66,MGM_W65,MGM_W64);
   not MGM_G85(MGM_W67,ssb_delay);
   and MGM_G86(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W67,MGM_W66);
   not MGM_G87(MGM_W68,clk_delay);
   and MGM_G88(MGM_W69,d_delay,MGM_W68);
   not MGM_G89(MGM_W70,si_delay);
   and MGM_G90(MGM_W71,MGM_W70,MGM_W69);
   and MGM_G91(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W71);
   not MGM_G92(MGM_W72,clk_delay);
   and MGM_G93(MGM_W73,d_delay,MGM_W72);
   and MGM_G94(MGM_W74,si_delay,MGM_W73);
   not MGM_G95(MGM_W75,ssb_delay);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G97(MGM_W76,clk_delay);
   and MGM_G98(MGM_W77,d_delay,MGM_W76);
   and MGM_G99(MGM_W78,si_delay,MGM_W77);
   and MGM_G100(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W78);
   not MGM_G101(MGM_W79,d_delay);
   and MGM_G102(MGM_W80,MGM_W79,clk_delay);
   not MGM_G103(MGM_W81,si_delay);
   and MGM_G104(MGM_W82,MGM_W81,MGM_W80);
   not MGM_G105(MGM_W83,ssb_delay);
   and MGM_G106(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W83,MGM_W82);
   not MGM_G107(MGM_W84,d_delay);
   and MGM_G108(MGM_W85,MGM_W84,clk_delay);
   not MGM_G109(MGM_W86,si_delay);
   and MGM_G110(MGM_W87,MGM_W86,MGM_W85);
   and MGM_G111(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W87);
   not MGM_G112(MGM_W88,d_delay);
   and MGM_G113(MGM_W89,MGM_W88,clk_delay);
   and MGM_G114(MGM_W90,si_delay,MGM_W89);
   not MGM_G115(MGM_W91,ssb_delay);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W91,MGM_W90);
   not MGM_G117(MGM_W92,d_delay);
   and MGM_G118(MGM_W93,MGM_W92,clk_delay);
   and MGM_G119(MGM_W94,si_delay,MGM_W93);
   and MGM_G120(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W94);
   and MGM_G121(MGM_W95,d_delay,clk_delay);
   not MGM_G122(MGM_W96,si_delay);
   and MGM_G123(MGM_W97,MGM_W96,MGM_W95);
   not MGM_G124(MGM_W98,ssb_delay);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W98,MGM_W97);
   and MGM_G126(MGM_W99,d_delay,clk_delay);
   not MGM_G127(MGM_W100,si_delay);
   and MGM_G128(MGM_W101,MGM_W100,MGM_W99);
   and MGM_G129(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W101);
   and MGM_G130(MGM_W102,d_delay,clk_delay);
   and MGM_G131(MGM_W103,si_delay,MGM_W102);
   not MGM_G132(MGM_W104,ssb_delay);
   and MGM_G133(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W104,MGM_W103);
   and MGM_G134(MGM_W105,d_delay,clk_delay);
   and MGM_G135(MGM_W106,si_delay,MGM_W105);
   and MGM_G136(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W106);
   not MGM_G137(MGM_W107,d_delay);
   and MGM_G138(MGM_W108,psb_delay,MGM_W107);
   not MGM_G139(MGM_W109,ssb_delay);
   and MGM_G140(ENABLE_NOT_d_AND_psb_AND_NOT_ssb,MGM_W109,MGM_W108);
   and MGM_G141(MGM_W110,psb_delay,d_delay);
   not MGM_G142(MGM_W111,ssb_delay);
   and MGM_G143(ENABLE_d_AND_psb_AND_NOT_ssb,MGM_W111,MGM_W110);
   not MGM_G144(MGM_W112,d_delay);
   and MGM_G145(MGM_W113,psb_delay,MGM_W112);
   and MGM_G146(ENABLE_NOT_d_AND_psb_AND_si,si_delay,MGM_W113);
   and MGM_G147(MGM_W114,psb_delay,d_delay);
   not MGM_G148(MGM_W115,si_delay);
   and MGM_G149(ENABLE_d_AND_psb_AND_NOT_si,MGM_W115,MGM_W114);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy00cah1n16x5( clk, d, o, psb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00cah_func b15fqy00cah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00cah_func b15fqy00cah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00cah_func b15fqy00cah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00cah_func b15fqy00cah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   not MGM_G2(MGM_W2,si_delay);
   and MGM_G3(MGM_W3,MGM_W2,MGM_W1);
   not MGM_G4(MGM_W4,ssb_delay);
   and MGM_G5(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W5,d_delay);
   and MGM_G7(MGM_W6,psb_delay,MGM_W5);
   not MGM_G8(MGM_W7,si_delay);
   and MGM_G9(MGM_W8,MGM_W7,MGM_W6);
   and MGM_G10(ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W8);
   not MGM_G11(MGM_W9,d_delay);
   and MGM_G12(MGM_W10,psb_delay,MGM_W9);
   and MGM_G13(MGM_W11,si_delay,MGM_W10);
   not MGM_G14(MGM_W12,ssb_delay);
   and MGM_G15(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G16(MGM_W13,d_delay);
   and MGM_G17(MGM_W14,psb_delay,MGM_W13);
   and MGM_G18(MGM_W15,si_delay,MGM_W14);
   and MGM_G19(ENABLE_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W15);
   and MGM_G20(MGM_W16,psb_delay,d_delay);
   not MGM_G21(MGM_W17,si_delay);
   and MGM_G22(MGM_W18,MGM_W17,MGM_W16);
   not MGM_G23(MGM_W19,ssb_delay);
   and MGM_G24(ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W19,MGM_W18);
   and MGM_G25(MGM_W20,psb_delay,d_delay);
   not MGM_G26(MGM_W21,si_delay);
   and MGM_G27(MGM_W22,MGM_W21,MGM_W20);
   and MGM_G28(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W22);
   and MGM_G29(MGM_W23,psb_delay,d_delay);
   and MGM_G30(MGM_W24,si_delay,MGM_W23);
   not MGM_G31(MGM_W25,ssb_delay);
   and MGM_G32(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W25,MGM_W24);
   and MGM_G33(MGM_W26,psb_delay,d_delay);
   and MGM_G34(MGM_W27,si_delay,MGM_W26);
   and MGM_G35(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W27);
   not MGM_G36(MGM_W28,si_delay);
   and MGM_G37(MGM_W29,MGM_W28,psb_delay);
   and MGM_G38(ENABLE_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W29);
   and MGM_G39(MGM_W30,si_delay,psb_delay);
   and MGM_G40(ENABLE_psb_AND_si_AND_ssb,ssb_delay,MGM_W30);
   not MGM_G41(MGM_W31,d_delay);
   not MGM_G42(MGM_W32,si_delay);
   and MGM_G43(MGM_W33,MGM_W32,MGM_W31);
   not MGM_G44(MGM_W34,ssb_delay);
   and MGM_G45(ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W34,MGM_W33);
   not MGM_G46(MGM_W35,d_delay);
   not MGM_G47(MGM_W36,si_delay);
   and MGM_G48(MGM_W37,MGM_W36,MGM_W35);
   and MGM_G49(ENABLE_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W37);
   not MGM_G50(MGM_W38,d_delay);
   and MGM_G51(MGM_W39,si_delay,MGM_W38);
   and MGM_G52(ENABLE_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W39);
   not MGM_G53(MGM_W40,si_delay);
   and MGM_G54(MGM_W41,MGM_W40,d_delay);
   not MGM_G55(MGM_W42,ssb_delay);
   and MGM_G56(ENABLE_d_AND_NOT_si_AND_NOT_ssb,MGM_W42,MGM_W41);
   not MGM_G57(MGM_W43,clk_delay);
   not MGM_G58(MGM_W44,d_delay);
   and MGM_G59(MGM_W45,MGM_W44,MGM_W43);
   not MGM_G60(MGM_W46,si_delay);
   and MGM_G61(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G62(MGM_W48,ssb_delay);
   and MGM_G63(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   not MGM_G64(MGM_W49,clk_delay);
   not MGM_G65(MGM_W50,d_delay);
   and MGM_G66(MGM_W51,MGM_W50,MGM_W49);
   not MGM_G67(MGM_W52,si_delay);
   and MGM_G68(MGM_W53,MGM_W52,MGM_W51);
   and MGM_G69(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W53);
   not MGM_G70(MGM_W54,clk_delay);
   not MGM_G71(MGM_W55,d_delay);
   and MGM_G72(MGM_W56,MGM_W55,MGM_W54);
   and MGM_G73(MGM_W57,si_delay,MGM_W56);
   not MGM_G74(MGM_W58,ssb_delay);
   and MGM_G75(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W58,MGM_W57);
   not MGM_G76(MGM_W59,clk_delay);
   not MGM_G77(MGM_W60,d_delay);
   and MGM_G78(MGM_W61,MGM_W60,MGM_W59);
   and MGM_G79(MGM_W62,si_delay,MGM_W61);
   and MGM_G80(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W62);
   not MGM_G81(MGM_W63,clk_delay);
   and MGM_G82(MGM_W64,d_delay,MGM_W63);
   not MGM_G83(MGM_W65,si_delay);
   and MGM_G84(MGM_W66,MGM_W65,MGM_W64);
   not MGM_G85(MGM_W67,ssb_delay);
   and MGM_G86(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W67,MGM_W66);
   not MGM_G87(MGM_W68,clk_delay);
   and MGM_G88(MGM_W69,d_delay,MGM_W68);
   not MGM_G89(MGM_W70,si_delay);
   and MGM_G90(MGM_W71,MGM_W70,MGM_W69);
   and MGM_G91(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W71);
   not MGM_G92(MGM_W72,clk_delay);
   and MGM_G93(MGM_W73,d_delay,MGM_W72);
   and MGM_G94(MGM_W74,si_delay,MGM_W73);
   not MGM_G95(MGM_W75,ssb_delay);
   and MGM_G96(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G97(MGM_W76,clk_delay);
   and MGM_G98(MGM_W77,d_delay,MGM_W76);
   and MGM_G99(MGM_W78,si_delay,MGM_W77);
   and MGM_G100(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W78);
   not MGM_G101(MGM_W79,d_delay);
   and MGM_G102(MGM_W80,MGM_W79,clk_delay);
   not MGM_G103(MGM_W81,si_delay);
   and MGM_G104(MGM_W82,MGM_W81,MGM_W80);
   not MGM_G105(MGM_W83,ssb_delay);
   and MGM_G106(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W83,MGM_W82);
   not MGM_G107(MGM_W84,d_delay);
   and MGM_G108(MGM_W85,MGM_W84,clk_delay);
   not MGM_G109(MGM_W86,si_delay);
   and MGM_G110(MGM_W87,MGM_W86,MGM_W85);
   and MGM_G111(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W87);
   not MGM_G112(MGM_W88,d_delay);
   and MGM_G113(MGM_W89,MGM_W88,clk_delay);
   and MGM_G114(MGM_W90,si_delay,MGM_W89);
   not MGM_G115(MGM_W91,ssb_delay);
   and MGM_G116(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W91,MGM_W90);
   not MGM_G117(MGM_W92,d_delay);
   and MGM_G118(MGM_W93,MGM_W92,clk_delay);
   and MGM_G119(MGM_W94,si_delay,MGM_W93);
   and MGM_G120(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W94);
   and MGM_G121(MGM_W95,d_delay,clk_delay);
   not MGM_G122(MGM_W96,si_delay);
   and MGM_G123(MGM_W97,MGM_W96,MGM_W95);
   not MGM_G124(MGM_W98,ssb_delay);
   and MGM_G125(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W98,MGM_W97);
   and MGM_G126(MGM_W99,d_delay,clk_delay);
   not MGM_G127(MGM_W100,si_delay);
   and MGM_G128(MGM_W101,MGM_W100,MGM_W99);
   and MGM_G129(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W101);
   and MGM_G130(MGM_W102,d_delay,clk_delay);
   and MGM_G131(MGM_W103,si_delay,MGM_W102);
   not MGM_G132(MGM_W104,ssb_delay);
   and MGM_G133(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W104,MGM_W103);
   and MGM_G134(MGM_W105,d_delay,clk_delay);
   and MGM_G135(MGM_W106,si_delay,MGM_W105);
   and MGM_G136(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W106);
   not MGM_G137(MGM_W107,d_delay);
   and MGM_G138(MGM_W108,psb_delay,MGM_W107);
   not MGM_G139(MGM_W109,ssb_delay);
   and MGM_G140(ENABLE_NOT_d_AND_psb_AND_NOT_ssb,MGM_W109,MGM_W108);
   and MGM_G141(MGM_W110,psb_delay,d_delay);
   not MGM_G142(MGM_W111,ssb_delay);
   and MGM_G143(ENABLE_d_AND_psb_AND_NOT_ssb,MGM_W111,MGM_W110);
   not MGM_G144(MGM_W112,d_delay);
   and MGM_G145(MGM_W113,psb_delay,MGM_W112);
   and MGM_G146(ENABLE_NOT_d_AND_psb_AND_si,si_delay,MGM_W113);
   and MGM_G147(MGM_W114,psb_delay,d_delay);
   not MGM_G148(MGM_W115,si_delay);
   and MGM_G149(ENABLE_d_AND_psb_AND_NOT_si,MGM_W115,MGM_W114);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fqy00fah_func( clk, d, o, psb, rb, si, ssb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb, si, ssb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_P0, psb, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_fqn00fah_LN_IQ_FF_UDP( IQ, MGM_C0, MGM_P0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_P0, psb );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_fqn00fah_LN_IQ_FF_UDP( IQ, MGM_C0, MGM_P0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fqy00fah1n02x5( clk, d, o, psb, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00fah_func b15fqy00fah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00fah_func b15fqy00fah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00fah_func b15fqy00fah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00fah_func b15fqy00fah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(MGM_W2,rb_delay,MGM_W1);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   and MGM_G8(MGM_W7,psb_delay,MGM_W6);
   and MGM_G9(MGM_W8,rb_delay,MGM_W7);
   not MGM_G10(MGM_W9,si_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G12(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W10);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,psb_delay,MGM_W11);
   and MGM_G15(MGM_W13,rb_delay,MGM_W12);
   and MGM_G16(MGM_W14,si_delay,MGM_W13);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,psb_delay,MGM_W16);
   and MGM_G21(MGM_W18,rb_delay,MGM_W17);
   and MGM_G22(MGM_W19,si_delay,MGM_W18);
   and MGM_G23(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W19);
   and MGM_G24(MGM_W20,psb_delay,d_delay);
   and MGM_G25(MGM_W21,rb_delay,MGM_W20);
   not MGM_G26(MGM_W22,si_delay);
   and MGM_G27(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G28(MGM_W24,ssb_delay);
   and MGM_G29(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W24,MGM_W23);
   and MGM_G30(MGM_W25,psb_delay,d_delay);
   and MGM_G31(MGM_W26,rb_delay,MGM_W25);
   not MGM_G32(MGM_W27,si_delay);
   and MGM_G33(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G34(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W28);
   and MGM_G35(MGM_W29,psb_delay,d_delay);
   and MGM_G36(MGM_W30,rb_delay,MGM_W29);
   and MGM_G37(MGM_W31,si_delay,MGM_W30);
   not MGM_G38(MGM_W32,ssb_delay);
   and MGM_G39(ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W32,MGM_W31);
   and MGM_G40(MGM_W33,psb_delay,d_delay);
   and MGM_G41(MGM_W34,rb_delay,MGM_W33);
   and MGM_G42(MGM_W35,si_delay,MGM_W34);
   and MGM_G43(ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G44(MGM_W36,rb_delay,psb_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   and MGM_G47(ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W38);
   and MGM_G48(MGM_W39,rb_delay,psb_delay);
   and MGM_G49(MGM_W40,si_delay,MGM_W39);
   and MGM_G50(ENABLE_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G51(MGM_W41,d_delay);
   and MGM_G52(MGM_W42,rb_delay,MGM_W41);
   not MGM_G53(MGM_W43,si_delay);
   and MGM_G54(MGM_W44,MGM_W43,MGM_W42);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   not MGM_G57(MGM_W46,d_delay);
   and MGM_G58(MGM_W47,rb_delay,MGM_W46);
   not MGM_G59(MGM_W48,si_delay);
   and MGM_G60(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G61(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G62(MGM_W50,d_delay);
   and MGM_G63(MGM_W51,rb_delay,MGM_W50);
   and MGM_G64(MGM_W52,si_delay,MGM_W51);
   and MGM_G65(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G66(MGM_W53,rb_delay,d_delay);
   not MGM_G67(MGM_W54,si_delay);
   and MGM_G68(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G69(MGM_W56,ssb_delay);
   and MGM_G70(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   not MGM_G71(MGM_W57,clk_delay);
   not MGM_G72(MGM_W58,d_delay);
   and MGM_G73(MGM_W59,MGM_W58,MGM_W57);
   and MGM_G74(MGM_W60,rb_delay,MGM_W59);
   not MGM_G75(MGM_W61,si_delay);
   and MGM_G76(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G77(MGM_W63,ssb_delay);
   and MGM_G78(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G79(MGM_W64,clk_delay);
   not MGM_G80(MGM_W65,d_delay);
   and MGM_G81(MGM_W66,MGM_W65,MGM_W64);
   and MGM_G82(MGM_W67,rb_delay,MGM_W66);
   not MGM_G83(MGM_W68,si_delay);
   and MGM_G84(MGM_W69,MGM_W68,MGM_W67);
   and MGM_G85(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W69);
   not MGM_G86(MGM_W70,clk_delay);
   not MGM_G87(MGM_W71,d_delay);
   and MGM_G88(MGM_W72,MGM_W71,MGM_W70);
   and MGM_G89(MGM_W73,rb_delay,MGM_W72);
   and MGM_G90(MGM_W74,si_delay,MGM_W73);
   not MGM_G91(MGM_W75,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G93(MGM_W76,clk_delay);
   not MGM_G94(MGM_W77,d_delay);
   and MGM_G95(MGM_W78,MGM_W77,MGM_W76);
   and MGM_G96(MGM_W79,rb_delay,MGM_W78);
   and MGM_G97(MGM_W80,si_delay,MGM_W79);
   and MGM_G98(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W80);
   not MGM_G99(MGM_W81,clk_delay);
   and MGM_G100(MGM_W82,d_delay,MGM_W81);
   and MGM_G101(MGM_W83,rb_delay,MGM_W82);
   not MGM_G102(MGM_W84,si_delay);
   and MGM_G103(MGM_W85,MGM_W84,MGM_W83);
   not MGM_G104(MGM_W86,ssb_delay);
   and MGM_G105(ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W86,MGM_W85);
   not MGM_G106(MGM_W87,clk_delay);
   and MGM_G107(MGM_W88,d_delay,MGM_W87);
   and MGM_G108(MGM_W89,rb_delay,MGM_W88);
   not MGM_G109(MGM_W90,si_delay);
   and MGM_G110(MGM_W91,MGM_W90,MGM_W89);
   and MGM_G111(ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W91);
   not MGM_G112(MGM_W92,clk_delay);
   and MGM_G113(MGM_W93,d_delay,MGM_W92);
   and MGM_G114(MGM_W94,rb_delay,MGM_W93);
   and MGM_G115(MGM_W95,si_delay,MGM_W94);
   not MGM_G116(MGM_W96,ssb_delay);
   and MGM_G117(ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W96,MGM_W95);
   not MGM_G118(MGM_W97,clk_delay);
   and MGM_G119(MGM_W98,d_delay,MGM_W97);
   and MGM_G120(MGM_W99,rb_delay,MGM_W98);
   and MGM_G121(MGM_W100,si_delay,MGM_W99);
   and MGM_G122(ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W100);
   not MGM_G123(MGM_W101,d_delay);
   and MGM_G124(MGM_W102,MGM_W101,clk_delay);
   and MGM_G125(MGM_W103,rb_delay,MGM_W102);
   not MGM_G126(MGM_W104,si_delay);
   and MGM_G127(MGM_W105,MGM_W104,MGM_W103);
   not MGM_G128(MGM_W106,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W106,MGM_W105);
   not MGM_G130(MGM_W107,d_delay);
   and MGM_G131(MGM_W108,MGM_W107,clk_delay);
   and MGM_G132(MGM_W109,rb_delay,MGM_W108);
   not MGM_G133(MGM_W110,si_delay);
   and MGM_G134(MGM_W111,MGM_W110,MGM_W109);
   and MGM_G135(ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W111);
   not MGM_G136(MGM_W112,d_delay);
   and MGM_G137(MGM_W113,MGM_W112,clk_delay);
   and MGM_G138(MGM_W114,rb_delay,MGM_W113);
   and MGM_G139(MGM_W115,si_delay,MGM_W114);
   not MGM_G140(MGM_W116,ssb_delay);
   and MGM_G141(ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W116,MGM_W115);
   not MGM_G142(MGM_W117,d_delay);
   and MGM_G143(MGM_W118,MGM_W117,clk_delay);
   and MGM_G144(MGM_W119,rb_delay,MGM_W118);
   and MGM_G145(MGM_W120,si_delay,MGM_W119);
   and MGM_G146(ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W120);
   and MGM_G147(MGM_W121,d_delay,clk_delay);
   and MGM_G148(MGM_W122,rb_delay,MGM_W121);
   not MGM_G149(MGM_W123,si_delay);
   and MGM_G150(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G151(MGM_W125,ssb_delay);
   and MGM_G152(ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W125,MGM_W124);
   and MGM_G153(MGM_W126,d_delay,clk_delay);
   and MGM_G154(MGM_W127,rb_delay,MGM_W126);
   not MGM_G155(MGM_W128,si_delay);
   and MGM_G156(MGM_W129,MGM_W128,MGM_W127);
   and MGM_G157(ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W129);
   and MGM_G158(MGM_W130,d_delay,clk_delay);
   and MGM_G159(MGM_W131,rb_delay,MGM_W130);
   and MGM_G160(MGM_W132,si_delay,MGM_W131);
   not MGM_G161(MGM_W133,ssb_delay);
   and MGM_G162(ENABLE_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W133,MGM_W132);
   and MGM_G163(MGM_W134,d_delay,clk_delay);
   and MGM_G164(MGM_W135,rb_delay,MGM_W134);
   and MGM_G165(MGM_W136,si_delay,MGM_W135);
   and MGM_G166(ENABLE_clk_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W136);
   not MGM_G167(MGM_W137,clk_delay);
   not MGM_G168(MGM_W138,d_delay);
   and MGM_G169(MGM_W139,MGM_W138,MGM_W137);
   not MGM_G170(MGM_W140,si_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   not MGM_G172(MGM_W142,ssb_delay);
   and MGM_G173(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W142,MGM_W141);
   not MGM_G174(MGM_W143,clk_delay);
   not MGM_G175(MGM_W144,d_delay);
   and MGM_G176(MGM_W145,MGM_W144,MGM_W143);
   not MGM_G177(MGM_W146,si_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W147);
   not MGM_G180(MGM_W148,clk_delay);
   not MGM_G181(MGM_W149,d_delay);
   and MGM_G182(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G183(MGM_W151,si_delay,MGM_W150);
   not MGM_G184(MGM_W152,ssb_delay);
   and MGM_G185(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W153,clk_delay);
   not MGM_G187(MGM_W154,d_delay);
   and MGM_G188(MGM_W155,MGM_W154,MGM_W153);
   and MGM_G189(MGM_W156,si_delay,MGM_W155);
   and MGM_G190(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W156);
   not MGM_G191(MGM_W157,clk_delay);
   and MGM_G192(MGM_W158,d_delay,MGM_W157);
   not MGM_G193(MGM_W159,si_delay);
   and MGM_G194(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G195(MGM_W161,ssb_delay);
   and MGM_G196(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W161,MGM_W160);
   not MGM_G197(MGM_W162,clk_delay);
   and MGM_G198(MGM_W163,d_delay,MGM_W162);
   not MGM_G199(MGM_W164,si_delay);
   and MGM_G200(MGM_W165,MGM_W164,MGM_W163);
   and MGM_G201(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W165);
   not MGM_G202(MGM_W166,clk_delay);
   and MGM_G203(MGM_W167,d_delay,MGM_W166);
   and MGM_G204(MGM_W168,si_delay,MGM_W167);
   not MGM_G205(MGM_W169,ssb_delay);
   and MGM_G206(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W169,MGM_W168);
   not MGM_G207(MGM_W170,clk_delay);
   and MGM_G208(MGM_W171,d_delay,MGM_W170);
   and MGM_G209(MGM_W172,si_delay,MGM_W171);
   and MGM_G210(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W172);
   not MGM_G211(MGM_W173,d_delay);
   and MGM_G212(MGM_W174,MGM_W173,clk_delay);
   not MGM_G213(MGM_W175,si_delay);
   and MGM_G214(MGM_W176,MGM_W175,MGM_W174);
   not MGM_G215(MGM_W177,ssb_delay);
   and MGM_G216(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W177,MGM_W176);
   not MGM_G217(MGM_W178,d_delay);
   and MGM_G218(MGM_W179,MGM_W178,clk_delay);
   not MGM_G219(MGM_W180,si_delay);
   and MGM_G220(MGM_W181,MGM_W180,MGM_W179);
   and MGM_G221(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W181);
   not MGM_G222(MGM_W182,d_delay);
   and MGM_G223(MGM_W183,MGM_W182,clk_delay);
   and MGM_G224(MGM_W184,si_delay,MGM_W183);
   not MGM_G225(MGM_W185,ssb_delay);
   and MGM_G226(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W185,MGM_W184);
   not MGM_G227(MGM_W186,d_delay);
   and MGM_G228(MGM_W187,MGM_W186,clk_delay);
   and MGM_G229(MGM_W188,si_delay,MGM_W187);
   and MGM_G230(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W188);
   and MGM_G231(MGM_W189,d_delay,clk_delay);
   not MGM_G232(MGM_W190,si_delay);
   and MGM_G233(MGM_W191,MGM_W190,MGM_W189);
   not MGM_G234(MGM_W192,ssb_delay);
   and MGM_G235(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W192,MGM_W191);
   and MGM_G236(MGM_W193,d_delay,clk_delay);
   not MGM_G237(MGM_W194,si_delay);
   and MGM_G238(MGM_W195,MGM_W194,MGM_W193);
   and MGM_G239(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W195);
   and MGM_G240(MGM_W196,d_delay,clk_delay);
   and MGM_G241(MGM_W197,si_delay,MGM_W196);
   not MGM_G242(MGM_W198,ssb_delay);
   and MGM_G243(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W198,MGM_W197);
   and MGM_G244(MGM_W199,d_delay,clk_delay);
   and MGM_G245(MGM_W200,si_delay,MGM_W199);
   and MGM_G246(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W200);
   not MGM_G247(MGM_W201,d_delay);
   and MGM_G248(MGM_W202,psb_delay,MGM_W201);
   and MGM_G249(MGM_W203,si_delay,MGM_W202);
   not MGM_G250(MGM_W204,ssb_delay);
   and MGM_G251(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W204,MGM_W203);
   and MGM_G252(MGM_W205,psb_delay,d_delay);
   not MGM_G253(MGM_W206,si_delay);
   and MGM_G254(MGM_W207,MGM_W206,MGM_W205);
   and MGM_G255(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W207);
   and MGM_G256(MGM_W208,psb_delay,d_delay);
   and MGM_G257(MGM_W209,si_delay,MGM_W208);
   not MGM_G258(MGM_W210,ssb_delay);
   and MGM_G259(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W210,MGM_W209);
   and MGM_G260(MGM_W211,psb_delay,d_delay);
   and MGM_G261(MGM_W212,si_delay,MGM_W211);
   and MGM_G262(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W212);
   not MGM_G263(MGM_W213,clk_delay);
   not MGM_G264(MGM_W214,d_delay);
   and MGM_G265(MGM_W215,MGM_W214,MGM_W213);
   and MGM_G266(MGM_W216,psb_delay,MGM_W215);
   not MGM_G267(MGM_W217,si_delay);
   and MGM_G268(MGM_W218,MGM_W217,MGM_W216);
   not MGM_G269(MGM_W219,ssb_delay);
   and MGM_G270(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W219,MGM_W218);
   not MGM_G271(MGM_W220,clk_delay);
   not MGM_G272(MGM_W221,d_delay);
   and MGM_G273(MGM_W222,MGM_W221,MGM_W220);
   and MGM_G274(MGM_W223,psb_delay,MGM_W222);
   not MGM_G275(MGM_W224,si_delay);
   and MGM_G276(MGM_W225,MGM_W224,MGM_W223);
   and MGM_G277(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W225);
   not MGM_G278(MGM_W226,clk_delay);
   not MGM_G279(MGM_W227,d_delay);
   and MGM_G280(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G281(MGM_W229,psb_delay,MGM_W228);
   and MGM_G282(MGM_W230,si_delay,MGM_W229);
   not MGM_G283(MGM_W231,ssb_delay);
   and MGM_G284(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W231,MGM_W230);
   not MGM_G285(MGM_W232,clk_delay);
   not MGM_G286(MGM_W233,d_delay);
   and MGM_G287(MGM_W234,MGM_W233,MGM_W232);
   and MGM_G288(MGM_W235,psb_delay,MGM_W234);
   and MGM_G289(MGM_W236,si_delay,MGM_W235);
   and MGM_G290(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W236);
   not MGM_G291(MGM_W237,clk_delay);
   and MGM_G292(MGM_W238,d_delay,MGM_W237);
   and MGM_G293(MGM_W239,psb_delay,MGM_W238);
   not MGM_G294(MGM_W240,si_delay);
   and MGM_G295(MGM_W241,MGM_W240,MGM_W239);
   not MGM_G296(MGM_W242,ssb_delay);
   and MGM_G297(ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W242,MGM_W241);
   not MGM_G298(MGM_W243,clk_delay);
   and MGM_G299(MGM_W244,d_delay,MGM_W243);
   and MGM_G300(MGM_W245,psb_delay,MGM_W244);
   not MGM_G301(MGM_W246,si_delay);
   and MGM_G302(MGM_W247,MGM_W246,MGM_W245);
   and MGM_G303(ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W247);
   not MGM_G304(MGM_W248,clk_delay);
   and MGM_G305(MGM_W249,d_delay,MGM_W248);
   and MGM_G306(MGM_W250,psb_delay,MGM_W249);
   and MGM_G307(MGM_W251,si_delay,MGM_W250);
   not MGM_G308(MGM_W252,ssb_delay);
   and MGM_G309(ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W252,MGM_W251);
   not MGM_G310(MGM_W253,clk_delay);
   and MGM_G311(MGM_W254,d_delay,MGM_W253);
   and MGM_G312(MGM_W255,psb_delay,MGM_W254);
   and MGM_G313(MGM_W256,si_delay,MGM_W255);
   and MGM_G314(ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W256);
   not MGM_G315(MGM_W257,d_delay);
   and MGM_G316(MGM_W258,MGM_W257,clk_delay);
   and MGM_G317(MGM_W259,psb_delay,MGM_W258);
   not MGM_G318(MGM_W260,si_delay);
   and MGM_G319(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G320(MGM_W262,ssb_delay);
   and MGM_G321(ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   not MGM_G322(MGM_W263,d_delay);
   and MGM_G323(MGM_W264,MGM_W263,clk_delay);
   and MGM_G324(MGM_W265,psb_delay,MGM_W264);
   not MGM_G325(MGM_W266,si_delay);
   and MGM_G326(MGM_W267,MGM_W266,MGM_W265);
   and MGM_G327(ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W267);
   not MGM_G328(MGM_W268,d_delay);
   and MGM_G329(MGM_W269,MGM_W268,clk_delay);
   and MGM_G330(MGM_W270,psb_delay,MGM_W269);
   and MGM_G331(MGM_W271,si_delay,MGM_W270);
   not MGM_G332(MGM_W272,ssb_delay);
   and MGM_G333(ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W272,MGM_W271);
   not MGM_G334(MGM_W273,d_delay);
   and MGM_G335(MGM_W274,MGM_W273,clk_delay);
   and MGM_G336(MGM_W275,psb_delay,MGM_W274);
   and MGM_G337(MGM_W276,si_delay,MGM_W275);
   and MGM_G338(ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W276);
   and MGM_G339(MGM_W277,d_delay,clk_delay);
   and MGM_G340(MGM_W278,psb_delay,MGM_W277);
   not MGM_G341(MGM_W279,si_delay);
   and MGM_G342(MGM_W280,MGM_W279,MGM_W278);
   not MGM_G343(MGM_W281,ssb_delay);
   and MGM_G344(ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W281,MGM_W280);
   and MGM_G345(MGM_W282,d_delay,clk_delay);
   and MGM_G346(MGM_W283,psb_delay,MGM_W282);
   not MGM_G347(MGM_W284,si_delay);
   and MGM_G348(MGM_W285,MGM_W284,MGM_W283);
   and MGM_G349(ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W285);
   and MGM_G350(MGM_W286,d_delay,clk_delay);
   and MGM_G351(MGM_W287,psb_delay,MGM_W286);
   and MGM_G352(MGM_W288,si_delay,MGM_W287);
   not MGM_G353(MGM_W289,ssb_delay);
   and MGM_G354(ENABLE_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W289,MGM_W288);
   and MGM_G355(MGM_W290,d_delay,clk_delay);
   and MGM_G356(MGM_W291,psb_delay,MGM_W290);
   and MGM_G357(MGM_W292,si_delay,MGM_W291);
   and MGM_G358(ENABLE_clk_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W292);
   not MGM_G359(MGM_W293,d_delay);
   and MGM_G360(MGM_W294,psb_delay,MGM_W293);
   and MGM_G361(MGM_W295,rb_delay,MGM_W294);
   not MGM_G362(MGM_W296,ssb_delay);
   and MGM_G363(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W296,MGM_W295);
   and MGM_G364(MGM_W297,psb_delay,d_delay);
   and MGM_G365(MGM_W298,rb_delay,MGM_W297);
   not MGM_G366(MGM_W299,ssb_delay);
   and MGM_G367(ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W299,MGM_W298);
   not MGM_G368(MGM_W300,d_delay);
   and MGM_G369(MGM_W301,psb_delay,MGM_W300);
   and MGM_G370(MGM_W302,rb_delay,MGM_W301);
   and MGM_G371(ENABLE_NOT_d_AND_psb_AND_rb_AND_si,si_delay,MGM_W302);
   and MGM_G372(MGM_W303,psb_delay,d_delay);
   and MGM_G373(MGM_W304,rb_delay,MGM_W303);
   not MGM_G374(MGM_W305,si_delay);
   and MGM_G375(ENABLE_d_AND_psb_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy00fah1n03x5( clk, d, o, psb, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00fah_func b15fqy00fah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00fah_func b15fqy00fah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00fah_func b15fqy00fah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00fah_func b15fqy00fah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(MGM_W2,rb_delay,MGM_W1);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   and MGM_G8(MGM_W7,psb_delay,MGM_W6);
   and MGM_G9(MGM_W8,rb_delay,MGM_W7);
   not MGM_G10(MGM_W9,si_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G12(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W10);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,psb_delay,MGM_W11);
   and MGM_G15(MGM_W13,rb_delay,MGM_W12);
   and MGM_G16(MGM_W14,si_delay,MGM_W13);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,psb_delay,MGM_W16);
   and MGM_G21(MGM_W18,rb_delay,MGM_W17);
   and MGM_G22(MGM_W19,si_delay,MGM_W18);
   and MGM_G23(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W19);
   and MGM_G24(MGM_W20,psb_delay,d_delay);
   and MGM_G25(MGM_W21,rb_delay,MGM_W20);
   not MGM_G26(MGM_W22,si_delay);
   and MGM_G27(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G28(MGM_W24,ssb_delay);
   and MGM_G29(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W24,MGM_W23);
   and MGM_G30(MGM_W25,psb_delay,d_delay);
   and MGM_G31(MGM_W26,rb_delay,MGM_W25);
   not MGM_G32(MGM_W27,si_delay);
   and MGM_G33(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G34(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W28);
   and MGM_G35(MGM_W29,psb_delay,d_delay);
   and MGM_G36(MGM_W30,rb_delay,MGM_W29);
   and MGM_G37(MGM_W31,si_delay,MGM_W30);
   not MGM_G38(MGM_W32,ssb_delay);
   and MGM_G39(ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W32,MGM_W31);
   and MGM_G40(MGM_W33,psb_delay,d_delay);
   and MGM_G41(MGM_W34,rb_delay,MGM_W33);
   and MGM_G42(MGM_W35,si_delay,MGM_W34);
   and MGM_G43(ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G44(MGM_W36,rb_delay,psb_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   and MGM_G47(ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W38);
   and MGM_G48(MGM_W39,rb_delay,psb_delay);
   and MGM_G49(MGM_W40,si_delay,MGM_W39);
   and MGM_G50(ENABLE_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G51(MGM_W41,d_delay);
   and MGM_G52(MGM_W42,rb_delay,MGM_W41);
   not MGM_G53(MGM_W43,si_delay);
   and MGM_G54(MGM_W44,MGM_W43,MGM_W42);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   not MGM_G57(MGM_W46,d_delay);
   and MGM_G58(MGM_W47,rb_delay,MGM_W46);
   not MGM_G59(MGM_W48,si_delay);
   and MGM_G60(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G61(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G62(MGM_W50,d_delay);
   and MGM_G63(MGM_W51,rb_delay,MGM_W50);
   and MGM_G64(MGM_W52,si_delay,MGM_W51);
   and MGM_G65(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G66(MGM_W53,rb_delay,d_delay);
   not MGM_G67(MGM_W54,si_delay);
   and MGM_G68(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G69(MGM_W56,ssb_delay);
   and MGM_G70(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   not MGM_G71(MGM_W57,clk_delay);
   not MGM_G72(MGM_W58,d_delay);
   and MGM_G73(MGM_W59,MGM_W58,MGM_W57);
   and MGM_G74(MGM_W60,rb_delay,MGM_W59);
   not MGM_G75(MGM_W61,si_delay);
   and MGM_G76(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G77(MGM_W63,ssb_delay);
   and MGM_G78(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G79(MGM_W64,clk_delay);
   not MGM_G80(MGM_W65,d_delay);
   and MGM_G81(MGM_W66,MGM_W65,MGM_W64);
   and MGM_G82(MGM_W67,rb_delay,MGM_W66);
   not MGM_G83(MGM_W68,si_delay);
   and MGM_G84(MGM_W69,MGM_W68,MGM_W67);
   and MGM_G85(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W69);
   not MGM_G86(MGM_W70,clk_delay);
   not MGM_G87(MGM_W71,d_delay);
   and MGM_G88(MGM_W72,MGM_W71,MGM_W70);
   and MGM_G89(MGM_W73,rb_delay,MGM_W72);
   and MGM_G90(MGM_W74,si_delay,MGM_W73);
   not MGM_G91(MGM_W75,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G93(MGM_W76,clk_delay);
   not MGM_G94(MGM_W77,d_delay);
   and MGM_G95(MGM_W78,MGM_W77,MGM_W76);
   and MGM_G96(MGM_W79,rb_delay,MGM_W78);
   and MGM_G97(MGM_W80,si_delay,MGM_W79);
   and MGM_G98(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W80);
   not MGM_G99(MGM_W81,clk_delay);
   and MGM_G100(MGM_W82,d_delay,MGM_W81);
   and MGM_G101(MGM_W83,rb_delay,MGM_W82);
   not MGM_G102(MGM_W84,si_delay);
   and MGM_G103(MGM_W85,MGM_W84,MGM_W83);
   not MGM_G104(MGM_W86,ssb_delay);
   and MGM_G105(ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W86,MGM_W85);
   not MGM_G106(MGM_W87,clk_delay);
   and MGM_G107(MGM_W88,d_delay,MGM_W87);
   and MGM_G108(MGM_W89,rb_delay,MGM_W88);
   not MGM_G109(MGM_W90,si_delay);
   and MGM_G110(MGM_W91,MGM_W90,MGM_W89);
   and MGM_G111(ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W91);
   not MGM_G112(MGM_W92,clk_delay);
   and MGM_G113(MGM_W93,d_delay,MGM_W92);
   and MGM_G114(MGM_W94,rb_delay,MGM_W93);
   and MGM_G115(MGM_W95,si_delay,MGM_W94);
   not MGM_G116(MGM_W96,ssb_delay);
   and MGM_G117(ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W96,MGM_W95);
   not MGM_G118(MGM_W97,clk_delay);
   and MGM_G119(MGM_W98,d_delay,MGM_W97);
   and MGM_G120(MGM_W99,rb_delay,MGM_W98);
   and MGM_G121(MGM_W100,si_delay,MGM_W99);
   and MGM_G122(ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W100);
   not MGM_G123(MGM_W101,d_delay);
   and MGM_G124(MGM_W102,MGM_W101,clk_delay);
   and MGM_G125(MGM_W103,rb_delay,MGM_W102);
   not MGM_G126(MGM_W104,si_delay);
   and MGM_G127(MGM_W105,MGM_W104,MGM_W103);
   not MGM_G128(MGM_W106,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W106,MGM_W105);
   not MGM_G130(MGM_W107,d_delay);
   and MGM_G131(MGM_W108,MGM_W107,clk_delay);
   and MGM_G132(MGM_W109,rb_delay,MGM_W108);
   not MGM_G133(MGM_W110,si_delay);
   and MGM_G134(MGM_W111,MGM_W110,MGM_W109);
   and MGM_G135(ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W111);
   not MGM_G136(MGM_W112,d_delay);
   and MGM_G137(MGM_W113,MGM_W112,clk_delay);
   and MGM_G138(MGM_W114,rb_delay,MGM_W113);
   and MGM_G139(MGM_W115,si_delay,MGM_W114);
   not MGM_G140(MGM_W116,ssb_delay);
   and MGM_G141(ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W116,MGM_W115);
   not MGM_G142(MGM_W117,d_delay);
   and MGM_G143(MGM_W118,MGM_W117,clk_delay);
   and MGM_G144(MGM_W119,rb_delay,MGM_W118);
   and MGM_G145(MGM_W120,si_delay,MGM_W119);
   and MGM_G146(ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W120);
   and MGM_G147(MGM_W121,d_delay,clk_delay);
   and MGM_G148(MGM_W122,rb_delay,MGM_W121);
   not MGM_G149(MGM_W123,si_delay);
   and MGM_G150(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G151(MGM_W125,ssb_delay);
   and MGM_G152(ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W125,MGM_W124);
   and MGM_G153(MGM_W126,d_delay,clk_delay);
   and MGM_G154(MGM_W127,rb_delay,MGM_W126);
   not MGM_G155(MGM_W128,si_delay);
   and MGM_G156(MGM_W129,MGM_W128,MGM_W127);
   and MGM_G157(ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W129);
   and MGM_G158(MGM_W130,d_delay,clk_delay);
   and MGM_G159(MGM_W131,rb_delay,MGM_W130);
   and MGM_G160(MGM_W132,si_delay,MGM_W131);
   not MGM_G161(MGM_W133,ssb_delay);
   and MGM_G162(ENABLE_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W133,MGM_W132);
   and MGM_G163(MGM_W134,d_delay,clk_delay);
   and MGM_G164(MGM_W135,rb_delay,MGM_W134);
   and MGM_G165(MGM_W136,si_delay,MGM_W135);
   and MGM_G166(ENABLE_clk_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W136);
   not MGM_G167(MGM_W137,clk_delay);
   not MGM_G168(MGM_W138,d_delay);
   and MGM_G169(MGM_W139,MGM_W138,MGM_W137);
   not MGM_G170(MGM_W140,si_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   not MGM_G172(MGM_W142,ssb_delay);
   and MGM_G173(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W142,MGM_W141);
   not MGM_G174(MGM_W143,clk_delay);
   not MGM_G175(MGM_W144,d_delay);
   and MGM_G176(MGM_W145,MGM_W144,MGM_W143);
   not MGM_G177(MGM_W146,si_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W147);
   not MGM_G180(MGM_W148,clk_delay);
   not MGM_G181(MGM_W149,d_delay);
   and MGM_G182(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G183(MGM_W151,si_delay,MGM_W150);
   not MGM_G184(MGM_W152,ssb_delay);
   and MGM_G185(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W153,clk_delay);
   not MGM_G187(MGM_W154,d_delay);
   and MGM_G188(MGM_W155,MGM_W154,MGM_W153);
   and MGM_G189(MGM_W156,si_delay,MGM_W155);
   and MGM_G190(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W156);
   not MGM_G191(MGM_W157,clk_delay);
   and MGM_G192(MGM_W158,d_delay,MGM_W157);
   not MGM_G193(MGM_W159,si_delay);
   and MGM_G194(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G195(MGM_W161,ssb_delay);
   and MGM_G196(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W161,MGM_W160);
   not MGM_G197(MGM_W162,clk_delay);
   and MGM_G198(MGM_W163,d_delay,MGM_W162);
   not MGM_G199(MGM_W164,si_delay);
   and MGM_G200(MGM_W165,MGM_W164,MGM_W163);
   and MGM_G201(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W165);
   not MGM_G202(MGM_W166,clk_delay);
   and MGM_G203(MGM_W167,d_delay,MGM_W166);
   and MGM_G204(MGM_W168,si_delay,MGM_W167);
   not MGM_G205(MGM_W169,ssb_delay);
   and MGM_G206(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W169,MGM_W168);
   not MGM_G207(MGM_W170,clk_delay);
   and MGM_G208(MGM_W171,d_delay,MGM_W170);
   and MGM_G209(MGM_W172,si_delay,MGM_W171);
   and MGM_G210(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W172);
   not MGM_G211(MGM_W173,d_delay);
   and MGM_G212(MGM_W174,MGM_W173,clk_delay);
   not MGM_G213(MGM_W175,si_delay);
   and MGM_G214(MGM_W176,MGM_W175,MGM_W174);
   not MGM_G215(MGM_W177,ssb_delay);
   and MGM_G216(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W177,MGM_W176);
   not MGM_G217(MGM_W178,d_delay);
   and MGM_G218(MGM_W179,MGM_W178,clk_delay);
   not MGM_G219(MGM_W180,si_delay);
   and MGM_G220(MGM_W181,MGM_W180,MGM_W179);
   and MGM_G221(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W181);
   not MGM_G222(MGM_W182,d_delay);
   and MGM_G223(MGM_W183,MGM_W182,clk_delay);
   and MGM_G224(MGM_W184,si_delay,MGM_W183);
   not MGM_G225(MGM_W185,ssb_delay);
   and MGM_G226(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W185,MGM_W184);
   not MGM_G227(MGM_W186,d_delay);
   and MGM_G228(MGM_W187,MGM_W186,clk_delay);
   and MGM_G229(MGM_W188,si_delay,MGM_W187);
   and MGM_G230(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W188);
   and MGM_G231(MGM_W189,d_delay,clk_delay);
   not MGM_G232(MGM_W190,si_delay);
   and MGM_G233(MGM_W191,MGM_W190,MGM_W189);
   not MGM_G234(MGM_W192,ssb_delay);
   and MGM_G235(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W192,MGM_W191);
   and MGM_G236(MGM_W193,d_delay,clk_delay);
   not MGM_G237(MGM_W194,si_delay);
   and MGM_G238(MGM_W195,MGM_W194,MGM_W193);
   and MGM_G239(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W195);
   and MGM_G240(MGM_W196,d_delay,clk_delay);
   and MGM_G241(MGM_W197,si_delay,MGM_W196);
   not MGM_G242(MGM_W198,ssb_delay);
   and MGM_G243(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W198,MGM_W197);
   and MGM_G244(MGM_W199,d_delay,clk_delay);
   and MGM_G245(MGM_W200,si_delay,MGM_W199);
   and MGM_G246(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W200);
   not MGM_G247(MGM_W201,d_delay);
   and MGM_G248(MGM_W202,psb_delay,MGM_W201);
   and MGM_G249(MGM_W203,si_delay,MGM_W202);
   not MGM_G250(MGM_W204,ssb_delay);
   and MGM_G251(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W204,MGM_W203);
   and MGM_G252(MGM_W205,psb_delay,d_delay);
   not MGM_G253(MGM_W206,si_delay);
   and MGM_G254(MGM_W207,MGM_W206,MGM_W205);
   and MGM_G255(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W207);
   and MGM_G256(MGM_W208,psb_delay,d_delay);
   and MGM_G257(MGM_W209,si_delay,MGM_W208);
   not MGM_G258(MGM_W210,ssb_delay);
   and MGM_G259(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W210,MGM_W209);
   and MGM_G260(MGM_W211,psb_delay,d_delay);
   and MGM_G261(MGM_W212,si_delay,MGM_W211);
   and MGM_G262(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W212);
   not MGM_G263(MGM_W213,clk_delay);
   not MGM_G264(MGM_W214,d_delay);
   and MGM_G265(MGM_W215,MGM_W214,MGM_W213);
   and MGM_G266(MGM_W216,psb_delay,MGM_W215);
   not MGM_G267(MGM_W217,si_delay);
   and MGM_G268(MGM_W218,MGM_W217,MGM_W216);
   not MGM_G269(MGM_W219,ssb_delay);
   and MGM_G270(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W219,MGM_W218);
   not MGM_G271(MGM_W220,clk_delay);
   not MGM_G272(MGM_W221,d_delay);
   and MGM_G273(MGM_W222,MGM_W221,MGM_W220);
   and MGM_G274(MGM_W223,psb_delay,MGM_W222);
   not MGM_G275(MGM_W224,si_delay);
   and MGM_G276(MGM_W225,MGM_W224,MGM_W223);
   and MGM_G277(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W225);
   not MGM_G278(MGM_W226,clk_delay);
   not MGM_G279(MGM_W227,d_delay);
   and MGM_G280(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G281(MGM_W229,psb_delay,MGM_W228);
   and MGM_G282(MGM_W230,si_delay,MGM_W229);
   not MGM_G283(MGM_W231,ssb_delay);
   and MGM_G284(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W231,MGM_W230);
   not MGM_G285(MGM_W232,clk_delay);
   not MGM_G286(MGM_W233,d_delay);
   and MGM_G287(MGM_W234,MGM_W233,MGM_W232);
   and MGM_G288(MGM_W235,psb_delay,MGM_W234);
   and MGM_G289(MGM_W236,si_delay,MGM_W235);
   and MGM_G290(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W236);
   not MGM_G291(MGM_W237,clk_delay);
   and MGM_G292(MGM_W238,d_delay,MGM_W237);
   and MGM_G293(MGM_W239,psb_delay,MGM_W238);
   not MGM_G294(MGM_W240,si_delay);
   and MGM_G295(MGM_W241,MGM_W240,MGM_W239);
   not MGM_G296(MGM_W242,ssb_delay);
   and MGM_G297(ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W242,MGM_W241);
   not MGM_G298(MGM_W243,clk_delay);
   and MGM_G299(MGM_W244,d_delay,MGM_W243);
   and MGM_G300(MGM_W245,psb_delay,MGM_W244);
   not MGM_G301(MGM_W246,si_delay);
   and MGM_G302(MGM_W247,MGM_W246,MGM_W245);
   and MGM_G303(ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W247);
   not MGM_G304(MGM_W248,clk_delay);
   and MGM_G305(MGM_W249,d_delay,MGM_W248);
   and MGM_G306(MGM_W250,psb_delay,MGM_W249);
   and MGM_G307(MGM_W251,si_delay,MGM_W250);
   not MGM_G308(MGM_W252,ssb_delay);
   and MGM_G309(ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W252,MGM_W251);
   not MGM_G310(MGM_W253,clk_delay);
   and MGM_G311(MGM_W254,d_delay,MGM_W253);
   and MGM_G312(MGM_W255,psb_delay,MGM_W254);
   and MGM_G313(MGM_W256,si_delay,MGM_W255);
   and MGM_G314(ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W256);
   not MGM_G315(MGM_W257,d_delay);
   and MGM_G316(MGM_W258,MGM_W257,clk_delay);
   and MGM_G317(MGM_W259,psb_delay,MGM_W258);
   not MGM_G318(MGM_W260,si_delay);
   and MGM_G319(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G320(MGM_W262,ssb_delay);
   and MGM_G321(ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   not MGM_G322(MGM_W263,d_delay);
   and MGM_G323(MGM_W264,MGM_W263,clk_delay);
   and MGM_G324(MGM_W265,psb_delay,MGM_W264);
   not MGM_G325(MGM_W266,si_delay);
   and MGM_G326(MGM_W267,MGM_W266,MGM_W265);
   and MGM_G327(ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W267);
   not MGM_G328(MGM_W268,d_delay);
   and MGM_G329(MGM_W269,MGM_W268,clk_delay);
   and MGM_G330(MGM_W270,psb_delay,MGM_W269);
   and MGM_G331(MGM_W271,si_delay,MGM_W270);
   not MGM_G332(MGM_W272,ssb_delay);
   and MGM_G333(ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W272,MGM_W271);
   not MGM_G334(MGM_W273,d_delay);
   and MGM_G335(MGM_W274,MGM_W273,clk_delay);
   and MGM_G336(MGM_W275,psb_delay,MGM_W274);
   and MGM_G337(MGM_W276,si_delay,MGM_W275);
   and MGM_G338(ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W276);
   and MGM_G339(MGM_W277,d_delay,clk_delay);
   and MGM_G340(MGM_W278,psb_delay,MGM_W277);
   not MGM_G341(MGM_W279,si_delay);
   and MGM_G342(MGM_W280,MGM_W279,MGM_W278);
   not MGM_G343(MGM_W281,ssb_delay);
   and MGM_G344(ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W281,MGM_W280);
   and MGM_G345(MGM_W282,d_delay,clk_delay);
   and MGM_G346(MGM_W283,psb_delay,MGM_W282);
   not MGM_G347(MGM_W284,si_delay);
   and MGM_G348(MGM_W285,MGM_W284,MGM_W283);
   and MGM_G349(ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W285);
   and MGM_G350(MGM_W286,d_delay,clk_delay);
   and MGM_G351(MGM_W287,psb_delay,MGM_W286);
   and MGM_G352(MGM_W288,si_delay,MGM_W287);
   not MGM_G353(MGM_W289,ssb_delay);
   and MGM_G354(ENABLE_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W289,MGM_W288);
   and MGM_G355(MGM_W290,d_delay,clk_delay);
   and MGM_G356(MGM_W291,psb_delay,MGM_W290);
   and MGM_G357(MGM_W292,si_delay,MGM_W291);
   and MGM_G358(ENABLE_clk_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W292);
   not MGM_G359(MGM_W293,d_delay);
   and MGM_G360(MGM_W294,psb_delay,MGM_W293);
   and MGM_G361(MGM_W295,rb_delay,MGM_W294);
   not MGM_G362(MGM_W296,ssb_delay);
   and MGM_G363(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W296,MGM_W295);
   and MGM_G364(MGM_W297,psb_delay,d_delay);
   and MGM_G365(MGM_W298,rb_delay,MGM_W297);
   not MGM_G366(MGM_W299,ssb_delay);
   and MGM_G367(ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W299,MGM_W298);
   not MGM_G368(MGM_W300,d_delay);
   and MGM_G369(MGM_W301,psb_delay,MGM_W300);
   and MGM_G370(MGM_W302,rb_delay,MGM_W301);
   and MGM_G371(ENABLE_NOT_d_AND_psb_AND_rb_AND_si,si_delay,MGM_W302);
   and MGM_G372(MGM_W303,psb_delay,d_delay);
   and MGM_G373(MGM_W304,rb_delay,MGM_W303);
   not MGM_G374(MGM_W305,si_delay);
   and MGM_G375(ENABLE_d_AND_psb_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy00fah1n04x5( clk, d, o, psb, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00fah_func b15fqy00fah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00fah_func b15fqy00fah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00fah_func b15fqy00fah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00fah_func b15fqy00fah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(MGM_W2,rb_delay,MGM_W1);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   and MGM_G8(MGM_W7,psb_delay,MGM_W6);
   and MGM_G9(MGM_W8,rb_delay,MGM_W7);
   not MGM_G10(MGM_W9,si_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G12(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W10);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,psb_delay,MGM_W11);
   and MGM_G15(MGM_W13,rb_delay,MGM_W12);
   and MGM_G16(MGM_W14,si_delay,MGM_W13);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,psb_delay,MGM_W16);
   and MGM_G21(MGM_W18,rb_delay,MGM_W17);
   and MGM_G22(MGM_W19,si_delay,MGM_W18);
   and MGM_G23(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W19);
   and MGM_G24(MGM_W20,psb_delay,d_delay);
   and MGM_G25(MGM_W21,rb_delay,MGM_W20);
   not MGM_G26(MGM_W22,si_delay);
   and MGM_G27(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G28(MGM_W24,ssb_delay);
   and MGM_G29(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W24,MGM_W23);
   and MGM_G30(MGM_W25,psb_delay,d_delay);
   and MGM_G31(MGM_W26,rb_delay,MGM_W25);
   not MGM_G32(MGM_W27,si_delay);
   and MGM_G33(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G34(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W28);
   and MGM_G35(MGM_W29,psb_delay,d_delay);
   and MGM_G36(MGM_W30,rb_delay,MGM_W29);
   and MGM_G37(MGM_W31,si_delay,MGM_W30);
   not MGM_G38(MGM_W32,ssb_delay);
   and MGM_G39(ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W32,MGM_W31);
   and MGM_G40(MGM_W33,psb_delay,d_delay);
   and MGM_G41(MGM_W34,rb_delay,MGM_W33);
   and MGM_G42(MGM_W35,si_delay,MGM_W34);
   and MGM_G43(ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G44(MGM_W36,rb_delay,psb_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   and MGM_G47(ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W38);
   and MGM_G48(MGM_W39,rb_delay,psb_delay);
   and MGM_G49(MGM_W40,si_delay,MGM_W39);
   and MGM_G50(ENABLE_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G51(MGM_W41,d_delay);
   and MGM_G52(MGM_W42,rb_delay,MGM_W41);
   not MGM_G53(MGM_W43,si_delay);
   and MGM_G54(MGM_W44,MGM_W43,MGM_W42);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   not MGM_G57(MGM_W46,d_delay);
   and MGM_G58(MGM_W47,rb_delay,MGM_W46);
   not MGM_G59(MGM_W48,si_delay);
   and MGM_G60(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G61(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G62(MGM_W50,d_delay);
   and MGM_G63(MGM_W51,rb_delay,MGM_W50);
   and MGM_G64(MGM_W52,si_delay,MGM_W51);
   and MGM_G65(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G66(MGM_W53,rb_delay,d_delay);
   not MGM_G67(MGM_W54,si_delay);
   and MGM_G68(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G69(MGM_W56,ssb_delay);
   and MGM_G70(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   not MGM_G71(MGM_W57,clk_delay);
   not MGM_G72(MGM_W58,d_delay);
   and MGM_G73(MGM_W59,MGM_W58,MGM_W57);
   and MGM_G74(MGM_W60,rb_delay,MGM_W59);
   not MGM_G75(MGM_W61,si_delay);
   and MGM_G76(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G77(MGM_W63,ssb_delay);
   and MGM_G78(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G79(MGM_W64,clk_delay);
   not MGM_G80(MGM_W65,d_delay);
   and MGM_G81(MGM_W66,MGM_W65,MGM_W64);
   and MGM_G82(MGM_W67,rb_delay,MGM_W66);
   not MGM_G83(MGM_W68,si_delay);
   and MGM_G84(MGM_W69,MGM_W68,MGM_W67);
   and MGM_G85(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W69);
   not MGM_G86(MGM_W70,clk_delay);
   not MGM_G87(MGM_W71,d_delay);
   and MGM_G88(MGM_W72,MGM_W71,MGM_W70);
   and MGM_G89(MGM_W73,rb_delay,MGM_W72);
   and MGM_G90(MGM_W74,si_delay,MGM_W73);
   not MGM_G91(MGM_W75,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G93(MGM_W76,clk_delay);
   not MGM_G94(MGM_W77,d_delay);
   and MGM_G95(MGM_W78,MGM_W77,MGM_W76);
   and MGM_G96(MGM_W79,rb_delay,MGM_W78);
   and MGM_G97(MGM_W80,si_delay,MGM_W79);
   and MGM_G98(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W80);
   not MGM_G99(MGM_W81,clk_delay);
   and MGM_G100(MGM_W82,d_delay,MGM_W81);
   and MGM_G101(MGM_W83,rb_delay,MGM_W82);
   not MGM_G102(MGM_W84,si_delay);
   and MGM_G103(MGM_W85,MGM_W84,MGM_W83);
   not MGM_G104(MGM_W86,ssb_delay);
   and MGM_G105(ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W86,MGM_W85);
   not MGM_G106(MGM_W87,clk_delay);
   and MGM_G107(MGM_W88,d_delay,MGM_W87);
   and MGM_G108(MGM_W89,rb_delay,MGM_W88);
   not MGM_G109(MGM_W90,si_delay);
   and MGM_G110(MGM_W91,MGM_W90,MGM_W89);
   and MGM_G111(ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W91);
   not MGM_G112(MGM_W92,clk_delay);
   and MGM_G113(MGM_W93,d_delay,MGM_W92);
   and MGM_G114(MGM_W94,rb_delay,MGM_W93);
   and MGM_G115(MGM_W95,si_delay,MGM_W94);
   not MGM_G116(MGM_W96,ssb_delay);
   and MGM_G117(ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W96,MGM_W95);
   not MGM_G118(MGM_W97,clk_delay);
   and MGM_G119(MGM_W98,d_delay,MGM_W97);
   and MGM_G120(MGM_W99,rb_delay,MGM_W98);
   and MGM_G121(MGM_W100,si_delay,MGM_W99);
   and MGM_G122(ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W100);
   not MGM_G123(MGM_W101,d_delay);
   and MGM_G124(MGM_W102,MGM_W101,clk_delay);
   and MGM_G125(MGM_W103,rb_delay,MGM_W102);
   not MGM_G126(MGM_W104,si_delay);
   and MGM_G127(MGM_W105,MGM_W104,MGM_W103);
   not MGM_G128(MGM_W106,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W106,MGM_W105);
   not MGM_G130(MGM_W107,d_delay);
   and MGM_G131(MGM_W108,MGM_W107,clk_delay);
   and MGM_G132(MGM_W109,rb_delay,MGM_W108);
   not MGM_G133(MGM_W110,si_delay);
   and MGM_G134(MGM_W111,MGM_W110,MGM_W109);
   and MGM_G135(ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W111);
   not MGM_G136(MGM_W112,d_delay);
   and MGM_G137(MGM_W113,MGM_W112,clk_delay);
   and MGM_G138(MGM_W114,rb_delay,MGM_W113);
   and MGM_G139(MGM_W115,si_delay,MGM_W114);
   not MGM_G140(MGM_W116,ssb_delay);
   and MGM_G141(ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W116,MGM_W115);
   not MGM_G142(MGM_W117,d_delay);
   and MGM_G143(MGM_W118,MGM_W117,clk_delay);
   and MGM_G144(MGM_W119,rb_delay,MGM_W118);
   and MGM_G145(MGM_W120,si_delay,MGM_W119);
   and MGM_G146(ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W120);
   and MGM_G147(MGM_W121,d_delay,clk_delay);
   and MGM_G148(MGM_W122,rb_delay,MGM_W121);
   not MGM_G149(MGM_W123,si_delay);
   and MGM_G150(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G151(MGM_W125,ssb_delay);
   and MGM_G152(ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W125,MGM_W124);
   and MGM_G153(MGM_W126,d_delay,clk_delay);
   and MGM_G154(MGM_W127,rb_delay,MGM_W126);
   not MGM_G155(MGM_W128,si_delay);
   and MGM_G156(MGM_W129,MGM_W128,MGM_W127);
   and MGM_G157(ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W129);
   and MGM_G158(MGM_W130,d_delay,clk_delay);
   and MGM_G159(MGM_W131,rb_delay,MGM_W130);
   and MGM_G160(MGM_W132,si_delay,MGM_W131);
   not MGM_G161(MGM_W133,ssb_delay);
   and MGM_G162(ENABLE_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W133,MGM_W132);
   and MGM_G163(MGM_W134,d_delay,clk_delay);
   and MGM_G164(MGM_W135,rb_delay,MGM_W134);
   and MGM_G165(MGM_W136,si_delay,MGM_W135);
   and MGM_G166(ENABLE_clk_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W136);
   not MGM_G167(MGM_W137,clk_delay);
   not MGM_G168(MGM_W138,d_delay);
   and MGM_G169(MGM_W139,MGM_W138,MGM_W137);
   not MGM_G170(MGM_W140,si_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   not MGM_G172(MGM_W142,ssb_delay);
   and MGM_G173(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W142,MGM_W141);
   not MGM_G174(MGM_W143,clk_delay);
   not MGM_G175(MGM_W144,d_delay);
   and MGM_G176(MGM_W145,MGM_W144,MGM_W143);
   not MGM_G177(MGM_W146,si_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W147);
   not MGM_G180(MGM_W148,clk_delay);
   not MGM_G181(MGM_W149,d_delay);
   and MGM_G182(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G183(MGM_W151,si_delay,MGM_W150);
   not MGM_G184(MGM_W152,ssb_delay);
   and MGM_G185(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W153,clk_delay);
   not MGM_G187(MGM_W154,d_delay);
   and MGM_G188(MGM_W155,MGM_W154,MGM_W153);
   and MGM_G189(MGM_W156,si_delay,MGM_W155);
   and MGM_G190(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W156);
   not MGM_G191(MGM_W157,clk_delay);
   and MGM_G192(MGM_W158,d_delay,MGM_W157);
   not MGM_G193(MGM_W159,si_delay);
   and MGM_G194(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G195(MGM_W161,ssb_delay);
   and MGM_G196(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W161,MGM_W160);
   not MGM_G197(MGM_W162,clk_delay);
   and MGM_G198(MGM_W163,d_delay,MGM_W162);
   not MGM_G199(MGM_W164,si_delay);
   and MGM_G200(MGM_W165,MGM_W164,MGM_W163);
   and MGM_G201(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W165);
   not MGM_G202(MGM_W166,clk_delay);
   and MGM_G203(MGM_W167,d_delay,MGM_W166);
   and MGM_G204(MGM_W168,si_delay,MGM_W167);
   not MGM_G205(MGM_W169,ssb_delay);
   and MGM_G206(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W169,MGM_W168);
   not MGM_G207(MGM_W170,clk_delay);
   and MGM_G208(MGM_W171,d_delay,MGM_W170);
   and MGM_G209(MGM_W172,si_delay,MGM_W171);
   and MGM_G210(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W172);
   not MGM_G211(MGM_W173,d_delay);
   and MGM_G212(MGM_W174,MGM_W173,clk_delay);
   not MGM_G213(MGM_W175,si_delay);
   and MGM_G214(MGM_W176,MGM_W175,MGM_W174);
   not MGM_G215(MGM_W177,ssb_delay);
   and MGM_G216(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W177,MGM_W176);
   not MGM_G217(MGM_W178,d_delay);
   and MGM_G218(MGM_W179,MGM_W178,clk_delay);
   not MGM_G219(MGM_W180,si_delay);
   and MGM_G220(MGM_W181,MGM_W180,MGM_W179);
   and MGM_G221(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W181);
   not MGM_G222(MGM_W182,d_delay);
   and MGM_G223(MGM_W183,MGM_W182,clk_delay);
   and MGM_G224(MGM_W184,si_delay,MGM_W183);
   not MGM_G225(MGM_W185,ssb_delay);
   and MGM_G226(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W185,MGM_W184);
   not MGM_G227(MGM_W186,d_delay);
   and MGM_G228(MGM_W187,MGM_W186,clk_delay);
   and MGM_G229(MGM_W188,si_delay,MGM_W187);
   and MGM_G230(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W188);
   and MGM_G231(MGM_W189,d_delay,clk_delay);
   not MGM_G232(MGM_W190,si_delay);
   and MGM_G233(MGM_W191,MGM_W190,MGM_W189);
   not MGM_G234(MGM_W192,ssb_delay);
   and MGM_G235(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W192,MGM_W191);
   and MGM_G236(MGM_W193,d_delay,clk_delay);
   not MGM_G237(MGM_W194,si_delay);
   and MGM_G238(MGM_W195,MGM_W194,MGM_W193);
   and MGM_G239(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W195);
   and MGM_G240(MGM_W196,d_delay,clk_delay);
   and MGM_G241(MGM_W197,si_delay,MGM_W196);
   not MGM_G242(MGM_W198,ssb_delay);
   and MGM_G243(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W198,MGM_W197);
   and MGM_G244(MGM_W199,d_delay,clk_delay);
   and MGM_G245(MGM_W200,si_delay,MGM_W199);
   and MGM_G246(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W200);
   not MGM_G247(MGM_W201,d_delay);
   and MGM_G248(MGM_W202,psb_delay,MGM_W201);
   and MGM_G249(MGM_W203,si_delay,MGM_W202);
   not MGM_G250(MGM_W204,ssb_delay);
   and MGM_G251(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W204,MGM_W203);
   and MGM_G252(MGM_W205,psb_delay,d_delay);
   not MGM_G253(MGM_W206,si_delay);
   and MGM_G254(MGM_W207,MGM_W206,MGM_W205);
   and MGM_G255(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W207);
   and MGM_G256(MGM_W208,psb_delay,d_delay);
   and MGM_G257(MGM_W209,si_delay,MGM_W208);
   not MGM_G258(MGM_W210,ssb_delay);
   and MGM_G259(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W210,MGM_W209);
   and MGM_G260(MGM_W211,psb_delay,d_delay);
   and MGM_G261(MGM_W212,si_delay,MGM_W211);
   and MGM_G262(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W212);
   not MGM_G263(MGM_W213,clk_delay);
   not MGM_G264(MGM_W214,d_delay);
   and MGM_G265(MGM_W215,MGM_W214,MGM_W213);
   and MGM_G266(MGM_W216,psb_delay,MGM_W215);
   not MGM_G267(MGM_W217,si_delay);
   and MGM_G268(MGM_W218,MGM_W217,MGM_W216);
   not MGM_G269(MGM_W219,ssb_delay);
   and MGM_G270(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W219,MGM_W218);
   not MGM_G271(MGM_W220,clk_delay);
   not MGM_G272(MGM_W221,d_delay);
   and MGM_G273(MGM_W222,MGM_W221,MGM_W220);
   and MGM_G274(MGM_W223,psb_delay,MGM_W222);
   not MGM_G275(MGM_W224,si_delay);
   and MGM_G276(MGM_W225,MGM_W224,MGM_W223);
   and MGM_G277(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W225);
   not MGM_G278(MGM_W226,clk_delay);
   not MGM_G279(MGM_W227,d_delay);
   and MGM_G280(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G281(MGM_W229,psb_delay,MGM_W228);
   and MGM_G282(MGM_W230,si_delay,MGM_W229);
   not MGM_G283(MGM_W231,ssb_delay);
   and MGM_G284(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W231,MGM_W230);
   not MGM_G285(MGM_W232,clk_delay);
   not MGM_G286(MGM_W233,d_delay);
   and MGM_G287(MGM_W234,MGM_W233,MGM_W232);
   and MGM_G288(MGM_W235,psb_delay,MGM_W234);
   and MGM_G289(MGM_W236,si_delay,MGM_W235);
   and MGM_G290(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W236);
   not MGM_G291(MGM_W237,clk_delay);
   and MGM_G292(MGM_W238,d_delay,MGM_W237);
   and MGM_G293(MGM_W239,psb_delay,MGM_W238);
   not MGM_G294(MGM_W240,si_delay);
   and MGM_G295(MGM_W241,MGM_W240,MGM_W239);
   not MGM_G296(MGM_W242,ssb_delay);
   and MGM_G297(ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W242,MGM_W241);
   not MGM_G298(MGM_W243,clk_delay);
   and MGM_G299(MGM_W244,d_delay,MGM_W243);
   and MGM_G300(MGM_W245,psb_delay,MGM_W244);
   not MGM_G301(MGM_W246,si_delay);
   and MGM_G302(MGM_W247,MGM_W246,MGM_W245);
   and MGM_G303(ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W247);
   not MGM_G304(MGM_W248,clk_delay);
   and MGM_G305(MGM_W249,d_delay,MGM_W248);
   and MGM_G306(MGM_W250,psb_delay,MGM_W249);
   and MGM_G307(MGM_W251,si_delay,MGM_W250);
   not MGM_G308(MGM_W252,ssb_delay);
   and MGM_G309(ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W252,MGM_W251);
   not MGM_G310(MGM_W253,clk_delay);
   and MGM_G311(MGM_W254,d_delay,MGM_W253);
   and MGM_G312(MGM_W255,psb_delay,MGM_W254);
   and MGM_G313(MGM_W256,si_delay,MGM_W255);
   and MGM_G314(ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W256);
   not MGM_G315(MGM_W257,d_delay);
   and MGM_G316(MGM_W258,MGM_W257,clk_delay);
   and MGM_G317(MGM_W259,psb_delay,MGM_W258);
   not MGM_G318(MGM_W260,si_delay);
   and MGM_G319(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G320(MGM_W262,ssb_delay);
   and MGM_G321(ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   not MGM_G322(MGM_W263,d_delay);
   and MGM_G323(MGM_W264,MGM_W263,clk_delay);
   and MGM_G324(MGM_W265,psb_delay,MGM_W264);
   not MGM_G325(MGM_W266,si_delay);
   and MGM_G326(MGM_W267,MGM_W266,MGM_W265);
   and MGM_G327(ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W267);
   not MGM_G328(MGM_W268,d_delay);
   and MGM_G329(MGM_W269,MGM_W268,clk_delay);
   and MGM_G330(MGM_W270,psb_delay,MGM_W269);
   and MGM_G331(MGM_W271,si_delay,MGM_W270);
   not MGM_G332(MGM_W272,ssb_delay);
   and MGM_G333(ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W272,MGM_W271);
   not MGM_G334(MGM_W273,d_delay);
   and MGM_G335(MGM_W274,MGM_W273,clk_delay);
   and MGM_G336(MGM_W275,psb_delay,MGM_W274);
   and MGM_G337(MGM_W276,si_delay,MGM_W275);
   and MGM_G338(ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W276);
   and MGM_G339(MGM_W277,d_delay,clk_delay);
   and MGM_G340(MGM_W278,psb_delay,MGM_W277);
   not MGM_G341(MGM_W279,si_delay);
   and MGM_G342(MGM_W280,MGM_W279,MGM_W278);
   not MGM_G343(MGM_W281,ssb_delay);
   and MGM_G344(ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W281,MGM_W280);
   and MGM_G345(MGM_W282,d_delay,clk_delay);
   and MGM_G346(MGM_W283,psb_delay,MGM_W282);
   not MGM_G347(MGM_W284,si_delay);
   and MGM_G348(MGM_W285,MGM_W284,MGM_W283);
   and MGM_G349(ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W285);
   and MGM_G350(MGM_W286,d_delay,clk_delay);
   and MGM_G351(MGM_W287,psb_delay,MGM_W286);
   and MGM_G352(MGM_W288,si_delay,MGM_W287);
   not MGM_G353(MGM_W289,ssb_delay);
   and MGM_G354(ENABLE_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W289,MGM_W288);
   and MGM_G355(MGM_W290,d_delay,clk_delay);
   and MGM_G356(MGM_W291,psb_delay,MGM_W290);
   and MGM_G357(MGM_W292,si_delay,MGM_W291);
   and MGM_G358(ENABLE_clk_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W292);
   not MGM_G359(MGM_W293,d_delay);
   and MGM_G360(MGM_W294,psb_delay,MGM_W293);
   and MGM_G361(MGM_W295,rb_delay,MGM_W294);
   not MGM_G362(MGM_W296,ssb_delay);
   and MGM_G363(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W296,MGM_W295);
   and MGM_G364(MGM_W297,psb_delay,d_delay);
   and MGM_G365(MGM_W298,rb_delay,MGM_W297);
   not MGM_G366(MGM_W299,ssb_delay);
   and MGM_G367(ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W299,MGM_W298);
   not MGM_G368(MGM_W300,d_delay);
   and MGM_G369(MGM_W301,psb_delay,MGM_W300);
   and MGM_G370(MGM_W302,rb_delay,MGM_W301);
   and MGM_G371(ENABLE_NOT_d_AND_psb_AND_rb_AND_si,si_delay,MGM_W302);
   and MGM_G372(MGM_W303,psb_delay,d_delay);
   and MGM_G373(MGM_W304,rb_delay,MGM_W303);
   not MGM_G374(MGM_W305,si_delay);
   and MGM_G375(ENABLE_d_AND_psb_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy00fah1n06x5( clk, d, o, psb, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00fah_func b15fqy00fah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00fah_func b15fqy00fah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00fah_func b15fqy00fah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00fah_func b15fqy00fah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(MGM_W2,rb_delay,MGM_W1);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   and MGM_G8(MGM_W7,psb_delay,MGM_W6);
   and MGM_G9(MGM_W8,rb_delay,MGM_W7);
   not MGM_G10(MGM_W9,si_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G12(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W10);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,psb_delay,MGM_W11);
   and MGM_G15(MGM_W13,rb_delay,MGM_W12);
   and MGM_G16(MGM_W14,si_delay,MGM_W13);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,psb_delay,MGM_W16);
   and MGM_G21(MGM_W18,rb_delay,MGM_W17);
   and MGM_G22(MGM_W19,si_delay,MGM_W18);
   and MGM_G23(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W19);
   and MGM_G24(MGM_W20,psb_delay,d_delay);
   and MGM_G25(MGM_W21,rb_delay,MGM_W20);
   not MGM_G26(MGM_W22,si_delay);
   and MGM_G27(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G28(MGM_W24,ssb_delay);
   and MGM_G29(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W24,MGM_W23);
   and MGM_G30(MGM_W25,psb_delay,d_delay);
   and MGM_G31(MGM_W26,rb_delay,MGM_W25);
   not MGM_G32(MGM_W27,si_delay);
   and MGM_G33(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G34(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W28);
   and MGM_G35(MGM_W29,psb_delay,d_delay);
   and MGM_G36(MGM_W30,rb_delay,MGM_W29);
   and MGM_G37(MGM_W31,si_delay,MGM_W30);
   not MGM_G38(MGM_W32,ssb_delay);
   and MGM_G39(ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W32,MGM_W31);
   and MGM_G40(MGM_W33,psb_delay,d_delay);
   and MGM_G41(MGM_W34,rb_delay,MGM_W33);
   and MGM_G42(MGM_W35,si_delay,MGM_W34);
   and MGM_G43(ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G44(MGM_W36,rb_delay,psb_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   and MGM_G47(ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W38);
   and MGM_G48(MGM_W39,rb_delay,psb_delay);
   and MGM_G49(MGM_W40,si_delay,MGM_W39);
   and MGM_G50(ENABLE_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G51(MGM_W41,d_delay);
   and MGM_G52(MGM_W42,rb_delay,MGM_W41);
   not MGM_G53(MGM_W43,si_delay);
   and MGM_G54(MGM_W44,MGM_W43,MGM_W42);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   not MGM_G57(MGM_W46,d_delay);
   and MGM_G58(MGM_W47,rb_delay,MGM_W46);
   not MGM_G59(MGM_W48,si_delay);
   and MGM_G60(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G61(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G62(MGM_W50,d_delay);
   and MGM_G63(MGM_W51,rb_delay,MGM_W50);
   and MGM_G64(MGM_W52,si_delay,MGM_W51);
   and MGM_G65(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G66(MGM_W53,rb_delay,d_delay);
   not MGM_G67(MGM_W54,si_delay);
   and MGM_G68(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G69(MGM_W56,ssb_delay);
   and MGM_G70(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   not MGM_G71(MGM_W57,clk_delay);
   not MGM_G72(MGM_W58,d_delay);
   and MGM_G73(MGM_W59,MGM_W58,MGM_W57);
   and MGM_G74(MGM_W60,rb_delay,MGM_W59);
   not MGM_G75(MGM_W61,si_delay);
   and MGM_G76(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G77(MGM_W63,ssb_delay);
   and MGM_G78(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G79(MGM_W64,clk_delay);
   not MGM_G80(MGM_W65,d_delay);
   and MGM_G81(MGM_W66,MGM_W65,MGM_W64);
   and MGM_G82(MGM_W67,rb_delay,MGM_W66);
   not MGM_G83(MGM_W68,si_delay);
   and MGM_G84(MGM_W69,MGM_W68,MGM_W67);
   and MGM_G85(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W69);
   not MGM_G86(MGM_W70,clk_delay);
   not MGM_G87(MGM_W71,d_delay);
   and MGM_G88(MGM_W72,MGM_W71,MGM_W70);
   and MGM_G89(MGM_W73,rb_delay,MGM_W72);
   and MGM_G90(MGM_W74,si_delay,MGM_W73);
   not MGM_G91(MGM_W75,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G93(MGM_W76,clk_delay);
   not MGM_G94(MGM_W77,d_delay);
   and MGM_G95(MGM_W78,MGM_W77,MGM_W76);
   and MGM_G96(MGM_W79,rb_delay,MGM_W78);
   and MGM_G97(MGM_W80,si_delay,MGM_W79);
   and MGM_G98(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W80);
   not MGM_G99(MGM_W81,clk_delay);
   and MGM_G100(MGM_W82,d_delay,MGM_W81);
   and MGM_G101(MGM_W83,rb_delay,MGM_W82);
   not MGM_G102(MGM_W84,si_delay);
   and MGM_G103(MGM_W85,MGM_W84,MGM_W83);
   not MGM_G104(MGM_W86,ssb_delay);
   and MGM_G105(ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W86,MGM_W85);
   not MGM_G106(MGM_W87,clk_delay);
   and MGM_G107(MGM_W88,d_delay,MGM_W87);
   and MGM_G108(MGM_W89,rb_delay,MGM_W88);
   not MGM_G109(MGM_W90,si_delay);
   and MGM_G110(MGM_W91,MGM_W90,MGM_W89);
   and MGM_G111(ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W91);
   not MGM_G112(MGM_W92,clk_delay);
   and MGM_G113(MGM_W93,d_delay,MGM_W92);
   and MGM_G114(MGM_W94,rb_delay,MGM_W93);
   and MGM_G115(MGM_W95,si_delay,MGM_W94);
   not MGM_G116(MGM_W96,ssb_delay);
   and MGM_G117(ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W96,MGM_W95);
   not MGM_G118(MGM_W97,clk_delay);
   and MGM_G119(MGM_W98,d_delay,MGM_W97);
   and MGM_G120(MGM_W99,rb_delay,MGM_W98);
   and MGM_G121(MGM_W100,si_delay,MGM_W99);
   and MGM_G122(ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W100);
   not MGM_G123(MGM_W101,d_delay);
   and MGM_G124(MGM_W102,MGM_W101,clk_delay);
   and MGM_G125(MGM_W103,rb_delay,MGM_W102);
   not MGM_G126(MGM_W104,si_delay);
   and MGM_G127(MGM_W105,MGM_W104,MGM_W103);
   not MGM_G128(MGM_W106,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W106,MGM_W105);
   not MGM_G130(MGM_W107,d_delay);
   and MGM_G131(MGM_W108,MGM_W107,clk_delay);
   and MGM_G132(MGM_W109,rb_delay,MGM_W108);
   not MGM_G133(MGM_W110,si_delay);
   and MGM_G134(MGM_W111,MGM_W110,MGM_W109);
   and MGM_G135(ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W111);
   not MGM_G136(MGM_W112,d_delay);
   and MGM_G137(MGM_W113,MGM_W112,clk_delay);
   and MGM_G138(MGM_W114,rb_delay,MGM_W113);
   and MGM_G139(MGM_W115,si_delay,MGM_W114);
   not MGM_G140(MGM_W116,ssb_delay);
   and MGM_G141(ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W116,MGM_W115);
   not MGM_G142(MGM_W117,d_delay);
   and MGM_G143(MGM_W118,MGM_W117,clk_delay);
   and MGM_G144(MGM_W119,rb_delay,MGM_W118);
   and MGM_G145(MGM_W120,si_delay,MGM_W119);
   and MGM_G146(ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W120);
   and MGM_G147(MGM_W121,d_delay,clk_delay);
   and MGM_G148(MGM_W122,rb_delay,MGM_W121);
   not MGM_G149(MGM_W123,si_delay);
   and MGM_G150(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G151(MGM_W125,ssb_delay);
   and MGM_G152(ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W125,MGM_W124);
   and MGM_G153(MGM_W126,d_delay,clk_delay);
   and MGM_G154(MGM_W127,rb_delay,MGM_W126);
   not MGM_G155(MGM_W128,si_delay);
   and MGM_G156(MGM_W129,MGM_W128,MGM_W127);
   and MGM_G157(ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W129);
   and MGM_G158(MGM_W130,d_delay,clk_delay);
   and MGM_G159(MGM_W131,rb_delay,MGM_W130);
   and MGM_G160(MGM_W132,si_delay,MGM_W131);
   not MGM_G161(MGM_W133,ssb_delay);
   and MGM_G162(ENABLE_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W133,MGM_W132);
   and MGM_G163(MGM_W134,d_delay,clk_delay);
   and MGM_G164(MGM_W135,rb_delay,MGM_W134);
   and MGM_G165(MGM_W136,si_delay,MGM_W135);
   and MGM_G166(ENABLE_clk_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W136);
   not MGM_G167(MGM_W137,clk_delay);
   not MGM_G168(MGM_W138,d_delay);
   and MGM_G169(MGM_W139,MGM_W138,MGM_W137);
   not MGM_G170(MGM_W140,si_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   not MGM_G172(MGM_W142,ssb_delay);
   and MGM_G173(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W142,MGM_W141);
   not MGM_G174(MGM_W143,clk_delay);
   not MGM_G175(MGM_W144,d_delay);
   and MGM_G176(MGM_W145,MGM_W144,MGM_W143);
   not MGM_G177(MGM_W146,si_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W147);
   not MGM_G180(MGM_W148,clk_delay);
   not MGM_G181(MGM_W149,d_delay);
   and MGM_G182(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G183(MGM_W151,si_delay,MGM_W150);
   not MGM_G184(MGM_W152,ssb_delay);
   and MGM_G185(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W153,clk_delay);
   not MGM_G187(MGM_W154,d_delay);
   and MGM_G188(MGM_W155,MGM_W154,MGM_W153);
   and MGM_G189(MGM_W156,si_delay,MGM_W155);
   and MGM_G190(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W156);
   not MGM_G191(MGM_W157,clk_delay);
   and MGM_G192(MGM_W158,d_delay,MGM_W157);
   not MGM_G193(MGM_W159,si_delay);
   and MGM_G194(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G195(MGM_W161,ssb_delay);
   and MGM_G196(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W161,MGM_W160);
   not MGM_G197(MGM_W162,clk_delay);
   and MGM_G198(MGM_W163,d_delay,MGM_W162);
   not MGM_G199(MGM_W164,si_delay);
   and MGM_G200(MGM_W165,MGM_W164,MGM_W163);
   and MGM_G201(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W165);
   not MGM_G202(MGM_W166,clk_delay);
   and MGM_G203(MGM_W167,d_delay,MGM_W166);
   and MGM_G204(MGM_W168,si_delay,MGM_W167);
   not MGM_G205(MGM_W169,ssb_delay);
   and MGM_G206(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W169,MGM_W168);
   not MGM_G207(MGM_W170,clk_delay);
   and MGM_G208(MGM_W171,d_delay,MGM_W170);
   and MGM_G209(MGM_W172,si_delay,MGM_W171);
   and MGM_G210(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W172);
   not MGM_G211(MGM_W173,d_delay);
   and MGM_G212(MGM_W174,MGM_W173,clk_delay);
   not MGM_G213(MGM_W175,si_delay);
   and MGM_G214(MGM_W176,MGM_W175,MGM_W174);
   not MGM_G215(MGM_W177,ssb_delay);
   and MGM_G216(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W177,MGM_W176);
   not MGM_G217(MGM_W178,d_delay);
   and MGM_G218(MGM_W179,MGM_W178,clk_delay);
   not MGM_G219(MGM_W180,si_delay);
   and MGM_G220(MGM_W181,MGM_W180,MGM_W179);
   and MGM_G221(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W181);
   not MGM_G222(MGM_W182,d_delay);
   and MGM_G223(MGM_W183,MGM_W182,clk_delay);
   and MGM_G224(MGM_W184,si_delay,MGM_W183);
   not MGM_G225(MGM_W185,ssb_delay);
   and MGM_G226(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W185,MGM_W184);
   not MGM_G227(MGM_W186,d_delay);
   and MGM_G228(MGM_W187,MGM_W186,clk_delay);
   and MGM_G229(MGM_W188,si_delay,MGM_W187);
   and MGM_G230(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W188);
   and MGM_G231(MGM_W189,d_delay,clk_delay);
   not MGM_G232(MGM_W190,si_delay);
   and MGM_G233(MGM_W191,MGM_W190,MGM_W189);
   not MGM_G234(MGM_W192,ssb_delay);
   and MGM_G235(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W192,MGM_W191);
   and MGM_G236(MGM_W193,d_delay,clk_delay);
   not MGM_G237(MGM_W194,si_delay);
   and MGM_G238(MGM_W195,MGM_W194,MGM_W193);
   and MGM_G239(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W195);
   and MGM_G240(MGM_W196,d_delay,clk_delay);
   and MGM_G241(MGM_W197,si_delay,MGM_W196);
   not MGM_G242(MGM_W198,ssb_delay);
   and MGM_G243(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W198,MGM_W197);
   and MGM_G244(MGM_W199,d_delay,clk_delay);
   and MGM_G245(MGM_W200,si_delay,MGM_W199);
   and MGM_G246(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W200);
   not MGM_G247(MGM_W201,d_delay);
   and MGM_G248(MGM_W202,psb_delay,MGM_W201);
   and MGM_G249(MGM_W203,si_delay,MGM_W202);
   not MGM_G250(MGM_W204,ssb_delay);
   and MGM_G251(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W204,MGM_W203);
   and MGM_G252(MGM_W205,psb_delay,d_delay);
   not MGM_G253(MGM_W206,si_delay);
   and MGM_G254(MGM_W207,MGM_W206,MGM_W205);
   and MGM_G255(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W207);
   and MGM_G256(MGM_W208,psb_delay,d_delay);
   and MGM_G257(MGM_W209,si_delay,MGM_W208);
   not MGM_G258(MGM_W210,ssb_delay);
   and MGM_G259(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W210,MGM_W209);
   and MGM_G260(MGM_W211,psb_delay,d_delay);
   and MGM_G261(MGM_W212,si_delay,MGM_W211);
   and MGM_G262(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W212);
   not MGM_G263(MGM_W213,clk_delay);
   not MGM_G264(MGM_W214,d_delay);
   and MGM_G265(MGM_W215,MGM_W214,MGM_W213);
   and MGM_G266(MGM_W216,psb_delay,MGM_W215);
   not MGM_G267(MGM_W217,si_delay);
   and MGM_G268(MGM_W218,MGM_W217,MGM_W216);
   not MGM_G269(MGM_W219,ssb_delay);
   and MGM_G270(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W219,MGM_W218);
   not MGM_G271(MGM_W220,clk_delay);
   not MGM_G272(MGM_W221,d_delay);
   and MGM_G273(MGM_W222,MGM_W221,MGM_W220);
   and MGM_G274(MGM_W223,psb_delay,MGM_W222);
   not MGM_G275(MGM_W224,si_delay);
   and MGM_G276(MGM_W225,MGM_W224,MGM_W223);
   and MGM_G277(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W225);
   not MGM_G278(MGM_W226,clk_delay);
   not MGM_G279(MGM_W227,d_delay);
   and MGM_G280(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G281(MGM_W229,psb_delay,MGM_W228);
   and MGM_G282(MGM_W230,si_delay,MGM_W229);
   not MGM_G283(MGM_W231,ssb_delay);
   and MGM_G284(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W231,MGM_W230);
   not MGM_G285(MGM_W232,clk_delay);
   not MGM_G286(MGM_W233,d_delay);
   and MGM_G287(MGM_W234,MGM_W233,MGM_W232);
   and MGM_G288(MGM_W235,psb_delay,MGM_W234);
   and MGM_G289(MGM_W236,si_delay,MGM_W235);
   and MGM_G290(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W236);
   not MGM_G291(MGM_W237,clk_delay);
   and MGM_G292(MGM_W238,d_delay,MGM_W237);
   and MGM_G293(MGM_W239,psb_delay,MGM_W238);
   not MGM_G294(MGM_W240,si_delay);
   and MGM_G295(MGM_W241,MGM_W240,MGM_W239);
   not MGM_G296(MGM_W242,ssb_delay);
   and MGM_G297(ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W242,MGM_W241);
   not MGM_G298(MGM_W243,clk_delay);
   and MGM_G299(MGM_W244,d_delay,MGM_W243);
   and MGM_G300(MGM_W245,psb_delay,MGM_W244);
   not MGM_G301(MGM_W246,si_delay);
   and MGM_G302(MGM_W247,MGM_W246,MGM_W245);
   and MGM_G303(ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W247);
   not MGM_G304(MGM_W248,clk_delay);
   and MGM_G305(MGM_W249,d_delay,MGM_W248);
   and MGM_G306(MGM_W250,psb_delay,MGM_W249);
   and MGM_G307(MGM_W251,si_delay,MGM_W250);
   not MGM_G308(MGM_W252,ssb_delay);
   and MGM_G309(ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W252,MGM_W251);
   not MGM_G310(MGM_W253,clk_delay);
   and MGM_G311(MGM_W254,d_delay,MGM_W253);
   and MGM_G312(MGM_W255,psb_delay,MGM_W254);
   and MGM_G313(MGM_W256,si_delay,MGM_W255);
   and MGM_G314(ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W256);
   not MGM_G315(MGM_W257,d_delay);
   and MGM_G316(MGM_W258,MGM_W257,clk_delay);
   and MGM_G317(MGM_W259,psb_delay,MGM_W258);
   not MGM_G318(MGM_W260,si_delay);
   and MGM_G319(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G320(MGM_W262,ssb_delay);
   and MGM_G321(ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   not MGM_G322(MGM_W263,d_delay);
   and MGM_G323(MGM_W264,MGM_W263,clk_delay);
   and MGM_G324(MGM_W265,psb_delay,MGM_W264);
   not MGM_G325(MGM_W266,si_delay);
   and MGM_G326(MGM_W267,MGM_W266,MGM_W265);
   and MGM_G327(ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W267);
   not MGM_G328(MGM_W268,d_delay);
   and MGM_G329(MGM_W269,MGM_W268,clk_delay);
   and MGM_G330(MGM_W270,psb_delay,MGM_W269);
   and MGM_G331(MGM_W271,si_delay,MGM_W270);
   not MGM_G332(MGM_W272,ssb_delay);
   and MGM_G333(ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W272,MGM_W271);
   not MGM_G334(MGM_W273,d_delay);
   and MGM_G335(MGM_W274,MGM_W273,clk_delay);
   and MGM_G336(MGM_W275,psb_delay,MGM_W274);
   and MGM_G337(MGM_W276,si_delay,MGM_W275);
   and MGM_G338(ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W276);
   and MGM_G339(MGM_W277,d_delay,clk_delay);
   and MGM_G340(MGM_W278,psb_delay,MGM_W277);
   not MGM_G341(MGM_W279,si_delay);
   and MGM_G342(MGM_W280,MGM_W279,MGM_W278);
   not MGM_G343(MGM_W281,ssb_delay);
   and MGM_G344(ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W281,MGM_W280);
   and MGM_G345(MGM_W282,d_delay,clk_delay);
   and MGM_G346(MGM_W283,psb_delay,MGM_W282);
   not MGM_G347(MGM_W284,si_delay);
   and MGM_G348(MGM_W285,MGM_W284,MGM_W283);
   and MGM_G349(ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W285);
   and MGM_G350(MGM_W286,d_delay,clk_delay);
   and MGM_G351(MGM_W287,psb_delay,MGM_W286);
   and MGM_G352(MGM_W288,si_delay,MGM_W287);
   not MGM_G353(MGM_W289,ssb_delay);
   and MGM_G354(ENABLE_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W289,MGM_W288);
   and MGM_G355(MGM_W290,d_delay,clk_delay);
   and MGM_G356(MGM_W291,psb_delay,MGM_W290);
   and MGM_G357(MGM_W292,si_delay,MGM_W291);
   and MGM_G358(ENABLE_clk_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W292);
   not MGM_G359(MGM_W293,d_delay);
   and MGM_G360(MGM_W294,psb_delay,MGM_W293);
   and MGM_G361(MGM_W295,rb_delay,MGM_W294);
   not MGM_G362(MGM_W296,ssb_delay);
   and MGM_G363(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W296,MGM_W295);
   and MGM_G364(MGM_W297,psb_delay,d_delay);
   and MGM_G365(MGM_W298,rb_delay,MGM_W297);
   not MGM_G366(MGM_W299,ssb_delay);
   and MGM_G367(ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W299,MGM_W298);
   not MGM_G368(MGM_W300,d_delay);
   and MGM_G369(MGM_W301,psb_delay,MGM_W300);
   and MGM_G370(MGM_W302,rb_delay,MGM_W301);
   and MGM_G371(ENABLE_NOT_d_AND_psb_AND_rb_AND_si,si_delay,MGM_W302);
   and MGM_G372(MGM_W303,psb_delay,d_delay);
   and MGM_G373(MGM_W304,rb_delay,MGM_W303);
   not MGM_G374(MGM_W305,si_delay);
   and MGM_G375(ENABLE_d_AND_psb_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy00fah1n08x5( clk, d, o, psb, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00fah_func b15fqy00fah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00fah_func b15fqy00fah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00fah_func b15fqy00fah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00fah_func b15fqy00fah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(MGM_W2,rb_delay,MGM_W1);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   and MGM_G8(MGM_W7,psb_delay,MGM_W6);
   and MGM_G9(MGM_W8,rb_delay,MGM_W7);
   not MGM_G10(MGM_W9,si_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G12(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W10);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,psb_delay,MGM_W11);
   and MGM_G15(MGM_W13,rb_delay,MGM_W12);
   and MGM_G16(MGM_W14,si_delay,MGM_W13);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,psb_delay,MGM_W16);
   and MGM_G21(MGM_W18,rb_delay,MGM_W17);
   and MGM_G22(MGM_W19,si_delay,MGM_W18);
   and MGM_G23(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W19);
   and MGM_G24(MGM_W20,psb_delay,d_delay);
   and MGM_G25(MGM_W21,rb_delay,MGM_W20);
   not MGM_G26(MGM_W22,si_delay);
   and MGM_G27(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G28(MGM_W24,ssb_delay);
   and MGM_G29(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W24,MGM_W23);
   and MGM_G30(MGM_W25,psb_delay,d_delay);
   and MGM_G31(MGM_W26,rb_delay,MGM_W25);
   not MGM_G32(MGM_W27,si_delay);
   and MGM_G33(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G34(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W28);
   and MGM_G35(MGM_W29,psb_delay,d_delay);
   and MGM_G36(MGM_W30,rb_delay,MGM_W29);
   and MGM_G37(MGM_W31,si_delay,MGM_W30);
   not MGM_G38(MGM_W32,ssb_delay);
   and MGM_G39(ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W32,MGM_W31);
   and MGM_G40(MGM_W33,psb_delay,d_delay);
   and MGM_G41(MGM_W34,rb_delay,MGM_W33);
   and MGM_G42(MGM_W35,si_delay,MGM_W34);
   and MGM_G43(ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G44(MGM_W36,rb_delay,psb_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   and MGM_G47(ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W38);
   and MGM_G48(MGM_W39,rb_delay,psb_delay);
   and MGM_G49(MGM_W40,si_delay,MGM_W39);
   and MGM_G50(ENABLE_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G51(MGM_W41,d_delay);
   and MGM_G52(MGM_W42,rb_delay,MGM_W41);
   not MGM_G53(MGM_W43,si_delay);
   and MGM_G54(MGM_W44,MGM_W43,MGM_W42);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   not MGM_G57(MGM_W46,d_delay);
   and MGM_G58(MGM_W47,rb_delay,MGM_W46);
   not MGM_G59(MGM_W48,si_delay);
   and MGM_G60(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G61(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G62(MGM_W50,d_delay);
   and MGM_G63(MGM_W51,rb_delay,MGM_W50);
   and MGM_G64(MGM_W52,si_delay,MGM_W51);
   and MGM_G65(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G66(MGM_W53,rb_delay,d_delay);
   not MGM_G67(MGM_W54,si_delay);
   and MGM_G68(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G69(MGM_W56,ssb_delay);
   and MGM_G70(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   not MGM_G71(MGM_W57,clk_delay);
   not MGM_G72(MGM_W58,d_delay);
   and MGM_G73(MGM_W59,MGM_W58,MGM_W57);
   and MGM_G74(MGM_W60,rb_delay,MGM_W59);
   not MGM_G75(MGM_W61,si_delay);
   and MGM_G76(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G77(MGM_W63,ssb_delay);
   and MGM_G78(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G79(MGM_W64,clk_delay);
   not MGM_G80(MGM_W65,d_delay);
   and MGM_G81(MGM_W66,MGM_W65,MGM_W64);
   and MGM_G82(MGM_W67,rb_delay,MGM_W66);
   not MGM_G83(MGM_W68,si_delay);
   and MGM_G84(MGM_W69,MGM_W68,MGM_W67);
   and MGM_G85(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W69);
   not MGM_G86(MGM_W70,clk_delay);
   not MGM_G87(MGM_W71,d_delay);
   and MGM_G88(MGM_W72,MGM_W71,MGM_W70);
   and MGM_G89(MGM_W73,rb_delay,MGM_W72);
   and MGM_G90(MGM_W74,si_delay,MGM_W73);
   not MGM_G91(MGM_W75,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G93(MGM_W76,clk_delay);
   not MGM_G94(MGM_W77,d_delay);
   and MGM_G95(MGM_W78,MGM_W77,MGM_W76);
   and MGM_G96(MGM_W79,rb_delay,MGM_W78);
   and MGM_G97(MGM_W80,si_delay,MGM_W79);
   and MGM_G98(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W80);
   not MGM_G99(MGM_W81,clk_delay);
   and MGM_G100(MGM_W82,d_delay,MGM_W81);
   and MGM_G101(MGM_W83,rb_delay,MGM_W82);
   not MGM_G102(MGM_W84,si_delay);
   and MGM_G103(MGM_W85,MGM_W84,MGM_W83);
   not MGM_G104(MGM_W86,ssb_delay);
   and MGM_G105(ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W86,MGM_W85);
   not MGM_G106(MGM_W87,clk_delay);
   and MGM_G107(MGM_W88,d_delay,MGM_W87);
   and MGM_G108(MGM_W89,rb_delay,MGM_W88);
   not MGM_G109(MGM_W90,si_delay);
   and MGM_G110(MGM_W91,MGM_W90,MGM_W89);
   and MGM_G111(ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W91);
   not MGM_G112(MGM_W92,clk_delay);
   and MGM_G113(MGM_W93,d_delay,MGM_W92);
   and MGM_G114(MGM_W94,rb_delay,MGM_W93);
   and MGM_G115(MGM_W95,si_delay,MGM_W94);
   not MGM_G116(MGM_W96,ssb_delay);
   and MGM_G117(ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W96,MGM_W95);
   not MGM_G118(MGM_W97,clk_delay);
   and MGM_G119(MGM_W98,d_delay,MGM_W97);
   and MGM_G120(MGM_W99,rb_delay,MGM_W98);
   and MGM_G121(MGM_W100,si_delay,MGM_W99);
   and MGM_G122(ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W100);
   not MGM_G123(MGM_W101,d_delay);
   and MGM_G124(MGM_W102,MGM_W101,clk_delay);
   and MGM_G125(MGM_W103,rb_delay,MGM_W102);
   not MGM_G126(MGM_W104,si_delay);
   and MGM_G127(MGM_W105,MGM_W104,MGM_W103);
   not MGM_G128(MGM_W106,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W106,MGM_W105);
   not MGM_G130(MGM_W107,d_delay);
   and MGM_G131(MGM_W108,MGM_W107,clk_delay);
   and MGM_G132(MGM_W109,rb_delay,MGM_W108);
   not MGM_G133(MGM_W110,si_delay);
   and MGM_G134(MGM_W111,MGM_W110,MGM_W109);
   and MGM_G135(ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W111);
   not MGM_G136(MGM_W112,d_delay);
   and MGM_G137(MGM_W113,MGM_W112,clk_delay);
   and MGM_G138(MGM_W114,rb_delay,MGM_W113);
   and MGM_G139(MGM_W115,si_delay,MGM_W114);
   not MGM_G140(MGM_W116,ssb_delay);
   and MGM_G141(ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W116,MGM_W115);
   not MGM_G142(MGM_W117,d_delay);
   and MGM_G143(MGM_W118,MGM_W117,clk_delay);
   and MGM_G144(MGM_W119,rb_delay,MGM_W118);
   and MGM_G145(MGM_W120,si_delay,MGM_W119);
   and MGM_G146(ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W120);
   and MGM_G147(MGM_W121,d_delay,clk_delay);
   and MGM_G148(MGM_W122,rb_delay,MGM_W121);
   not MGM_G149(MGM_W123,si_delay);
   and MGM_G150(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G151(MGM_W125,ssb_delay);
   and MGM_G152(ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W125,MGM_W124);
   and MGM_G153(MGM_W126,d_delay,clk_delay);
   and MGM_G154(MGM_W127,rb_delay,MGM_W126);
   not MGM_G155(MGM_W128,si_delay);
   and MGM_G156(MGM_W129,MGM_W128,MGM_W127);
   and MGM_G157(ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W129);
   and MGM_G158(MGM_W130,d_delay,clk_delay);
   and MGM_G159(MGM_W131,rb_delay,MGM_W130);
   and MGM_G160(MGM_W132,si_delay,MGM_W131);
   not MGM_G161(MGM_W133,ssb_delay);
   and MGM_G162(ENABLE_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W133,MGM_W132);
   and MGM_G163(MGM_W134,d_delay,clk_delay);
   and MGM_G164(MGM_W135,rb_delay,MGM_W134);
   and MGM_G165(MGM_W136,si_delay,MGM_W135);
   and MGM_G166(ENABLE_clk_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W136);
   not MGM_G167(MGM_W137,clk_delay);
   not MGM_G168(MGM_W138,d_delay);
   and MGM_G169(MGM_W139,MGM_W138,MGM_W137);
   not MGM_G170(MGM_W140,si_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   not MGM_G172(MGM_W142,ssb_delay);
   and MGM_G173(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W142,MGM_W141);
   not MGM_G174(MGM_W143,clk_delay);
   not MGM_G175(MGM_W144,d_delay);
   and MGM_G176(MGM_W145,MGM_W144,MGM_W143);
   not MGM_G177(MGM_W146,si_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W147);
   not MGM_G180(MGM_W148,clk_delay);
   not MGM_G181(MGM_W149,d_delay);
   and MGM_G182(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G183(MGM_W151,si_delay,MGM_W150);
   not MGM_G184(MGM_W152,ssb_delay);
   and MGM_G185(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W153,clk_delay);
   not MGM_G187(MGM_W154,d_delay);
   and MGM_G188(MGM_W155,MGM_W154,MGM_W153);
   and MGM_G189(MGM_W156,si_delay,MGM_W155);
   and MGM_G190(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W156);
   not MGM_G191(MGM_W157,clk_delay);
   and MGM_G192(MGM_W158,d_delay,MGM_W157);
   not MGM_G193(MGM_W159,si_delay);
   and MGM_G194(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G195(MGM_W161,ssb_delay);
   and MGM_G196(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W161,MGM_W160);
   not MGM_G197(MGM_W162,clk_delay);
   and MGM_G198(MGM_W163,d_delay,MGM_W162);
   not MGM_G199(MGM_W164,si_delay);
   and MGM_G200(MGM_W165,MGM_W164,MGM_W163);
   and MGM_G201(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W165);
   not MGM_G202(MGM_W166,clk_delay);
   and MGM_G203(MGM_W167,d_delay,MGM_W166);
   and MGM_G204(MGM_W168,si_delay,MGM_W167);
   not MGM_G205(MGM_W169,ssb_delay);
   and MGM_G206(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W169,MGM_W168);
   not MGM_G207(MGM_W170,clk_delay);
   and MGM_G208(MGM_W171,d_delay,MGM_W170);
   and MGM_G209(MGM_W172,si_delay,MGM_W171);
   and MGM_G210(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W172);
   not MGM_G211(MGM_W173,d_delay);
   and MGM_G212(MGM_W174,MGM_W173,clk_delay);
   not MGM_G213(MGM_W175,si_delay);
   and MGM_G214(MGM_W176,MGM_W175,MGM_W174);
   not MGM_G215(MGM_W177,ssb_delay);
   and MGM_G216(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W177,MGM_W176);
   not MGM_G217(MGM_W178,d_delay);
   and MGM_G218(MGM_W179,MGM_W178,clk_delay);
   not MGM_G219(MGM_W180,si_delay);
   and MGM_G220(MGM_W181,MGM_W180,MGM_W179);
   and MGM_G221(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W181);
   not MGM_G222(MGM_W182,d_delay);
   and MGM_G223(MGM_W183,MGM_W182,clk_delay);
   and MGM_G224(MGM_W184,si_delay,MGM_W183);
   not MGM_G225(MGM_W185,ssb_delay);
   and MGM_G226(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W185,MGM_W184);
   not MGM_G227(MGM_W186,d_delay);
   and MGM_G228(MGM_W187,MGM_W186,clk_delay);
   and MGM_G229(MGM_W188,si_delay,MGM_W187);
   and MGM_G230(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W188);
   and MGM_G231(MGM_W189,d_delay,clk_delay);
   not MGM_G232(MGM_W190,si_delay);
   and MGM_G233(MGM_W191,MGM_W190,MGM_W189);
   not MGM_G234(MGM_W192,ssb_delay);
   and MGM_G235(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W192,MGM_W191);
   and MGM_G236(MGM_W193,d_delay,clk_delay);
   not MGM_G237(MGM_W194,si_delay);
   and MGM_G238(MGM_W195,MGM_W194,MGM_W193);
   and MGM_G239(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W195);
   and MGM_G240(MGM_W196,d_delay,clk_delay);
   and MGM_G241(MGM_W197,si_delay,MGM_W196);
   not MGM_G242(MGM_W198,ssb_delay);
   and MGM_G243(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W198,MGM_W197);
   and MGM_G244(MGM_W199,d_delay,clk_delay);
   and MGM_G245(MGM_W200,si_delay,MGM_W199);
   and MGM_G246(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W200);
   not MGM_G247(MGM_W201,d_delay);
   and MGM_G248(MGM_W202,psb_delay,MGM_W201);
   and MGM_G249(MGM_W203,si_delay,MGM_W202);
   not MGM_G250(MGM_W204,ssb_delay);
   and MGM_G251(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W204,MGM_W203);
   and MGM_G252(MGM_W205,psb_delay,d_delay);
   not MGM_G253(MGM_W206,si_delay);
   and MGM_G254(MGM_W207,MGM_W206,MGM_W205);
   and MGM_G255(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W207);
   and MGM_G256(MGM_W208,psb_delay,d_delay);
   and MGM_G257(MGM_W209,si_delay,MGM_W208);
   not MGM_G258(MGM_W210,ssb_delay);
   and MGM_G259(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W210,MGM_W209);
   and MGM_G260(MGM_W211,psb_delay,d_delay);
   and MGM_G261(MGM_W212,si_delay,MGM_W211);
   and MGM_G262(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W212);
   not MGM_G263(MGM_W213,clk_delay);
   not MGM_G264(MGM_W214,d_delay);
   and MGM_G265(MGM_W215,MGM_W214,MGM_W213);
   and MGM_G266(MGM_W216,psb_delay,MGM_W215);
   not MGM_G267(MGM_W217,si_delay);
   and MGM_G268(MGM_W218,MGM_W217,MGM_W216);
   not MGM_G269(MGM_W219,ssb_delay);
   and MGM_G270(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W219,MGM_W218);
   not MGM_G271(MGM_W220,clk_delay);
   not MGM_G272(MGM_W221,d_delay);
   and MGM_G273(MGM_W222,MGM_W221,MGM_W220);
   and MGM_G274(MGM_W223,psb_delay,MGM_W222);
   not MGM_G275(MGM_W224,si_delay);
   and MGM_G276(MGM_W225,MGM_W224,MGM_W223);
   and MGM_G277(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W225);
   not MGM_G278(MGM_W226,clk_delay);
   not MGM_G279(MGM_W227,d_delay);
   and MGM_G280(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G281(MGM_W229,psb_delay,MGM_W228);
   and MGM_G282(MGM_W230,si_delay,MGM_W229);
   not MGM_G283(MGM_W231,ssb_delay);
   and MGM_G284(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W231,MGM_W230);
   not MGM_G285(MGM_W232,clk_delay);
   not MGM_G286(MGM_W233,d_delay);
   and MGM_G287(MGM_W234,MGM_W233,MGM_W232);
   and MGM_G288(MGM_W235,psb_delay,MGM_W234);
   and MGM_G289(MGM_W236,si_delay,MGM_W235);
   and MGM_G290(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W236);
   not MGM_G291(MGM_W237,clk_delay);
   and MGM_G292(MGM_W238,d_delay,MGM_W237);
   and MGM_G293(MGM_W239,psb_delay,MGM_W238);
   not MGM_G294(MGM_W240,si_delay);
   and MGM_G295(MGM_W241,MGM_W240,MGM_W239);
   not MGM_G296(MGM_W242,ssb_delay);
   and MGM_G297(ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W242,MGM_W241);
   not MGM_G298(MGM_W243,clk_delay);
   and MGM_G299(MGM_W244,d_delay,MGM_W243);
   and MGM_G300(MGM_W245,psb_delay,MGM_W244);
   not MGM_G301(MGM_W246,si_delay);
   and MGM_G302(MGM_W247,MGM_W246,MGM_W245);
   and MGM_G303(ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W247);
   not MGM_G304(MGM_W248,clk_delay);
   and MGM_G305(MGM_W249,d_delay,MGM_W248);
   and MGM_G306(MGM_W250,psb_delay,MGM_W249);
   and MGM_G307(MGM_W251,si_delay,MGM_W250);
   not MGM_G308(MGM_W252,ssb_delay);
   and MGM_G309(ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W252,MGM_W251);
   not MGM_G310(MGM_W253,clk_delay);
   and MGM_G311(MGM_W254,d_delay,MGM_W253);
   and MGM_G312(MGM_W255,psb_delay,MGM_W254);
   and MGM_G313(MGM_W256,si_delay,MGM_W255);
   and MGM_G314(ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W256);
   not MGM_G315(MGM_W257,d_delay);
   and MGM_G316(MGM_W258,MGM_W257,clk_delay);
   and MGM_G317(MGM_W259,psb_delay,MGM_W258);
   not MGM_G318(MGM_W260,si_delay);
   and MGM_G319(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G320(MGM_W262,ssb_delay);
   and MGM_G321(ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   not MGM_G322(MGM_W263,d_delay);
   and MGM_G323(MGM_W264,MGM_W263,clk_delay);
   and MGM_G324(MGM_W265,psb_delay,MGM_W264);
   not MGM_G325(MGM_W266,si_delay);
   and MGM_G326(MGM_W267,MGM_W266,MGM_W265);
   and MGM_G327(ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W267);
   not MGM_G328(MGM_W268,d_delay);
   and MGM_G329(MGM_W269,MGM_W268,clk_delay);
   and MGM_G330(MGM_W270,psb_delay,MGM_W269);
   and MGM_G331(MGM_W271,si_delay,MGM_W270);
   not MGM_G332(MGM_W272,ssb_delay);
   and MGM_G333(ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W272,MGM_W271);
   not MGM_G334(MGM_W273,d_delay);
   and MGM_G335(MGM_W274,MGM_W273,clk_delay);
   and MGM_G336(MGM_W275,psb_delay,MGM_W274);
   and MGM_G337(MGM_W276,si_delay,MGM_W275);
   and MGM_G338(ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W276);
   and MGM_G339(MGM_W277,d_delay,clk_delay);
   and MGM_G340(MGM_W278,psb_delay,MGM_W277);
   not MGM_G341(MGM_W279,si_delay);
   and MGM_G342(MGM_W280,MGM_W279,MGM_W278);
   not MGM_G343(MGM_W281,ssb_delay);
   and MGM_G344(ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W281,MGM_W280);
   and MGM_G345(MGM_W282,d_delay,clk_delay);
   and MGM_G346(MGM_W283,psb_delay,MGM_W282);
   not MGM_G347(MGM_W284,si_delay);
   and MGM_G348(MGM_W285,MGM_W284,MGM_W283);
   and MGM_G349(ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W285);
   and MGM_G350(MGM_W286,d_delay,clk_delay);
   and MGM_G351(MGM_W287,psb_delay,MGM_W286);
   and MGM_G352(MGM_W288,si_delay,MGM_W287);
   not MGM_G353(MGM_W289,ssb_delay);
   and MGM_G354(ENABLE_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W289,MGM_W288);
   and MGM_G355(MGM_W290,d_delay,clk_delay);
   and MGM_G356(MGM_W291,psb_delay,MGM_W290);
   and MGM_G357(MGM_W292,si_delay,MGM_W291);
   and MGM_G358(ENABLE_clk_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W292);
   not MGM_G359(MGM_W293,d_delay);
   and MGM_G360(MGM_W294,psb_delay,MGM_W293);
   and MGM_G361(MGM_W295,rb_delay,MGM_W294);
   not MGM_G362(MGM_W296,ssb_delay);
   and MGM_G363(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W296,MGM_W295);
   and MGM_G364(MGM_W297,psb_delay,d_delay);
   and MGM_G365(MGM_W298,rb_delay,MGM_W297);
   not MGM_G366(MGM_W299,ssb_delay);
   and MGM_G367(ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W299,MGM_W298);
   not MGM_G368(MGM_W300,d_delay);
   and MGM_G369(MGM_W301,psb_delay,MGM_W300);
   and MGM_G370(MGM_W302,rb_delay,MGM_W301);
   and MGM_G371(ENABLE_NOT_d_AND_psb_AND_rb_AND_si,si_delay,MGM_W302);
   and MGM_G372(MGM_W303,psb_delay,d_delay);
   and MGM_G373(MGM_W304,rb_delay,MGM_W303);
   not MGM_G374(MGM_W305,si_delay);
   and MGM_G375(ENABLE_d_AND_psb_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy00fah1n12x5( clk, d, o, psb, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00fah_func b15fqy00fah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00fah_func b15fqy00fah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00fah_func b15fqy00fah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00fah_func b15fqy00fah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(MGM_W2,rb_delay,MGM_W1);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   and MGM_G8(MGM_W7,psb_delay,MGM_W6);
   and MGM_G9(MGM_W8,rb_delay,MGM_W7);
   not MGM_G10(MGM_W9,si_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G12(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W10);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,psb_delay,MGM_W11);
   and MGM_G15(MGM_W13,rb_delay,MGM_W12);
   and MGM_G16(MGM_W14,si_delay,MGM_W13);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,psb_delay,MGM_W16);
   and MGM_G21(MGM_W18,rb_delay,MGM_W17);
   and MGM_G22(MGM_W19,si_delay,MGM_W18);
   and MGM_G23(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W19);
   and MGM_G24(MGM_W20,psb_delay,d_delay);
   and MGM_G25(MGM_W21,rb_delay,MGM_W20);
   not MGM_G26(MGM_W22,si_delay);
   and MGM_G27(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G28(MGM_W24,ssb_delay);
   and MGM_G29(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W24,MGM_W23);
   and MGM_G30(MGM_W25,psb_delay,d_delay);
   and MGM_G31(MGM_W26,rb_delay,MGM_W25);
   not MGM_G32(MGM_W27,si_delay);
   and MGM_G33(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G34(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W28);
   and MGM_G35(MGM_W29,psb_delay,d_delay);
   and MGM_G36(MGM_W30,rb_delay,MGM_W29);
   and MGM_G37(MGM_W31,si_delay,MGM_W30);
   not MGM_G38(MGM_W32,ssb_delay);
   and MGM_G39(ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W32,MGM_W31);
   and MGM_G40(MGM_W33,psb_delay,d_delay);
   and MGM_G41(MGM_W34,rb_delay,MGM_W33);
   and MGM_G42(MGM_W35,si_delay,MGM_W34);
   and MGM_G43(ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G44(MGM_W36,rb_delay,psb_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   and MGM_G47(ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W38);
   and MGM_G48(MGM_W39,rb_delay,psb_delay);
   and MGM_G49(MGM_W40,si_delay,MGM_W39);
   and MGM_G50(ENABLE_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G51(MGM_W41,d_delay);
   and MGM_G52(MGM_W42,rb_delay,MGM_W41);
   not MGM_G53(MGM_W43,si_delay);
   and MGM_G54(MGM_W44,MGM_W43,MGM_W42);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   not MGM_G57(MGM_W46,d_delay);
   and MGM_G58(MGM_W47,rb_delay,MGM_W46);
   not MGM_G59(MGM_W48,si_delay);
   and MGM_G60(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G61(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G62(MGM_W50,d_delay);
   and MGM_G63(MGM_W51,rb_delay,MGM_W50);
   and MGM_G64(MGM_W52,si_delay,MGM_W51);
   and MGM_G65(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G66(MGM_W53,rb_delay,d_delay);
   not MGM_G67(MGM_W54,si_delay);
   and MGM_G68(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G69(MGM_W56,ssb_delay);
   and MGM_G70(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   not MGM_G71(MGM_W57,clk_delay);
   not MGM_G72(MGM_W58,d_delay);
   and MGM_G73(MGM_W59,MGM_W58,MGM_W57);
   and MGM_G74(MGM_W60,rb_delay,MGM_W59);
   not MGM_G75(MGM_W61,si_delay);
   and MGM_G76(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G77(MGM_W63,ssb_delay);
   and MGM_G78(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G79(MGM_W64,clk_delay);
   not MGM_G80(MGM_W65,d_delay);
   and MGM_G81(MGM_W66,MGM_W65,MGM_W64);
   and MGM_G82(MGM_W67,rb_delay,MGM_W66);
   not MGM_G83(MGM_W68,si_delay);
   and MGM_G84(MGM_W69,MGM_W68,MGM_W67);
   and MGM_G85(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W69);
   not MGM_G86(MGM_W70,clk_delay);
   not MGM_G87(MGM_W71,d_delay);
   and MGM_G88(MGM_W72,MGM_W71,MGM_W70);
   and MGM_G89(MGM_W73,rb_delay,MGM_W72);
   and MGM_G90(MGM_W74,si_delay,MGM_W73);
   not MGM_G91(MGM_W75,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G93(MGM_W76,clk_delay);
   not MGM_G94(MGM_W77,d_delay);
   and MGM_G95(MGM_W78,MGM_W77,MGM_W76);
   and MGM_G96(MGM_W79,rb_delay,MGM_W78);
   and MGM_G97(MGM_W80,si_delay,MGM_W79);
   and MGM_G98(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W80);
   not MGM_G99(MGM_W81,clk_delay);
   and MGM_G100(MGM_W82,d_delay,MGM_W81);
   and MGM_G101(MGM_W83,rb_delay,MGM_W82);
   not MGM_G102(MGM_W84,si_delay);
   and MGM_G103(MGM_W85,MGM_W84,MGM_W83);
   not MGM_G104(MGM_W86,ssb_delay);
   and MGM_G105(ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W86,MGM_W85);
   not MGM_G106(MGM_W87,clk_delay);
   and MGM_G107(MGM_W88,d_delay,MGM_W87);
   and MGM_G108(MGM_W89,rb_delay,MGM_W88);
   not MGM_G109(MGM_W90,si_delay);
   and MGM_G110(MGM_W91,MGM_W90,MGM_W89);
   and MGM_G111(ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W91);
   not MGM_G112(MGM_W92,clk_delay);
   and MGM_G113(MGM_W93,d_delay,MGM_W92);
   and MGM_G114(MGM_W94,rb_delay,MGM_W93);
   and MGM_G115(MGM_W95,si_delay,MGM_W94);
   not MGM_G116(MGM_W96,ssb_delay);
   and MGM_G117(ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W96,MGM_W95);
   not MGM_G118(MGM_W97,clk_delay);
   and MGM_G119(MGM_W98,d_delay,MGM_W97);
   and MGM_G120(MGM_W99,rb_delay,MGM_W98);
   and MGM_G121(MGM_W100,si_delay,MGM_W99);
   and MGM_G122(ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W100);
   not MGM_G123(MGM_W101,d_delay);
   and MGM_G124(MGM_W102,MGM_W101,clk_delay);
   and MGM_G125(MGM_W103,rb_delay,MGM_W102);
   not MGM_G126(MGM_W104,si_delay);
   and MGM_G127(MGM_W105,MGM_W104,MGM_W103);
   not MGM_G128(MGM_W106,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W106,MGM_W105);
   not MGM_G130(MGM_W107,d_delay);
   and MGM_G131(MGM_W108,MGM_W107,clk_delay);
   and MGM_G132(MGM_W109,rb_delay,MGM_W108);
   not MGM_G133(MGM_W110,si_delay);
   and MGM_G134(MGM_W111,MGM_W110,MGM_W109);
   and MGM_G135(ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W111);
   not MGM_G136(MGM_W112,d_delay);
   and MGM_G137(MGM_W113,MGM_W112,clk_delay);
   and MGM_G138(MGM_W114,rb_delay,MGM_W113);
   and MGM_G139(MGM_W115,si_delay,MGM_W114);
   not MGM_G140(MGM_W116,ssb_delay);
   and MGM_G141(ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W116,MGM_W115);
   not MGM_G142(MGM_W117,d_delay);
   and MGM_G143(MGM_W118,MGM_W117,clk_delay);
   and MGM_G144(MGM_W119,rb_delay,MGM_W118);
   and MGM_G145(MGM_W120,si_delay,MGM_W119);
   and MGM_G146(ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W120);
   and MGM_G147(MGM_W121,d_delay,clk_delay);
   and MGM_G148(MGM_W122,rb_delay,MGM_W121);
   not MGM_G149(MGM_W123,si_delay);
   and MGM_G150(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G151(MGM_W125,ssb_delay);
   and MGM_G152(ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W125,MGM_W124);
   and MGM_G153(MGM_W126,d_delay,clk_delay);
   and MGM_G154(MGM_W127,rb_delay,MGM_W126);
   not MGM_G155(MGM_W128,si_delay);
   and MGM_G156(MGM_W129,MGM_W128,MGM_W127);
   and MGM_G157(ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W129);
   and MGM_G158(MGM_W130,d_delay,clk_delay);
   and MGM_G159(MGM_W131,rb_delay,MGM_W130);
   and MGM_G160(MGM_W132,si_delay,MGM_W131);
   not MGM_G161(MGM_W133,ssb_delay);
   and MGM_G162(ENABLE_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W133,MGM_W132);
   and MGM_G163(MGM_W134,d_delay,clk_delay);
   and MGM_G164(MGM_W135,rb_delay,MGM_W134);
   and MGM_G165(MGM_W136,si_delay,MGM_W135);
   and MGM_G166(ENABLE_clk_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W136);
   not MGM_G167(MGM_W137,clk_delay);
   not MGM_G168(MGM_W138,d_delay);
   and MGM_G169(MGM_W139,MGM_W138,MGM_W137);
   not MGM_G170(MGM_W140,si_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   not MGM_G172(MGM_W142,ssb_delay);
   and MGM_G173(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W142,MGM_W141);
   not MGM_G174(MGM_W143,clk_delay);
   not MGM_G175(MGM_W144,d_delay);
   and MGM_G176(MGM_W145,MGM_W144,MGM_W143);
   not MGM_G177(MGM_W146,si_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W147);
   not MGM_G180(MGM_W148,clk_delay);
   not MGM_G181(MGM_W149,d_delay);
   and MGM_G182(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G183(MGM_W151,si_delay,MGM_W150);
   not MGM_G184(MGM_W152,ssb_delay);
   and MGM_G185(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W153,clk_delay);
   not MGM_G187(MGM_W154,d_delay);
   and MGM_G188(MGM_W155,MGM_W154,MGM_W153);
   and MGM_G189(MGM_W156,si_delay,MGM_W155);
   and MGM_G190(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W156);
   not MGM_G191(MGM_W157,clk_delay);
   and MGM_G192(MGM_W158,d_delay,MGM_W157);
   not MGM_G193(MGM_W159,si_delay);
   and MGM_G194(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G195(MGM_W161,ssb_delay);
   and MGM_G196(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W161,MGM_W160);
   not MGM_G197(MGM_W162,clk_delay);
   and MGM_G198(MGM_W163,d_delay,MGM_W162);
   not MGM_G199(MGM_W164,si_delay);
   and MGM_G200(MGM_W165,MGM_W164,MGM_W163);
   and MGM_G201(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W165);
   not MGM_G202(MGM_W166,clk_delay);
   and MGM_G203(MGM_W167,d_delay,MGM_W166);
   and MGM_G204(MGM_W168,si_delay,MGM_W167);
   not MGM_G205(MGM_W169,ssb_delay);
   and MGM_G206(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W169,MGM_W168);
   not MGM_G207(MGM_W170,clk_delay);
   and MGM_G208(MGM_W171,d_delay,MGM_W170);
   and MGM_G209(MGM_W172,si_delay,MGM_W171);
   and MGM_G210(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W172);
   not MGM_G211(MGM_W173,d_delay);
   and MGM_G212(MGM_W174,MGM_W173,clk_delay);
   not MGM_G213(MGM_W175,si_delay);
   and MGM_G214(MGM_W176,MGM_W175,MGM_W174);
   not MGM_G215(MGM_W177,ssb_delay);
   and MGM_G216(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W177,MGM_W176);
   not MGM_G217(MGM_W178,d_delay);
   and MGM_G218(MGM_W179,MGM_W178,clk_delay);
   not MGM_G219(MGM_W180,si_delay);
   and MGM_G220(MGM_W181,MGM_W180,MGM_W179);
   and MGM_G221(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W181);
   not MGM_G222(MGM_W182,d_delay);
   and MGM_G223(MGM_W183,MGM_W182,clk_delay);
   and MGM_G224(MGM_W184,si_delay,MGM_W183);
   not MGM_G225(MGM_W185,ssb_delay);
   and MGM_G226(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W185,MGM_W184);
   not MGM_G227(MGM_W186,d_delay);
   and MGM_G228(MGM_W187,MGM_W186,clk_delay);
   and MGM_G229(MGM_W188,si_delay,MGM_W187);
   and MGM_G230(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W188);
   and MGM_G231(MGM_W189,d_delay,clk_delay);
   not MGM_G232(MGM_W190,si_delay);
   and MGM_G233(MGM_W191,MGM_W190,MGM_W189);
   not MGM_G234(MGM_W192,ssb_delay);
   and MGM_G235(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W192,MGM_W191);
   and MGM_G236(MGM_W193,d_delay,clk_delay);
   not MGM_G237(MGM_W194,si_delay);
   and MGM_G238(MGM_W195,MGM_W194,MGM_W193);
   and MGM_G239(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W195);
   and MGM_G240(MGM_W196,d_delay,clk_delay);
   and MGM_G241(MGM_W197,si_delay,MGM_W196);
   not MGM_G242(MGM_W198,ssb_delay);
   and MGM_G243(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W198,MGM_W197);
   and MGM_G244(MGM_W199,d_delay,clk_delay);
   and MGM_G245(MGM_W200,si_delay,MGM_W199);
   and MGM_G246(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W200);
   not MGM_G247(MGM_W201,d_delay);
   and MGM_G248(MGM_W202,psb_delay,MGM_W201);
   and MGM_G249(MGM_W203,si_delay,MGM_W202);
   not MGM_G250(MGM_W204,ssb_delay);
   and MGM_G251(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W204,MGM_W203);
   and MGM_G252(MGM_W205,psb_delay,d_delay);
   not MGM_G253(MGM_W206,si_delay);
   and MGM_G254(MGM_W207,MGM_W206,MGM_W205);
   and MGM_G255(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W207);
   and MGM_G256(MGM_W208,psb_delay,d_delay);
   and MGM_G257(MGM_W209,si_delay,MGM_W208);
   not MGM_G258(MGM_W210,ssb_delay);
   and MGM_G259(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W210,MGM_W209);
   and MGM_G260(MGM_W211,psb_delay,d_delay);
   and MGM_G261(MGM_W212,si_delay,MGM_W211);
   and MGM_G262(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W212);
   not MGM_G263(MGM_W213,clk_delay);
   not MGM_G264(MGM_W214,d_delay);
   and MGM_G265(MGM_W215,MGM_W214,MGM_W213);
   and MGM_G266(MGM_W216,psb_delay,MGM_W215);
   not MGM_G267(MGM_W217,si_delay);
   and MGM_G268(MGM_W218,MGM_W217,MGM_W216);
   not MGM_G269(MGM_W219,ssb_delay);
   and MGM_G270(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W219,MGM_W218);
   not MGM_G271(MGM_W220,clk_delay);
   not MGM_G272(MGM_W221,d_delay);
   and MGM_G273(MGM_W222,MGM_W221,MGM_W220);
   and MGM_G274(MGM_W223,psb_delay,MGM_W222);
   not MGM_G275(MGM_W224,si_delay);
   and MGM_G276(MGM_W225,MGM_W224,MGM_W223);
   and MGM_G277(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W225);
   not MGM_G278(MGM_W226,clk_delay);
   not MGM_G279(MGM_W227,d_delay);
   and MGM_G280(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G281(MGM_W229,psb_delay,MGM_W228);
   and MGM_G282(MGM_W230,si_delay,MGM_W229);
   not MGM_G283(MGM_W231,ssb_delay);
   and MGM_G284(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W231,MGM_W230);
   not MGM_G285(MGM_W232,clk_delay);
   not MGM_G286(MGM_W233,d_delay);
   and MGM_G287(MGM_W234,MGM_W233,MGM_W232);
   and MGM_G288(MGM_W235,psb_delay,MGM_W234);
   and MGM_G289(MGM_W236,si_delay,MGM_W235);
   and MGM_G290(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W236);
   not MGM_G291(MGM_W237,clk_delay);
   and MGM_G292(MGM_W238,d_delay,MGM_W237);
   and MGM_G293(MGM_W239,psb_delay,MGM_W238);
   not MGM_G294(MGM_W240,si_delay);
   and MGM_G295(MGM_W241,MGM_W240,MGM_W239);
   not MGM_G296(MGM_W242,ssb_delay);
   and MGM_G297(ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W242,MGM_W241);
   not MGM_G298(MGM_W243,clk_delay);
   and MGM_G299(MGM_W244,d_delay,MGM_W243);
   and MGM_G300(MGM_W245,psb_delay,MGM_W244);
   not MGM_G301(MGM_W246,si_delay);
   and MGM_G302(MGM_W247,MGM_W246,MGM_W245);
   and MGM_G303(ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W247);
   not MGM_G304(MGM_W248,clk_delay);
   and MGM_G305(MGM_W249,d_delay,MGM_W248);
   and MGM_G306(MGM_W250,psb_delay,MGM_W249);
   and MGM_G307(MGM_W251,si_delay,MGM_W250);
   not MGM_G308(MGM_W252,ssb_delay);
   and MGM_G309(ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W252,MGM_W251);
   not MGM_G310(MGM_W253,clk_delay);
   and MGM_G311(MGM_W254,d_delay,MGM_W253);
   and MGM_G312(MGM_W255,psb_delay,MGM_W254);
   and MGM_G313(MGM_W256,si_delay,MGM_W255);
   and MGM_G314(ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W256);
   not MGM_G315(MGM_W257,d_delay);
   and MGM_G316(MGM_W258,MGM_W257,clk_delay);
   and MGM_G317(MGM_W259,psb_delay,MGM_W258);
   not MGM_G318(MGM_W260,si_delay);
   and MGM_G319(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G320(MGM_W262,ssb_delay);
   and MGM_G321(ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   not MGM_G322(MGM_W263,d_delay);
   and MGM_G323(MGM_W264,MGM_W263,clk_delay);
   and MGM_G324(MGM_W265,psb_delay,MGM_W264);
   not MGM_G325(MGM_W266,si_delay);
   and MGM_G326(MGM_W267,MGM_W266,MGM_W265);
   and MGM_G327(ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W267);
   not MGM_G328(MGM_W268,d_delay);
   and MGM_G329(MGM_W269,MGM_W268,clk_delay);
   and MGM_G330(MGM_W270,psb_delay,MGM_W269);
   and MGM_G331(MGM_W271,si_delay,MGM_W270);
   not MGM_G332(MGM_W272,ssb_delay);
   and MGM_G333(ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W272,MGM_W271);
   not MGM_G334(MGM_W273,d_delay);
   and MGM_G335(MGM_W274,MGM_W273,clk_delay);
   and MGM_G336(MGM_W275,psb_delay,MGM_W274);
   and MGM_G337(MGM_W276,si_delay,MGM_W275);
   and MGM_G338(ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W276);
   and MGM_G339(MGM_W277,d_delay,clk_delay);
   and MGM_G340(MGM_W278,psb_delay,MGM_W277);
   not MGM_G341(MGM_W279,si_delay);
   and MGM_G342(MGM_W280,MGM_W279,MGM_W278);
   not MGM_G343(MGM_W281,ssb_delay);
   and MGM_G344(ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W281,MGM_W280);
   and MGM_G345(MGM_W282,d_delay,clk_delay);
   and MGM_G346(MGM_W283,psb_delay,MGM_W282);
   not MGM_G347(MGM_W284,si_delay);
   and MGM_G348(MGM_W285,MGM_W284,MGM_W283);
   and MGM_G349(ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W285);
   and MGM_G350(MGM_W286,d_delay,clk_delay);
   and MGM_G351(MGM_W287,psb_delay,MGM_W286);
   and MGM_G352(MGM_W288,si_delay,MGM_W287);
   not MGM_G353(MGM_W289,ssb_delay);
   and MGM_G354(ENABLE_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W289,MGM_W288);
   and MGM_G355(MGM_W290,d_delay,clk_delay);
   and MGM_G356(MGM_W291,psb_delay,MGM_W290);
   and MGM_G357(MGM_W292,si_delay,MGM_W291);
   and MGM_G358(ENABLE_clk_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W292);
   not MGM_G359(MGM_W293,d_delay);
   and MGM_G360(MGM_W294,psb_delay,MGM_W293);
   and MGM_G361(MGM_W295,rb_delay,MGM_W294);
   not MGM_G362(MGM_W296,ssb_delay);
   and MGM_G363(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W296,MGM_W295);
   and MGM_G364(MGM_W297,psb_delay,d_delay);
   and MGM_G365(MGM_W298,rb_delay,MGM_W297);
   not MGM_G366(MGM_W299,ssb_delay);
   and MGM_G367(ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W299,MGM_W298);
   not MGM_G368(MGM_W300,d_delay);
   and MGM_G369(MGM_W301,psb_delay,MGM_W300);
   and MGM_G370(MGM_W302,rb_delay,MGM_W301);
   and MGM_G371(ENABLE_NOT_d_AND_psb_AND_rb_AND_si,si_delay,MGM_W302);
   and MGM_G372(MGM_W303,psb_delay,d_delay);
   and MGM_G373(MGM_W304,rb_delay,MGM_W303);
   not MGM_G374(MGM_W305,si_delay);
   and MGM_G375(ENABLE_d_AND_psb_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy00fah1n16x5( clk, d, o, psb, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00fah_func b15fqy00fah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00fah_func b15fqy00fah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy00fah_func b15fqy00fah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy00fah_func b15fqy00fah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(MGM_W2,rb_delay,MGM_W1);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   and MGM_G8(MGM_W7,psb_delay,MGM_W6);
   and MGM_G9(MGM_W8,rb_delay,MGM_W7);
   not MGM_G10(MGM_W9,si_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G12(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W10);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,psb_delay,MGM_W11);
   and MGM_G15(MGM_W13,rb_delay,MGM_W12);
   and MGM_G16(MGM_W14,si_delay,MGM_W13);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,psb_delay,MGM_W16);
   and MGM_G21(MGM_W18,rb_delay,MGM_W17);
   and MGM_G22(MGM_W19,si_delay,MGM_W18);
   and MGM_G23(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W19);
   and MGM_G24(MGM_W20,psb_delay,d_delay);
   and MGM_G25(MGM_W21,rb_delay,MGM_W20);
   not MGM_G26(MGM_W22,si_delay);
   and MGM_G27(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G28(MGM_W24,ssb_delay);
   and MGM_G29(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W24,MGM_W23);
   and MGM_G30(MGM_W25,psb_delay,d_delay);
   and MGM_G31(MGM_W26,rb_delay,MGM_W25);
   not MGM_G32(MGM_W27,si_delay);
   and MGM_G33(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G34(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W28);
   and MGM_G35(MGM_W29,psb_delay,d_delay);
   and MGM_G36(MGM_W30,rb_delay,MGM_W29);
   and MGM_G37(MGM_W31,si_delay,MGM_W30);
   not MGM_G38(MGM_W32,ssb_delay);
   and MGM_G39(ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W32,MGM_W31);
   and MGM_G40(MGM_W33,psb_delay,d_delay);
   and MGM_G41(MGM_W34,rb_delay,MGM_W33);
   and MGM_G42(MGM_W35,si_delay,MGM_W34);
   and MGM_G43(ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G44(MGM_W36,rb_delay,psb_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   and MGM_G47(ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W38);
   and MGM_G48(MGM_W39,rb_delay,psb_delay);
   and MGM_G49(MGM_W40,si_delay,MGM_W39);
   and MGM_G50(ENABLE_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G51(MGM_W41,d_delay);
   and MGM_G52(MGM_W42,rb_delay,MGM_W41);
   not MGM_G53(MGM_W43,si_delay);
   and MGM_G54(MGM_W44,MGM_W43,MGM_W42);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   not MGM_G57(MGM_W46,d_delay);
   and MGM_G58(MGM_W47,rb_delay,MGM_W46);
   not MGM_G59(MGM_W48,si_delay);
   and MGM_G60(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G61(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G62(MGM_W50,d_delay);
   and MGM_G63(MGM_W51,rb_delay,MGM_W50);
   and MGM_G64(MGM_W52,si_delay,MGM_W51);
   and MGM_G65(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G66(MGM_W53,rb_delay,d_delay);
   not MGM_G67(MGM_W54,si_delay);
   and MGM_G68(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G69(MGM_W56,ssb_delay);
   and MGM_G70(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   not MGM_G71(MGM_W57,clk_delay);
   not MGM_G72(MGM_W58,d_delay);
   and MGM_G73(MGM_W59,MGM_W58,MGM_W57);
   and MGM_G74(MGM_W60,rb_delay,MGM_W59);
   not MGM_G75(MGM_W61,si_delay);
   and MGM_G76(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G77(MGM_W63,ssb_delay);
   and MGM_G78(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G79(MGM_W64,clk_delay);
   not MGM_G80(MGM_W65,d_delay);
   and MGM_G81(MGM_W66,MGM_W65,MGM_W64);
   and MGM_G82(MGM_W67,rb_delay,MGM_W66);
   not MGM_G83(MGM_W68,si_delay);
   and MGM_G84(MGM_W69,MGM_W68,MGM_W67);
   and MGM_G85(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W69);
   not MGM_G86(MGM_W70,clk_delay);
   not MGM_G87(MGM_W71,d_delay);
   and MGM_G88(MGM_W72,MGM_W71,MGM_W70);
   and MGM_G89(MGM_W73,rb_delay,MGM_W72);
   and MGM_G90(MGM_W74,si_delay,MGM_W73);
   not MGM_G91(MGM_W75,ssb_delay);
   and MGM_G92(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G93(MGM_W76,clk_delay);
   not MGM_G94(MGM_W77,d_delay);
   and MGM_G95(MGM_W78,MGM_W77,MGM_W76);
   and MGM_G96(MGM_W79,rb_delay,MGM_W78);
   and MGM_G97(MGM_W80,si_delay,MGM_W79);
   and MGM_G98(ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W80);
   not MGM_G99(MGM_W81,clk_delay);
   and MGM_G100(MGM_W82,d_delay,MGM_W81);
   and MGM_G101(MGM_W83,rb_delay,MGM_W82);
   not MGM_G102(MGM_W84,si_delay);
   and MGM_G103(MGM_W85,MGM_W84,MGM_W83);
   not MGM_G104(MGM_W86,ssb_delay);
   and MGM_G105(ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W86,MGM_W85);
   not MGM_G106(MGM_W87,clk_delay);
   and MGM_G107(MGM_W88,d_delay,MGM_W87);
   and MGM_G108(MGM_W89,rb_delay,MGM_W88);
   not MGM_G109(MGM_W90,si_delay);
   and MGM_G110(MGM_W91,MGM_W90,MGM_W89);
   and MGM_G111(ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W91);
   not MGM_G112(MGM_W92,clk_delay);
   and MGM_G113(MGM_W93,d_delay,MGM_W92);
   and MGM_G114(MGM_W94,rb_delay,MGM_W93);
   and MGM_G115(MGM_W95,si_delay,MGM_W94);
   not MGM_G116(MGM_W96,ssb_delay);
   and MGM_G117(ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W96,MGM_W95);
   not MGM_G118(MGM_W97,clk_delay);
   and MGM_G119(MGM_W98,d_delay,MGM_W97);
   and MGM_G120(MGM_W99,rb_delay,MGM_W98);
   and MGM_G121(MGM_W100,si_delay,MGM_W99);
   and MGM_G122(ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W100);
   not MGM_G123(MGM_W101,d_delay);
   and MGM_G124(MGM_W102,MGM_W101,clk_delay);
   and MGM_G125(MGM_W103,rb_delay,MGM_W102);
   not MGM_G126(MGM_W104,si_delay);
   and MGM_G127(MGM_W105,MGM_W104,MGM_W103);
   not MGM_G128(MGM_W106,ssb_delay);
   and MGM_G129(ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W106,MGM_W105);
   not MGM_G130(MGM_W107,d_delay);
   and MGM_G131(MGM_W108,MGM_W107,clk_delay);
   and MGM_G132(MGM_W109,rb_delay,MGM_W108);
   not MGM_G133(MGM_W110,si_delay);
   and MGM_G134(MGM_W111,MGM_W110,MGM_W109);
   and MGM_G135(ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W111);
   not MGM_G136(MGM_W112,d_delay);
   and MGM_G137(MGM_W113,MGM_W112,clk_delay);
   and MGM_G138(MGM_W114,rb_delay,MGM_W113);
   and MGM_G139(MGM_W115,si_delay,MGM_W114);
   not MGM_G140(MGM_W116,ssb_delay);
   and MGM_G141(ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W116,MGM_W115);
   not MGM_G142(MGM_W117,d_delay);
   and MGM_G143(MGM_W118,MGM_W117,clk_delay);
   and MGM_G144(MGM_W119,rb_delay,MGM_W118);
   and MGM_G145(MGM_W120,si_delay,MGM_W119);
   and MGM_G146(ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W120);
   and MGM_G147(MGM_W121,d_delay,clk_delay);
   and MGM_G148(MGM_W122,rb_delay,MGM_W121);
   not MGM_G149(MGM_W123,si_delay);
   and MGM_G150(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G151(MGM_W125,ssb_delay);
   and MGM_G152(ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W125,MGM_W124);
   and MGM_G153(MGM_W126,d_delay,clk_delay);
   and MGM_G154(MGM_W127,rb_delay,MGM_W126);
   not MGM_G155(MGM_W128,si_delay);
   and MGM_G156(MGM_W129,MGM_W128,MGM_W127);
   and MGM_G157(ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W129);
   and MGM_G158(MGM_W130,d_delay,clk_delay);
   and MGM_G159(MGM_W131,rb_delay,MGM_W130);
   and MGM_G160(MGM_W132,si_delay,MGM_W131);
   not MGM_G161(MGM_W133,ssb_delay);
   and MGM_G162(ENABLE_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W133,MGM_W132);
   and MGM_G163(MGM_W134,d_delay,clk_delay);
   and MGM_G164(MGM_W135,rb_delay,MGM_W134);
   and MGM_G165(MGM_W136,si_delay,MGM_W135);
   and MGM_G166(ENABLE_clk_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W136);
   not MGM_G167(MGM_W137,clk_delay);
   not MGM_G168(MGM_W138,d_delay);
   and MGM_G169(MGM_W139,MGM_W138,MGM_W137);
   not MGM_G170(MGM_W140,si_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   not MGM_G172(MGM_W142,ssb_delay);
   and MGM_G173(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W142,MGM_W141);
   not MGM_G174(MGM_W143,clk_delay);
   not MGM_G175(MGM_W144,d_delay);
   and MGM_G176(MGM_W145,MGM_W144,MGM_W143);
   not MGM_G177(MGM_W146,si_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W147);
   not MGM_G180(MGM_W148,clk_delay);
   not MGM_G181(MGM_W149,d_delay);
   and MGM_G182(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G183(MGM_W151,si_delay,MGM_W150);
   not MGM_G184(MGM_W152,ssb_delay);
   and MGM_G185(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W153,clk_delay);
   not MGM_G187(MGM_W154,d_delay);
   and MGM_G188(MGM_W155,MGM_W154,MGM_W153);
   and MGM_G189(MGM_W156,si_delay,MGM_W155);
   and MGM_G190(ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W156);
   not MGM_G191(MGM_W157,clk_delay);
   and MGM_G192(MGM_W158,d_delay,MGM_W157);
   not MGM_G193(MGM_W159,si_delay);
   and MGM_G194(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G195(MGM_W161,ssb_delay);
   and MGM_G196(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W161,MGM_W160);
   not MGM_G197(MGM_W162,clk_delay);
   and MGM_G198(MGM_W163,d_delay,MGM_W162);
   not MGM_G199(MGM_W164,si_delay);
   and MGM_G200(MGM_W165,MGM_W164,MGM_W163);
   and MGM_G201(ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W165);
   not MGM_G202(MGM_W166,clk_delay);
   and MGM_G203(MGM_W167,d_delay,MGM_W166);
   and MGM_G204(MGM_W168,si_delay,MGM_W167);
   not MGM_G205(MGM_W169,ssb_delay);
   and MGM_G206(ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W169,MGM_W168);
   not MGM_G207(MGM_W170,clk_delay);
   and MGM_G208(MGM_W171,d_delay,MGM_W170);
   and MGM_G209(MGM_W172,si_delay,MGM_W171);
   and MGM_G210(ENABLE_NOT_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W172);
   not MGM_G211(MGM_W173,d_delay);
   and MGM_G212(MGM_W174,MGM_W173,clk_delay);
   not MGM_G213(MGM_W175,si_delay);
   and MGM_G214(MGM_W176,MGM_W175,MGM_W174);
   not MGM_G215(MGM_W177,ssb_delay);
   and MGM_G216(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W177,MGM_W176);
   not MGM_G217(MGM_W178,d_delay);
   and MGM_G218(MGM_W179,MGM_W178,clk_delay);
   not MGM_G219(MGM_W180,si_delay);
   and MGM_G220(MGM_W181,MGM_W180,MGM_W179);
   and MGM_G221(ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W181);
   not MGM_G222(MGM_W182,d_delay);
   and MGM_G223(MGM_W183,MGM_W182,clk_delay);
   and MGM_G224(MGM_W184,si_delay,MGM_W183);
   not MGM_G225(MGM_W185,ssb_delay);
   and MGM_G226(ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W185,MGM_W184);
   not MGM_G227(MGM_W186,d_delay);
   and MGM_G228(MGM_W187,MGM_W186,clk_delay);
   and MGM_G229(MGM_W188,si_delay,MGM_W187);
   and MGM_G230(ENABLE_clk_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W188);
   and MGM_G231(MGM_W189,d_delay,clk_delay);
   not MGM_G232(MGM_W190,si_delay);
   and MGM_G233(MGM_W191,MGM_W190,MGM_W189);
   not MGM_G234(MGM_W192,ssb_delay);
   and MGM_G235(ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W192,MGM_W191);
   and MGM_G236(MGM_W193,d_delay,clk_delay);
   not MGM_G237(MGM_W194,si_delay);
   and MGM_G238(MGM_W195,MGM_W194,MGM_W193);
   and MGM_G239(ENABLE_clk_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W195);
   and MGM_G240(MGM_W196,d_delay,clk_delay);
   and MGM_G241(MGM_W197,si_delay,MGM_W196);
   not MGM_G242(MGM_W198,ssb_delay);
   and MGM_G243(ENABLE_clk_AND_d_AND_si_AND_NOT_ssb,MGM_W198,MGM_W197);
   and MGM_G244(MGM_W199,d_delay,clk_delay);
   and MGM_G245(MGM_W200,si_delay,MGM_W199);
   and MGM_G246(ENABLE_clk_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W200);
   not MGM_G247(MGM_W201,d_delay);
   and MGM_G248(MGM_W202,psb_delay,MGM_W201);
   and MGM_G249(MGM_W203,si_delay,MGM_W202);
   not MGM_G250(MGM_W204,ssb_delay);
   and MGM_G251(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W204,MGM_W203);
   and MGM_G252(MGM_W205,psb_delay,d_delay);
   not MGM_G253(MGM_W206,si_delay);
   and MGM_G254(MGM_W207,MGM_W206,MGM_W205);
   and MGM_G255(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W207);
   and MGM_G256(MGM_W208,psb_delay,d_delay);
   and MGM_G257(MGM_W209,si_delay,MGM_W208);
   not MGM_G258(MGM_W210,ssb_delay);
   and MGM_G259(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W210,MGM_W209);
   and MGM_G260(MGM_W211,psb_delay,d_delay);
   and MGM_G261(MGM_W212,si_delay,MGM_W211);
   and MGM_G262(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W212);
   not MGM_G263(MGM_W213,clk_delay);
   not MGM_G264(MGM_W214,d_delay);
   and MGM_G265(MGM_W215,MGM_W214,MGM_W213);
   and MGM_G266(MGM_W216,psb_delay,MGM_W215);
   not MGM_G267(MGM_W217,si_delay);
   and MGM_G268(MGM_W218,MGM_W217,MGM_W216);
   not MGM_G269(MGM_W219,ssb_delay);
   and MGM_G270(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W219,MGM_W218);
   not MGM_G271(MGM_W220,clk_delay);
   not MGM_G272(MGM_W221,d_delay);
   and MGM_G273(MGM_W222,MGM_W221,MGM_W220);
   and MGM_G274(MGM_W223,psb_delay,MGM_W222);
   not MGM_G275(MGM_W224,si_delay);
   and MGM_G276(MGM_W225,MGM_W224,MGM_W223);
   and MGM_G277(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W225);
   not MGM_G278(MGM_W226,clk_delay);
   not MGM_G279(MGM_W227,d_delay);
   and MGM_G280(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G281(MGM_W229,psb_delay,MGM_W228);
   and MGM_G282(MGM_W230,si_delay,MGM_W229);
   not MGM_G283(MGM_W231,ssb_delay);
   and MGM_G284(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W231,MGM_W230);
   not MGM_G285(MGM_W232,clk_delay);
   not MGM_G286(MGM_W233,d_delay);
   and MGM_G287(MGM_W234,MGM_W233,MGM_W232);
   and MGM_G288(MGM_W235,psb_delay,MGM_W234);
   and MGM_G289(MGM_W236,si_delay,MGM_W235);
   and MGM_G290(ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W236);
   not MGM_G291(MGM_W237,clk_delay);
   and MGM_G292(MGM_W238,d_delay,MGM_W237);
   and MGM_G293(MGM_W239,psb_delay,MGM_W238);
   not MGM_G294(MGM_W240,si_delay);
   and MGM_G295(MGM_W241,MGM_W240,MGM_W239);
   not MGM_G296(MGM_W242,ssb_delay);
   and MGM_G297(ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W242,MGM_W241);
   not MGM_G298(MGM_W243,clk_delay);
   and MGM_G299(MGM_W244,d_delay,MGM_W243);
   and MGM_G300(MGM_W245,psb_delay,MGM_W244);
   not MGM_G301(MGM_W246,si_delay);
   and MGM_G302(MGM_W247,MGM_W246,MGM_W245);
   and MGM_G303(ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W247);
   not MGM_G304(MGM_W248,clk_delay);
   and MGM_G305(MGM_W249,d_delay,MGM_W248);
   and MGM_G306(MGM_W250,psb_delay,MGM_W249);
   and MGM_G307(MGM_W251,si_delay,MGM_W250);
   not MGM_G308(MGM_W252,ssb_delay);
   and MGM_G309(ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W252,MGM_W251);
   not MGM_G310(MGM_W253,clk_delay);
   and MGM_G311(MGM_W254,d_delay,MGM_W253);
   and MGM_G312(MGM_W255,psb_delay,MGM_W254);
   and MGM_G313(MGM_W256,si_delay,MGM_W255);
   and MGM_G314(ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W256);
   not MGM_G315(MGM_W257,d_delay);
   and MGM_G316(MGM_W258,MGM_W257,clk_delay);
   and MGM_G317(MGM_W259,psb_delay,MGM_W258);
   not MGM_G318(MGM_W260,si_delay);
   and MGM_G319(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G320(MGM_W262,ssb_delay);
   and MGM_G321(ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   not MGM_G322(MGM_W263,d_delay);
   and MGM_G323(MGM_W264,MGM_W263,clk_delay);
   and MGM_G324(MGM_W265,psb_delay,MGM_W264);
   not MGM_G325(MGM_W266,si_delay);
   and MGM_G326(MGM_W267,MGM_W266,MGM_W265);
   and MGM_G327(ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W267);
   not MGM_G328(MGM_W268,d_delay);
   and MGM_G329(MGM_W269,MGM_W268,clk_delay);
   and MGM_G330(MGM_W270,psb_delay,MGM_W269);
   and MGM_G331(MGM_W271,si_delay,MGM_W270);
   not MGM_G332(MGM_W272,ssb_delay);
   and MGM_G333(ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W272,MGM_W271);
   not MGM_G334(MGM_W273,d_delay);
   and MGM_G335(MGM_W274,MGM_W273,clk_delay);
   and MGM_G336(MGM_W275,psb_delay,MGM_W274);
   and MGM_G337(MGM_W276,si_delay,MGM_W275);
   and MGM_G338(ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W276);
   and MGM_G339(MGM_W277,d_delay,clk_delay);
   and MGM_G340(MGM_W278,psb_delay,MGM_W277);
   not MGM_G341(MGM_W279,si_delay);
   and MGM_G342(MGM_W280,MGM_W279,MGM_W278);
   not MGM_G343(MGM_W281,ssb_delay);
   and MGM_G344(ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W281,MGM_W280);
   and MGM_G345(MGM_W282,d_delay,clk_delay);
   and MGM_G346(MGM_W283,psb_delay,MGM_W282);
   not MGM_G347(MGM_W284,si_delay);
   and MGM_G348(MGM_W285,MGM_W284,MGM_W283);
   and MGM_G349(ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W285);
   and MGM_G350(MGM_W286,d_delay,clk_delay);
   and MGM_G351(MGM_W287,psb_delay,MGM_W286);
   and MGM_G352(MGM_W288,si_delay,MGM_W287);
   not MGM_G353(MGM_W289,ssb_delay);
   and MGM_G354(ENABLE_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W289,MGM_W288);
   and MGM_G355(MGM_W290,d_delay,clk_delay);
   and MGM_G356(MGM_W291,psb_delay,MGM_W290);
   and MGM_G357(MGM_W292,si_delay,MGM_W291);
   and MGM_G358(ENABLE_clk_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W292);
   not MGM_G359(MGM_W293,d_delay);
   and MGM_G360(MGM_W294,psb_delay,MGM_W293);
   and MGM_G361(MGM_W295,rb_delay,MGM_W294);
   not MGM_G362(MGM_W296,ssb_delay);
   and MGM_G363(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W296,MGM_W295);
   and MGM_G364(MGM_W297,psb_delay,d_delay);
   and MGM_G365(MGM_W298,rb_delay,MGM_W297);
   not MGM_G366(MGM_W299,ssb_delay);
   and MGM_G367(ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W299,MGM_W298);
   not MGM_G368(MGM_W300,d_delay);
   and MGM_G369(MGM_W301,psb_delay,MGM_W300);
   and MGM_G370(MGM_W302,rb_delay,MGM_W301);
   and MGM_G371(ENABLE_NOT_d_AND_psb_AND_rb_AND_si,si_delay,MGM_W302);
   and MGM_G372(MGM_W303,psb_delay,d_delay);
   and MGM_G373(MGM_W304,rb_delay,MGM_W303);
   not MGM_G374(MGM_W305,si_delay);
   and MGM_G375(ENABLE_d_AND_psb_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      // recrem psb-clk-posedge
      $recrem(posedge psb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clk_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clk_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fqy043ah_func( clk, d, den, o, rb, si, ssb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb, si, ssb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, int2, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_fpn040ah_6( int1, IQ, d, den, vcc, vssx );
   INTCseq_fdw003ah_5( int2, int1, si, ssb, vcc, vssx );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_cdiar2ah_0( MGM_D0, int2 );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_fpn040ah_6( int1, IQ, d, den );
   INTCseq_fdw003ah_5( int2, int1, si, ssb );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fqy043ah1n02x5( clk, d, den, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy043ah_func b15fqy043ah1n02x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy043ah_func b15fqy043ah1n02x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy043ah_func b15fqy043ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy043ah_func b15fqy043ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,den_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   and MGM_G3(MGM_W3,rb_delay,MGM_W2);
   not MGM_G4(MGM_W4,si_delay);
   and MGM_G5(MGM_W5,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W6,ssb_delay);
   and MGM_G7(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W6,MGM_W5);
   not MGM_G8(MGM_W7,d_delay);
   not MGM_G9(MGM_W8,den_delay);
   and MGM_G10(MGM_W9,MGM_W8,MGM_W7);
   and MGM_G11(MGM_W10,rb_delay,MGM_W9);
   and MGM_G12(MGM_W11,si_delay,MGM_W10);
   not MGM_G13(MGM_W12,ssb_delay);
   and MGM_G14(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G15(MGM_W13,d_delay);
   and MGM_G16(MGM_W14,den_delay,MGM_W13);
   and MGM_G17(MGM_W15,rb_delay,MGM_W14);
   not MGM_G18(MGM_W16,si_delay);
   and MGM_G19(MGM_W17,MGM_W16,MGM_W15);
   not MGM_G20(MGM_W18,ssb_delay);
   and MGM_G21(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   not MGM_G22(MGM_W19,d_delay);
   and MGM_G23(MGM_W20,den_delay,MGM_W19);
   and MGM_G24(MGM_W21,rb_delay,MGM_W20);
   not MGM_G25(MGM_W22,si_delay);
   and MGM_G26(MGM_W23,MGM_W22,MGM_W21);
   and MGM_G27(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W23);
   not MGM_G28(MGM_W24,d_delay);
   and MGM_G29(MGM_W25,den_delay,MGM_W24);
   and MGM_G30(MGM_W26,rb_delay,MGM_W25);
   and MGM_G31(MGM_W27,si_delay,MGM_W26);
   not MGM_G32(MGM_W28,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W28,MGM_W27);
   not MGM_G34(MGM_W29,d_delay);
   and MGM_G35(MGM_W30,den_delay,MGM_W29);
   and MGM_G36(MGM_W31,rb_delay,MGM_W30);
   and MGM_G37(MGM_W32,si_delay,MGM_W31);
   and MGM_G38(ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W32);
   not MGM_G39(MGM_W33,den_delay);
   and MGM_G40(MGM_W34,MGM_W33,d_delay);
   and MGM_G41(MGM_W35,rb_delay,MGM_W34);
   not MGM_G42(MGM_W36,si_delay);
   and MGM_G43(MGM_W37,MGM_W36,MGM_W35);
   not MGM_G44(MGM_W38,ssb_delay);
   and MGM_G45(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W38,MGM_W37);
   not MGM_G46(MGM_W39,den_delay);
   and MGM_G47(MGM_W40,MGM_W39,d_delay);
   and MGM_G48(MGM_W41,rb_delay,MGM_W40);
   and MGM_G49(MGM_W42,si_delay,MGM_W41);
   not MGM_G50(MGM_W43,ssb_delay);
   and MGM_G51(ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W43,MGM_W42);
   and MGM_G52(MGM_W44,den_delay,d_delay);
   and MGM_G53(MGM_W45,rb_delay,MGM_W44);
   not MGM_G54(MGM_W46,si_delay);
   and MGM_G55(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G56(MGM_W48,ssb_delay);
   and MGM_G57(ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   and MGM_G58(MGM_W49,den_delay,d_delay);
   and MGM_G59(MGM_W50,rb_delay,MGM_W49);
   not MGM_G60(MGM_W51,si_delay);
   and MGM_G61(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G62(ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G63(MGM_W53,den_delay,d_delay);
   and MGM_G64(MGM_W54,rb_delay,MGM_W53);
   and MGM_G65(MGM_W55,si_delay,MGM_W54);
   not MGM_G66(MGM_W56,ssb_delay);
   and MGM_G67(ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   and MGM_G68(MGM_W57,den_delay,d_delay);
   and MGM_G69(MGM_W58,rb_delay,MGM_W57);
   and MGM_G70(MGM_W59,si_delay,MGM_W58);
   and MGM_G71(ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W59);
   and MGM_G72(MGM_W60,rb_delay,den_delay);
   not MGM_G73(MGM_W61,si_delay);
   and MGM_G74(MGM_W62,MGM_W61,MGM_W60);
   and MGM_G75(ENABLE_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W62);
   and MGM_G76(MGM_W63,rb_delay,den_delay);
   and MGM_G77(MGM_W64,si_delay,MGM_W63);
   and MGM_G78(ENABLE_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W64);
   not MGM_G79(MGM_W65,d_delay);
   and MGM_G80(MGM_W66,rb_delay,MGM_W65);
   not MGM_G81(MGM_W67,si_delay);
   and MGM_G82(MGM_W68,MGM_W67,MGM_W66);
   and MGM_G83(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W68);
   not MGM_G84(MGM_W69,d_delay);
   and MGM_G85(MGM_W70,rb_delay,MGM_W69);
   and MGM_G86(MGM_W71,si_delay,MGM_W70);
   and MGM_G87(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W71);
   and MGM_G88(MGM_W72,rb_delay,d_delay);
   not MGM_G89(MGM_W73,si_delay);
   and MGM_G90(MGM_W74,MGM_W73,MGM_W72);
   and MGM_G91(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W74);
   and MGM_G92(MGM_W75,rb_delay,d_delay);
   and MGM_G93(MGM_W76,si_delay,MGM_W75);
   and MGM_G94(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W76);
   not MGM_G95(MGM_W77,d_delay);
   not MGM_G96(MGM_W78,den_delay);
   and MGM_G97(MGM_W79,MGM_W78,MGM_W77);
   and MGM_G98(MGM_W80,si_delay,MGM_W79);
   not MGM_G99(MGM_W81,ssb_delay);
   and MGM_G100(ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W81,MGM_W80);
   not MGM_G101(MGM_W82,d_delay);
   and MGM_G102(MGM_W83,den_delay,MGM_W82);
   and MGM_G103(MGM_W84,si_delay,MGM_W83);
   not MGM_G104(MGM_W85,ssb_delay);
   and MGM_G105(ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W85,MGM_W84);
   not MGM_G106(MGM_W86,den_delay);
   and MGM_G107(MGM_W87,MGM_W86,d_delay);
   and MGM_G108(MGM_W88,si_delay,MGM_W87);
   not MGM_G109(MGM_W89,ssb_delay);
   and MGM_G110(ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W89,MGM_W88);
   and MGM_G111(MGM_W90,den_delay,d_delay);
   not MGM_G112(MGM_W91,si_delay);
   and MGM_G113(MGM_W92,MGM_W91,MGM_W90);
   and MGM_G114(ENABLE_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W92);
   and MGM_G115(MGM_W93,den_delay,d_delay);
   and MGM_G116(MGM_W94,si_delay,MGM_W93);
   not MGM_G117(MGM_W95,ssb_delay);
   and MGM_G118(ENABLE_d_AND_den_AND_si_AND_NOT_ssb,MGM_W95,MGM_W94);
   and MGM_G119(MGM_W96,den_delay,d_delay);
   and MGM_G120(MGM_W97,si_delay,MGM_W96);
   and MGM_G121(ENABLE_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W97);
   not MGM_G122(MGM_W98,clk_delay);
   not MGM_G123(MGM_W99,d_delay);
   and MGM_G124(MGM_W100,MGM_W99,MGM_W98);
   not MGM_G125(MGM_W101,den_delay);
   and MGM_G126(MGM_W102,MGM_W101,MGM_W100);
   not MGM_G127(MGM_W103,si_delay);
   and MGM_G128(MGM_W104,MGM_W103,MGM_W102);
   not MGM_G129(MGM_W105,ssb_delay);
   and MGM_G130(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W105,MGM_W104);
   not MGM_G131(MGM_W106,clk_delay);
   not MGM_G132(MGM_W107,d_delay);
   and MGM_G133(MGM_W108,MGM_W107,MGM_W106);
   not MGM_G134(MGM_W109,den_delay);
   and MGM_G135(MGM_W110,MGM_W109,MGM_W108);
   not MGM_G136(MGM_W111,si_delay);
   and MGM_G137(MGM_W112,MGM_W111,MGM_W110);
   and MGM_G138(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W112);
   not MGM_G139(MGM_W113,clk_delay);
   not MGM_G140(MGM_W114,d_delay);
   and MGM_G141(MGM_W115,MGM_W114,MGM_W113);
   not MGM_G142(MGM_W116,den_delay);
   and MGM_G143(MGM_W117,MGM_W116,MGM_W115);
   and MGM_G144(MGM_W118,si_delay,MGM_W117);
   not MGM_G145(MGM_W119,ssb_delay);
   and MGM_G146(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W119,MGM_W118);
   not MGM_G147(MGM_W120,clk_delay);
   not MGM_G148(MGM_W121,d_delay);
   and MGM_G149(MGM_W122,MGM_W121,MGM_W120);
   not MGM_G150(MGM_W123,den_delay);
   and MGM_G151(MGM_W124,MGM_W123,MGM_W122);
   and MGM_G152(MGM_W125,si_delay,MGM_W124);
   and MGM_G153(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W125);
   not MGM_G154(MGM_W126,clk_delay);
   not MGM_G155(MGM_W127,d_delay);
   and MGM_G156(MGM_W128,MGM_W127,MGM_W126);
   and MGM_G157(MGM_W129,den_delay,MGM_W128);
   not MGM_G158(MGM_W130,si_delay);
   and MGM_G159(MGM_W131,MGM_W130,MGM_W129);
   not MGM_G160(MGM_W132,ssb_delay);
   and MGM_G161(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W132,MGM_W131);
   not MGM_G162(MGM_W133,clk_delay);
   not MGM_G163(MGM_W134,d_delay);
   and MGM_G164(MGM_W135,MGM_W134,MGM_W133);
   and MGM_G165(MGM_W136,den_delay,MGM_W135);
   not MGM_G166(MGM_W137,si_delay);
   and MGM_G167(MGM_W138,MGM_W137,MGM_W136);
   and MGM_G168(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W138);
   not MGM_G169(MGM_W139,clk_delay);
   not MGM_G170(MGM_W140,d_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   and MGM_G172(MGM_W142,den_delay,MGM_W141);
   and MGM_G173(MGM_W143,si_delay,MGM_W142);
   not MGM_G174(MGM_W144,ssb_delay);
   and MGM_G175(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W144,MGM_W143);
   not MGM_G176(MGM_W145,clk_delay);
   not MGM_G177(MGM_W146,d_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(MGM_W148,den_delay,MGM_W147);
   and MGM_G180(MGM_W149,si_delay,MGM_W148);
   and MGM_G181(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W149);
   not MGM_G182(MGM_W150,clk_delay);
   and MGM_G183(MGM_W151,d_delay,MGM_W150);
   not MGM_G184(MGM_W152,den_delay);
   and MGM_G185(MGM_W153,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W154,si_delay);
   and MGM_G187(MGM_W155,MGM_W154,MGM_W153);
   not MGM_G188(MGM_W156,ssb_delay);
   and MGM_G189(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W156,MGM_W155);
   not MGM_G190(MGM_W157,clk_delay);
   and MGM_G191(MGM_W158,d_delay,MGM_W157);
   not MGM_G192(MGM_W159,den_delay);
   and MGM_G193(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G194(MGM_W161,si_delay);
   and MGM_G195(MGM_W162,MGM_W161,MGM_W160);
   and MGM_G196(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W162);
   not MGM_G197(MGM_W163,clk_delay);
   and MGM_G198(MGM_W164,d_delay,MGM_W163);
   not MGM_G199(MGM_W165,den_delay);
   and MGM_G200(MGM_W166,MGM_W165,MGM_W164);
   and MGM_G201(MGM_W167,si_delay,MGM_W166);
   not MGM_G202(MGM_W168,ssb_delay);
   and MGM_G203(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W168,MGM_W167);
   not MGM_G204(MGM_W169,clk_delay);
   and MGM_G205(MGM_W170,d_delay,MGM_W169);
   not MGM_G206(MGM_W171,den_delay);
   and MGM_G207(MGM_W172,MGM_W171,MGM_W170);
   and MGM_G208(MGM_W173,si_delay,MGM_W172);
   and MGM_G209(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W173);
   not MGM_G210(MGM_W174,clk_delay);
   and MGM_G211(MGM_W175,d_delay,MGM_W174);
   and MGM_G212(MGM_W176,den_delay,MGM_W175);
   not MGM_G213(MGM_W177,si_delay);
   and MGM_G214(MGM_W178,MGM_W177,MGM_W176);
   not MGM_G215(MGM_W179,ssb_delay);
   and MGM_G216(ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W179,MGM_W178);
   not MGM_G217(MGM_W180,clk_delay);
   and MGM_G218(MGM_W181,d_delay,MGM_W180);
   and MGM_G219(MGM_W182,den_delay,MGM_W181);
   not MGM_G220(MGM_W183,si_delay);
   and MGM_G221(MGM_W184,MGM_W183,MGM_W182);
   and MGM_G222(ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W184);
   not MGM_G223(MGM_W185,clk_delay);
   and MGM_G224(MGM_W186,d_delay,MGM_W185);
   and MGM_G225(MGM_W187,den_delay,MGM_W186);
   and MGM_G226(MGM_W188,si_delay,MGM_W187);
   not MGM_G227(MGM_W189,ssb_delay);
   and MGM_G228(ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_NOT_ssb,MGM_W189,MGM_W188);
   not MGM_G229(MGM_W190,clk_delay);
   and MGM_G230(MGM_W191,d_delay,MGM_W190);
   and MGM_G231(MGM_W192,den_delay,MGM_W191);
   and MGM_G232(MGM_W193,si_delay,MGM_W192);
   and MGM_G233(ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W193);
   not MGM_G234(MGM_W194,d_delay);
   and MGM_G235(MGM_W195,MGM_W194,clk_delay);
   not MGM_G236(MGM_W196,den_delay);
   and MGM_G237(MGM_W197,MGM_W196,MGM_W195);
   not MGM_G238(MGM_W198,si_delay);
   and MGM_G239(MGM_W199,MGM_W198,MGM_W197);
   not MGM_G240(MGM_W200,ssb_delay);
   and MGM_G241(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W200,MGM_W199);
   not MGM_G242(MGM_W201,d_delay);
   and MGM_G243(MGM_W202,MGM_W201,clk_delay);
   not MGM_G244(MGM_W203,den_delay);
   and MGM_G245(MGM_W204,MGM_W203,MGM_W202);
   not MGM_G246(MGM_W205,si_delay);
   and MGM_G247(MGM_W206,MGM_W205,MGM_W204);
   and MGM_G248(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W206);
   not MGM_G249(MGM_W207,d_delay);
   and MGM_G250(MGM_W208,MGM_W207,clk_delay);
   not MGM_G251(MGM_W209,den_delay);
   and MGM_G252(MGM_W210,MGM_W209,MGM_W208);
   and MGM_G253(MGM_W211,si_delay,MGM_W210);
   not MGM_G254(MGM_W212,ssb_delay);
   and MGM_G255(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W212,MGM_W211);
   not MGM_G256(MGM_W213,d_delay);
   and MGM_G257(MGM_W214,MGM_W213,clk_delay);
   not MGM_G258(MGM_W215,den_delay);
   and MGM_G259(MGM_W216,MGM_W215,MGM_W214);
   and MGM_G260(MGM_W217,si_delay,MGM_W216);
   and MGM_G261(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W217);
   not MGM_G262(MGM_W218,d_delay);
   and MGM_G263(MGM_W219,MGM_W218,clk_delay);
   and MGM_G264(MGM_W220,den_delay,MGM_W219);
   not MGM_G265(MGM_W221,si_delay);
   and MGM_G266(MGM_W222,MGM_W221,MGM_W220);
   not MGM_G267(MGM_W223,ssb_delay);
   and MGM_G268(ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W223,MGM_W222);
   not MGM_G269(MGM_W224,d_delay);
   and MGM_G270(MGM_W225,MGM_W224,clk_delay);
   and MGM_G271(MGM_W226,den_delay,MGM_W225);
   not MGM_G272(MGM_W227,si_delay);
   and MGM_G273(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G274(ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W228);
   not MGM_G275(MGM_W229,d_delay);
   and MGM_G276(MGM_W230,MGM_W229,clk_delay);
   and MGM_G277(MGM_W231,den_delay,MGM_W230);
   and MGM_G278(MGM_W232,si_delay,MGM_W231);
   not MGM_G279(MGM_W233,ssb_delay);
   and MGM_G280(ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W233,MGM_W232);
   not MGM_G281(MGM_W234,d_delay);
   and MGM_G282(MGM_W235,MGM_W234,clk_delay);
   and MGM_G283(MGM_W236,den_delay,MGM_W235);
   and MGM_G284(MGM_W237,si_delay,MGM_W236);
   and MGM_G285(ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W237);
   and MGM_G286(MGM_W238,d_delay,clk_delay);
   not MGM_G287(MGM_W239,den_delay);
   and MGM_G288(MGM_W240,MGM_W239,MGM_W238);
   not MGM_G289(MGM_W241,si_delay);
   and MGM_G290(MGM_W242,MGM_W241,MGM_W240);
   not MGM_G291(MGM_W243,ssb_delay);
   and MGM_G292(ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W243,MGM_W242);
   and MGM_G293(MGM_W244,d_delay,clk_delay);
   not MGM_G294(MGM_W245,den_delay);
   and MGM_G295(MGM_W246,MGM_W245,MGM_W244);
   not MGM_G296(MGM_W247,si_delay);
   and MGM_G297(MGM_W248,MGM_W247,MGM_W246);
   and MGM_G298(ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W248);
   and MGM_G299(MGM_W249,d_delay,clk_delay);
   not MGM_G300(MGM_W250,den_delay);
   and MGM_G301(MGM_W251,MGM_W250,MGM_W249);
   and MGM_G302(MGM_W252,si_delay,MGM_W251);
   not MGM_G303(MGM_W253,ssb_delay);
   and MGM_G304(ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W253,MGM_W252);
   and MGM_G305(MGM_W254,d_delay,clk_delay);
   not MGM_G306(MGM_W255,den_delay);
   and MGM_G307(MGM_W256,MGM_W255,MGM_W254);
   and MGM_G308(MGM_W257,si_delay,MGM_W256);
   and MGM_G309(ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W257);
   and MGM_G310(MGM_W258,d_delay,clk_delay);
   and MGM_G311(MGM_W259,den_delay,MGM_W258);
   not MGM_G312(MGM_W260,si_delay);
   and MGM_G313(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G314(MGM_W262,ssb_delay);
   and MGM_G315(ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   and MGM_G316(MGM_W263,d_delay,clk_delay);
   and MGM_G317(MGM_W264,den_delay,MGM_W263);
   not MGM_G318(MGM_W265,si_delay);
   and MGM_G319(MGM_W266,MGM_W265,MGM_W264);
   and MGM_G320(ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W266);
   and MGM_G321(MGM_W267,d_delay,clk_delay);
   and MGM_G322(MGM_W268,den_delay,MGM_W267);
   and MGM_G323(MGM_W269,si_delay,MGM_W268);
   not MGM_G324(MGM_W270,ssb_delay);
   and MGM_G325(ENABLE_clk_AND_d_AND_den_AND_si_AND_NOT_ssb,MGM_W270,MGM_W269);
   and MGM_G326(MGM_W271,d_delay,clk_delay);
   and MGM_G327(MGM_W272,den_delay,MGM_W271);
   and MGM_G328(MGM_W273,si_delay,MGM_W272);
   and MGM_G329(ENABLE_clk_AND_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W273);
   not MGM_G330(MGM_W274,d_delay);
   not MGM_G331(MGM_W275,den_delay);
   and MGM_G332(MGM_W276,MGM_W275,MGM_W274);
   and MGM_G333(MGM_W277,rb_delay,MGM_W276);
   not MGM_G334(MGM_W278,ssb_delay);
   and MGM_G335(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb,MGM_W278,MGM_W277);
   not MGM_G336(MGM_W279,d_delay);
   and MGM_G337(MGM_W280,den_delay,MGM_W279);
   and MGM_G338(MGM_W281,rb_delay,MGM_W280);
   not MGM_G339(MGM_W282,ssb_delay);
   and MGM_G340(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb,MGM_W282,MGM_W281);
   not MGM_G341(MGM_W283,den_delay);
   and MGM_G342(MGM_W284,MGM_W283,d_delay);
   and MGM_G343(MGM_W285,rb_delay,MGM_W284);
   not MGM_G344(MGM_W286,ssb_delay);
   and MGM_G345(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb,MGM_W286,MGM_W285);
   and MGM_G346(MGM_W287,den_delay,d_delay);
   and MGM_G347(MGM_W288,rb_delay,MGM_W287);
   not MGM_G348(MGM_W289,ssb_delay);
   and MGM_G349(ENABLE_d_AND_den_AND_rb_AND_NOT_ssb,MGM_W289,MGM_W288);
   not MGM_G350(MGM_W290,d_delay);
   not MGM_G351(MGM_W291,den_delay);
   and MGM_G352(MGM_W292,MGM_W291,MGM_W290);
   and MGM_G353(MGM_W293,rb_delay,MGM_W292);
   not MGM_G354(MGM_W294,si_delay);
   and MGM_G355(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si,MGM_W294,MGM_W293);
   not MGM_G356(MGM_W295,d_delay);
   not MGM_G357(MGM_W296,den_delay);
   and MGM_G358(MGM_W297,MGM_W296,MGM_W295);
   and MGM_G359(MGM_W298,rb_delay,MGM_W297);
   and MGM_G360(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si,si_delay,MGM_W298);
   not MGM_G361(MGM_W299,d_delay);
   and MGM_G362(MGM_W300,den_delay,MGM_W299);
   and MGM_G363(MGM_W301,rb_delay,MGM_W300);
   and MGM_G364(ENABLE_NOT_d_AND_den_AND_rb_AND_si,si_delay,MGM_W301);
   not MGM_G365(MGM_W302,den_delay);
   and MGM_G366(MGM_W303,MGM_W302,d_delay);
   and MGM_G367(MGM_W304,rb_delay,MGM_W303);
   not MGM_G368(MGM_W305,si_delay);
   and MGM_G369(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   not MGM_G370(MGM_W306,den_delay);
   and MGM_G371(MGM_W307,MGM_W306,d_delay);
   and MGM_G372(MGM_W308,rb_delay,MGM_W307);
   and MGM_G373(ENABLE_d_AND_NOT_den_AND_rb_AND_si,si_delay,MGM_W308);
   and MGM_G374(MGM_W309,den_delay,d_delay);
   and MGM_G375(MGM_W310,rb_delay,MGM_W309);
   not MGM_G376(MGM_W311,si_delay);
   and MGM_G377(ENABLE_d_AND_den_AND_rb_AND_NOT_si,MGM_W311,MGM_W310);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy043ah1n03x5( clk, d, den, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy043ah_func b15fqy043ah1n03x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy043ah_func b15fqy043ah1n03x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy043ah_func b15fqy043ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy043ah_func b15fqy043ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,den_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   and MGM_G3(MGM_W3,rb_delay,MGM_W2);
   not MGM_G4(MGM_W4,si_delay);
   and MGM_G5(MGM_W5,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W6,ssb_delay);
   and MGM_G7(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W6,MGM_W5);
   not MGM_G8(MGM_W7,d_delay);
   not MGM_G9(MGM_W8,den_delay);
   and MGM_G10(MGM_W9,MGM_W8,MGM_W7);
   and MGM_G11(MGM_W10,rb_delay,MGM_W9);
   and MGM_G12(MGM_W11,si_delay,MGM_W10);
   not MGM_G13(MGM_W12,ssb_delay);
   and MGM_G14(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G15(MGM_W13,d_delay);
   and MGM_G16(MGM_W14,den_delay,MGM_W13);
   and MGM_G17(MGM_W15,rb_delay,MGM_W14);
   not MGM_G18(MGM_W16,si_delay);
   and MGM_G19(MGM_W17,MGM_W16,MGM_W15);
   not MGM_G20(MGM_W18,ssb_delay);
   and MGM_G21(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   not MGM_G22(MGM_W19,d_delay);
   and MGM_G23(MGM_W20,den_delay,MGM_W19);
   and MGM_G24(MGM_W21,rb_delay,MGM_W20);
   not MGM_G25(MGM_W22,si_delay);
   and MGM_G26(MGM_W23,MGM_W22,MGM_W21);
   and MGM_G27(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W23);
   not MGM_G28(MGM_W24,d_delay);
   and MGM_G29(MGM_W25,den_delay,MGM_W24);
   and MGM_G30(MGM_W26,rb_delay,MGM_W25);
   and MGM_G31(MGM_W27,si_delay,MGM_W26);
   not MGM_G32(MGM_W28,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W28,MGM_W27);
   not MGM_G34(MGM_W29,d_delay);
   and MGM_G35(MGM_W30,den_delay,MGM_W29);
   and MGM_G36(MGM_W31,rb_delay,MGM_W30);
   and MGM_G37(MGM_W32,si_delay,MGM_W31);
   and MGM_G38(ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W32);
   not MGM_G39(MGM_W33,den_delay);
   and MGM_G40(MGM_W34,MGM_W33,d_delay);
   and MGM_G41(MGM_W35,rb_delay,MGM_W34);
   not MGM_G42(MGM_W36,si_delay);
   and MGM_G43(MGM_W37,MGM_W36,MGM_W35);
   not MGM_G44(MGM_W38,ssb_delay);
   and MGM_G45(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W38,MGM_W37);
   not MGM_G46(MGM_W39,den_delay);
   and MGM_G47(MGM_W40,MGM_W39,d_delay);
   and MGM_G48(MGM_W41,rb_delay,MGM_W40);
   and MGM_G49(MGM_W42,si_delay,MGM_W41);
   not MGM_G50(MGM_W43,ssb_delay);
   and MGM_G51(ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W43,MGM_W42);
   and MGM_G52(MGM_W44,den_delay,d_delay);
   and MGM_G53(MGM_W45,rb_delay,MGM_W44);
   not MGM_G54(MGM_W46,si_delay);
   and MGM_G55(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G56(MGM_W48,ssb_delay);
   and MGM_G57(ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   and MGM_G58(MGM_W49,den_delay,d_delay);
   and MGM_G59(MGM_W50,rb_delay,MGM_W49);
   not MGM_G60(MGM_W51,si_delay);
   and MGM_G61(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G62(ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G63(MGM_W53,den_delay,d_delay);
   and MGM_G64(MGM_W54,rb_delay,MGM_W53);
   and MGM_G65(MGM_W55,si_delay,MGM_W54);
   not MGM_G66(MGM_W56,ssb_delay);
   and MGM_G67(ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   and MGM_G68(MGM_W57,den_delay,d_delay);
   and MGM_G69(MGM_W58,rb_delay,MGM_W57);
   and MGM_G70(MGM_W59,si_delay,MGM_W58);
   and MGM_G71(ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W59);
   and MGM_G72(MGM_W60,rb_delay,den_delay);
   not MGM_G73(MGM_W61,si_delay);
   and MGM_G74(MGM_W62,MGM_W61,MGM_W60);
   and MGM_G75(ENABLE_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W62);
   and MGM_G76(MGM_W63,rb_delay,den_delay);
   and MGM_G77(MGM_W64,si_delay,MGM_W63);
   and MGM_G78(ENABLE_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W64);
   not MGM_G79(MGM_W65,d_delay);
   and MGM_G80(MGM_W66,rb_delay,MGM_W65);
   not MGM_G81(MGM_W67,si_delay);
   and MGM_G82(MGM_W68,MGM_W67,MGM_W66);
   and MGM_G83(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W68);
   not MGM_G84(MGM_W69,d_delay);
   and MGM_G85(MGM_W70,rb_delay,MGM_W69);
   and MGM_G86(MGM_W71,si_delay,MGM_W70);
   and MGM_G87(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W71);
   and MGM_G88(MGM_W72,rb_delay,d_delay);
   not MGM_G89(MGM_W73,si_delay);
   and MGM_G90(MGM_W74,MGM_W73,MGM_W72);
   and MGM_G91(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W74);
   and MGM_G92(MGM_W75,rb_delay,d_delay);
   and MGM_G93(MGM_W76,si_delay,MGM_W75);
   and MGM_G94(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W76);
   not MGM_G95(MGM_W77,d_delay);
   not MGM_G96(MGM_W78,den_delay);
   and MGM_G97(MGM_W79,MGM_W78,MGM_W77);
   and MGM_G98(MGM_W80,si_delay,MGM_W79);
   not MGM_G99(MGM_W81,ssb_delay);
   and MGM_G100(ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W81,MGM_W80);
   not MGM_G101(MGM_W82,d_delay);
   and MGM_G102(MGM_W83,den_delay,MGM_W82);
   and MGM_G103(MGM_W84,si_delay,MGM_W83);
   not MGM_G104(MGM_W85,ssb_delay);
   and MGM_G105(ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W85,MGM_W84);
   not MGM_G106(MGM_W86,den_delay);
   and MGM_G107(MGM_W87,MGM_W86,d_delay);
   and MGM_G108(MGM_W88,si_delay,MGM_W87);
   not MGM_G109(MGM_W89,ssb_delay);
   and MGM_G110(ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W89,MGM_W88);
   and MGM_G111(MGM_W90,den_delay,d_delay);
   not MGM_G112(MGM_W91,si_delay);
   and MGM_G113(MGM_W92,MGM_W91,MGM_W90);
   and MGM_G114(ENABLE_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W92);
   and MGM_G115(MGM_W93,den_delay,d_delay);
   and MGM_G116(MGM_W94,si_delay,MGM_W93);
   not MGM_G117(MGM_W95,ssb_delay);
   and MGM_G118(ENABLE_d_AND_den_AND_si_AND_NOT_ssb,MGM_W95,MGM_W94);
   and MGM_G119(MGM_W96,den_delay,d_delay);
   and MGM_G120(MGM_W97,si_delay,MGM_W96);
   and MGM_G121(ENABLE_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W97);
   not MGM_G122(MGM_W98,clk_delay);
   not MGM_G123(MGM_W99,d_delay);
   and MGM_G124(MGM_W100,MGM_W99,MGM_W98);
   not MGM_G125(MGM_W101,den_delay);
   and MGM_G126(MGM_W102,MGM_W101,MGM_W100);
   not MGM_G127(MGM_W103,si_delay);
   and MGM_G128(MGM_W104,MGM_W103,MGM_W102);
   not MGM_G129(MGM_W105,ssb_delay);
   and MGM_G130(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W105,MGM_W104);
   not MGM_G131(MGM_W106,clk_delay);
   not MGM_G132(MGM_W107,d_delay);
   and MGM_G133(MGM_W108,MGM_W107,MGM_W106);
   not MGM_G134(MGM_W109,den_delay);
   and MGM_G135(MGM_W110,MGM_W109,MGM_W108);
   not MGM_G136(MGM_W111,si_delay);
   and MGM_G137(MGM_W112,MGM_W111,MGM_W110);
   and MGM_G138(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W112);
   not MGM_G139(MGM_W113,clk_delay);
   not MGM_G140(MGM_W114,d_delay);
   and MGM_G141(MGM_W115,MGM_W114,MGM_W113);
   not MGM_G142(MGM_W116,den_delay);
   and MGM_G143(MGM_W117,MGM_W116,MGM_W115);
   and MGM_G144(MGM_W118,si_delay,MGM_W117);
   not MGM_G145(MGM_W119,ssb_delay);
   and MGM_G146(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W119,MGM_W118);
   not MGM_G147(MGM_W120,clk_delay);
   not MGM_G148(MGM_W121,d_delay);
   and MGM_G149(MGM_W122,MGM_W121,MGM_W120);
   not MGM_G150(MGM_W123,den_delay);
   and MGM_G151(MGM_W124,MGM_W123,MGM_W122);
   and MGM_G152(MGM_W125,si_delay,MGM_W124);
   and MGM_G153(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W125);
   not MGM_G154(MGM_W126,clk_delay);
   not MGM_G155(MGM_W127,d_delay);
   and MGM_G156(MGM_W128,MGM_W127,MGM_W126);
   and MGM_G157(MGM_W129,den_delay,MGM_W128);
   not MGM_G158(MGM_W130,si_delay);
   and MGM_G159(MGM_W131,MGM_W130,MGM_W129);
   not MGM_G160(MGM_W132,ssb_delay);
   and MGM_G161(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W132,MGM_W131);
   not MGM_G162(MGM_W133,clk_delay);
   not MGM_G163(MGM_W134,d_delay);
   and MGM_G164(MGM_W135,MGM_W134,MGM_W133);
   and MGM_G165(MGM_W136,den_delay,MGM_W135);
   not MGM_G166(MGM_W137,si_delay);
   and MGM_G167(MGM_W138,MGM_W137,MGM_W136);
   and MGM_G168(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W138);
   not MGM_G169(MGM_W139,clk_delay);
   not MGM_G170(MGM_W140,d_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   and MGM_G172(MGM_W142,den_delay,MGM_W141);
   and MGM_G173(MGM_W143,si_delay,MGM_W142);
   not MGM_G174(MGM_W144,ssb_delay);
   and MGM_G175(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W144,MGM_W143);
   not MGM_G176(MGM_W145,clk_delay);
   not MGM_G177(MGM_W146,d_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(MGM_W148,den_delay,MGM_W147);
   and MGM_G180(MGM_W149,si_delay,MGM_W148);
   and MGM_G181(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W149);
   not MGM_G182(MGM_W150,clk_delay);
   and MGM_G183(MGM_W151,d_delay,MGM_W150);
   not MGM_G184(MGM_W152,den_delay);
   and MGM_G185(MGM_W153,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W154,si_delay);
   and MGM_G187(MGM_W155,MGM_W154,MGM_W153);
   not MGM_G188(MGM_W156,ssb_delay);
   and MGM_G189(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W156,MGM_W155);
   not MGM_G190(MGM_W157,clk_delay);
   and MGM_G191(MGM_W158,d_delay,MGM_W157);
   not MGM_G192(MGM_W159,den_delay);
   and MGM_G193(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G194(MGM_W161,si_delay);
   and MGM_G195(MGM_W162,MGM_W161,MGM_W160);
   and MGM_G196(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W162);
   not MGM_G197(MGM_W163,clk_delay);
   and MGM_G198(MGM_W164,d_delay,MGM_W163);
   not MGM_G199(MGM_W165,den_delay);
   and MGM_G200(MGM_W166,MGM_W165,MGM_W164);
   and MGM_G201(MGM_W167,si_delay,MGM_W166);
   not MGM_G202(MGM_W168,ssb_delay);
   and MGM_G203(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W168,MGM_W167);
   not MGM_G204(MGM_W169,clk_delay);
   and MGM_G205(MGM_W170,d_delay,MGM_W169);
   not MGM_G206(MGM_W171,den_delay);
   and MGM_G207(MGM_W172,MGM_W171,MGM_W170);
   and MGM_G208(MGM_W173,si_delay,MGM_W172);
   and MGM_G209(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W173);
   not MGM_G210(MGM_W174,clk_delay);
   and MGM_G211(MGM_W175,d_delay,MGM_W174);
   and MGM_G212(MGM_W176,den_delay,MGM_W175);
   not MGM_G213(MGM_W177,si_delay);
   and MGM_G214(MGM_W178,MGM_W177,MGM_W176);
   not MGM_G215(MGM_W179,ssb_delay);
   and MGM_G216(ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W179,MGM_W178);
   not MGM_G217(MGM_W180,clk_delay);
   and MGM_G218(MGM_W181,d_delay,MGM_W180);
   and MGM_G219(MGM_W182,den_delay,MGM_W181);
   not MGM_G220(MGM_W183,si_delay);
   and MGM_G221(MGM_W184,MGM_W183,MGM_W182);
   and MGM_G222(ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W184);
   not MGM_G223(MGM_W185,clk_delay);
   and MGM_G224(MGM_W186,d_delay,MGM_W185);
   and MGM_G225(MGM_W187,den_delay,MGM_W186);
   and MGM_G226(MGM_W188,si_delay,MGM_W187);
   not MGM_G227(MGM_W189,ssb_delay);
   and MGM_G228(ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_NOT_ssb,MGM_W189,MGM_W188);
   not MGM_G229(MGM_W190,clk_delay);
   and MGM_G230(MGM_W191,d_delay,MGM_W190);
   and MGM_G231(MGM_W192,den_delay,MGM_W191);
   and MGM_G232(MGM_W193,si_delay,MGM_W192);
   and MGM_G233(ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W193);
   not MGM_G234(MGM_W194,d_delay);
   and MGM_G235(MGM_W195,MGM_W194,clk_delay);
   not MGM_G236(MGM_W196,den_delay);
   and MGM_G237(MGM_W197,MGM_W196,MGM_W195);
   not MGM_G238(MGM_W198,si_delay);
   and MGM_G239(MGM_W199,MGM_W198,MGM_W197);
   not MGM_G240(MGM_W200,ssb_delay);
   and MGM_G241(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W200,MGM_W199);
   not MGM_G242(MGM_W201,d_delay);
   and MGM_G243(MGM_W202,MGM_W201,clk_delay);
   not MGM_G244(MGM_W203,den_delay);
   and MGM_G245(MGM_W204,MGM_W203,MGM_W202);
   not MGM_G246(MGM_W205,si_delay);
   and MGM_G247(MGM_W206,MGM_W205,MGM_W204);
   and MGM_G248(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W206);
   not MGM_G249(MGM_W207,d_delay);
   and MGM_G250(MGM_W208,MGM_W207,clk_delay);
   not MGM_G251(MGM_W209,den_delay);
   and MGM_G252(MGM_W210,MGM_W209,MGM_W208);
   and MGM_G253(MGM_W211,si_delay,MGM_W210);
   not MGM_G254(MGM_W212,ssb_delay);
   and MGM_G255(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W212,MGM_W211);
   not MGM_G256(MGM_W213,d_delay);
   and MGM_G257(MGM_W214,MGM_W213,clk_delay);
   not MGM_G258(MGM_W215,den_delay);
   and MGM_G259(MGM_W216,MGM_W215,MGM_W214);
   and MGM_G260(MGM_W217,si_delay,MGM_W216);
   and MGM_G261(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W217);
   not MGM_G262(MGM_W218,d_delay);
   and MGM_G263(MGM_W219,MGM_W218,clk_delay);
   and MGM_G264(MGM_W220,den_delay,MGM_W219);
   not MGM_G265(MGM_W221,si_delay);
   and MGM_G266(MGM_W222,MGM_W221,MGM_W220);
   not MGM_G267(MGM_W223,ssb_delay);
   and MGM_G268(ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W223,MGM_W222);
   not MGM_G269(MGM_W224,d_delay);
   and MGM_G270(MGM_W225,MGM_W224,clk_delay);
   and MGM_G271(MGM_W226,den_delay,MGM_W225);
   not MGM_G272(MGM_W227,si_delay);
   and MGM_G273(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G274(ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W228);
   not MGM_G275(MGM_W229,d_delay);
   and MGM_G276(MGM_W230,MGM_W229,clk_delay);
   and MGM_G277(MGM_W231,den_delay,MGM_W230);
   and MGM_G278(MGM_W232,si_delay,MGM_W231);
   not MGM_G279(MGM_W233,ssb_delay);
   and MGM_G280(ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W233,MGM_W232);
   not MGM_G281(MGM_W234,d_delay);
   and MGM_G282(MGM_W235,MGM_W234,clk_delay);
   and MGM_G283(MGM_W236,den_delay,MGM_W235);
   and MGM_G284(MGM_W237,si_delay,MGM_W236);
   and MGM_G285(ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W237);
   and MGM_G286(MGM_W238,d_delay,clk_delay);
   not MGM_G287(MGM_W239,den_delay);
   and MGM_G288(MGM_W240,MGM_W239,MGM_W238);
   not MGM_G289(MGM_W241,si_delay);
   and MGM_G290(MGM_W242,MGM_W241,MGM_W240);
   not MGM_G291(MGM_W243,ssb_delay);
   and MGM_G292(ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W243,MGM_W242);
   and MGM_G293(MGM_W244,d_delay,clk_delay);
   not MGM_G294(MGM_W245,den_delay);
   and MGM_G295(MGM_W246,MGM_W245,MGM_W244);
   not MGM_G296(MGM_W247,si_delay);
   and MGM_G297(MGM_W248,MGM_W247,MGM_W246);
   and MGM_G298(ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W248);
   and MGM_G299(MGM_W249,d_delay,clk_delay);
   not MGM_G300(MGM_W250,den_delay);
   and MGM_G301(MGM_W251,MGM_W250,MGM_W249);
   and MGM_G302(MGM_W252,si_delay,MGM_W251);
   not MGM_G303(MGM_W253,ssb_delay);
   and MGM_G304(ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W253,MGM_W252);
   and MGM_G305(MGM_W254,d_delay,clk_delay);
   not MGM_G306(MGM_W255,den_delay);
   and MGM_G307(MGM_W256,MGM_W255,MGM_W254);
   and MGM_G308(MGM_W257,si_delay,MGM_W256);
   and MGM_G309(ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W257);
   and MGM_G310(MGM_W258,d_delay,clk_delay);
   and MGM_G311(MGM_W259,den_delay,MGM_W258);
   not MGM_G312(MGM_W260,si_delay);
   and MGM_G313(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G314(MGM_W262,ssb_delay);
   and MGM_G315(ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   and MGM_G316(MGM_W263,d_delay,clk_delay);
   and MGM_G317(MGM_W264,den_delay,MGM_W263);
   not MGM_G318(MGM_W265,si_delay);
   and MGM_G319(MGM_W266,MGM_W265,MGM_W264);
   and MGM_G320(ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W266);
   and MGM_G321(MGM_W267,d_delay,clk_delay);
   and MGM_G322(MGM_W268,den_delay,MGM_W267);
   and MGM_G323(MGM_W269,si_delay,MGM_W268);
   not MGM_G324(MGM_W270,ssb_delay);
   and MGM_G325(ENABLE_clk_AND_d_AND_den_AND_si_AND_NOT_ssb,MGM_W270,MGM_W269);
   and MGM_G326(MGM_W271,d_delay,clk_delay);
   and MGM_G327(MGM_W272,den_delay,MGM_W271);
   and MGM_G328(MGM_W273,si_delay,MGM_W272);
   and MGM_G329(ENABLE_clk_AND_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W273);
   not MGM_G330(MGM_W274,d_delay);
   not MGM_G331(MGM_W275,den_delay);
   and MGM_G332(MGM_W276,MGM_W275,MGM_W274);
   and MGM_G333(MGM_W277,rb_delay,MGM_W276);
   not MGM_G334(MGM_W278,ssb_delay);
   and MGM_G335(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb,MGM_W278,MGM_W277);
   not MGM_G336(MGM_W279,d_delay);
   and MGM_G337(MGM_W280,den_delay,MGM_W279);
   and MGM_G338(MGM_W281,rb_delay,MGM_W280);
   not MGM_G339(MGM_W282,ssb_delay);
   and MGM_G340(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb,MGM_W282,MGM_W281);
   not MGM_G341(MGM_W283,den_delay);
   and MGM_G342(MGM_W284,MGM_W283,d_delay);
   and MGM_G343(MGM_W285,rb_delay,MGM_W284);
   not MGM_G344(MGM_W286,ssb_delay);
   and MGM_G345(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb,MGM_W286,MGM_W285);
   and MGM_G346(MGM_W287,den_delay,d_delay);
   and MGM_G347(MGM_W288,rb_delay,MGM_W287);
   not MGM_G348(MGM_W289,ssb_delay);
   and MGM_G349(ENABLE_d_AND_den_AND_rb_AND_NOT_ssb,MGM_W289,MGM_W288);
   not MGM_G350(MGM_W290,d_delay);
   not MGM_G351(MGM_W291,den_delay);
   and MGM_G352(MGM_W292,MGM_W291,MGM_W290);
   and MGM_G353(MGM_W293,rb_delay,MGM_W292);
   not MGM_G354(MGM_W294,si_delay);
   and MGM_G355(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si,MGM_W294,MGM_W293);
   not MGM_G356(MGM_W295,d_delay);
   not MGM_G357(MGM_W296,den_delay);
   and MGM_G358(MGM_W297,MGM_W296,MGM_W295);
   and MGM_G359(MGM_W298,rb_delay,MGM_W297);
   and MGM_G360(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si,si_delay,MGM_W298);
   not MGM_G361(MGM_W299,d_delay);
   and MGM_G362(MGM_W300,den_delay,MGM_W299);
   and MGM_G363(MGM_W301,rb_delay,MGM_W300);
   and MGM_G364(ENABLE_NOT_d_AND_den_AND_rb_AND_si,si_delay,MGM_W301);
   not MGM_G365(MGM_W302,den_delay);
   and MGM_G366(MGM_W303,MGM_W302,d_delay);
   and MGM_G367(MGM_W304,rb_delay,MGM_W303);
   not MGM_G368(MGM_W305,si_delay);
   and MGM_G369(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   not MGM_G370(MGM_W306,den_delay);
   and MGM_G371(MGM_W307,MGM_W306,d_delay);
   and MGM_G372(MGM_W308,rb_delay,MGM_W307);
   and MGM_G373(ENABLE_d_AND_NOT_den_AND_rb_AND_si,si_delay,MGM_W308);
   and MGM_G374(MGM_W309,den_delay,d_delay);
   and MGM_G375(MGM_W310,rb_delay,MGM_W309);
   not MGM_G376(MGM_W311,si_delay);
   and MGM_G377(ENABLE_d_AND_den_AND_rb_AND_NOT_si,MGM_W311,MGM_W310);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy043ah1n04x5( clk, d, den, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy043ah_func b15fqy043ah1n04x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy043ah_func b15fqy043ah1n04x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy043ah_func b15fqy043ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy043ah_func b15fqy043ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,den_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   and MGM_G3(MGM_W3,rb_delay,MGM_W2);
   not MGM_G4(MGM_W4,si_delay);
   and MGM_G5(MGM_W5,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W6,ssb_delay);
   and MGM_G7(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W6,MGM_W5);
   not MGM_G8(MGM_W7,d_delay);
   not MGM_G9(MGM_W8,den_delay);
   and MGM_G10(MGM_W9,MGM_W8,MGM_W7);
   and MGM_G11(MGM_W10,rb_delay,MGM_W9);
   and MGM_G12(MGM_W11,si_delay,MGM_W10);
   not MGM_G13(MGM_W12,ssb_delay);
   and MGM_G14(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G15(MGM_W13,d_delay);
   and MGM_G16(MGM_W14,den_delay,MGM_W13);
   and MGM_G17(MGM_W15,rb_delay,MGM_W14);
   not MGM_G18(MGM_W16,si_delay);
   and MGM_G19(MGM_W17,MGM_W16,MGM_W15);
   not MGM_G20(MGM_W18,ssb_delay);
   and MGM_G21(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   not MGM_G22(MGM_W19,d_delay);
   and MGM_G23(MGM_W20,den_delay,MGM_W19);
   and MGM_G24(MGM_W21,rb_delay,MGM_W20);
   not MGM_G25(MGM_W22,si_delay);
   and MGM_G26(MGM_W23,MGM_W22,MGM_W21);
   and MGM_G27(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W23);
   not MGM_G28(MGM_W24,d_delay);
   and MGM_G29(MGM_W25,den_delay,MGM_W24);
   and MGM_G30(MGM_W26,rb_delay,MGM_W25);
   and MGM_G31(MGM_W27,si_delay,MGM_W26);
   not MGM_G32(MGM_W28,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W28,MGM_W27);
   not MGM_G34(MGM_W29,d_delay);
   and MGM_G35(MGM_W30,den_delay,MGM_W29);
   and MGM_G36(MGM_W31,rb_delay,MGM_W30);
   and MGM_G37(MGM_W32,si_delay,MGM_W31);
   and MGM_G38(ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W32);
   not MGM_G39(MGM_W33,den_delay);
   and MGM_G40(MGM_W34,MGM_W33,d_delay);
   and MGM_G41(MGM_W35,rb_delay,MGM_W34);
   not MGM_G42(MGM_W36,si_delay);
   and MGM_G43(MGM_W37,MGM_W36,MGM_W35);
   not MGM_G44(MGM_W38,ssb_delay);
   and MGM_G45(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W38,MGM_W37);
   not MGM_G46(MGM_W39,den_delay);
   and MGM_G47(MGM_W40,MGM_W39,d_delay);
   and MGM_G48(MGM_W41,rb_delay,MGM_W40);
   and MGM_G49(MGM_W42,si_delay,MGM_W41);
   not MGM_G50(MGM_W43,ssb_delay);
   and MGM_G51(ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W43,MGM_W42);
   and MGM_G52(MGM_W44,den_delay,d_delay);
   and MGM_G53(MGM_W45,rb_delay,MGM_W44);
   not MGM_G54(MGM_W46,si_delay);
   and MGM_G55(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G56(MGM_W48,ssb_delay);
   and MGM_G57(ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   and MGM_G58(MGM_W49,den_delay,d_delay);
   and MGM_G59(MGM_W50,rb_delay,MGM_W49);
   not MGM_G60(MGM_W51,si_delay);
   and MGM_G61(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G62(ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G63(MGM_W53,den_delay,d_delay);
   and MGM_G64(MGM_W54,rb_delay,MGM_W53);
   and MGM_G65(MGM_W55,si_delay,MGM_W54);
   not MGM_G66(MGM_W56,ssb_delay);
   and MGM_G67(ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   and MGM_G68(MGM_W57,den_delay,d_delay);
   and MGM_G69(MGM_W58,rb_delay,MGM_W57);
   and MGM_G70(MGM_W59,si_delay,MGM_W58);
   and MGM_G71(ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W59);
   and MGM_G72(MGM_W60,rb_delay,den_delay);
   not MGM_G73(MGM_W61,si_delay);
   and MGM_G74(MGM_W62,MGM_W61,MGM_W60);
   and MGM_G75(ENABLE_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W62);
   and MGM_G76(MGM_W63,rb_delay,den_delay);
   and MGM_G77(MGM_W64,si_delay,MGM_W63);
   and MGM_G78(ENABLE_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W64);
   not MGM_G79(MGM_W65,d_delay);
   and MGM_G80(MGM_W66,rb_delay,MGM_W65);
   not MGM_G81(MGM_W67,si_delay);
   and MGM_G82(MGM_W68,MGM_W67,MGM_W66);
   and MGM_G83(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W68);
   not MGM_G84(MGM_W69,d_delay);
   and MGM_G85(MGM_W70,rb_delay,MGM_W69);
   and MGM_G86(MGM_W71,si_delay,MGM_W70);
   and MGM_G87(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W71);
   and MGM_G88(MGM_W72,rb_delay,d_delay);
   not MGM_G89(MGM_W73,si_delay);
   and MGM_G90(MGM_W74,MGM_W73,MGM_W72);
   and MGM_G91(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W74);
   and MGM_G92(MGM_W75,rb_delay,d_delay);
   and MGM_G93(MGM_W76,si_delay,MGM_W75);
   and MGM_G94(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W76);
   not MGM_G95(MGM_W77,d_delay);
   not MGM_G96(MGM_W78,den_delay);
   and MGM_G97(MGM_W79,MGM_W78,MGM_W77);
   and MGM_G98(MGM_W80,si_delay,MGM_W79);
   not MGM_G99(MGM_W81,ssb_delay);
   and MGM_G100(ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W81,MGM_W80);
   not MGM_G101(MGM_W82,d_delay);
   and MGM_G102(MGM_W83,den_delay,MGM_W82);
   and MGM_G103(MGM_W84,si_delay,MGM_W83);
   not MGM_G104(MGM_W85,ssb_delay);
   and MGM_G105(ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W85,MGM_W84);
   not MGM_G106(MGM_W86,den_delay);
   and MGM_G107(MGM_W87,MGM_W86,d_delay);
   and MGM_G108(MGM_W88,si_delay,MGM_W87);
   not MGM_G109(MGM_W89,ssb_delay);
   and MGM_G110(ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W89,MGM_W88);
   and MGM_G111(MGM_W90,den_delay,d_delay);
   not MGM_G112(MGM_W91,si_delay);
   and MGM_G113(MGM_W92,MGM_W91,MGM_W90);
   and MGM_G114(ENABLE_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W92);
   and MGM_G115(MGM_W93,den_delay,d_delay);
   and MGM_G116(MGM_W94,si_delay,MGM_W93);
   not MGM_G117(MGM_W95,ssb_delay);
   and MGM_G118(ENABLE_d_AND_den_AND_si_AND_NOT_ssb,MGM_W95,MGM_W94);
   and MGM_G119(MGM_W96,den_delay,d_delay);
   and MGM_G120(MGM_W97,si_delay,MGM_W96);
   and MGM_G121(ENABLE_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W97);
   not MGM_G122(MGM_W98,clk_delay);
   not MGM_G123(MGM_W99,d_delay);
   and MGM_G124(MGM_W100,MGM_W99,MGM_W98);
   not MGM_G125(MGM_W101,den_delay);
   and MGM_G126(MGM_W102,MGM_W101,MGM_W100);
   not MGM_G127(MGM_W103,si_delay);
   and MGM_G128(MGM_W104,MGM_W103,MGM_W102);
   not MGM_G129(MGM_W105,ssb_delay);
   and MGM_G130(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W105,MGM_W104);
   not MGM_G131(MGM_W106,clk_delay);
   not MGM_G132(MGM_W107,d_delay);
   and MGM_G133(MGM_W108,MGM_W107,MGM_W106);
   not MGM_G134(MGM_W109,den_delay);
   and MGM_G135(MGM_W110,MGM_W109,MGM_W108);
   not MGM_G136(MGM_W111,si_delay);
   and MGM_G137(MGM_W112,MGM_W111,MGM_W110);
   and MGM_G138(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W112);
   not MGM_G139(MGM_W113,clk_delay);
   not MGM_G140(MGM_W114,d_delay);
   and MGM_G141(MGM_W115,MGM_W114,MGM_W113);
   not MGM_G142(MGM_W116,den_delay);
   and MGM_G143(MGM_W117,MGM_W116,MGM_W115);
   and MGM_G144(MGM_W118,si_delay,MGM_W117);
   not MGM_G145(MGM_W119,ssb_delay);
   and MGM_G146(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W119,MGM_W118);
   not MGM_G147(MGM_W120,clk_delay);
   not MGM_G148(MGM_W121,d_delay);
   and MGM_G149(MGM_W122,MGM_W121,MGM_W120);
   not MGM_G150(MGM_W123,den_delay);
   and MGM_G151(MGM_W124,MGM_W123,MGM_W122);
   and MGM_G152(MGM_W125,si_delay,MGM_W124);
   and MGM_G153(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W125);
   not MGM_G154(MGM_W126,clk_delay);
   not MGM_G155(MGM_W127,d_delay);
   and MGM_G156(MGM_W128,MGM_W127,MGM_W126);
   and MGM_G157(MGM_W129,den_delay,MGM_W128);
   not MGM_G158(MGM_W130,si_delay);
   and MGM_G159(MGM_W131,MGM_W130,MGM_W129);
   not MGM_G160(MGM_W132,ssb_delay);
   and MGM_G161(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W132,MGM_W131);
   not MGM_G162(MGM_W133,clk_delay);
   not MGM_G163(MGM_W134,d_delay);
   and MGM_G164(MGM_W135,MGM_W134,MGM_W133);
   and MGM_G165(MGM_W136,den_delay,MGM_W135);
   not MGM_G166(MGM_W137,si_delay);
   and MGM_G167(MGM_W138,MGM_W137,MGM_W136);
   and MGM_G168(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W138);
   not MGM_G169(MGM_W139,clk_delay);
   not MGM_G170(MGM_W140,d_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   and MGM_G172(MGM_W142,den_delay,MGM_W141);
   and MGM_G173(MGM_W143,si_delay,MGM_W142);
   not MGM_G174(MGM_W144,ssb_delay);
   and MGM_G175(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W144,MGM_W143);
   not MGM_G176(MGM_W145,clk_delay);
   not MGM_G177(MGM_W146,d_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(MGM_W148,den_delay,MGM_W147);
   and MGM_G180(MGM_W149,si_delay,MGM_W148);
   and MGM_G181(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W149);
   not MGM_G182(MGM_W150,clk_delay);
   and MGM_G183(MGM_W151,d_delay,MGM_W150);
   not MGM_G184(MGM_W152,den_delay);
   and MGM_G185(MGM_W153,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W154,si_delay);
   and MGM_G187(MGM_W155,MGM_W154,MGM_W153);
   not MGM_G188(MGM_W156,ssb_delay);
   and MGM_G189(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W156,MGM_W155);
   not MGM_G190(MGM_W157,clk_delay);
   and MGM_G191(MGM_W158,d_delay,MGM_W157);
   not MGM_G192(MGM_W159,den_delay);
   and MGM_G193(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G194(MGM_W161,si_delay);
   and MGM_G195(MGM_W162,MGM_W161,MGM_W160);
   and MGM_G196(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W162);
   not MGM_G197(MGM_W163,clk_delay);
   and MGM_G198(MGM_W164,d_delay,MGM_W163);
   not MGM_G199(MGM_W165,den_delay);
   and MGM_G200(MGM_W166,MGM_W165,MGM_W164);
   and MGM_G201(MGM_W167,si_delay,MGM_W166);
   not MGM_G202(MGM_W168,ssb_delay);
   and MGM_G203(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W168,MGM_W167);
   not MGM_G204(MGM_W169,clk_delay);
   and MGM_G205(MGM_W170,d_delay,MGM_W169);
   not MGM_G206(MGM_W171,den_delay);
   and MGM_G207(MGM_W172,MGM_W171,MGM_W170);
   and MGM_G208(MGM_W173,si_delay,MGM_W172);
   and MGM_G209(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W173);
   not MGM_G210(MGM_W174,clk_delay);
   and MGM_G211(MGM_W175,d_delay,MGM_W174);
   and MGM_G212(MGM_W176,den_delay,MGM_W175);
   not MGM_G213(MGM_W177,si_delay);
   and MGM_G214(MGM_W178,MGM_W177,MGM_W176);
   not MGM_G215(MGM_W179,ssb_delay);
   and MGM_G216(ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W179,MGM_W178);
   not MGM_G217(MGM_W180,clk_delay);
   and MGM_G218(MGM_W181,d_delay,MGM_W180);
   and MGM_G219(MGM_W182,den_delay,MGM_W181);
   not MGM_G220(MGM_W183,si_delay);
   and MGM_G221(MGM_W184,MGM_W183,MGM_W182);
   and MGM_G222(ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W184);
   not MGM_G223(MGM_W185,clk_delay);
   and MGM_G224(MGM_W186,d_delay,MGM_W185);
   and MGM_G225(MGM_W187,den_delay,MGM_W186);
   and MGM_G226(MGM_W188,si_delay,MGM_W187);
   not MGM_G227(MGM_W189,ssb_delay);
   and MGM_G228(ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_NOT_ssb,MGM_W189,MGM_W188);
   not MGM_G229(MGM_W190,clk_delay);
   and MGM_G230(MGM_W191,d_delay,MGM_W190);
   and MGM_G231(MGM_W192,den_delay,MGM_W191);
   and MGM_G232(MGM_W193,si_delay,MGM_W192);
   and MGM_G233(ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W193);
   not MGM_G234(MGM_W194,d_delay);
   and MGM_G235(MGM_W195,MGM_W194,clk_delay);
   not MGM_G236(MGM_W196,den_delay);
   and MGM_G237(MGM_W197,MGM_W196,MGM_W195);
   not MGM_G238(MGM_W198,si_delay);
   and MGM_G239(MGM_W199,MGM_W198,MGM_W197);
   not MGM_G240(MGM_W200,ssb_delay);
   and MGM_G241(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W200,MGM_W199);
   not MGM_G242(MGM_W201,d_delay);
   and MGM_G243(MGM_W202,MGM_W201,clk_delay);
   not MGM_G244(MGM_W203,den_delay);
   and MGM_G245(MGM_W204,MGM_W203,MGM_W202);
   not MGM_G246(MGM_W205,si_delay);
   and MGM_G247(MGM_W206,MGM_W205,MGM_W204);
   and MGM_G248(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W206);
   not MGM_G249(MGM_W207,d_delay);
   and MGM_G250(MGM_W208,MGM_W207,clk_delay);
   not MGM_G251(MGM_W209,den_delay);
   and MGM_G252(MGM_W210,MGM_W209,MGM_W208);
   and MGM_G253(MGM_W211,si_delay,MGM_W210);
   not MGM_G254(MGM_W212,ssb_delay);
   and MGM_G255(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W212,MGM_W211);
   not MGM_G256(MGM_W213,d_delay);
   and MGM_G257(MGM_W214,MGM_W213,clk_delay);
   not MGM_G258(MGM_W215,den_delay);
   and MGM_G259(MGM_W216,MGM_W215,MGM_W214);
   and MGM_G260(MGM_W217,si_delay,MGM_W216);
   and MGM_G261(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W217);
   not MGM_G262(MGM_W218,d_delay);
   and MGM_G263(MGM_W219,MGM_W218,clk_delay);
   and MGM_G264(MGM_W220,den_delay,MGM_W219);
   not MGM_G265(MGM_W221,si_delay);
   and MGM_G266(MGM_W222,MGM_W221,MGM_W220);
   not MGM_G267(MGM_W223,ssb_delay);
   and MGM_G268(ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W223,MGM_W222);
   not MGM_G269(MGM_W224,d_delay);
   and MGM_G270(MGM_W225,MGM_W224,clk_delay);
   and MGM_G271(MGM_W226,den_delay,MGM_W225);
   not MGM_G272(MGM_W227,si_delay);
   and MGM_G273(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G274(ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W228);
   not MGM_G275(MGM_W229,d_delay);
   and MGM_G276(MGM_W230,MGM_W229,clk_delay);
   and MGM_G277(MGM_W231,den_delay,MGM_W230);
   and MGM_G278(MGM_W232,si_delay,MGM_W231);
   not MGM_G279(MGM_W233,ssb_delay);
   and MGM_G280(ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W233,MGM_W232);
   not MGM_G281(MGM_W234,d_delay);
   and MGM_G282(MGM_W235,MGM_W234,clk_delay);
   and MGM_G283(MGM_W236,den_delay,MGM_W235);
   and MGM_G284(MGM_W237,si_delay,MGM_W236);
   and MGM_G285(ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W237);
   and MGM_G286(MGM_W238,d_delay,clk_delay);
   not MGM_G287(MGM_W239,den_delay);
   and MGM_G288(MGM_W240,MGM_W239,MGM_W238);
   not MGM_G289(MGM_W241,si_delay);
   and MGM_G290(MGM_W242,MGM_W241,MGM_W240);
   not MGM_G291(MGM_W243,ssb_delay);
   and MGM_G292(ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W243,MGM_W242);
   and MGM_G293(MGM_W244,d_delay,clk_delay);
   not MGM_G294(MGM_W245,den_delay);
   and MGM_G295(MGM_W246,MGM_W245,MGM_W244);
   not MGM_G296(MGM_W247,si_delay);
   and MGM_G297(MGM_W248,MGM_W247,MGM_W246);
   and MGM_G298(ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W248);
   and MGM_G299(MGM_W249,d_delay,clk_delay);
   not MGM_G300(MGM_W250,den_delay);
   and MGM_G301(MGM_W251,MGM_W250,MGM_W249);
   and MGM_G302(MGM_W252,si_delay,MGM_W251);
   not MGM_G303(MGM_W253,ssb_delay);
   and MGM_G304(ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W253,MGM_W252);
   and MGM_G305(MGM_W254,d_delay,clk_delay);
   not MGM_G306(MGM_W255,den_delay);
   and MGM_G307(MGM_W256,MGM_W255,MGM_W254);
   and MGM_G308(MGM_W257,si_delay,MGM_W256);
   and MGM_G309(ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W257);
   and MGM_G310(MGM_W258,d_delay,clk_delay);
   and MGM_G311(MGM_W259,den_delay,MGM_W258);
   not MGM_G312(MGM_W260,si_delay);
   and MGM_G313(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G314(MGM_W262,ssb_delay);
   and MGM_G315(ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   and MGM_G316(MGM_W263,d_delay,clk_delay);
   and MGM_G317(MGM_W264,den_delay,MGM_W263);
   not MGM_G318(MGM_W265,si_delay);
   and MGM_G319(MGM_W266,MGM_W265,MGM_W264);
   and MGM_G320(ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W266);
   and MGM_G321(MGM_W267,d_delay,clk_delay);
   and MGM_G322(MGM_W268,den_delay,MGM_W267);
   and MGM_G323(MGM_W269,si_delay,MGM_W268);
   not MGM_G324(MGM_W270,ssb_delay);
   and MGM_G325(ENABLE_clk_AND_d_AND_den_AND_si_AND_NOT_ssb,MGM_W270,MGM_W269);
   and MGM_G326(MGM_W271,d_delay,clk_delay);
   and MGM_G327(MGM_W272,den_delay,MGM_W271);
   and MGM_G328(MGM_W273,si_delay,MGM_W272);
   and MGM_G329(ENABLE_clk_AND_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W273);
   not MGM_G330(MGM_W274,d_delay);
   not MGM_G331(MGM_W275,den_delay);
   and MGM_G332(MGM_W276,MGM_W275,MGM_W274);
   and MGM_G333(MGM_W277,rb_delay,MGM_W276);
   not MGM_G334(MGM_W278,ssb_delay);
   and MGM_G335(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb,MGM_W278,MGM_W277);
   not MGM_G336(MGM_W279,d_delay);
   and MGM_G337(MGM_W280,den_delay,MGM_W279);
   and MGM_G338(MGM_W281,rb_delay,MGM_W280);
   not MGM_G339(MGM_W282,ssb_delay);
   and MGM_G340(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb,MGM_W282,MGM_W281);
   not MGM_G341(MGM_W283,den_delay);
   and MGM_G342(MGM_W284,MGM_W283,d_delay);
   and MGM_G343(MGM_W285,rb_delay,MGM_W284);
   not MGM_G344(MGM_W286,ssb_delay);
   and MGM_G345(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb,MGM_W286,MGM_W285);
   and MGM_G346(MGM_W287,den_delay,d_delay);
   and MGM_G347(MGM_W288,rb_delay,MGM_W287);
   not MGM_G348(MGM_W289,ssb_delay);
   and MGM_G349(ENABLE_d_AND_den_AND_rb_AND_NOT_ssb,MGM_W289,MGM_W288);
   not MGM_G350(MGM_W290,d_delay);
   not MGM_G351(MGM_W291,den_delay);
   and MGM_G352(MGM_W292,MGM_W291,MGM_W290);
   and MGM_G353(MGM_W293,rb_delay,MGM_W292);
   not MGM_G354(MGM_W294,si_delay);
   and MGM_G355(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si,MGM_W294,MGM_W293);
   not MGM_G356(MGM_W295,d_delay);
   not MGM_G357(MGM_W296,den_delay);
   and MGM_G358(MGM_W297,MGM_W296,MGM_W295);
   and MGM_G359(MGM_W298,rb_delay,MGM_W297);
   and MGM_G360(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si,si_delay,MGM_W298);
   not MGM_G361(MGM_W299,d_delay);
   and MGM_G362(MGM_W300,den_delay,MGM_W299);
   and MGM_G363(MGM_W301,rb_delay,MGM_W300);
   and MGM_G364(ENABLE_NOT_d_AND_den_AND_rb_AND_si,si_delay,MGM_W301);
   not MGM_G365(MGM_W302,den_delay);
   and MGM_G366(MGM_W303,MGM_W302,d_delay);
   and MGM_G367(MGM_W304,rb_delay,MGM_W303);
   not MGM_G368(MGM_W305,si_delay);
   and MGM_G369(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   not MGM_G370(MGM_W306,den_delay);
   and MGM_G371(MGM_W307,MGM_W306,d_delay);
   and MGM_G372(MGM_W308,rb_delay,MGM_W307);
   and MGM_G373(ENABLE_d_AND_NOT_den_AND_rb_AND_si,si_delay,MGM_W308);
   and MGM_G374(MGM_W309,den_delay,d_delay);
   and MGM_G375(MGM_W310,rb_delay,MGM_W309);
   not MGM_G376(MGM_W311,si_delay);
   and MGM_G377(ENABLE_d_AND_den_AND_rb_AND_NOT_si,MGM_W311,MGM_W310);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy043ah1n06x5( clk, d, den, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy043ah_func b15fqy043ah1n06x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy043ah_func b15fqy043ah1n06x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy043ah_func b15fqy043ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy043ah_func b15fqy043ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,den_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   and MGM_G3(MGM_W3,rb_delay,MGM_W2);
   not MGM_G4(MGM_W4,si_delay);
   and MGM_G5(MGM_W5,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W6,ssb_delay);
   and MGM_G7(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W6,MGM_W5);
   not MGM_G8(MGM_W7,d_delay);
   not MGM_G9(MGM_W8,den_delay);
   and MGM_G10(MGM_W9,MGM_W8,MGM_W7);
   and MGM_G11(MGM_W10,rb_delay,MGM_W9);
   and MGM_G12(MGM_W11,si_delay,MGM_W10);
   not MGM_G13(MGM_W12,ssb_delay);
   and MGM_G14(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G15(MGM_W13,d_delay);
   and MGM_G16(MGM_W14,den_delay,MGM_W13);
   and MGM_G17(MGM_W15,rb_delay,MGM_W14);
   not MGM_G18(MGM_W16,si_delay);
   and MGM_G19(MGM_W17,MGM_W16,MGM_W15);
   not MGM_G20(MGM_W18,ssb_delay);
   and MGM_G21(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   not MGM_G22(MGM_W19,d_delay);
   and MGM_G23(MGM_W20,den_delay,MGM_W19);
   and MGM_G24(MGM_W21,rb_delay,MGM_W20);
   not MGM_G25(MGM_W22,si_delay);
   and MGM_G26(MGM_W23,MGM_W22,MGM_W21);
   and MGM_G27(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W23);
   not MGM_G28(MGM_W24,d_delay);
   and MGM_G29(MGM_W25,den_delay,MGM_W24);
   and MGM_G30(MGM_W26,rb_delay,MGM_W25);
   and MGM_G31(MGM_W27,si_delay,MGM_W26);
   not MGM_G32(MGM_W28,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W28,MGM_W27);
   not MGM_G34(MGM_W29,d_delay);
   and MGM_G35(MGM_W30,den_delay,MGM_W29);
   and MGM_G36(MGM_W31,rb_delay,MGM_W30);
   and MGM_G37(MGM_W32,si_delay,MGM_W31);
   and MGM_G38(ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W32);
   not MGM_G39(MGM_W33,den_delay);
   and MGM_G40(MGM_W34,MGM_W33,d_delay);
   and MGM_G41(MGM_W35,rb_delay,MGM_W34);
   not MGM_G42(MGM_W36,si_delay);
   and MGM_G43(MGM_W37,MGM_W36,MGM_W35);
   not MGM_G44(MGM_W38,ssb_delay);
   and MGM_G45(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W38,MGM_W37);
   not MGM_G46(MGM_W39,den_delay);
   and MGM_G47(MGM_W40,MGM_W39,d_delay);
   and MGM_G48(MGM_W41,rb_delay,MGM_W40);
   and MGM_G49(MGM_W42,si_delay,MGM_W41);
   not MGM_G50(MGM_W43,ssb_delay);
   and MGM_G51(ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W43,MGM_W42);
   and MGM_G52(MGM_W44,den_delay,d_delay);
   and MGM_G53(MGM_W45,rb_delay,MGM_W44);
   not MGM_G54(MGM_W46,si_delay);
   and MGM_G55(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G56(MGM_W48,ssb_delay);
   and MGM_G57(ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   and MGM_G58(MGM_W49,den_delay,d_delay);
   and MGM_G59(MGM_W50,rb_delay,MGM_W49);
   not MGM_G60(MGM_W51,si_delay);
   and MGM_G61(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G62(ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G63(MGM_W53,den_delay,d_delay);
   and MGM_G64(MGM_W54,rb_delay,MGM_W53);
   and MGM_G65(MGM_W55,si_delay,MGM_W54);
   not MGM_G66(MGM_W56,ssb_delay);
   and MGM_G67(ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   and MGM_G68(MGM_W57,den_delay,d_delay);
   and MGM_G69(MGM_W58,rb_delay,MGM_W57);
   and MGM_G70(MGM_W59,si_delay,MGM_W58);
   and MGM_G71(ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W59);
   and MGM_G72(MGM_W60,rb_delay,den_delay);
   not MGM_G73(MGM_W61,si_delay);
   and MGM_G74(MGM_W62,MGM_W61,MGM_W60);
   and MGM_G75(ENABLE_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W62);
   and MGM_G76(MGM_W63,rb_delay,den_delay);
   and MGM_G77(MGM_W64,si_delay,MGM_W63);
   and MGM_G78(ENABLE_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W64);
   not MGM_G79(MGM_W65,d_delay);
   and MGM_G80(MGM_W66,rb_delay,MGM_W65);
   not MGM_G81(MGM_W67,si_delay);
   and MGM_G82(MGM_W68,MGM_W67,MGM_W66);
   and MGM_G83(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W68);
   not MGM_G84(MGM_W69,d_delay);
   and MGM_G85(MGM_W70,rb_delay,MGM_W69);
   and MGM_G86(MGM_W71,si_delay,MGM_W70);
   and MGM_G87(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W71);
   and MGM_G88(MGM_W72,rb_delay,d_delay);
   not MGM_G89(MGM_W73,si_delay);
   and MGM_G90(MGM_W74,MGM_W73,MGM_W72);
   and MGM_G91(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W74);
   and MGM_G92(MGM_W75,rb_delay,d_delay);
   and MGM_G93(MGM_W76,si_delay,MGM_W75);
   and MGM_G94(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W76);
   not MGM_G95(MGM_W77,d_delay);
   not MGM_G96(MGM_W78,den_delay);
   and MGM_G97(MGM_W79,MGM_W78,MGM_W77);
   and MGM_G98(MGM_W80,si_delay,MGM_W79);
   not MGM_G99(MGM_W81,ssb_delay);
   and MGM_G100(ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W81,MGM_W80);
   not MGM_G101(MGM_W82,d_delay);
   and MGM_G102(MGM_W83,den_delay,MGM_W82);
   and MGM_G103(MGM_W84,si_delay,MGM_W83);
   not MGM_G104(MGM_W85,ssb_delay);
   and MGM_G105(ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W85,MGM_W84);
   not MGM_G106(MGM_W86,den_delay);
   and MGM_G107(MGM_W87,MGM_W86,d_delay);
   and MGM_G108(MGM_W88,si_delay,MGM_W87);
   not MGM_G109(MGM_W89,ssb_delay);
   and MGM_G110(ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W89,MGM_W88);
   and MGM_G111(MGM_W90,den_delay,d_delay);
   not MGM_G112(MGM_W91,si_delay);
   and MGM_G113(MGM_W92,MGM_W91,MGM_W90);
   and MGM_G114(ENABLE_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W92);
   and MGM_G115(MGM_W93,den_delay,d_delay);
   and MGM_G116(MGM_W94,si_delay,MGM_W93);
   not MGM_G117(MGM_W95,ssb_delay);
   and MGM_G118(ENABLE_d_AND_den_AND_si_AND_NOT_ssb,MGM_W95,MGM_W94);
   and MGM_G119(MGM_W96,den_delay,d_delay);
   and MGM_G120(MGM_W97,si_delay,MGM_W96);
   and MGM_G121(ENABLE_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W97);
   not MGM_G122(MGM_W98,clk_delay);
   not MGM_G123(MGM_W99,d_delay);
   and MGM_G124(MGM_W100,MGM_W99,MGM_W98);
   not MGM_G125(MGM_W101,den_delay);
   and MGM_G126(MGM_W102,MGM_W101,MGM_W100);
   not MGM_G127(MGM_W103,si_delay);
   and MGM_G128(MGM_W104,MGM_W103,MGM_W102);
   not MGM_G129(MGM_W105,ssb_delay);
   and MGM_G130(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W105,MGM_W104);
   not MGM_G131(MGM_W106,clk_delay);
   not MGM_G132(MGM_W107,d_delay);
   and MGM_G133(MGM_W108,MGM_W107,MGM_W106);
   not MGM_G134(MGM_W109,den_delay);
   and MGM_G135(MGM_W110,MGM_W109,MGM_W108);
   not MGM_G136(MGM_W111,si_delay);
   and MGM_G137(MGM_W112,MGM_W111,MGM_W110);
   and MGM_G138(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W112);
   not MGM_G139(MGM_W113,clk_delay);
   not MGM_G140(MGM_W114,d_delay);
   and MGM_G141(MGM_W115,MGM_W114,MGM_W113);
   not MGM_G142(MGM_W116,den_delay);
   and MGM_G143(MGM_W117,MGM_W116,MGM_W115);
   and MGM_G144(MGM_W118,si_delay,MGM_W117);
   not MGM_G145(MGM_W119,ssb_delay);
   and MGM_G146(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W119,MGM_W118);
   not MGM_G147(MGM_W120,clk_delay);
   not MGM_G148(MGM_W121,d_delay);
   and MGM_G149(MGM_W122,MGM_W121,MGM_W120);
   not MGM_G150(MGM_W123,den_delay);
   and MGM_G151(MGM_W124,MGM_W123,MGM_W122);
   and MGM_G152(MGM_W125,si_delay,MGM_W124);
   and MGM_G153(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W125);
   not MGM_G154(MGM_W126,clk_delay);
   not MGM_G155(MGM_W127,d_delay);
   and MGM_G156(MGM_W128,MGM_W127,MGM_W126);
   and MGM_G157(MGM_W129,den_delay,MGM_W128);
   not MGM_G158(MGM_W130,si_delay);
   and MGM_G159(MGM_W131,MGM_W130,MGM_W129);
   not MGM_G160(MGM_W132,ssb_delay);
   and MGM_G161(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W132,MGM_W131);
   not MGM_G162(MGM_W133,clk_delay);
   not MGM_G163(MGM_W134,d_delay);
   and MGM_G164(MGM_W135,MGM_W134,MGM_W133);
   and MGM_G165(MGM_W136,den_delay,MGM_W135);
   not MGM_G166(MGM_W137,si_delay);
   and MGM_G167(MGM_W138,MGM_W137,MGM_W136);
   and MGM_G168(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W138);
   not MGM_G169(MGM_W139,clk_delay);
   not MGM_G170(MGM_W140,d_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   and MGM_G172(MGM_W142,den_delay,MGM_W141);
   and MGM_G173(MGM_W143,si_delay,MGM_W142);
   not MGM_G174(MGM_W144,ssb_delay);
   and MGM_G175(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W144,MGM_W143);
   not MGM_G176(MGM_W145,clk_delay);
   not MGM_G177(MGM_W146,d_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(MGM_W148,den_delay,MGM_W147);
   and MGM_G180(MGM_W149,si_delay,MGM_W148);
   and MGM_G181(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W149);
   not MGM_G182(MGM_W150,clk_delay);
   and MGM_G183(MGM_W151,d_delay,MGM_W150);
   not MGM_G184(MGM_W152,den_delay);
   and MGM_G185(MGM_W153,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W154,si_delay);
   and MGM_G187(MGM_W155,MGM_W154,MGM_W153);
   not MGM_G188(MGM_W156,ssb_delay);
   and MGM_G189(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W156,MGM_W155);
   not MGM_G190(MGM_W157,clk_delay);
   and MGM_G191(MGM_W158,d_delay,MGM_W157);
   not MGM_G192(MGM_W159,den_delay);
   and MGM_G193(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G194(MGM_W161,si_delay);
   and MGM_G195(MGM_W162,MGM_W161,MGM_W160);
   and MGM_G196(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W162);
   not MGM_G197(MGM_W163,clk_delay);
   and MGM_G198(MGM_W164,d_delay,MGM_W163);
   not MGM_G199(MGM_W165,den_delay);
   and MGM_G200(MGM_W166,MGM_W165,MGM_W164);
   and MGM_G201(MGM_W167,si_delay,MGM_W166);
   not MGM_G202(MGM_W168,ssb_delay);
   and MGM_G203(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W168,MGM_W167);
   not MGM_G204(MGM_W169,clk_delay);
   and MGM_G205(MGM_W170,d_delay,MGM_W169);
   not MGM_G206(MGM_W171,den_delay);
   and MGM_G207(MGM_W172,MGM_W171,MGM_W170);
   and MGM_G208(MGM_W173,si_delay,MGM_W172);
   and MGM_G209(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W173);
   not MGM_G210(MGM_W174,clk_delay);
   and MGM_G211(MGM_W175,d_delay,MGM_W174);
   and MGM_G212(MGM_W176,den_delay,MGM_W175);
   not MGM_G213(MGM_W177,si_delay);
   and MGM_G214(MGM_W178,MGM_W177,MGM_W176);
   not MGM_G215(MGM_W179,ssb_delay);
   and MGM_G216(ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W179,MGM_W178);
   not MGM_G217(MGM_W180,clk_delay);
   and MGM_G218(MGM_W181,d_delay,MGM_W180);
   and MGM_G219(MGM_W182,den_delay,MGM_W181);
   not MGM_G220(MGM_W183,si_delay);
   and MGM_G221(MGM_W184,MGM_W183,MGM_W182);
   and MGM_G222(ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W184);
   not MGM_G223(MGM_W185,clk_delay);
   and MGM_G224(MGM_W186,d_delay,MGM_W185);
   and MGM_G225(MGM_W187,den_delay,MGM_W186);
   and MGM_G226(MGM_W188,si_delay,MGM_W187);
   not MGM_G227(MGM_W189,ssb_delay);
   and MGM_G228(ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_NOT_ssb,MGM_W189,MGM_W188);
   not MGM_G229(MGM_W190,clk_delay);
   and MGM_G230(MGM_W191,d_delay,MGM_W190);
   and MGM_G231(MGM_W192,den_delay,MGM_W191);
   and MGM_G232(MGM_W193,si_delay,MGM_W192);
   and MGM_G233(ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W193);
   not MGM_G234(MGM_W194,d_delay);
   and MGM_G235(MGM_W195,MGM_W194,clk_delay);
   not MGM_G236(MGM_W196,den_delay);
   and MGM_G237(MGM_W197,MGM_W196,MGM_W195);
   not MGM_G238(MGM_W198,si_delay);
   and MGM_G239(MGM_W199,MGM_W198,MGM_W197);
   not MGM_G240(MGM_W200,ssb_delay);
   and MGM_G241(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W200,MGM_W199);
   not MGM_G242(MGM_W201,d_delay);
   and MGM_G243(MGM_W202,MGM_W201,clk_delay);
   not MGM_G244(MGM_W203,den_delay);
   and MGM_G245(MGM_W204,MGM_W203,MGM_W202);
   not MGM_G246(MGM_W205,si_delay);
   and MGM_G247(MGM_W206,MGM_W205,MGM_W204);
   and MGM_G248(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W206);
   not MGM_G249(MGM_W207,d_delay);
   and MGM_G250(MGM_W208,MGM_W207,clk_delay);
   not MGM_G251(MGM_W209,den_delay);
   and MGM_G252(MGM_W210,MGM_W209,MGM_W208);
   and MGM_G253(MGM_W211,si_delay,MGM_W210);
   not MGM_G254(MGM_W212,ssb_delay);
   and MGM_G255(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W212,MGM_W211);
   not MGM_G256(MGM_W213,d_delay);
   and MGM_G257(MGM_W214,MGM_W213,clk_delay);
   not MGM_G258(MGM_W215,den_delay);
   and MGM_G259(MGM_W216,MGM_W215,MGM_W214);
   and MGM_G260(MGM_W217,si_delay,MGM_W216);
   and MGM_G261(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W217);
   not MGM_G262(MGM_W218,d_delay);
   and MGM_G263(MGM_W219,MGM_W218,clk_delay);
   and MGM_G264(MGM_W220,den_delay,MGM_W219);
   not MGM_G265(MGM_W221,si_delay);
   and MGM_G266(MGM_W222,MGM_W221,MGM_W220);
   not MGM_G267(MGM_W223,ssb_delay);
   and MGM_G268(ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W223,MGM_W222);
   not MGM_G269(MGM_W224,d_delay);
   and MGM_G270(MGM_W225,MGM_W224,clk_delay);
   and MGM_G271(MGM_W226,den_delay,MGM_W225);
   not MGM_G272(MGM_W227,si_delay);
   and MGM_G273(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G274(ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W228);
   not MGM_G275(MGM_W229,d_delay);
   and MGM_G276(MGM_W230,MGM_W229,clk_delay);
   and MGM_G277(MGM_W231,den_delay,MGM_W230);
   and MGM_G278(MGM_W232,si_delay,MGM_W231);
   not MGM_G279(MGM_W233,ssb_delay);
   and MGM_G280(ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W233,MGM_W232);
   not MGM_G281(MGM_W234,d_delay);
   and MGM_G282(MGM_W235,MGM_W234,clk_delay);
   and MGM_G283(MGM_W236,den_delay,MGM_W235);
   and MGM_G284(MGM_W237,si_delay,MGM_W236);
   and MGM_G285(ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W237);
   and MGM_G286(MGM_W238,d_delay,clk_delay);
   not MGM_G287(MGM_W239,den_delay);
   and MGM_G288(MGM_W240,MGM_W239,MGM_W238);
   not MGM_G289(MGM_W241,si_delay);
   and MGM_G290(MGM_W242,MGM_W241,MGM_W240);
   not MGM_G291(MGM_W243,ssb_delay);
   and MGM_G292(ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W243,MGM_W242);
   and MGM_G293(MGM_W244,d_delay,clk_delay);
   not MGM_G294(MGM_W245,den_delay);
   and MGM_G295(MGM_W246,MGM_W245,MGM_W244);
   not MGM_G296(MGM_W247,si_delay);
   and MGM_G297(MGM_W248,MGM_W247,MGM_W246);
   and MGM_G298(ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W248);
   and MGM_G299(MGM_W249,d_delay,clk_delay);
   not MGM_G300(MGM_W250,den_delay);
   and MGM_G301(MGM_W251,MGM_W250,MGM_W249);
   and MGM_G302(MGM_W252,si_delay,MGM_W251);
   not MGM_G303(MGM_W253,ssb_delay);
   and MGM_G304(ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W253,MGM_W252);
   and MGM_G305(MGM_W254,d_delay,clk_delay);
   not MGM_G306(MGM_W255,den_delay);
   and MGM_G307(MGM_W256,MGM_W255,MGM_W254);
   and MGM_G308(MGM_W257,si_delay,MGM_W256);
   and MGM_G309(ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W257);
   and MGM_G310(MGM_W258,d_delay,clk_delay);
   and MGM_G311(MGM_W259,den_delay,MGM_W258);
   not MGM_G312(MGM_W260,si_delay);
   and MGM_G313(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G314(MGM_W262,ssb_delay);
   and MGM_G315(ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   and MGM_G316(MGM_W263,d_delay,clk_delay);
   and MGM_G317(MGM_W264,den_delay,MGM_W263);
   not MGM_G318(MGM_W265,si_delay);
   and MGM_G319(MGM_W266,MGM_W265,MGM_W264);
   and MGM_G320(ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W266);
   and MGM_G321(MGM_W267,d_delay,clk_delay);
   and MGM_G322(MGM_W268,den_delay,MGM_W267);
   and MGM_G323(MGM_W269,si_delay,MGM_W268);
   not MGM_G324(MGM_W270,ssb_delay);
   and MGM_G325(ENABLE_clk_AND_d_AND_den_AND_si_AND_NOT_ssb,MGM_W270,MGM_W269);
   and MGM_G326(MGM_W271,d_delay,clk_delay);
   and MGM_G327(MGM_W272,den_delay,MGM_W271);
   and MGM_G328(MGM_W273,si_delay,MGM_W272);
   and MGM_G329(ENABLE_clk_AND_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W273);
   not MGM_G330(MGM_W274,d_delay);
   not MGM_G331(MGM_W275,den_delay);
   and MGM_G332(MGM_W276,MGM_W275,MGM_W274);
   and MGM_G333(MGM_W277,rb_delay,MGM_W276);
   not MGM_G334(MGM_W278,ssb_delay);
   and MGM_G335(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb,MGM_W278,MGM_W277);
   not MGM_G336(MGM_W279,d_delay);
   and MGM_G337(MGM_W280,den_delay,MGM_W279);
   and MGM_G338(MGM_W281,rb_delay,MGM_W280);
   not MGM_G339(MGM_W282,ssb_delay);
   and MGM_G340(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb,MGM_W282,MGM_W281);
   not MGM_G341(MGM_W283,den_delay);
   and MGM_G342(MGM_W284,MGM_W283,d_delay);
   and MGM_G343(MGM_W285,rb_delay,MGM_W284);
   not MGM_G344(MGM_W286,ssb_delay);
   and MGM_G345(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb,MGM_W286,MGM_W285);
   and MGM_G346(MGM_W287,den_delay,d_delay);
   and MGM_G347(MGM_W288,rb_delay,MGM_W287);
   not MGM_G348(MGM_W289,ssb_delay);
   and MGM_G349(ENABLE_d_AND_den_AND_rb_AND_NOT_ssb,MGM_W289,MGM_W288);
   not MGM_G350(MGM_W290,d_delay);
   not MGM_G351(MGM_W291,den_delay);
   and MGM_G352(MGM_W292,MGM_W291,MGM_W290);
   and MGM_G353(MGM_W293,rb_delay,MGM_W292);
   not MGM_G354(MGM_W294,si_delay);
   and MGM_G355(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si,MGM_W294,MGM_W293);
   not MGM_G356(MGM_W295,d_delay);
   not MGM_G357(MGM_W296,den_delay);
   and MGM_G358(MGM_W297,MGM_W296,MGM_W295);
   and MGM_G359(MGM_W298,rb_delay,MGM_W297);
   and MGM_G360(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si,si_delay,MGM_W298);
   not MGM_G361(MGM_W299,d_delay);
   and MGM_G362(MGM_W300,den_delay,MGM_W299);
   and MGM_G363(MGM_W301,rb_delay,MGM_W300);
   and MGM_G364(ENABLE_NOT_d_AND_den_AND_rb_AND_si,si_delay,MGM_W301);
   not MGM_G365(MGM_W302,den_delay);
   and MGM_G366(MGM_W303,MGM_W302,d_delay);
   and MGM_G367(MGM_W304,rb_delay,MGM_W303);
   not MGM_G368(MGM_W305,si_delay);
   and MGM_G369(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   not MGM_G370(MGM_W306,den_delay);
   and MGM_G371(MGM_W307,MGM_W306,d_delay);
   and MGM_G372(MGM_W308,rb_delay,MGM_W307);
   and MGM_G373(ENABLE_d_AND_NOT_den_AND_rb_AND_si,si_delay,MGM_W308);
   and MGM_G374(MGM_W309,den_delay,d_delay);
   and MGM_G375(MGM_W310,rb_delay,MGM_W309);
   not MGM_G376(MGM_W311,si_delay);
   and MGM_G377(ENABLE_d_AND_den_AND_rb_AND_NOT_si,MGM_W311,MGM_W310);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy043ah1n08x5( clk, d, den, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy043ah_func b15fqy043ah1n08x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy043ah_func b15fqy043ah1n08x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy043ah_func b15fqy043ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy043ah_func b15fqy043ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,den_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   and MGM_G3(MGM_W3,rb_delay,MGM_W2);
   not MGM_G4(MGM_W4,si_delay);
   and MGM_G5(MGM_W5,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W6,ssb_delay);
   and MGM_G7(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W6,MGM_W5);
   not MGM_G8(MGM_W7,d_delay);
   not MGM_G9(MGM_W8,den_delay);
   and MGM_G10(MGM_W9,MGM_W8,MGM_W7);
   and MGM_G11(MGM_W10,rb_delay,MGM_W9);
   and MGM_G12(MGM_W11,si_delay,MGM_W10);
   not MGM_G13(MGM_W12,ssb_delay);
   and MGM_G14(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G15(MGM_W13,d_delay);
   and MGM_G16(MGM_W14,den_delay,MGM_W13);
   and MGM_G17(MGM_W15,rb_delay,MGM_W14);
   not MGM_G18(MGM_W16,si_delay);
   and MGM_G19(MGM_W17,MGM_W16,MGM_W15);
   not MGM_G20(MGM_W18,ssb_delay);
   and MGM_G21(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   not MGM_G22(MGM_W19,d_delay);
   and MGM_G23(MGM_W20,den_delay,MGM_W19);
   and MGM_G24(MGM_W21,rb_delay,MGM_W20);
   not MGM_G25(MGM_W22,si_delay);
   and MGM_G26(MGM_W23,MGM_W22,MGM_W21);
   and MGM_G27(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W23);
   not MGM_G28(MGM_W24,d_delay);
   and MGM_G29(MGM_W25,den_delay,MGM_W24);
   and MGM_G30(MGM_W26,rb_delay,MGM_W25);
   and MGM_G31(MGM_W27,si_delay,MGM_W26);
   not MGM_G32(MGM_W28,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W28,MGM_W27);
   not MGM_G34(MGM_W29,d_delay);
   and MGM_G35(MGM_W30,den_delay,MGM_W29);
   and MGM_G36(MGM_W31,rb_delay,MGM_W30);
   and MGM_G37(MGM_W32,si_delay,MGM_W31);
   and MGM_G38(ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W32);
   not MGM_G39(MGM_W33,den_delay);
   and MGM_G40(MGM_W34,MGM_W33,d_delay);
   and MGM_G41(MGM_W35,rb_delay,MGM_W34);
   not MGM_G42(MGM_W36,si_delay);
   and MGM_G43(MGM_W37,MGM_W36,MGM_W35);
   not MGM_G44(MGM_W38,ssb_delay);
   and MGM_G45(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W38,MGM_W37);
   not MGM_G46(MGM_W39,den_delay);
   and MGM_G47(MGM_W40,MGM_W39,d_delay);
   and MGM_G48(MGM_W41,rb_delay,MGM_W40);
   and MGM_G49(MGM_W42,si_delay,MGM_W41);
   not MGM_G50(MGM_W43,ssb_delay);
   and MGM_G51(ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W43,MGM_W42);
   and MGM_G52(MGM_W44,den_delay,d_delay);
   and MGM_G53(MGM_W45,rb_delay,MGM_W44);
   not MGM_G54(MGM_W46,si_delay);
   and MGM_G55(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G56(MGM_W48,ssb_delay);
   and MGM_G57(ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   and MGM_G58(MGM_W49,den_delay,d_delay);
   and MGM_G59(MGM_W50,rb_delay,MGM_W49);
   not MGM_G60(MGM_W51,si_delay);
   and MGM_G61(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G62(ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G63(MGM_W53,den_delay,d_delay);
   and MGM_G64(MGM_W54,rb_delay,MGM_W53);
   and MGM_G65(MGM_W55,si_delay,MGM_W54);
   not MGM_G66(MGM_W56,ssb_delay);
   and MGM_G67(ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   and MGM_G68(MGM_W57,den_delay,d_delay);
   and MGM_G69(MGM_W58,rb_delay,MGM_W57);
   and MGM_G70(MGM_W59,si_delay,MGM_W58);
   and MGM_G71(ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W59);
   and MGM_G72(MGM_W60,rb_delay,den_delay);
   not MGM_G73(MGM_W61,si_delay);
   and MGM_G74(MGM_W62,MGM_W61,MGM_W60);
   and MGM_G75(ENABLE_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W62);
   and MGM_G76(MGM_W63,rb_delay,den_delay);
   and MGM_G77(MGM_W64,si_delay,MGM_W63);
   and MGM_G78(ENABLE_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W64);
   not MGM_G79(MGM_W65,d_delay);
   and MGM_G80(MGM_W66,rb_delay,MGM_W65);
   not MGM_G81(MGM_W67,si_delay);
   and MGM_G82(MGM_W68,MGM_W67,MGM_W66);
   and MGM_G83(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W68);
   not MGM_G84(MGM_W69,d_delay);
   and MGM_G85(MGM_W70,rb_delay,MGM_W69);
   and MGM_G86(MGM_W71,si_delay,MGM_W70);
   and MGM_G87(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W71);
   and MGM_G88(MGM_W72,rb_delay,d_delay);
   not MGM_G89(MGM_W73,si_delay);
   and MGM_G90(MGM_W74,MGM_W73,MGM_W72);
   and MGM_G91(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W74);
   and MGM_G92(MGM_W75,rb_delay,d_delay);
   and MGM_G93(MGM_W76,si_delay,MGM_W75);
   and MGM_G94(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W76);
   not MGM_G95(MGM_W77,d_delay);
   not MGM_G96(MGM_W78,den_delay);
   and MGM_G97(MGM_W79,MGM_W78,MGM_W77);
   and MGM_G98(MGM_W80,si_delay,MGM_W79);
   not MGM_G99(MGM_W81,ssb_delay);
   and MGM_G100(ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W81,MGM_W80);
   not MGM_G101(MGM_W82,d_delay);
   and MGM_G102(MGM_W83,den_delay,MGM_W82);
   and MGM_G103(MGM_W84,si_delay,MGM_W83);
   not MGM_G104(MGM_W85,ssb_delay);
   and MGM_G105(ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W85,MGM_W84);
   not MGM_G106(MGM_W86,den_delay);
   and MGM_G107(MGM_W87,MGM_W86,d_delay);
   and MGM_G108(MGM_W88,si_delay,MGM_W87);
   not MGM_G109(MGM_W89,ssb_delay);
   and MGM_G110(ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W89,MGM_W88);
   and MGM_G111(MGM_W90,den_delay,d_delay);
   not MGM_G112(MGM_W91,si_delay);
   and MGM_G113(MGM_W92,MGM_W91,MGM_W90);
   and MGM_G114(ENABLE_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W92);
   and MGM_G115(MGM_W93,den_delay,d_delay);
   and MGM_G116(MGM_W94,si_delay,MGM_W93);
   not MGM_G117(MGM_W95,ssb_delay);
   and MGM_G118(ENABLE_d_AND_den_AND_si_AND_NOT_ssb,MGM_W95,MGM_W94);
   and MGM_G119(MGM_W96,den_delay,d_delay);
   and MGM_G120(MGM_W97,si_delay,MGM_W96);
   and MGM_G121(ENABLE_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W97);
   not MGM_G122(MGM_W98,clk_delay);
   not MGM_G123(MGM_W99,d_delay);
   and MGM_G124(MGM_W100,MGM_W99,MGM_W98);
   not MGM_G125(MGM_W101,den_delay);
   and MGM_G126(MGM_W102,MGM_W101,MGM_W100);
   not MGM_G127(MGM_W103,si_delay);
   and MGM_G128(MGM_W104,MGM_W103,MGM_W102);
   not MGM_G129(MGM_W105,ssb_delay);
   and MGM_G130(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W105,MGM_W104);
   not MGM_G131(MGM_W106,clk_delay);
   not MGM_G132(MGM_W107,d_delay);
   and MGM_G133(MGM_W108,MGM_W107,MGM_W106);
   not MGM_G134(MGM_W109,den_delay);
   and MGM_G135(MGM_W110,MGM_W109,MGM_W108);
   not MGM_G136(MGM_W111,si_delay);
   and MGM_G137(MGM_W112,MGM_W111,MGM_W110);
   and MGM_G138(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W112);
   not MGM_G139(MGM_W113,clk_delay);
   not MGM_G140(MGM_W114,d_delay);
   and MGM_G141(MGM_W115,MGM_W114,MGM_W113);
   not MGM_G142(MGM_W116,den_delay);
   and MGM_G143(MGM_W117,MGM_W116,MGM_W115);
   and MGM_G144(MGM_W118,si_delay,MGM_W117);
   not MGM_G145(MGM_W119,ssb_delay);
   and MGM_G146(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W119,MGM_W118);
   not MGM_G147(MGM_W120,clk_delay);
   not MGM_G148(MGM_W121,d_delay);
   and MGM_G149(MGM_W122,MGM_W121,MGM_W120);
   not MGM_G150(MGM_W123,den_delay);
   and MGM_G151(MGM_W124,MGM_W123,MGM_W122);
   and MGM_G152(MGM_W125,si_delay,MGM_W124);
   and MGM_G153(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W125);
   not MGM_G154(MGM_W126,clk_delay);
   not MGM_G155(MGM_W127,d_delay);
   and MGM_G156(MGM_W128,MGM_W127,MGM_W126);
   and MGM_G157(MGM_W129,den_delay,MGM_W128);
   not MGM_G158(MGM_W130,si_delay);
   and MGM_G159(MGM_W131,MGM_W130,MGM_W129);
   not MGM_G160(MGM_W132,ssb_delay);
   and MGM_G161(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W132,MGM_W131);
   not MGM_G162(MGM_W133,clk_delay);
   not MGM_G163(MGM_W134,d_delay);
   and MGM_G164(MGM_W135,MGM_W134,MGM_W133);
   and MGM_G165(MGM_W136,den_delay,MGM_W135);
   not MGM_G166(MGM_W137,si_delay);
   and MGM_G167(MGM_W138,MGM_W137,MGM_W136);
   and MGM_G168(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W138);
   not MGM_G169(MGM_W139,clk_delay);
   not MGM_G170(MGM_W140,d_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   and MGM_G172(MGM_W142,den_delay,MGM_W141);
   and MGM_G173(MGM_W143,si_delay,MGM_W142);
   not MGM_G174(MGM_W144,ssb_delay);
   and MGM_G175(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W144,MGM_W143);
   not MGM_G176(MGM_W145,clk_delay);
   not MGM_G177(MGM_W146,d_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(MGM_W148,den_delay,MGM_W147);
   and MGM_G180(MGM_W149,si_delay,MGM_W148);
   and MGM_G181(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W149);
   not MGM_G182(MGM_W150,clk_delay);
   and MGM_G183(MGM_W151,d_delay,MGM_W150);
   not MGM_G184(MGM_W152,den_delay);
   and MGM_G185(MGM_W153,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W154,si_delay);
   and MGM_G187(MGM_W155,MGM_W154,MGM_W153);
   not MGM_G188(MGM_W156,ssb_delay);
   and MGM_G189(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W156,MGM_W155);
   not MGM_G190(MGM_W157,clk_delay);
   and MGM_G191(MGM_W158,d_delay,MGM_W157);
   not MGM_G192(MGM_W159,den_delay);
   and MGM_G193(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G194(MGM_W161,si_delay);
   and MGM_G195(MGM_W162,MGM_W161,MGM_W160);
   and MGM_G196(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W162);
   not MGM_G197(MGM_W163,clk_delay);
   and MGM_G198(MGM_W164,d_delay,MGM_W163);
   not MGM_G199(MGM_W165,den_delay);
   and MGM_G200(MGM_W166,MGM_W165,MGM_W164);
   and MGM_G201(MGM_W167,si_delay,MGM_W166);
   not MGM_G202(MGM_W168,ssb_delay);
   and MGM_G203(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W168,MGM_W167);
   not MGM_G204(MGM_W169,clk_delay);
   and MGM_G205(MGM_W170,d_delay,MGM_W169);
   not MGM_G206(MGM_W171,den_delay);
   and MGM_G207(MGM_W172,MGM_W171,MGM_W170);
   and MGM_G208(MGM_W173,si_delay,MGM_W172);
   and MGM_G209(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W173);
   not MGM_G210(MGM_W174,clk_delay);
   and MGM_G211(MGM_W175,d_delay,MGM_W174);
   and MGM_G212(MGM_W176,den_delay,MGM_W175);
   not MGM_G213(MGM_W177,si_delay);
   and MGM_G214(MGM_W178,MGM_W177,MGM_W176);
   not MGM_G215(MGM_W179,ssb_delay);
   and MGM_G216(ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W179,MGM_W178);
   not MGM_G217(MGM_W180,clk_delay);
   and MGM_G218(MGM_W181,d_delay,MGM_W180);
   and MGM_G219(MGM_W182,den_delay,MGM_W181);
   not MGM_G220(MGM_W183,si_delay);
   and MGM_G221(MGM_W184,MGM_W183,MGM_W182);
   and MGM_G222(ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W184);
   not MGM_G223(MGM_W185,clk_delay);
   and MGM_G224(MGM_W186,d_delay,MGM_W185);
   and MGM_G225(MGM_W187,den_delay,MGM_W186);
   and MGM_G226(MGM_W188,si_delay,MGM_W187);
   not MGM_G227(MGM_W189,ssb_delay);
   and MGM_G228(ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_NOT_ssb,MGM_W189,MGM_W188);
   not MGM_G229(MGM_W190,clk_delay);
   and MGM_G230(MGM_W191,d_delay,MGM_W190);
   and MGM_G231(MGM_W192,den_delay,MGM_W191);
   and MGM_G232(MGM_W193,si_delay,MGM_W192);
   and MGM_G233(ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W193);
   not MGM_G234(MGM_W194,d_delay);
   and MGM_G235(MGM_W195,MGM_W194,clk_delay);
   not MGM_G236(MGM_W196,den_delay);
   and MGM_G237(MGM_W197,MGM_W196,MGM_W195);
   not MGM_G238(MGM_W198,si_delay);
   and MGM_G239(MGM_W199,MGM_W198,MGM_W197);
   not MGM_G240(MGM_W200,ssb_delay);
   and MGM_G241(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W200,MGM_W199);
   not MGM_G242(MGM_W201,d_delay);
   and MGM_G243(MGM_W202,MGM_W201,clk_delay);
   not MGM_G244(MGM_W203,den_delay);
   and MGM_G245(MGM_W204,MGM_W203,MGM_W202);
   not MGM_G246(MGM_W205,si_delay);
   and MGM_G247(MGM_W206,MGM_W205,MGM_W204);
   and MGM_G248(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W206);
   not MGM_G249(MGM_W207,d_delay);
   and MGM_G250(MGM_W208,MGM_W207,clk_delay);
   not MGM_G251(MGM_W209,den_delay);
   and MGM_G252(MGM_W210,MGM_W209,MGM_W208);
   and MGM_G253(MGM_W211,si_delay,MGM_W210);
   not MGM_G254(MGM_W212,ssb_delay);
   and MGM_G255(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W212,MGM_W211);
   not MGM_G256(MGM_W213,d_delay);
   and MGM_G257(MGM_W214,MGM_W213,clk_delay);
   not MGM_G258(MGM_W215,den_delay);
   and MGM_G259(MGM_W216,MGM_W215,MGM_W214);
   and MGM_G260(MGM_W217,si_delay,MGM_W216);
   and MGM_G261(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W217);
   not MGM_G262(MGM_W218,d_delay);
   and MGM_G263(MGM_W219,MGM_W218,clk_delay);
   and MGM_G264(MGM_W220,den_delay,MGM_W219);
   not MGM_G265(MGM_W221,si_delay);
   and MGM_G266(MGM_W222,MGM_W221,MGM_W220);
   not MGM_G267(MGM_W223,ssb_delay);
   and MGM_G268(ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W223,MGM_W222);
   not MGM_G269(MGM_W224,d_delay);
   and MGM_G270(MGM_W225,MGM_W224,clk_delay);
   and MGM_G271(MGM_W226,den_delay,MGM_W225);
   not MGM_G272(MGM_W227,si_delay);
   and MGM_G273(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G274(ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W228);
   not MGM_G275(MGM_W229,d_delay);
   and MGM_G276(MGM_W230,MGM_W229,clk_delay);
   and MGM_G277(MGM_W231,den_delay,MGM_W230);
   and MGM_G278(MGM_W232,si_delay,MGM_W231);
   not MGM_G279(MGM_W233,ssb_delay);
   and MGM_G280(ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W233,MGM_W232);
   not MGM_G281(MGM_W234,d_delay);
   and MGM_G282(MGM_W235,MGM_W234,clk_delay);
   and MGM_G283(MGM_W236,den_delay,MGM_W235);
   and MGM_G284(MGM_W237,si_delay,MGM_W236);
   and MGM_G285(ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W237);
   and MGM_G286(MGM_W238,d_delay,clk_delay);
   not MGM_G287(MGM_W239,den_delay);
   and MGM_G288(MGM_W240,MGM_W239,MGM_W238);
   not MGM_G289(MGM_W241,si_delay);
   and MGM_G290(MGM_W242,MGM_W241,MGM_W240);
   not MGM_G291(MGM_W243,ssb_delay);
   and MGM_G292(ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W243,MGM_W242);
   and MGM_G293(MGM_W244,d_delay,clk_delay);
   not MGM_G294(MGM_W245,den_delay);
   and MGM_G295(MGM_W246,MGM_W245,MGM_W244);
   not MGM_G296(MGM_W247,si_delay);
   and MGM_G297(MGM_W248,MGM_W247,MGM_W246);
   and MGM_G298(ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W248);
   and MGM_G299(MGM_W249,d_delay,clk_delay);
   not MGM_G300(MGM_W250,den_delay);
   and MGM_G301(MGM_W251,MGM_W250,MGM_W249);
   and MGM_G302(MGM_W252,si_delay,MGM_W251);
   not MGM_G303(MGM_W253,ssb_delay);
   and MGM_G304(ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W253,MGM_W252);
   and MGM_G305(MGM_W254,d_delay,clk_delay);
   not MGM_G306(MGM_W255,den_delay);
   and MGM_G307(MGM_W256,MGM_W255,MGM_W254);
   and MGM_G308(MGM_W257,si_delay,MGM_W256);
   and MGM_G309(ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W257);
   and MGM_G310(MGM_W258,d_delay,clk_delay);
   and MGM_G311(MGM_W259,den_delay,MGM_W258);
   not MGM_G312(MGM_W260,si_delay);
   and MGM_G313(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G314(MGM_W262,ssb_delay);
   and MGM_G315(ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   and MGM_G316(MGM_W263,d_delay,clk_delay);
   and MGM_G317(MGM_W264,den_delay,MGM_W263);
   not MGM_G318(MGM_W265,si_delay);
   and MGM_G319(MGM_W266,MGM_W265,MGM_W264);
   and MGM_G320(ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W266);
   and MGM_G321(MGM_W267,d_delay,clk_delay);
   and MGM_G322(MGM_W268,den_delay,MGM_W267);
   and MGM_G323(MGM_W269,si_delay,MGM_W268);
   not MGM_G324(MGM_W270,ssb_delay);
   and MGM_G325(ENABLE_clk_AND_d_AND_den_AND_si_AND_NOT_ssb,MGM_W270,MGM_W269);
   and MGM_G326(MGM_W271,d_delay,clk_delay);
   and MGM_G327(MGM_W272,den_delay,MGM_W271);
   and MGM_G328(MGM_W273,si_delay,MGM_W272);
   and MGM_G329(ENABLE_clk_AND_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W273);
   not MGM_G330(MGM_W274,d_delay);
   not MGM_G331(MGM_W275,den_delay);
   and MGM_G332(MGM_W276,MGM_W275,MGM_W274);
   and MGM_G333(MGM_W277,rb_delay,MGM_W276);
   not MGM_G334(MGM_W278,ssb_delay);
   and MGM_G335(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb,MGM_W278,MGM_W277);
   not MGM_G336(MGM_W279,d_delay);
   and MGM_G337(MGM_W280,den_delay,MGM_W279);
   and MGM_G338(MGM_W281,rb_delay,MGM_W280);
   not MGM_G339(MGM_W282,ssb_delay);
   and MGM_G340(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb,MGM_W282,MGM_W281);
   not MGM_G341(MGM_W283,den_delay);
   and MGM_G342(MGM_W284,MGM_W283,d_delay);
   and MGM_G343(MGM_W285,rb_delay,MGM_W284);
   not MGM_G344(MGM_W286,ssb_delay);
   and MGM_G345(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb,MGM_W286,MGM_W285);
   and MGM_G346(MGM_W287,den_delay,d_delay);
   and MGM_G347(MGM_W288,rb_delay,MGM_W287);
   not MGM_G348(MGM_W289,ssb_delay);
   and MGM_G349(ENABLE_d_AND_den_AND_rb_AND_NOT_ssb,MGM_W289,MGM_W288);
   not MGM_G350(MGM_W290,d_delay);
   not MGM_G351(MGM_W291,den_delay);
   and MGM_G352(MGM_W292,MGM_W291,MGM_W290);
   and MGM_G353(MGM_W293,rb_delay,MGM_W292);
   not MGM_G354(MGM_W294,si_delay);
   and MGM_G355(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si,MGM_W294,MGM_W293);
   not MGM_G356(MGM_W295,d_delay);
   not MGM_G357(MGM_W296,den_delay);
   and MGM_G358(MGM_W297,MGM_W296,MGM_W295);
   and MGM_G359(MGM_W298,rb_delay,MGM_W297);
   and MGM_G360(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si,si_delay,MGM_W298);
   not MGM_G361(MGM_W299,d_delay);
   and MGM_G362(MGM_W300,den_delay,MGM_W299);
   and MGM_G363(MGM_W301,rb_delay,MGM_W300);
   and MGM_G364(ENABLE_NOT_d_AND_den_AND_rb_AND_si,si_delay,MGM_W301);
   not MGM_G365(MGM_W302,den_delay);
   and MGM_G366(MGM_W303,MGM_W302,d_delay);
   and MGM_G367(MGM_W304,rb_delay,MGM_W303);
   not MGM_G368(MGM_W305,si_delay);
   and MGM_G369(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   not MGM_G370(MGM_W306,den_delay);
   and MGM_G371(MGM_W307,MGM_W306,d_delay);
   and MGM_G372(MGM_W308,rb_delay,MGM_W307);
   and MGM_G373(ENABLE_d_AND_NOT_den_AND_rb_AND_si,si_delay,MGM_W308);
   and MGM_G374(MGM_W309,den_delay,d_delay);
   and MGM_G375(MGM_W310,rb_delay,MGM_W309);
   not MGM_G376(MGM_W311,si_delay);
   and MGM_G377(ENABLE_d_AND_den_AND_rb_AND_NOT_si,MGM_W311,MGM_W310);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy043ah1n12x5( clk, d, den, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy043ah_func b15fqy043ah1n12x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy043ah_func b15fqy043ah1n12x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy043ah_func b15fqy043ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy043ah_func b15fqy043ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,den_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   and MGM_G3(MGM_W3,rb_delay,MGM_W2);
   not MGM_G4(MGM_W4,si_delay);
   and MGM_G5(MGM_W5,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W6,ssb_delay);
   and MGM_G7(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W6,MGM_W5);
   not MGM_G8(MGM_W7,d_delay);
   not MGM_G9(MGM_W8,den_delay);
   and MGM_G10(MGM_W9,MGM_W8,MGM_W7);
   and MGM_G11(MGM_W10,rb_delay,MGM_W9);
   and MGM_G12(MGM_W11,si_delay,MGM_W10);
   not MGM_G13(MGM_W12,ssb_delay);
   and MGM_G14(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G15(MGM_W13,d_delay);
   and MGM_G16(MGM_W14,den_delay,MGM_W13);
   and MGM_G17(MGM_W15,rb_delay,MGM_W14);
   not MGM_G18(MGM_W16,si_delay);
   and MGM_G19(MGM_W17,MGM_W16,MGM_W15);
   not MGM_G20(MGM_W18,ssb_delay);
   and MGM_G21(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   not MGM_G22(MGM_W19,d_delay);
   and MGM_G23(MGM_W20,den_delay,MGM_W19);
   and MGM_G24(MGM_W21,rb_delay,MGM_W20);
   not MGM_G25(MGM_W22,si_delay);
   and MGM_G26(MGM_W23,MGM_W22,MGM_W21);
   and MGM_G27(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W23);
   not MGM_G28(MGM_W24,d_delay);
   and MGM_G29(MGM_W25,den_delay,MGM_W24);
   and MGM_G30(MGM_W26,rb_delay,MGM_W25);
   and MGM_G31(MGM_W27,si_delay,MGM_W26);
   not MGM_G32(MGM_W28,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W28,MGM_W27);
   not MGM_G34(MGM_W29,d_delay);
   and MGM_G35(MGM_W30,den_delay,MGM_W29);
   and MGM_G36(MGM_W31,rb_delay,MGM_W30);
   and MGM_G37(MGM_W32,si_delay,MGM_W31);
   and MGM_G38(ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W32);
   not MGM_G39(MGM_W33,den_delay);
   and MGM_G40(MGM_W34,MGM_W33,d_delay);
   and MGM_G41(MGM_W35,rb_delay,MGM_W34);
   not MGM_G42(MGM_W36,si_delay);
   and MGM_G43(MGM_W37,MGM_W36,MGM_W35);
   not MGM_G44(MGM_W38,ssb_delay);
   and MGM_G45(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W38,MGM_W37);
   not MGM_G46(MGM_W39,den_delay);
   and MGM_G47(MGM_W40,MGM_W39,d_delay);
   and MGM_G48(MGM_W41,rb_delay,MGM_W40);
   and MGM_G49(MGM_W42,si_delay,MGM_W41);
   not MGM_G50(MGM_W43,ssb_delay);
   and MGM_G51(ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W43,MGM_W42);
   and MGM_G52(MGM_W44,den_delay,d_delay);
   and MGM_G53(MGM_W45,rb_delay,MGM_W44);
   not MGM_G54(MGM_W46,si_delay);
   and MGM_G55(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G56(MGM_W48,ssb_delay);
   and MGM_G57(ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   and MGM_G58(MGM_W49,den_delay,d_delay);
   and MGM_G59(MGM_W50,rb_delay,MGM_W49);
   not MGM_G60(MGM_W51,si_delay);
   and MGM_G61(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G62(ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G63(MGM_W53,den_delay,d_delay);
   and MGM_G64(MGM_W54,rb_delay,MGM_W53);
   and MGM_G65(MGM_W55,si_delay,MGM_W54);
   not MGM_G66(MGM_W56,ssb_delay);
   and MGM_G67(ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   and MGM_G68(MGM_W57,den_delay,d_delay);
   and MGM_G69(MGM_W58,rb_delay,MGM_W57);
   and MGM_G70(MGM_W59,si_delay,MGM_W58);
   and MGM_G71(ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W59);
   and MGM_G72(MGM_W60,rb_delay,den_delay);
   not MGM_G73(MGM_W61,si_delay);
   and MGM_G74(MGM_W62,MGM_W61,MGM_W60);
   and MGM_G75(ENABLE_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W62);
   and MGM_G76(MGM_W63,rb_delay,den_delay);
   and MGM_G77(MGM_W64,si_delay,MGM_W63);
   and MGM_G78(ENABLE_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W64);
   not MGM_G79(MGM_W65,d_delay);
   and MGM_G80(MGM_W66,rb_delay,MGM_W65);
   not MGM_G81(MGM_W67,si_delay);
   and MGM_G82(MGM_W68,MGM_W67,MGM_W66);
   and MGM_G83(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W68);
   not MGM_G84(MGM_W69,d_delay);
   and MGM_G85(MGM_W70,rb_delay,MGM_W69);
   and MGM_G86(MGM_W71,si_delay,MGM_W70);
   and MGM_G87(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W71);
   and MGM_G88(MGM_W72,rb_delay,d_delay);
   not MGM_G89(MGM_W73,si_delay);
   and MGM_G90(MGM_W74,MGM_W73,MGM_W72);
   and MGM_G91(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W74);
   and MGM_G92(MGM_W75,rb_delay,d_delay);
   and MGM_G93(MGM_W76,si_delay,MGM_W75);
   and MGM_G94(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W76);
   not MGM_G95(MGM_W77,d_delay);
   not MGM_G96(MGM_W78,den_delay);
   and MGM_G97(MGM_W79,MGM_W78,MGM_W77);
   and MGM_G98(MGM_W80,si_delay,MGM_W79);
   not MGM_G99(MGM_W81,ssb_delay);
   and MGM_G100(ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W81,MGM_W80);
   not MGM_G101(MGM_W82,d_delay);
   and MGM_G102(MGM_W83,den_delay,MGM_W82);
   and MGM_G103(MGM_W84,si_delay,MGM_W83);
   not MGM_G104(MGM_W85,ssb_delay);
   and MGM_G105(ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W85,MGM_W84);
   not MGM_G106(MGM_W86,den_delay);
   and MGM_G107(MGM_W87,MGM_W86,d_delay);
   and MGM_G108(MGM_W88,si_delay,MGM_W87);
   not MGM_G109(MGM_W89,ssb_delay);
   and MGM_G110(ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W89,MGM_W88);
   and MGM_G111(MGM_W90,den_delay,d_delay);
   not MGM_G112(MGM_W91,si_delay);
   and MGM_G113(MGM_W92,MGM_W91,MGM_W90);
   and MGM_G114(ENABLE_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W92);
   and MGM_G115(MGM_W93,den_delay,d_delay);
   and MGM_G116(MGM_W94,si_delay,MGM_W93);
   not MGM_G117(MGM_W95,ssb_delay);
   and MGM_G118(ENABLE_d_AND_den_AND_si_AND_NOT_ssb,MGM_W95,MGM_W94);
   and MGM_G119(MGM_W96,den_delay,d_delay);
   and MGM_G120(MGM_W97,si_delay,MGM_W96);
   and MGM_G121(ENABLE_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W97);
   not MGM_G122(MGM_W98,clk_delay);
   not MGM_G123(MGM_W99,d_delay);
   and MGM_G124(MGM_W100,MGM_W99,MGM_W98);
   not MGM_G125(MGM_W101,den_delay);
   and MGM_G126(MGM_W102,MGM_W101,MGM_W100);
   not MGM_G127(MGM_W103,si_delay);
   and MGM_G128(MGM_W104,MGM_W103,MGM_W102);
   not MGM_G129(MGM_W105,ssb_delay);
   and MGM_G130(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W105,MGM_W104);
   not MGM_G131(MGM_W106,clk_delay);
   not MGM_G132(MGM_W107,d_delay);
   and MGM_G133(MGM_W108,MGM_W107,MGM_W106);
   not MGM_G134(MGM_W109,den_delay);
   and MGM_G135(MGM_W110,MGM_W109,MGM_W108);
   not MGM_G136(MGM_W111,si_delay);
   and MGM_G137(MGM_W112,MGM_W111,MGM_W110);
   and MGM_G138(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W112);
   not MGM_G139(MGM_W113,clk_delay);
   not MGM_G140(MGM_W114,d_delay);
   and MGM_G141(MGM_W115,MGM_W114,MGM_W113);
   not MGM_G142(MGM_W116,den_delay);
   and MGM_G143(MGM_W117,MGM_W116,MGM_W115);
   and MGM_G144(MGM_W118,si_delay,MGM_W117);
   not MGM_G145(MGM_W119,ssb_delay);
   and MGM_G146(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W119,MGM_W118);
   not MGM_G147(MGM_W120,clk_delay);
   not MGM_G148(MGM_W121,d_delay);
   and MGM_G149(MGM_W122,MGM_W121,MGM_W120);
   not MGM_G150(MGM_W123,den_delay);
   and MGM_G151(MGM_W124,MGM_W123,MGM_W122);
   and MGM_G152(MGM_W125,si_delay,MGM_W124);
   and MGM_G153(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W125);
   not MGM_G154(MGM_W126,clk_delay);
   not MGM_G155(MGM_W127,d_delay);
   and MGM_G156(MGM_W128,MGM_W127,MGM_W126);
   and MGM_G157(MGM_W129,den_delay,MGM_W128);
   not MGM_G158(MGM_W130,si_delay);
   and MGM_G159(MGM_W131,MGM_W130,MGM_W129);
   not MGM_G160(MGM_W132,ssb_delay);
   and MGM_G161(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W132,MGM_W131);
   not MGM_G162(MGM_W133,clk_delay);
   not MGM_G163(MGM_W134,d_delay);
   and MGM_G164(MGM_W135,MGM_W134,MGM_W133);
   and MGM_G165(MGM_W136,den_delay,MGM_W135);
   not MGM_G166(MGM_W137,si_delay);
   and MGM_G167(MGM_W138,MGM_W137,MGM_W136);
   and MGM_G168(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W138);
   not MGM_G169(MGM_W139,clk_delay);
   not MGM_G170(MGM_W140,d_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   and MGM_G172(MGM_W142,den_delay,MGM_W141);
   and MGM_G173(MGM_W143,si_delay,MGM_W142);
   not MGM_G174(MGM_W144,ssb_delay);
   and MGM_G175(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W144,MGM_W143);
   not MGM_G176(MGM_W145,clk_delay);
   not MGM_G177(MGM_W146,d_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(MGM_W148,den_delay,MGM_W147);
   and MGM_G180(MGM_W149,si_delay,MGM_W148);
   and MGM_G181(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W149);
   not MGM_G182(MGM_W150,clk_delay);
   and MGM_G183(MGM_W151,d_delay,MGM_W150);
   not MGM_G184(MGM_W152,den_delay);
   and MGM_G185(MGM_W153,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W154,si_delay);
   and MGM_G187(MGM_W155,MGM_W154,MGM_W153);
   not MGM_G188(MGM_W156,ssb_delay);
   and MGM_G189(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W156,MGM_W155);
   not MGM_G190(MGM_W157,clk_delay);
   and MGM_G191(MGM_W158,d_delay,MGM_W157);
   not MGM_G192(MGM_W159,den_delay);
   and MGM_G193(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G194(MGM_W161,si_delay);
   and MGM_G195(MGM_W162,MGM_W161,MGM_W160);
   and MGM_G196(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W162);
   not MGM_G197(MGM_W163,clk_delay);
   and MGM_G198(MGM_W164,d_delay,MGM_W163);
   not MGM_G199(MGM_W165,den_delay);
   and MGM_G200(MGM_W166,MGM_W165,MGM_W164);
   and MGM_G201(MGM_W167,si_delay,MGM_W166);
   not MGM_G202(MGM_W168,ssb_delay);
   and MGM_G203(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W168,MGM_W167);
   not MGM_G204(MGM_W169,clk_delay);
   and MGM_G205(MGM_W170,d_delay,MGM_W169);
   not MGM_G206(MGM_W171,den_delay);
   and MGM_G207(MGM_W172,MGM_W171,MGM_W170);
   and MGM_G208(MGM_W173,si_delay,MGM_W172);
   and MGM_G209(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W173);
   not MGM_G210(MGM_W174,clk_delay);
   and MGM_G211(MGM_W175,d_delay,MGM_W174);
   and MGM_G212(MGM_W176,den_delay,MGM_W175);
   not MGM_G213(MGM_W177,si_delay);
   and MGM_G214(MGM_W178,MGM_W177,MGM_W176);
   not MGM_G215(MGM_W179,ssb_delay);
   and MGM_G216(ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W179,MGM_W178);
   not MGM_G217(MGM_W180,clk_delay);
   and MGM_G218(MGM_W181,d_delay,MGM_W180);
   and MGM_G219(MGM_W182,den_delay,MGM_W181);
   not MGM_G220(MGM_W183,si_delay);
   and MGM_G221(MGM_W184,MGM_W183,MGM_W182);
   and MGM_G222(ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W184);
   not MGM_G223(MGM_W185,clk_delay);
   and MGM_G224(MGM_W186,d_delay,MGM_W185);
   and MGM_G225(MGM_W187,den_delay,MGM_W186);
   and MGM_G226(MGM_W188,si_delay,MGM_W187);
   not MGM_G227(MGM_W189,ssb_delay);
   and MGM_G228(ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_NOT_ssb,MGM_W189,MGM_W188);
   not MGM_G229(MGM_W190,clk_delay);
   and MGM_G230(MGM_W191,d_delay,MGM_W190);
   and MGM_G231(MGM_W192,den_delay,MGM_W191);
   and MGM_G232(MGM_W193,si_delay,MGM_W192);
   and MGM_G233(ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W193);
   not MGM_G234(MGM_W194,d_delay);
   and MGM_G235(MGM_W195,MGM_W194,clk_delay);
   not MGM_G236(MGM_W196,den_delay);
   and MGM_G237(MGM_W197,MGM_W196,MGM_W195);
   not MGM_G238(MGM_W198,si_delay);
   and MGM_G239(MGM_W199,MGM_W198,MGM_W197);
   not MGM_G240(MGM_W200,ssb_delay);
   and MGM_G241(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W200,MGM_W199);
   not MGM_G242(MGM_W201,d_delay);
   and MGM_G243(MGM_W202,MGM_W201,clk_delay);
   not MGM_G244(MGM_W203,den_delay);
   and MGM_G245(MGM_W204,MGM_W203,MGM_W202);
   not MGM_G246(MGM_W205,si_delay);
   and MGM_G247(MGM_W206,MGM_W205,MGM_W204);
   and MGM_G248(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W206);
   not MGM_G249(MGM_W207,d_delay);
   and MGM_G250(MGM_W208,MGM_W207,clk_delay);
   not MGM_G251(MGM_W209,den_delay);
   and MGM_G252(MGM_W210,MGM_W209,MGM_W208);
   and MGM_G253(MGM_W211,si_delay,MGM_W210);
   not MGM_G254(MGM_W212,ssb_delay);
   and MGM_G255(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W212,MGM_W211);
   not MGM_G256(MGM_W213,d_delay);
   and MGM_G257(MGM_W214,MGM_W213,clk_delay);
   not MGM_G258(MGM_W215,den_delay);
   and MGM_G259(MGM_W216,MGM_W215,MGM_W214);
   and MGM_G260(MGM_W217,si_delay,MGM_W216);
   and MGM_G261(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W217);
   not MGM_G262(MGM_W218,d_delay);
   and MGM_G263(MGM_W219,MGM_W218,clk_delay);
   and MGM_G264(MGM_W220,den_delay,MGM_W219);
   not MGM_G265(MGM_W221,si_delay);
   and MGM_G266(MGM_W222,MGM_W221,MGM_W220);
   not MGM_G267(MGM_W223,ssb_delay);
   and MGM_G268(ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W223,MGM_W222);
   not MGM_G269(MGM_W224,d_delay);
   and MGM_G270(MGM_W225,MGM_W224,clk_delay);
   and MGM_G271(MGM_W226,den_delay,MGM_W225);
   not MGM_G272(MGM_W227,si_delay);
   and MGM_G273(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G274(ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W228);
   not MGM_G275(MGM_W229,d_delay);
   and MGM_G276(MGM_W230,MGM_W229,clk_delay);
   and MGM_G277(MGM_W231,den_delay,MGM_W230);
   and MGM_G278(MGM_W232,si_delay,MGM_W231);
   not MGM_G279(MGM_W233,ssb_delay);
   and MGM_G280(ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W233,MGM_W232);
   not MGM_G281(MGM_W234,d_delay);
   and MGM_G282(MGM_W235,MGM_W234,clk_delay);
   and MGM_G283(MGM_W236,den_delay,MGM_W235);
   and MGM_G284(MGM_W237,si_delay,MGM_W236);
   and MGM_G285(ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W237);
   and MGM_G286(MGM_W238,d_delay,clk_delay);
   not MGM_G287(MGM_W239,den_delay);
   and MGM_G288(MGM_W240,MGM_W239,MGM_W238);
   not MGM_G289(MGM_W241,si_delay);
   and MGM_G290(MGM_W242,MGM_W241,MGM_W240);
   not MGM_G291(MGM_W243,ssb_delay);
   and MGM_G292(ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W243,MGM_W242);
   and MGM_G293(MGM_W244,d_delay,clk_delay);
   not MGM_G294(MGM_W245,den_delay);
   and MGM_G295(MGM_W246,MGM_W245,MGM_W244);
   not MGM_G296(MGM_W247,si_delay);
   and MGM_G297(MGM_W248,MGM_W247,MGM_W246);
   and MGM_G298(ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W248);
   and MGM_G299(MGM_W249,d_delay,clk_delay);
   not MGM_G300(MGM_W250,den_delay);
   and MGM_G301(MGM_W251,MGM_W250,MGM_W249);
   and MGM_G302(MGM_W252,si_delay,MGM_W251);
   not MGM_G303(MGM_W253,ssb_delay);
   and MGM_G304(ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W253,MGM_W252);
   and MGM_G305(MGM_W254,d_delay,clk_delay);
   not MGM_G306(MGM_W255,den_delay);
   and MGM_G307(MGM_W256,MGM_W255,MGM_W254);
   and MGM_G308(MGM_W257,si_delay,MGM_W256);
   and MGM_G309(ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W257);
   and MGM_G310(MGM_W258,d_delay,clk_delay);
   and MGM_G311(MGM_W259,den_delay,MGM_W258);
   not MGM_G312(MGM_W260,si_delay);
   and MGM_G313(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G314(MGM_W262,ssb_delay);
   and MGM_G315(ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   and MGM_G316(MGM_W263,d_delay,clk_delay);
   and MGM_G317(MGM_W264,den_delay,MGM_W263);
   not MGM_G318(MGM_W265,si_delay);
   and MGM_G319(MGM_W266,MGM_W265,MGM_W264);
   and MGM_G320(ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W266);
   and MGM_G321(MGM_W267,d_delay,clk_delay);
   and MGM_G322(MGM_W268,den_delay,MGM_W267);
   and MGM_G323(MGM_W269,si_delay,MGM_W268);
   not MGM_G324(MGM_W270,ssb_delay);
   and MGM_G325(ENABLE_clk_AND_d_AND_den_AND_si_AND_NOT_ssb,MGM_W270,MGM_W269);
   and MGM_G326(MGM_W271,d_delay,clk_delay);
   and MGM_G327(MGM_W272,den_delay,MGM_W271);
   and MGM_G328(MGM_W273,si_delay,MGM_W272);
   and MGM_G329(ENABLE_clk_AND_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W273);
   not MGM_G330(MGM_W274,d_delay);
   not MGM_G331(MGM_W275,den_delay);
   and MGM_G332(MGM_W276,MGM_W275,MGM_W274);
   and MGM_G333(MGM_W277,rb_delay,MGM_W276);
   not MGM_G334(MGM_W278,ssb_delay);
   and MGM_G335(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb,MGM_W278,MGM_W277);
   not MGM_G336(MGM_W279,d_delay);
   and MGM_G337(MGM_W280,den_delay,MGM_W279);
   and MGM_G338(MGM_W281,rb_delay,MGM_W280);
   not MGM_G339(MGM_W282,ssb_delay);
   and MGM_G340(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb,MGM_W282,MGM_W281);
   not MGM_G341(MGM_W283,den_delay);
   and MGM_G342(MGM_W284,MGM_W283,d_delay);
   and MGM_G343(MGM_W285,rb_delay,MGM_W284);
   not MGM_G344(MGM_W286,ssb_delay);
   and MGM_G345(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb,MGM_W286,MGM_W285);
   and MGM_G346(MGM_W287,den_delay,d_delay);
   and MGM_G347(MGM_W288,rb_delay,MGM_W287);
   not MGM_G348(MGM_W289,ssb_delay);
   and MGM_G349(ENABLE_d_AND_den_AND_rb_AND_NOT_ssb,MGM_W289,MGM_W288);
   not MGM_G350(MGM_W290,d_delay);
   not MGM_G351(MGM_W291,den_delay);
   and MGM_G352(MGM_W292,MGM_W291,MGM_W290);
   and MGM_G353(MGM_W293,rb_delay,MGM_W292);
   not MGM_G354(MGM_W294,si_delay);
   and MGM_G355(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si,MGM_W294,MGM_W293);
   not MGM_G356(MGM_W295,d_delay);
   not MGM_G357(MGM_W296,den_delay);
   and MGM_G358(MGM_W297,MGM_W296,MGM_W295);
   and MGM_G359(MGM_W298,rb_delay,MGM_W297);
   and MGM_G360(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si,si_delay,MGM_W298);
   not MGM_G361(MGM_W299,d_delay);
   and MGM_G362(MGM_W300,den_delay,MGM_W299);
   and MGM_G363(MGM_W301,rb_delay,MGM_W300);
   and MGM_G364(ENABLE_NOT_d_AND_den_AND_rb_AND_si,si_delay,MGM_W301);
   not MGM_G365(MGM_W302,den_delay);
   and MGM_G366(MGM_W303,MGM_W302,d_delay);
   and MGM_G367(MGM_W304,rb_delay,MGM_W303);
   not MGM_G368(MGM_W305,si_delay);
   and MGM_G369(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   not MGM_G370(MGM_W306,den_delay);
   and MGM_G371(MGM_W307,MGM_W306,d_delay);
   and MGM_G372(MGM_W308,rb_delay,MGM_W307);
   and MGM_G373(ENABLE_d_AND_NOT_den_AND_rb_AND_si,si_delay,MGM_W308);
   and MGM_G374(MGM_W309,den_delay,d_delay);
   and MGM_G375(MGM_W310,rb_delay,MGM_W309);
   not MGM_G376(MGM_W311,si_delay);
   and MGM_G377(ENABLE_d_AND_den_AND_rb_AND_NOT_si,MGM_W311,MGM_W310);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy043ah1n16x5( clk, d, den, o, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, den, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy043ah_func b15fqy043ah1n16x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy043ah_func b15fqy043ah1n16x5_behav_inst(.clk(clk),.d(d),.den(den),.o(o),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire den_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy043ah_func b15fqy043ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy043ah_func b15fqy043ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.den(den_delay),.o(o),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   not MGM_G1(MGM_W1,den_delay);
   and MGM_G2(MGM_W2,MGM_W1,MGM_W0);
   and MGM_G3(MGM_W3,rb_delay,MGM_W2);
   not MGM_G4(MGM_W4,si_delay);
   and MGM_G5(MGM_W5,MGM_W4,MGM_W3);
   not MGM_G6(MGM_W6,ssb_delay);
   and MGM_G7(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W6,MGM_W5);
   not MGM_G8(MGM_W7,d_delay);
   not MGM_G9(MGM_W8,den_delay);
   and MGM_G10(MGM_W9,MGM_W8,MGM_W7);
   and MGM_G11(MGM_W10,rb_delay,MGM_W9);
   and MGM_G12(MGM_W11,si_delay,MGM_W10);
   not MGM_G13(MGM_W12,ssb_delay);
   and MGM_G14(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W12,MGM_W11);
   not MGM_G15(MGM_W13,d_delay);
   and MGM_G16(MGM_W14,den_delay,MGM_W13);
   and MGM_G17(MGM_W15,rb_delay,MGM_W14);
   not MGM_G18(MGM_W16,si_delay);
   and MGM_G19(MGM_W17,MGM_W16,MGM_W15);
   not MGM_G20(MGM_W18,ssb_delay);
   and MGM_G21(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W18,MGM_W17);
   not MGM_G22(MGM_W19,d_delay);
   and MGM_G23(MGM_W20,den_delay,MGM_W19);
   and MGM_G24(MGM_W21,rb_delay,MGM_W20);
   not MGM_G25(MGM_W22,si_delay);
   and MGM_G26(MGM_W23,MGM_W22,MGM_W21);
   and MGM_G27(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W23);
   not MGM_G28(MGM_W24,d_delay);
   and MGM_G29(MGM_W25,den_delay,MGM_W24);
   and MGM_G30(MGM_W26,rb_delay,MGM_W25);
   and MGM_G31(MGM_W27,si_delay,MGM_W26);
   not MGM_G32(MGM_W28,ssb_delay);
   and MGM_G33(ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W28,MGM_W27);
   not MGM_G34(MGM_W29,d_delay);
   and MGM_G35(MGM_W30,den_delay,MGM_W29);
   and MGM_G36(MGM_W31,rb_delay,MGM_W30);
   and MGM_G37(MGM_W32,si_delay,MGM_W31);
   and MGM_G38(ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W32);
   not MGM_G39(MGM_W33,den_delay);
   and MGM_G40(MGM_W34,MGM_W33,d_delay);
   and MGM_G41(MGM_W35,rb_delay,MGM_W34);
   not MGM_G42(MGM_W36,si_delay);
   and MGM_G43(MGM_W37,MGM_W36,MGM_W35);
   not MGM_G44(MGM_W38,ssb_delay);
   and MGM_G45(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W38,MGM_W37);
   not MGM_G46(MGM_W39,den_delay);
   and MGM_G47(MGM_W40,MGM_W39,d_delay);
   and MGM_G48(MGM_W41,rb_delay,MGM_W40);
   and MGM_G49(MGM_W42,si_delay,MGM_W41);
   not MGM_G50(MGM_W43,ssb_delay);
   and MGM_G51(ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W43,MGM_W42);
   and MGM_G52(MGM_W44,den_delay,d_delay);
   and MGM_G53(MGM_W45,rb_delay,MGM_W44);
   not MGM_G54(MGM_W46,si_delay);
   and MGM_G55(MGM_W47,MGM_W46,MGM_W45);
   not MGM_G56(MGM_W48,ssb_delay);
   and MGM_G57(ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W48,MGM_W47);
   and MGM_G58(MGM_W49,den_delay,d_delay);
   and MGM_G59(MGM_W50,rb_delay,MGM_W49);
   not MGM_G60(MGM_W51,si_delay);
   and MGM_G61(MGM_W52,MGM_W51,MGM_W50);
   and MGM_G62(ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G63(MGM_W53,den_delay,d_delay);
   and MGM_G64(MGM_W54,rb_delay,MGM_W53);
   and MGM_G65(MGM_W55,si_delay,MGM_W54);
   not MGM_G66(MGM_W56,ssb_delay);
   and MGM_G67(ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   and MGM_G68(MGM_W57,den_delay,d_delay);
   and MGM_G69(MGM_W58,rb_delay,MGM_W57);
   and MGM_G70(MGM_W59,si_delay,MGM_W58);
   and MGM_G71(ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W59);
   and MGM_G72(MGM_W60,rb_delay,den_delay);
   not MGM_G73(MGM_W61,si_delay);
   and MGM_G74(MGM_W62,MGM_W61,MGM_W60);
   and MGM_G75(ENABLE_den_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W62);
   and MGM_G76(MGM_W63,rb_delay,den_delay);
   and MGM_G77(MGM_W64,si_delay,MGM_W63);
   and MGM_G78(ENABLE_den_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W64);
   not MGM_G79(MGM_W65,d_delay);
   and MGM_G80(MGM_W66,rb_delay,MGM_W65);
   not MGM_G81(MGM_W67,si_delay);
   and MGM_G82(MGM_W68,MGM_W67,MGM_W66);
   and MGM_G83(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W68);
   not MGM_G84(MGM_W69,d_delay);
   and MGM_G85(MGM_W70,rb_delay,MGM_W69);
   and MGM_G86(MGM_W71,si_delay,MGM_W70);
   and MGM_G87(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W71);
   and MGM_G88(MGM_W72,rb_delay,d_delay);
   not MGM_G89(MGM_W73,si_delay);
   and MGM_G90(MGM_W74,MGM_W73,MGM_W72);
   and MGM_G91(ENABLE_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W74);
   and MGM_G92(MGM_W75,rb_delay,d_delay);
   and MGM_G93(MGM_W76,si_delay,MGM_W75);
   and MGM_G94(ENABLE_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W76);
   not MGM_G95(MGM_W77,d_delay);
   not MGM_G96(MGM_W78,den_delay);
   and MGM_G97(MGM_W79,MGM_W78,MGM_W77);
   and MGM_G98(MGM_W80,si_delay,MGM_W79);
   not MGM_G99(MGM_W81,ssb_delay);
   and MGM_G100(ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W81,MGM_W80);
   not MGM_G101(MGM_W82,d_delay);
   and MGM_G102(MGM_W83,den_delay,MGM_W82);
   and MGM_G103(MGM_W84,si_delay,MGM_W83);
   not MGM_G104(MGM_W85,ssb_delay);
   and MGM_G105(ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W85,MGM_W84);
   not MGM_G106(MGM_W86,den_delay);
   and MGM_G107(MGM_W87,MGM_W86,d_delay);
   and MGM_G108(MGM_W88,si_delay,MGM_W87);
   not MGM_G109(MGM_W89,ssb_delay);
   and MGM_G110(ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W89,MGM_W88);
   and MGM_G111(MGM_W90,den_delay,d_delay);
   not MGM_G112(MGM_W91,si_delay);
   and MGM_G113(MGM_W92,MGM_W91,MGM_W90);
   and MGM_G114(ENABLE_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W92);
   and MGM_G115(MGM_W93,den_delay,d_delay);
   and MGM_G116(MGM_W94,si_delay,MGM_W93);
   not MGM_G117(MGM_W95,ssb_delay);
   and MGM_G118(ENABLE_d_AND_den_AND_si_AND_NOT_ssb,MGM_W95,MGM_W94);
   and MGM_G119(MGM_W96,den_delay,d_delay);
   and MGM_G120(MGM_W97,si_delay,MGM_W96);
   and MGM_G121(ENABLE_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W97);
   not MGM_G122(MGM_W98,clk_delay);
   not MGM_G123(MGM_W99,d_delay);
   and MGM_G124(MGM_W100,MGM_W99,MGM_W98);
   not MGM_G125(MGM_W101,den_delay);
   and MGM_G126(MGM_W102,MGM_W101,MGM_W100);
   not MGM_G127(MGM_W103,si_delay);
   and MGM_G128(MGM_W104,MGM_W103,MGM_W102);
   not MGM_G129(MGM_W105,ssb_delay);
   and MGM_G130(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W105,MGM_W104);
   not MGM_G131(MGM_W106,clk_delay);
   not MGM_G132(MGM_W107,d_delay);
   and MGM_G133(MGM_W108,MGM_W107,MGM_W106);
   not MGM_G134(MGM_W109,den_delay);
   and MGM_G135(MGM_W110,MGM_W109,MGM_W108);
   not MGM_G136(MGM_W111,si_delay);
   and MGM_G137(MGM_W112,MGM_W111,MGM_W110);
   and MGM_G138(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W112);
   not MGM_G139(MGM_W113,clk_delay);
   not MGM_G140(MGM_W114,d_delay);
   and MGM_G141(MGM_W115,MGM_W114,MGM_W113);
   not MGM_G142(MGM_W116,den_delay);
   and MGM_G143(MGM_W117,MGM_W116,MGM_W115);
   and MGM_G144(MGM_W118,si_delay,MGM_W117);
   not MGM_G145(MGM_W119,ssb_delay);
   and MGM_G146(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W119,MGM_W118);
   not MGM_G147(MGM_W120,clk_delay);
   not MGM_G148(MGM_W121,d_delay);
   and MGM_G149(MGM_W122,MGM_W121,MGM_W120);
   not MGM_G150(MGM_W123,den_delay);
   and MGM_G151(MGM_W124,MGM_W123,MGM_W122);
   and MGM_G152(MGM_W125,si_delay,MGM_W124);
   and MGM_G153(ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W125);
   not MGM_G154(MGM_W126,clk_delay);
   not MGM_G155(MGM_W127,d_delay);
   and MGM_G156(MGM_W128,MGM_W127,MGM_W126);
   and MGM_G157(MGM_W129,den_delay,MGM_W128);
   not MGM_G158(MGM_W130,si_delay);
   and MGM_G159(MGM_W131,MGM_W130,MGM_W129);
   not MGM_G160(MGM_W132,ssb_delay);
   and MGM_G161(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W132,MGM_W131);
   not MGM_G162(MGM_W133,clk_delay);
   not MGM_G163(MGM_W134,d_delay);
   and MGM_G164(MGM_W135,MGM_W134,MGM_W133);
   and MGM_G165(MGM_W136,den_delay,MGM_W135);
   not MGM_G166(MGM_W137,si_delay);
   and MGM_G167(MGM_W138,MGM_W137,MGM_W136);
   and MGM_G168(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W138);
   not MGM_G169(MGM_W139,clk_delay);
   not MGM_G170(MGM_W140,d_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   and MGM_G172(MGM_W142,den_delay,MGM_W141);
   and MGM_G173(MGM_W143,si_delay,MGM_W142);
   not MGM_G174(MGM_W144,ssb_delay);
   and MGM_G175(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W144,MGM_W143);
   not MGM_G176(MGM_W145,clk_delay);
   not MGM_G177(MGM_W146,d_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(MGM_W148,den_delay,MGM_W147);
   and MGM_G180(MGM_W149,si_delay,MGM_W148);
   and MGM_G181(ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W149);
   not MGM_G182(MGM_W150,clk_delay);
   and MGM_G183(MGM_W151,d_delay,MGM_W150);
   not MGM_G184(MGM_W152,den_delay);
   and MGM_G185(MGM_W153,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W154,si_delay);
   and MGM_G187(MGM_W155,MGM_W154,MGM_W153);
   not MGM_G188(MGM_W156,ssb_delay);
   and MGM_G189(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W156,MGM_W155);
   not MGM_G190(MGM_W157,clk_delay);
   and MGM_G191(MGM_W158,d_delay,MGM_W157);
   not MGM_G192(MGM_W159,den_delay);
   and MGM_G193(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G194(MGM_W161,si_delay);
   and MGM_G195(MGM_W162,MGM_W161,MGM_W160);
   and MGM_G196(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W162);
   not MGM_G197(MGM_W163,clk_delay);
   and MGM_G198(MGM_W164,d_delay,MGM_W163);
   not MGM_G199(MGM_W165,den_delay);
   and MGM_G200(MGM_W166,MGM_W165,MGM_W164);
   and MGM_G201(MGM_W167,si_delay,MGM_W166);
   not MGM_G202(MGM_W168,ssb_delay);
   and MGM_G203(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W168,MGM_W167);
   not MGM_G204(MGM_W169,clk_delay);
   and MGM_G205(MGM_W170,d_delay,MGM_W169);
   not MGM_G206(MGM_W171,den_delay);
   and MGM_G207(MGM_W172,MGM_W171,MGM_W170);
   and MGM_G208(MGM_W173,si_delay,MGM_W172);
   and MGM_G209(ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W173);
   not MGM_G210(MGM_W174,clk_delay);
   and MGM_G211(MGM_W175,d_delay,MGM_W174);
   and MGM_G212(MGM_W176,den_delay,MGM_W175);
   not MGM_G213(MGM_W177,si_delay);
   and MGM_G214(MGM_W178,MGM_W177,MGM_W176);
   not MGM_G215(MGM_W179,ssb_delay);
   and MGM_G216(ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W179,MGM_W178);
   not MGM_G217(MGM_W180,clk_delay);
   and MGM_G218(MGM_W181,d_delay,MGM_W180);
   and MGM_G219(MGM_W182,den_delay,MGM_W181);
   not MGM_G220(MGM_W183,si_delay);
   and MGM_G221(MGM_W184,MGM_W183,MGM_W182);
   and MGM_G222(ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W184);
   not MGM_G223(MGM_W185,clk_delay);
   and MGM_G224(MGM_W186,d_delay,MGM_W185);
   and MGM_G225(MGM_W187,den_delay,MGM_W186);
   and MGM_G226(MGM_W188,si_delay,MGM_W187);
   not MGM_G227(MGM_W189,ssb_delay);
   and MGM_G228(ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_NOT_ssb,MGM_W189,MGM_W188);
   not MGM_G229(MGM_W190,clk_delay);
   and MGM_G230(MGM_W191,d_delay,MGM_W190);
   and MGM_G231(MGM_W192,den_delay,MGM_W191);
   and MGM_G232(MGM_W193,si_delay,MGM_W192);
   and MGM_G233(ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W193);
   not MGM_G234(MGM_W194,d_delay);
   and MGM_G235(MGM_W195,MGM_W194,clk_delay);
   not MGM_G236(MGM_W196,den_delay);
   and MGM_G237(MGM_W197,MGM_W196,MGM_W195);
   not MGM_G238(MGM_W198,si_delay);
   and MGM_G239(MGM_W199,MGM_W198,MGM_W197);
   not MGM_G240(MGM_W200,ssb_delay);
   and MGM_G241(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W200,MGM_W199);
   not MGM_G242(MGM_W201,d_delay);
   and MGM_G243(MGM_W202,MGM_W201,clk_delay);
   not MGM_G244(MGM_W203,den_delay);
   and MGM_G245(MGM_W204,MGM_W203,MGM_W202);
   not MGM_G246(MGM_W205,si_delay);
   and MGM_G247(MGM_W206,MGM_W205,MGM_W204);
   and MGM_G248(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W206);
   not MGM_G249(MGM_W207,d_delay);
   and MGM_G250(MGM_W208,MGM_W207,clk_delay);
   not MGM_G251(MGM_W209,den_delay);
   and MGM_G252(MGM_W210,MGM_W209,MGM_W208);
   and MGM_G253(MGM_W211,si_delay,MGM_W210);
   not MGM_G254(MGM_W212,ssb_delay);
   and MGM_G255(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W212,MGM_W211);
   not MGM_G256(MGM_W213,d_delay);
   and MGM_G257(MGM_W214,MGM_W213,clk_delay);
   not MGM_G258(MGM_W215,den_delay);
   and MGM_G259(MGM_W216,MGM_W215,MGM_W214);
   and MGM_G260(MGM_W217,si_delay,MGM_W216);
   and MGM_G261(ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W217);
   not MGM_G262(MGM_W218,d_delay);
   and MGM_G263(MGM_W219,MGM_W218,clk_delay);
   and MGM_G264(MGM_W220,den_delay,MGM_W219);
   not MGM_G265(MGM_W221,si_delay);
   and MGM_G266(MGM_W222,MGM_W221,MGM_W220);
   not MGM_G267(MGM_W223,ssb_delay);
   and MGM_G268(ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W223,MGM_W222);
   not MGM_G269(MGM_W224,d_delay);
   and MGM_G270(MGM_W225,MGM_W224,clk_delay);
   and MGM_G271(MGM_W226,den_delay,MGM_W225);
   not MGM_G272(MGM_W227,si_delay);
   and MGM_G273(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G274(ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W228);
   not MGM_G275(MGM_W229,d_delay);
   and MGM_G276(MGM_W230,MGM_W229,clk_delay);
   and MGM_G277(MGM_W231,den_delay,MGM_W230);
   and MGM_G278(MGM_W232,si_delay,MGM_W231);
   not MGM_G279(MGM_W233,ssb_delay);
   and MGM_G280(ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb,MGM_W233,MGM_W232);
   not MGM_G281(MGM_W234,d_delay);
   and MGM_G282(MGM_W235,MGM_W234,clk_delay);
   and MGM_G283(MGM_W236,den_delay,MGM_W235);
   and MGM_G284(MGM_W237,si_delay,MGM_W236);
   and MGM_G285(ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W237);
   and MGM_G286(MGM_W238,d_delay,clk_delay);
   not MGM_G287(MGM_W239,den_delay);
   and MGM_G288(MGM_W240,MGM_W239,MGM_W238);
   not MGM_G289(MGM_W241,si_delay);
   and MGM_G290(MGM_W242,MGM_W241,MGM_W240);
   not MGM_G291(MGM_W243,ssb_delay);
   and MGM_G292(ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb,MGM_W243,MGM_W242);
   and MGM_G293(MGM_W244,d_delay,clk_delay);
   not MGM_G294(MGM_W245,den_delay);
   and MGM_G295(MGM_W246,MGM_W245,MGM_W244);
   not MGM_G296(MGM_W247,si_delay);
   and MGM_G297(MGM_W248,MGM_W247,MGM_W246);
   and MGM_G298(ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W248);
   and MGM_G299(MGM_W249,d_delay,clk_delay);
   not MGM_G300(MGM_W250,den_delay);
   and MGM_G301(MGM_W251,MGM_W250,MGM_W249);
   and MGM_G302(MGM_W252,si_delay,MGM_W251);
   not MGM_G303(MGM_W253,ssb_delay);
   and MGM_G304(ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb,MGM_W253,MGM_W252);
   and MGM_G305(MGM_W254,d_delay,clk_delay);
   not MGM_G306(MGM_W255,den_delay);
   and MGM_G307(MGM_W256,MGM_W255,MGM_W254);
   and MGM_G308(MGM_W257,si_delay,MGM_W256);
   and MGM_G309(ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_ssb,ssb_delay,MGM_W257);
   and MGM_G310(MGM_W258,d_delay,clk_delay);
   and MGM_G311(MGM_W259,den_delay,MGM_W258);
   not MGM_G312(MGM_W260,si_delay);
   and MGM_G313(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G314(MGM_W262,ssb_delay);
   and MGM_G315(ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   and MGM_G316(MGM_W263,d_delay,clk_delay);
   and MGM_G317(MGM_W264,den_delay,MGM_W263);
   not MGM_G318(MGM_W265,si_delay);
   and MGM_G319(MGM_W266,MGM_W265,MGM_W264);
   and MGM_G320(ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_ssb,ssb_delay,MGM_W266);
   and MGM_G321(MGM_W267,d_delay,clk_delay);
   and MGM_G322(MGM_W268,den_delay,MGM_W267);
   and MGM_G323(MGM_W269,si_delay,MGM_W268);
   not MGM_G324(MGM_W270,ssb_delay);
   and MGM_G325(ENABLE_clk_AND_d_AND_den_AND_si_AND_NOT_ssb,MGM_W270,MGM_W269);
   and MGM_G326(MGM_W271,d_delay,clk_delay);
   and MGM_G327(MGM_W272,den_delay,MGM_W271);
   and MGM_G328(MGM_W273,si_delay,MGM_W272);
   and MGM_G329(ENABLE_clk_AND_d_AND_den_AND_si_AND_ssb,ssb_delay,MGM_W273);
   not MGM_G330(MGM_W274,d_delay);
   not MGM_G331(MGM_W275,den_delay);
   and MGM_G332(MGM_W276,MGM_W275,MGM_W274);
   and MGM_G333(MGM_W277,rb_delay,MGM_W276);
   not MGM_G334(MGM_W278,ssb_delay);
   and MGM_G335(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb,MGM_W278,MGM_W277);
   not MGM_G336(MGM_W279,d_delay);
   and MGM_G337(MGM_W280,den_delay,MGM_W279);
   and MGM_G338(MGM_W281,rb_delay,MGM_W280);
   not MGM_G339(MGM_W282,ssb_delay);
   and MGM_G340(ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb,MGM_W282,MGM_W281);
   not MGM_G341(MGM_W283,den_delay);
   and MGM_G342(MGM_W284,MGM_W283,d_delay);
   and MGM_G343(MGM_W285,rb_delay,MGM_W284);
   not MGM_G344(MGM_W286,ssb_delay);
   and MGM_G345(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb,MGM_W286,MGM_W285);
   and MGM_G346(MGM_W287,den_delay,d_delay);
   and MGM_G347(MGM_W288,rb_delay,MGM_W287);
   not MGM_G348(MGM_W289,ssb_delay);
   and MGM_G349(ENABLE_d_AND_den_AND_rb_AND_NOT_ssb,MGM_W289,MGM_W288);
   not MGM_G350(MGM_W290,d_delay);
   not MGM_G351(MGM_W291,den_delay);
   and MGM_G352(MGM_W292,MGM_W291,MGM_W290);
   and MGM_G353(MGM_W293,rb_delay,MGM_W292);
   not MGM_G354(MGM_W294,si_delay);
   and MGM_G355(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si,MGM_W294,MGM_W293);
   not MGM_G356(MGM_W295,d_delay);
   not MGM_G357(MGM_W296,den_delay);
   and MGM_G358(MGM_W297,MGM_W296,MGM_W295);
   and MGM_G359(MGM_W298,rb_delay,MGM_W297);
   and MGM_G360(ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si,si_delay,MGM_W298);
   not MGM_G361(MGM_W299,d_delay);
   and MGM_G362(MGM_W300,den_delay,MGM_W299);
   and MGM_G363(MGM_W301,rb_delay,MGM_W300);
   and MGM_G364(ENABLE_NOT_d_AND_den_AND_rb_AND_si,si_delay,MGM_W301);
   not MGM_G365(MGM_W302,den_delay);
   and MGM_G366(MGM_W303,MGM_W302,d_delay);
   and MGM_G367(MGM_W304,rb_delay,MGM_W303);
   not MGM_G368(MGM_W305,si_delay);
   and MGM_G369(ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   not MGM_G370(MGM_W306,den_delay);
   and MGM_G371(MGM_W307,MGM_W306,d_delay);
   and MGM_G372(MGM_W308,rb_delay,MGM_W307);
   and MGM_G373(ENABLE_d_AND_NOT_den_AND_rb_AND_si,si_delay,MGM_W308);
   and MGM_G374(MGM_W309,den_delay,d_delay);
   and MGM_G375(MGM_W310,rb_delay,MGM_W309);
   not MGM_G376(MGM_W311,si_delay);
   and MGM_G377(ENABLE_d_AND_den_AND_rb_AND_NOT_si,MGM_W311,MGM_W310);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && den==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && den==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && den==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-LH
      $setuphold(posedge clk &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_den_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge den &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // setuphold den- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge den &&& (ENABLE_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,den_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d_AND_den_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_NOT_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d_AND_den_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold si- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,si_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_NOT_den_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_den_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fqy08fah_func( clkb, d, o, psb, rb, si, ssb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, psb, rb, si, ssb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_1( MGM_CLK0, clkb, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_P0, psb, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb, vcc, vssx );
   INTCseq_fqn00fah_LN_IQ_FF_UDP( IQ, MGM_C0, MGM_P0, MGM_CLK0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_1( MGM_CLK0, clkb );
   INTCseq_cdiar2ah_1( MGM_P0, psb );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_fdw003ah_5( MGM_D0, d, si, ssb );
   INTCseq_fqn00fah_LN_IQ_FF_UDP( IQ, MGM_C0, MGM_P0, MGM_CLK0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15fqy08fah1n02x5( clkb, d, o, psb, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, psb, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy08fah_func b15fqy08fah1n02x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy08fah_func b15fqy08fah1n02x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy08fah_func b15fqy08fah1n02x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy08fah_func b15fqy08fah1n02x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(MGM_W2,rb_delay,MGM_W1);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   and MGM_G8(MGM_W7,psb_delay,MGM_W6);
   and MGM_G9(MGM_W8,rb_delay,MGM_W7);
   not MGM_G10(MGM_W9,si_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G12(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W10);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,psb_delay,MGM_W11);
   and MGM_G15(MGM_W13,rb_delay,MGM_W12);
   and MGM_G16(MGM_W14,si_delay,MGM_W13);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,psb_delay,MGM_W16);
   and MGM_G21(MGM_W18,rb_delay,MGM_W17);
   and MGM_G22(MGM_W19,si_delay,MGM_W18);
   and MGM_G23(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W19);
   and MGM_G24(MGM_W20,psb_delay,d_delay);
   and MGM_G25(MGM_W21,rb_delay,MGM_W20);
   not MGM_G26(MGM_W22,si_delay);
   and MGM_G27(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G28(MGM_W24,ssb_delay);
   and MGM_G29(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W24,MGM_W23);
   and MGM_G30(MGM_W25,psb_delay,d_delay);
   and MGM_G31(MGM_W26,rb_delay,MGM_W25);
   not MGM_G32(MGM_W27,si_delay);
   and MGM_G33(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G34(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W28);
   and MGM_G35(MGM_W29,psb_delay,d_delay);
   and MGM_G36(MGM_W30,rb_delay,MGM_W29);
   and MGM_G37(MGM_W31,si_delay,MGM_W30);
   not MGM_G38(MGM_W32,ssb_delay);
   and MGM_G39(ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W32,MGM_W31);
   and MGM_G40(MGM_W33,psb_delay,d_delay);
   and MGM_G41(MGM_W34,rb_delay,MGM_W33);
   and MGM_G42(MGM_W35,si_delay,MGM_W34);
   and MGM_G43(ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G44(MGM_W36,rb_delay,psb_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   and MGM_G47(ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W38);
   and MGM_G48(MGM_W39,rb_delay,psb_delay);
   and MGM_G49(MGM_W40,si_delay,MGM_W39);
   and MGM_G50(ENABLE_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G51(MGM_W41,d_delay);
   and MGM_G52(MGM_W42,rb_delay,MGM_W41);
   not MGM_G53(MGM_W43,si_delay);
   and MGM_G54(MGM_W44,MGM_W43,MGM_W42);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   not MGM_G57(MGM_W46,d_delay);
   and MGM_G58(MGM_W47,rb_delay,MGM_W46);
   not MGM_G59(MGM_W48,si_delay);
   and MGM_G60(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G61(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G62(MGM_W50,d_delay);
   and MGM_G63(MGM_W51,rb_delay,MGM_W50);
   and MGM_G64(MGM_W52,si_delay,MGM_W51);
   and MGM_G65(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G66(MGM_W53,rb_delay,d_delay);
   not MGM_G67(MGM_W54,si_delay);
   and MGM_G68(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G69(MGM_W56,ssb_delay);
   and MGM_G70(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   not MGM_G71(MGM_W57,clkb_delay);
   not MGM_G72(MGM_W58,d_delay);
   and MGM_G73(MGM_W59,MGM_W58,MGM_W57);
   and MGM_G74(MGM_W60,rb_delay,MGM_W59);
   not MGM_G75(MGM_W61,si_delay);
   and MGM_G76(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G77(MGM_W63,ssb_delay);
   and MGM_G78(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G79(MGM_W64,clkb_delay);
   not MGM_G80(MGM_W65,d_delay);
   and MGM_G81(MGM_W66,MGM_W65,MGM_W64);
   and MGM_G82(MGM_W67,rb_delay,MGM_W66);
   not MGM_G83(MGM_W68,si_delay);
   and MGM_G84(MGM_W69,MGM_W68,MGM_W67);
   and MGM_G85(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W69);
   not MGM_G86(MGM_W70,clkb_delay);
   not MGM_G87(MGM_W71,d_delay);
   and MGM_G88(MGM_W72,MGM_W71,MGM_W70);
   and MGM_G89(MGM_W73,rb_delay,MGM_W72);
   and MGM_G90(MGM_W74,si_delay,MGM_W73);
   not MGM_G91(MGM_W75,ssb_delay);
   and MGM_G92(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G93(MGM_W76,clkb_delay);
   not MGM_G94(MGM_W77,d_delay);
   and MGM_G95(MGM_W78,MGM_W77,MGM_W76);
   and MGM_G96(MGM_W79,rb_delay,MGM_W78);
   and MGM_G97(MGM_W80,si_delay,MGM_W79);
   and MGM_G98(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W80);
   not MGM_G99(MGM_W81,clkb_delay);
   and MGM_G100(MGM_W82,d_delay,MGM_W81);
   and MGM_G101(MGM_W83,rb_delay,MGM_W82);
   not MGM_G102(MGM_W84,si_delay);
   and MGM_G103(MGM_W85,MGM_W84,MGM_W83);
   not MGM_G104(MGM_W86,ssb_delay);
   and MGM_G105(ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W86,MGM_W85);
   not MGM_G106(MGM_W87,clkb_delay);
   and MGM_G107(MGM_W88,d_delay,MGM_W87);
   and MGM_G108(MGM_W89,rb_delay,MGM_W88);
   not MGM_G109(MGM_W90,si_delay);
   and MGM_G110(MGM_W91,MGM_W90,MGM_W89);
   and MGM_G111(ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W91);
   not MGM_G112(MGM_W92,clkb_delay);
   and MGM_G113(MGM_W93,d_delay,MGM_W92);
   and MGM_G114(MGM_W94,rb_delay,MGM_W93);
   and MGM_G115(MGM_W95,si_delay,MGM_W94);
   not MGM_G116(MGM_W96,ssb_delay);
   and MGM_G117(ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W96,MGM_W95);
   not MGM_G118(MGM_W97,clkb_delay);
   and MGM_G119(MGM_W98,d_delay,MGM_W97);
   and MGM_G120(MGM_W99,rb_delay,MGM_W98);
   and MGM_G121(MGM_W100,si_delay,MGM_W99);
   and MGM_G122(ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W100);
   not MGM_G123(MGM_W101,d_delay);
   and MGM_G124(MGM_W102,MGM_W101,clkb_delay);
   and MGM_G125(MGM_W103,rb_delay,MGM_W102);
   not MGM_G126(MGM_W104,si_delay);
   and MGM_G127(MGM_W105,MGM_W104,MGM_W103);
   not MGM_G128(MGM_W106,ssb_delay);
   and MGM_G129(ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W106,MGM_W105);
   not MGM_G130(MGM_W107,d_delay);
   and MGM_G131(MGM_W108,MGM_W107,clkb_delay);
   and MGM_G132(MGM_W109,rb_delay,MGM_W108);
   not MGM_G133(MGM_W110,si_delay);
   and MGM_G134(MGM_W111,MGM_W110,MGM_W109);
   and MGM_G135(ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W111);
   not MGM_G136(MGM_W112,d_delay);
   and MGM_G137(MGM_W113,MGM_W112,clkb_delay);
   and MGM_G138(MGM_W114,rb_delay,MGM_W113);
   and MGM_G139(MGM_W115,si_delay,MGM_W114);
   not MGM_G140(MGM_W116,ssb_delay);
   and MGM_G141(ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W116,MGM_W115);
   not MGM_G142(MGM_W117,d_delay);
   and MGM_G143(MGM_W118,MGM_W117,clkb_delay);
   and MGM_G144(MGM_W119,rb_delay,MGM_W118);
   and MGM_G145(MGM_W120,si_delay,MGM_W119);
   and MGM_G146(ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W120);
   and MGM_G147(MGM_W121,d_delay,clkb_delay);
   and MGM_G148(MGM_W122,rb_delay,MGM_W121);
   not MGM_G149(MGM_W123,si_delay);
   and MGM_G150(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G151(MGM_W125,ssb_delay);
   and MGM_G152(ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W125,MGM_W124);
   and MGM_G153(MGM_W126,d_delay,clkb_delay);
   and MGM_G154(MGM_W127,rb_delay,MGM_W126);
   not MGM_G155(MGM_W128,si_delay);
   and MGM_G156(MGM_W129,MGM_W128,MGM_W127);
   and MGM_G157(ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W129);
   and MGM_G158(MGM_W130,d_delay,clkb_delay);
   and MGM_G159(MGM_W131,rb_delay,MGM_W130);
   and MGM_G160(MGM_W132,si_delay,MGM_W131);
   not MGM_G161(MGM_W133,ssb_delay);
   and MGM_G162(ENABLE_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W133,MGM_W132);
   and MGM_G163(MGM_W134,d_delay,clkb_delay);
   and MGM_G164(MGM_W135,rb_delay,MGM_W134);
   and MGM_G165(MGM_W136,si_delay,MGM_W135);
   and MGM_G166(ENABLE_clkb_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W136);
   not MGM_G167(MGM_W137,clkb_delay);
   not MGM_G168(MGM_W138,d_delay);
   and MGM_G169(MGM_W139,MGM_W138,MGM_W137);
   not MGM_G170(MGM_W140,si_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   not MGM_G172(MGM_W142,ssb_delay);
   and MGM_G173(ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W142,MGM_W141);
   not MGM_G174(MGM_W143,clkb_delay);
   not MGM_G175(MGM_W144,d_delay);
   and MGM_G176(MGM_W145,MGM_W144,MGM_W143);
   not MGM_G177(MGM_W146,si_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W147);
   not MGM_G180(MGM_W148,clkb_delay);
   not MGM_G181(MGM_W149,d_delay);
   and MGM_G182(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G183(MGM_W151,si_delay,MGM_W150);
   not MGM_G184(MGM_W152,ssb_delay);
   and MGM_G185(ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W153,clkb_delay);
   not MGM_G187(MGM_W154,d_delay);
   and MGM_G188(MGM_W155,MGM_W154,MGM_W153);
   and MGM_G189(MGM_W156,si_delay,MGM_W155);
   and MGM_G190(ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W156);
   not MGM_G191(MGM_W157,clkb_delay);
   and MGM_G192(MGM_W158,d_delay,MGM_W157);
   not MGM_G193(MGM_W159,si_delay);
   and MGM_G194(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G195(MGM_W161,ssb_delay);
   and MGM_G196(ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W161,MGM_W160);
   not MGM_G197(MGM_W162,clkb_delay);
   and MGM_G198(MGM_W163,d_delay,MGM_W162);
   not MGM_G199(MGM_W164,si_delay);
   and MGM_G200(MGM_W165,MGM_W164,MGM_W163);
   and MGM_G201(ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W165);
   not MGM_G202(MGM_W166,clkb_delay);
   and MGM_G203(MGM_W167,d_delay,MGM_W166);
   and MGM_G204(MGM_W168,si_delay,MGM_W167);
   not MGM_G205(MGM_W169,ssb_delay);
   and MGM_G206(ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb,MGM_W169,MGM_W168);
   not MGM_G207(MGM_W170,clkb_delay);
   and MGM_G208(MGM_W171,d_delay,MGM_W170);
   and MGM_G209(MGM_W172,si_delay,MGM_W171);
   and MGM_G210(ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W172);
   not MGM_G211(MGM_W173,d_delay);
   and MGM_G212(MGM_W174,MGM_W173,clkb_delay);
   not MGM_G213(MGM_W175,si_delay);
   and MGM_G214(MGM_W176,MGM_W175,MGM_W174);
   not MGM_G215(MGM_W177,ssb_delay);
   and MGM_G216(ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W177,MGM_W176);
   not MGM_G217(MGM_W178,d_delay);
   and MGM_G218(MGM_W179,MGM_W178,clkb_delay);
   not MGM_G219(MGM_W180,si_delay);
   and MGM_G220(MGM_W181,MGM_W180,MGM_W179);
   and MGM_G221(ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W181);
   not MGM_G222(MGM_W182,d_delay);
   and MGM_G223(MGM_W183,MGM_W182,clkb_delay);
   and MGM_G224(MGM_W184,si_delay,MGM_W183);
   not MGM_G225(MGM_W185,ssb_delay);
   and MGM_G226(ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W185,MGM_W184);
   not MGM_G227(MGM_W186,d_delay);
   and MGM_G228(MGM_W187,MGM_W186,clkb_delay);
   and MGM_G229(MGM_W188,si_delay,MGM_W187);
   and MGM_G230(ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W188);
   and MGM_G231(MGM_W189,d_delay,clkb_delay);
   not MGM_G232(MGM_W190,si_delay);
   and MGM_G233(MGM_W191,MGM_W190,MGM_W189);
   not MGM_G234(MGM_W192,ssb_delay);
   and MGM_G235(ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W192,MGM_W191);
   and MGM_G236(MGM_W193,d_delay,clkb_delay);
   not MGM_G237(MGM_W194,si_delay);
   and MGM_G238(MGM_W195,MGM_W194,MGM_W193);
   and MGM_G239(ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W195);
   and MGM_G240(MGM_W196,d_delay,clkb_delay);
   and MGM_G241(MGM_W197,si_delay,MGM_W196);
   not MGM_G242(MGM_W198,ssb_delay);
   and MGM_G243(ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb,MGM_W198,MGM_W197);
   and MGM_G244(MGM_W199,d_delay,clkb_delay);
   and MGM_G245(MGM_W200,si_delay,MGM_W199);
   and MGM_G246(ENABLE_clkb_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W200);
   not MGM_G247(MGM_W201,d_delay);
   and MGM_G248(MGM_W202,psb_delay,MGM_W201);
   and MGM_G249(MGM_W203,si_delay,MGM_W202);
   not MGM_G250(MGM_W204,ssb_delay);
   and MGM_G251(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W204,MGM_W203);
   and MGM_G252(MGM_W205,psb_delay,d_delay);
   not MGM_G253(MGM_W206,si_delay);
   and MGM_G254(MGM_W207,MGM_W206,MGM_W205);
   and MGM_G255(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W207);
   and MGM_G256(MGM_W208,psb_delay,d_delay);
   and MGM_G257(MGM_W209,si_delay,MGM_W208);
   not MGM_G258(MGM_W210,ssb_delay);
   and MGM_G259(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W210,MGM_W209);
   and MGM_G260(MGM_W211,psb_delay,d_delay);
   and MGM_G261(MGM_W212,si_delay,MGM_W211);
   and MGM_G262(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W212);
   not MGM_G263(MGM_W213,clkb_delay);
   not MGM_G264(MGM_W214,d_delay);
   and MGM_G265(MGM_W215,MGM_W214,MGM_W213);
   and MGM_G266(MGM_W216,psb_delay,MGM_W215);
   not MGM_G267(MGM_W217,si_delay);
   and MGM_G268(MGM_W218,MGM_W217,MGM_W216);
   not MGM_G269(MGM_W219,ssb_delay);
   and MGM_G270(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W219,MGM_W218);
   not MGM_G271(MGM_W220,clkb_delay);
   not MGM_G272(MGM_W221,d_delay);
   and MGM_G273(MGM_W222,MGM_W221,MGM_W220);
   and MGM_G274(MGM_W223,psb_delay,MGM_W222);
   not MGM_G275(MGM_W224,si_delay);
   and MGM_G276(MGM_W225,MGM_W224,MGM_W223);
   and MGM_G277(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W225);
   not MGM_G278(MGM_W226,clkb_delay);
   not MGM_G279(MGM_W227,d_delay);
   and MGM_G280(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G281(MGM_W229,psb_delay,MGM_W228);
   and MGM_G282(MGM_W230,si_delay,MGM_W229);
   not MGM_G283(MGM_W231,ssb_delay);
   and MGM_G284(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W231,MGM_W230);
   not MGM_G285(MGM_W232,clkb_delay);
   not MGM_G286(MGM_W233,d_delay);
   and MGM_G287(MGM_W234,MGM_W233,MGM_W232);
   and MGM_G288(MGM_W235,psb_delay,MGM_W234);
   and MGM_G289(MGM_W236,si_delay,MGM_W235);
   and MGM_G290(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W236);
   not MGM_G291(MGM_W237,clkb_delay);
   and MGM_G292(MGM_W238,d_delay,MGM_W237);
   and MGM_G293(MGM_W239,psb_delay,MGM_W238);
   not MGM_G294(MGM_W240,si_delay);
   and MGM_G295(MGM_W241,MGM_W240,MGM_W239);
   not MGM_G296(MGM_W242,ssb_delay);
   and MGM_G297(ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W242,MGM_W241);
   not MGM_G298(MGM_W243,clkb_delay);
   and MGM_G299(MGM_W244,d_delay,MGM_W243);
   and MGM_G300(MGM_W245,psb_delay,MGM_W244);
   not MGM_G301(MGM_W246,si_delay);
   and MGM_G302(MGM_W247,MGM_W246,MGM_W245);
   and MGM_G303(ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W247);
   not MGM_G304(MGM_W248,clkb_delay);
   and MGM_G305(MGM_W249,d_delay,MGM_W248);
   and MGM_G306(MGM_W250,psb_delay,MGM_W249);
   and MGM_G307(MGM_W251,si_delay,MGM_W250);
   not MGM_G308(MGM_W252,ssb_delay);
   and MGM_G309(ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W252,MGM_W251);
   not MGM_G310(MGM_W253,clkb_delay);
   and MGM_G311(MGM_W254,d_delay,MGM_W253);
   and MGM_G312(MGM_W255,psb_delay,MGM_W254);
   and MGM_G313(MGM_W256,si_delay,MGM_W255);
   and MGM_G314(ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W256);
   not MGM_G315(MGM_W257,d_delay);
   and MGM_G316(MGM_W258,MGM_W257,clkb_delay);
   and MGM_G317(MGM_W259,psb_delay,MGM_W258);
   not MGM_G318(MGM_W260,si_delay);
   and MGM_G319(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G320(MGM_W262,ssb_delay);
   and MGM_G321(ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   not MGM_G322(MGM_W263,d_delay);
   and MGM_G323(MGM_W264,MGM_W263,clkb_delay);
   and MGM_G324(MGM_W265,psb_delay,MGM_W264);
   not MGM_G325(MGM_W266,si_delay);
   and MGM_G326(MGM_W267,MGM_W266,MGM_W265);
   and MGM_G327(ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W267);
   not MGM_G328(MGM_W268,d_delay);
   and MGM_G329(MGM_W269,MGM_W268,clkb_delay);
   and MGM_G330(MGM_W270,psb_delay,MGM_W269);
   and MGM_G331(MGM_W271,si_delay,MGM_W270);
   not MGM_G332(MGM_W272,ssb_delay);
   and MGM_G333(ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W272,MGM_W271);
   not MGM_G334(MGM_W273,d_delay);
   and MGM_G335(MGM_W274,MGM_W273,clkb_delay);
   and MGM_G336(MGM_W275,psb_delay,MGM_W274);
   and MGM_G337(MGM_W276,si_delay,MGM_W275);
   and MGM_G338(ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W276);
   and MGM_G339(MGM_W277,d_delay,clkb_delay);
   and MGM_G340(MGM_W278,psb_delay,MGM_W277);
   not MGM_G341(MGM_W279,si_delay);
   and MGM_G342(MGM_W280,MGM_W279,MGM_W278);
   not MGM_G343(MGM_W281,ssb_delay);
   and MGM_G344(ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W281,MGM_W280);
   and MGM_G345(MGM_W282,d_delay,clkb_delay);
   and MGM_G346(MGM_W283,psb_delay,MGM_W282);
   not MGM_G347(MGM_W284,si_delay);
   and MGM_G348(MGM_W285,MGM_W284,MGM_W283);
   and MGM_G349(ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W285);
   and MGM_G350(MGM_W286,d_delay,clkb_delay);
   and MGM_G351(MGM_W287,psb_delay,MGM_W286);
   and MGM_G352(MGM_W288,si_delay,MGM_W287);
   not MGM_G353(MGM_W289,ssb_delay);
   and MGM_G354(ENABLE_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W289,MGM_W288);
   and MGM_G355(MGM_W290,d_delay,clkb_delay);
   and MGM_G356(MGM_W291,psb_delay,MGM_W290);
   and MGM_G357(MGM_W292,si_delay,MGM_W291);
   and MGM_G358(ENABLE_clkb_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W292);
   not MGM_G359(MGM_W293,d_delay);
   and MGM_G360(MGM_W294,psb_delay,MGM_W293);
   and MGM_G361(MGM_W295,rb_delay,MGM_W294);
   not MGM_G362(MGM_W296,ssb_delay);
   and MGM_G363(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W296,MGM_W295);
   and MGM_G364(MGM_W297,psb_delay,d_delay);
   and MGM_G365(MGM_W298,rb_delay,MGM_W297);
   not MGM_G366(MGM_W299,ssb_delay);
   and MGM_G367(ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W299,MGM_W298);
   not MGM_G368(MGM_W300,d_delay);
   and MGM_G369(MGM_W301,psb_delay,MGM_W300);
   and MGM_G370(MGM_W302,rb_delay,MGM_W301);
   and MGM_G371(ENABLE_NOT_d_AND_psb_AND_rb_AND_si,si_delay,MGM_W302);
   and MGM_G372(MGM_W303,psb_delay,d_delay);
   and MGM_G373(MGM_W304,rb_delay,MGM_W303);
   not MGM_G374(MGM_W305,si_delay);
   and MGM_G375(ENABLE_d_AND_psb_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy08fah1n04x5( clkb, d, o, psb, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, psb, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy08fah_func b15fqy08fah1n04x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy08fah_func b15fqy08fah1n04x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy08fah_func b15fqy08fah1n04x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy08fah_func b15fqy08fah1n04x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(MGM_W2,rb_delay,MGM_W1);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   and MGM_G8(MGM_W7,psb_delay,MGM_W6);
   and MGM_G9(MGM_W8,rb_delay,MGM_W7);
   not MGM_G10(MGM_W9,si_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G12(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W10);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,psb_delay,MGM_W11);
   and MGM_G15(MGM_W13,rb_delay,MGM_W12);
   and MGM_G16(MGM_W14,si_delay,MGM_W13);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,psb_delay,MGM_W16);
   and MGM_G21(MGM_W18,rb_delay,MGM_W17);
   and MGM_G22(MGM_W19,si_delay,MGM_W18);
   and MGM_G23(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W19);
   and MGM_G24(MGM_W20,psb_delay,d_delay);
   and MGM_G25(MGM_W21,rb_delay,MGM_W20);
   not MGM_G26(MGM_W22,si_delay);
   and MGM_G27(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G28(MGM_W24,ssb_delay);
   and MGM_G29(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W24,MGM_W23);
   and MGM_G30(MGM_W25,psb_delay,d_delay);
   and MGM_G31(MGM_W26,rb_delay,MGM_W25);
   not MGM_G32(MGM_W27,si_delay);
   and MGM_G33(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G34(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W28);
   and MGM_G35(MGM_W29,psb_delay,d_delay);
   and MGM_G36(MGM_W30,rb_delay,MGM_W29);
   and MGM_G37(MGM_W31,si_delay,MGM_W30);
   not MGM_G38(MGM_W32,ssb_delay);
   and MGM_G39(ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W32,MGM_W31);
   and MGM_G40(MGM_W33,psb_delay,d_delay);
   and MGM_G41(MGM_W34,rb_delay,MGM_W33);
   and MGM_G42(MGM_W35,si_delay,MGM_W34);
   and MGM_G43(ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G44(MGM_W36,rb_delay,psb_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   and MGM_G47(ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W38);
   and MGM_G48(MGM_W39,rb_delay,psb_delay);
   and MGM_G49(MGM_W40,si_delay,MGM_W39);
   and MGM_G50(ENABLE_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G51(MGM_W41,d_delay);
   and MGM_G52(MGM_W42,rb_delay,MGM_W41);
   not MGM_G53(MGM_W43,si_delay);
   and MGM_G54(MGM_W44,MGM_W43,MGM_W42);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   not MGM_G57(MGM_W46,d_delay);
   and MGM_G58(MGM_W47,rb_delay,MGM_W46);
   not MGM_G59(MGM_W48,si_delay);
   and MGM_G60(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G61(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G62(MGM_W50,d_delay);
   and MGM_G63(MGM_W51,rb_delay,MGM_W50);
   and MGM_G64(MGM_W52,si_delay,MGM_W51);
   and MGM_G65(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G66(MGM_W53,rb_delay,d_delay);
   not MGM_G67(MGM_W54,si_delay);
   and MGM_G68(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G69(MGM_W56,ssb_delay);
   and MGM_G70(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   not MGM_G71(MGM_W57,clkb_delay);
   not MGM_G72(MGM_W58,d_delay);
   and MGM_G73(MGM_W59,MGM_W58,MGM_W57);
   and MGM_G74(MGM_W60,rb_delay,MGM_W59);
   not MGM_G75(MGM_W61,si_delay);
   and MGM_G76(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G77(MGM_W63,ssb_delay);
   and MGM_G78(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G79(MGM_W64,clkb_delay);
   not MGM_G80(MGM_W65,d_delay);
   and MGM_G81(MGM_W66,MGM_W65,MGM_W64);
   and MGM_G82(MGM_W67,rb_delay,MGM_W66);
   not MGM_G83(MGM_W68,si_delay);
   and MGM_G84(MGM_W69,MGM_W68,MGM_W67);
   and MGM_G85(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W69);
   not MGM_G86(MGM_W70,clkb_delay);
   not MGM_G87(MGM_W71,d_delay);
   and MGM_G88(MGM_W72,MGM_W71,MGM_W70);
   and MGM_G89(MGM_W73,rb_delay,MGM_W72);
   and MGM_G90(MGM_W74,si_delay,MGM_W73);
   not MGM_G91(MGM_W75,ssb_delay);
   and MGM_G92(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G93(MGM_W76,clkb_delay);
   not MGM_G94(MGM_W77,d_delay);
   and MGM_G95(MGM_W78,MGM_W77,MGM_W76);
   and MGM_G96(MGM_W79,rb_delay,MGM_W78);
   and MGM_G97(MGM_W80,si_delay,MGM_W79);
   and MGM_G98(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W80);
   not MGM_G99(MGM_W81,clkb_delay);
   and MGM_G100(MGM_W82,d_delay,MGM_W81);
   and MGM_G101(MGM_W83,rb_delay,MGM_W82);
   not MGM_G102(MGM_W84,si_delay);
   and MGM_G103(MGM_W85,MGM_W84,MGM_W83);
   not MGM_G104(MGM_W86,ssb_delay);
   and MGM_G105(ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W86,MGM_W85);
   not MGM_G106(MGM_W87,clkb_delay);
   and MGM_G107(MGM_W88,d_delay,MGM_W87);
   and MGM_G108(MGM_W89,rb_delay,MGM_W88);
   not MGM_G109(MGM_W90,si_delay);
   and MGM_G110(MGM_W91,MGM_W90,MGM_W89);
   and MGM_G111(ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W91);
   not MGM_G112(MGM_W92,clkb_delay);
   and MGM_G113(MGM_W93,d_delay,MGM_W92);
   and MGM_G114(MGM_W94,rb_delay,MGM_W93);
   and MGM_G115(MGM_W95,si_delay,MGM_W94);
   not MGM_G116(MGM_W96,ssb_delay);
   and MGM_G117(ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W96,MGM_W95);
   not MGM_G118(MGM_W97,clkb_delay);
   and MGM_G119(MGM_W98,d_delay,MGM_W97);
   and MGM_G120(MGM_W99,rb_delay,MGM_W98);
   and MGM_G121(MGM_W100,si_delay,MGM_W99);
   and MGM_G122(ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W100);
   not MGM_G123(MGM_W101,d_delay);
   and MGM_G124(MGM_W102,MGM_W101,clkb_delay);
   and MGM_G125(MGM_W103,rb_delay,MGM_W102);
   not MGM_G126(MGM_W104,si_delay);
   and MGM_G127(MGM_W105,MGM_W104,MGM_W103);
   not MGM_G128(MGM_W106,ssb_delay);
   and MGM_G129(ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W106,MGM_W105);
   not MGM_G130(MGM_W107,d_delay);
   and MGM_G131(MGM_W108,MGM_W107,clkb_delay);
   and MGM_G132(MGM_W109,rb_delay,MGM_W108);
   not MGM_G133(MGM_W110,si_delay);
   and MGM_G134(MGM_W111,MGM_W110,MGM_W109);
   and MGM_G135(ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W111);
   not MGM_G136(MGM_W112,d_delay);
   and MGM_G137(MGM_W113,MGM_W112,clkb_delay);
   and MGM_G138(MGM_W114,rb_delay,MGM_W113);
   and MGM_G139(MGM_W115,si_delay,MGM_W114);
   not MGM_G140(MGM_W116,ssb_delay);
   and MGM_G141(ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W116,MGM_W115);
   not MGM_G142(MGM_W117,d_delay);
   and MGM_G143(MGM_W118,MGM_W117,clkb_delay);
   and MGM_G144(MGM_W119,rb_delay,MGM_W118);
   and MGM_G145(MGM_W120,si_delay,MGM_W119);
   and MGM_G146(ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W120);
   and MGM_G147(MGM_W121,d_delay,clkb_delay);
   and MGM_G148(MGM_W122,rb_delay,MGM_W121);
   not MGM_G149(MGM_W123,si_delay);
   and MGM_G150(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G151(MGM_W125,ssb_delay);
   and MGM_G152(ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W125,MGM_W124);
   and MGM_G153(MGM_W126,d_delay,clkb_delay);
   and MGM_G154(MGM_W127,rb_delay,MGM_W126);
   not MGM_G155(MGM_W128,si_delay);
   and MGM_G156(MGM_W129,MGM_W128,MGM_W127);
   and MGM_G157(ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W129);
   and MGM_G158(MGM_W130,d_delay,clkb_delay);
   and MGM_G159(MGM_W131,rb_delay,MGM_W130);
   and MGM_G160(MGM_W132,si_delay,MGM_W131);
   not MGM_G161(MGM_W133,ssb_delay);
   and MGM_G162(ENABLE_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W133,MGM_W132);
   and MGM_G163(MGM_W134,d_delay,clkb_delay);
   and MGM_G164(MGM_W135,rb_delay,MGM_W134);
   and MGM_G165(MGM_W136,si_delay,MGM_W135);
   and MGM_G166(ENABLE_clkb_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W136);
   not MGM_G167(MGM_W137,clkb_delay);
   not MGM_G168(MGM_W138,d_delay);
   and MGM_G169(MGM_W139,MGM_W138,MGM_W137);
   not MGM_G170(MGM_W140,si_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   not MGM_G172(MGM_W142,ssb_delay);
   and MGM_G173(ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W142,MGM_W141);
   not MGM_G174(MGM_W143,clkb_delay);
   not MGM_G175(MGM_W144,d_delay);
   and MGM_G176(MGM_W145,MGM_W144,MGM_W143);
   not MGM_G177(MGM_W146,si_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W147);
   not MGM_G180(MGM_W148,clkb_delay);
   not MGM_G181(MGM_W149,d_delay);
   and MGM_G182(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G183(MGM_W151,si_delay,MGM_W150);
   not MGM_G184(MGM_W152,ssb_delay);
   and MGM_G185(ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W153,clkb_delay);
   not MGM_G187(MGM_W154,d_delay);
   and MGM_G188(MGM_W155,MGM_W154,MGM_W153);
   and MGM_G189(MGM_W156,si_delay,MGM_W155);
   and MGM_G190(ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W156);
   not MGM_G191(MGM_W157,clkb_delay);
   and MGM_G192(MGM_W158,d_delay,MGM_W157);
   not MGM_G193(MGM_W159,si_delay);
   and MGM_G194(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G195(MGM_W161,ssb_delay);
   and MGM_G196(ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W161,MGM_W160);
   not MGM_G197(MGM_W162,clkb_delay);
   and MGM_G198(MGM_W163,d_delay,MGM_W162);
   not MGM_G199(MGM_W164,si_delay);
   and MGM_G200(MGM_W165,MGM_W164,MGM_W163);
   and MGM_G201(ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W165);
   not MGM_G202(MGM_W166,clkb_delay);
   and MGM_G203(MGM_W167,d_delay,MGM_W166);
   and MGM_G204(MGM_W168,si_delay,MGM_W167);
   not MGM_G205(MGM_W169,ssb_delay);
   and MGM_G206(ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb,MGM_W169,MGM_W168);
   not MGM_G207(MGM_W170,clkb_delay);
   and MGM_G208(MGM_W171,d_delay,MGM_W170);
   and MGM_G209(MGM_W172,si_delay,MGM_W171);
   and MGM_G210(ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W172);
   not MGM_G211(MGM_W173,d_delay);
   and MGM_G212(MGM_W174,MGM_W173,clkb_delay);
   not MGM_G213(MGM_W175,si_delay);
   and MGM_G214(MGM_W176,MGM_W175,MGM_W174);
   not MGM_G215(MGM_W177,ssb_delay);
   and MGM_G216(ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W177,MGM_W176);
   not MGM_G217(MGM_W178,d_delay);
   and MGM_G218(MGM_W179,MGM_W178,clkb_delay);
   not MGM_G219(MGM_W180,si_delay);
   and MGM_G220(MGM_W181,MGM_W180,MGM_W179);
   and MGM_G221(ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W181);
   not MGM_G222(MGM_W182,d_delay);
   and MGM_G223(MGM_W183,MGM_W182,clkb_delay);
   and MGM_G224(MGM_W184,si_delay,MGM_W183);
   not MGM_G225(MGM_W185,ssb_delay);
   and MGM_G226(ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W185,MGM_W184);
   not MGM_G227(MGM_W186,d_delay);
   and MGM_G228(MGM_W187,MGM_W186,clkb_delay);
   and MGM_G229(MGM_W188,si_delay,MGM_W187);
   and MGM_G230(ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W188);
   and MGM_G231(MGM_W189,d_delay,clkb_delay);
   not MGM_G232(MGM_W190,si_delay);
   and MGM_G233(MGM_W191,MGM_W190,MGM_W189);
   not MGM_G234(MGM_W192,ssb_delay);
   and MGM_G235(ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W192,MGM_W191);
   and MGM_G236(MGM_W193,d_delay,clkb_delay);
   not MGM_G237(MGM_W194,si_delay);
   and MGM_G238(MGM_W195,MGM_W194,MGM_W193);
   and MGM_G239(ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W195);
   and MGM_G240(MGM_W196,d_delay,clkb_delay);
   and MGM_G241(MGM_W197,si_delay,MGM_W196);
   not MGM_G242(MGM_W198,ssb_delay);
   and MGM_G243(ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb,MGM_W198,MGM_W197);
   and MGM_G244(MGM_W199,d_delay,clkb_delay);
   and MGM_G245(MGM_W200,si_delay,MGM_W199);
   and MGM_G246(ENABLE_clkb_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W200);
   not MGM_G247(MGM_W201,d_delay);
   and MGM_G248(MGM_W202,psb_delay,MGM_W201);
   and MGM_G249(MGM_W203,si_delay,MGM_W202);
   not MGM_G250(MGM_W204,ssb_delay);
   and MGM_G251(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W204,MGM_W203);
   and MGM_G252(MGM_W205,psb_delay,d_delay);
   not MGM_G253(MGM_W206,si_delay);
   and MGM_G254(MGM_W207,MGM_W206,MGM_W205);
   and MGM_G255(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W207);
   and MGM_G256(MGM_W208,psb_delay,d_delay);
   and MGM_G257(MGM_W209,si_delay,MGM_W208);
   not MGM_G258(MGM_W210,ssb_delay);
   and MGM_G259(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W210,MGM_W209);
   and MGM_G260(MGM_W211,psb_delay,d_delay);
   and MGM_G261(MGM_W212,si_delay,MGM_W211);
   and MGM_G262(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W212);
   not MGM_G263(MGM_W213,clkb_delay);
   not MGM_G264(MGM_W214,d_delay);
   and MGM_G265(MGM_W215,MGM_W214,MGM_W213);
   and MGM_G266(MGM_W216,psb_delay,MGM_W215);
   not MGM_G267(MGM_W217,si_delay);
   and MGM_G268(MGM_W218,MGM_W217,MGM_W216);
   not MGM_G269(MGM_W219,ssb_delay);
   and MGM_G270(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W219,MGM_W218);
   not MGM_G271(MGM_W220,clkb_delay);
   not MGM_G272(MGM_W221,d_delay);
   and MGM_G273(MGM_W222,MGM_W221,MGM_W220);
   and MGM_G274(MGM_W223,psb_delay,MGM_W222);
   not MGM_G275(MGM_W224,si_delay);
   and MGM_G276(MGM_W225,MGM_W224,MGM_W223);
   and MGM_G277(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W225);
   not MGM_G278(MGM_W226,clkb_delay);
   not MGM_G279(MGM_W227,d_delay);
   and MGM_G280(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G281(MGM_W229,psb_delay,MGM_W228);
   and MGM_G282(MGM_W230,si_delay,MGM_W229);
   not MGM_G283(MGM_W231,ssb_delay);
   and MGM_G284(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W231,MGM_W230);
   not MGM_G285(MGM_W232,clkb_delay);
   not MGM_G286(MGM_W233,d_delay);
   and MGM_G287(MGM_W234,MGM_W233,MGM_W232);
   and MGM_G288(MGM_W235,psb_delay,MGM_W234);
   and MGM_G289(MGM_W236,si_delay,MGM_W235);
   and MGM_G290(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W236);
   not MGM_G291(MGM_W237,clkb_delay);
   and MGM_G292(MGM_W238,d_delay,MGM_W237);
   and MGM_G293(MGM_W239,psb_delay,MGM_W238);
   not MGM_G294(MGM_W240,si_delay);
   and MGM_G295(MGM_W241,MGM_W240,MGM_W239);
   not MGM_G296(MGM_W242,ssb_delay);
   and MGM_G297(ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W242,MGM_W241);
   not MGM_G298(MGM_W243,clkb_delay);
   and MGM_G299(MGM_W244,d_delay,MGM_W243);
   and MGM_G300(MGM_W245,psb_delay,MGM_W244);
   not MGM_G301(MGM_W246,si_delay);
   and MGM_G302(MGM_W247,MGM_W246,MGM_W245);
   and MGM_G303(ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W247);
   not MGM_G304(MGM_W248,clkb_delay);
   and MGM_G305(MGM_W249,d_delay,MGM_W248);
   and MGM_G306(MGM_W250,psb_delay,MGM_W249);
   and MGM_G307(MGM_W251,si_delay,MGM_W250);
   not MGM_G308(MGM_W252,ssb_delay);
   and MGM_G309(ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W252,MGM_W251);
   not MGM_G310(MGM_W253,clkb_delay);
   and MGM_G311(MGM_W254,d_delay,MGM_W253);
   and MGM_G312(MGM_W255,psb_delay,MGM_W254);
   and MGM_G313(MGM_W256,si_delay,MGM_W255);
   and MGM_G314(ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W256);
   not MGM_G315(MGM_W257,d_delay);
   and MGM_G316(MGM_W258,MGM_W257,clkb_delay);
   and MGM_G317(MGM_W259,psb_delay,MGM_W258);
   not MGM_G318(MGM_W260,si_delay);
   and MGM_G319(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G320(MGM_W262,ssb_delay);
   and MGM_G321(ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   not MGM_G322(MGM_W263,d_delay);
   and MGM_G323(MGM_W264,MGM_W263,clkb_delay);
   and MGM_G324(MGM_W265,psb_delay,MGM_W264);
   not MGM_G325(MGM_W266,si_delay);
   and MGM_G326(MGM_W267,MGM_W266,MGM_W265);
   and MGM_G327(ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W267);
   not MGM_G328(MGM_W268,d_delay);
   and MGM_G329(MGM_W269,MGM_W268,clkb_delay);
   and MGM_G330(MGM_W270,psb_delay,MGM_W269);
   and MGM_G331(MGM_W271,si_delay,MGM_W270);
   not MGM_G332(MGM_W272,ssb_delay);
   and MGM_G333(ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W272,MGM_W271);
   not MGM_G334(MGM_W273,d_delay);
   and MGM_G335(MGM_W274,MGM_W273,clkb_delay);
   and MGM_G336(MGM_W275,psb_delay,MGM_W274);
   and MGM_G337(MGM_W276,si_delay,MGM_W275);
   and MGM_G338(ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W276);
   and MGM_G339(MGM_W277,d_delay,clkb_delay);
   and MGM_G340(MGM_W278,psb_delay,MGM_W277);
   not MGM_G341(MGM_W279,si_delay);
   and MGM_G342(MGM_W280,MGM_W279,MGM_W278);
   not MGM_G343(MGM_W281,ssb_delay);
   and MGM_G344(ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W281,MGM_W280);
   and MGM_G345(MGM_W282,d_delay,clkb_delay);
   and MGM_G346(MGM_W283,psb_delay,MGM_W282);
   not MGM_G347(MGM_W284,si_delay);
   and MGM_G348(MGM_W285,MGM_W284,MGM_W283);
   and MGM_G349(ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W285);
   and MGM_G350(MGM_W286,d_delay,clkb_delay);
   and MGM_G351(MGM_W287,psb_delay,MGM_W286);
   and MGM_G352(MGM_W288,si_delay,MGM_W287);
   not MGM_G353(MGM_W289,ssb_delay);
   and MGM_G354(ENABLE_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W289,MGM_W288);
   and MGM_G355(MGM_W290,d_delay,clkb_delay);
   and MGM_G356(MGM_W291,psb_delay,MGM_W290);
   and MGM_G357(MGM_W292,si_delay,MGM_W291);
   and MGM_G358(ENABLE_clkb_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W292);
   not MGM_G359(MGM_W293,d_delay);
   and MGM_G360(MGM_W294,psb_delay,MGM_W293);
   and MGM_G361(MGM_W295,rb_delay,MGM_W294);
   not MGM_G362(MGM_W296,ssb_delay);
   and MGM_G363(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W296,MGM_W295);
   and MGM_G364(MGM_W297,psb_delay,d_delay);
   and MGM_G365(MGM_W298,rb_delay,MGM_W297);
   not MGM_G366(MGM_W299,ssb_delay);
   and MGM_G367(ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W299,MGM_W298);
   not MGM_G368(MGM_W300,d_delay);
   and MGM_G369(MGM_W301,psb_delay,MGM_W300);
   and MGM_G370(MGM_W302,rb_delay,MGM_W301);
   and MGM_G371(ENABLE_NOT_d_AND_psb_AND_rb_AND_si,si_delay,MGM_W302);
   and MGM_G372(MGM_W303,psb_delay,d_delay);
   and MGM_G373(MGM_W304,rb_delay,MGM_W303);
   not MGM_G374(MGM_W305,si_delay);
   and MGM_G375(ENABLE_d_AND_psb_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy08fah1n08x5( clkb, d, o, psb, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, psb, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy08fah_func b15fqy08fah1n08x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy08fah_func b15fqy08fah1n08x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy08fah_func b15fqy08fah1n08x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy08fah_func b15fqy08fah1n08x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(MGM_W2,rb_delay,MGM_W1);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   and MGM_G8(MGM_W7,psb_delay,MGM_W6);
   and MGM_G9(MGM_W8,rb_delay,MGM_W7);
   not MGM_G10(MGM_W9,si_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G12(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W10);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,psb_delay,MGM_W11);
   and MGM_G15(MGM_W13,rb_delay,MGM_W12);
   and MGM_G16(MGM_W14,si_delay,MGM_W13);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,psb_delay,MGM_W16);
   and MGM_G21(MGM_W18,rb_delay,MGM_W17);
   and MGM_G22(MGM_W19,si_delay,MGM_W18);
   and MGM_G23(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W19);
   and MGM_G24(MGM_W20,psb_delay,d_delay);
   and MGM_G25(MGM_W21,rb_delay,MGM_W20);
   not MGM_G26(MGM_W22,si_delay);
   and MGM_G27(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G28(MGM_W24,ssb_delay);
   and MGM_G29(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W24,MGM_W23);
   and MGM_G30(MGM_W25,psb_delay,d_delay);
   and MGM_G31(MGM_W26,rb_delay,MGM_W25);
   not MGM_G32(MGM_W27,si_delay);
   and MGM_G33(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G34(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W28);
   and MGM_G35(MGM_W29,psb_delay,d_delay);
   and MGM_G36(MGM_W30,rb_delay,MGM_W29);
   and MGM_G37(MGM_W31,si_delay,MGM_W30);
   not MGM_G38(MGM_W32,ssb_delay);
   and MGM_G39(ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W32,MGM_W31);
   and MGM_G40(MGM_W33,psb_delay,d_delay);
   and MGM_G41(MGM_W34,rb_delay,MGM_W33);
   and MGM_G42(MGM_W35,si_delay,MGM_W34);
   and MGM_G43(ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G44(MGM_W36,rb_delay,psb_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   and MGM_G47(ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W38);
   and MGM_G48(MGM_W39,rb_delay,psb_delay);
   and MGM_G49(MGM_W40,si_delay,MGM_W39);
   and MGM_G50(ENABLE_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G51(MGM_W41,d_delay);
   and MGM_G52(MGM_W42,rb_delay,MGM_W41);
   not MGM_G53(MGM_W43,si_delay);
   and MGM_G54(MGM_W44,MGM_W43,MGM_W42);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   not MGM_G57(MGM_W46,d_delay);
   and MGM_G58(MGM_W47,rb_delay,MGM_W46);
   not MGM_G59(MGM_W48,si_delay);
   and MGM_G60(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G61(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G62(MGM_W50,d_delay);
   and MGM_G63(MGM_W51,rb_delay,MGM_W50);
   and MGM_G64(MGM_W52,si_delay,MGM_W51);
   and MGM_G65(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G66(MGM_W53,rb_delay,d_delay);
   not MGM_G67(MGM_W54,si_delay);
   and MGM_G68(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G69(MGM_W56,ssb_delay);
   and MGM_G70(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   not MGM_G71(MGM_W57,clkb_delay);
   not MGM_G72(MGM_W58,d_delay);
   and MGM_G73(MGM_W59,MGM_W58,MGM_W57);
   and MGM_G74(MGM_W60,rb_delay,MGM_W59);
   not MGM_G75(MGM_W61,si_delay);
   and MGM_G76(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G77(MGM_W63,ssb_delay);
   and MGM_G78(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G79(MGM_W64,clkb_delay);
   not MGM_G80(MGM_W65,d_delay);
   and MGM_G81(MGM_W66,MGM_W65,MGM_W64);
   and MGM_G82(MGM_W67,rb_delay,MGM_W66);
   not MGM_G83(MGM_W68,si_delay);
   and MGM_G84(MGM_W69,MGM_W68,MGM_W67);
   and MGM_G85(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W69);
   not MGM_G86(MGM_W70,clkb_delay);
   not MGM_G87(MGM_W71,d_delay);
   and MGM_G88(MGM_W72,MGM_W71,MGM_W70);
   and MGM_G89(MGM_W73,rb_delay,MGM_W72);
   and MGM_G90(MGM_W74,si_delay,MGM_W73);
   not MGM_G91(MGM_W75,ssb_delay);
   and MGM_G92(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G93(MGM_W76,clkb_delay);
   not MGM_G94(MGM_W77,d_delay);
   and MGM_G95(MGM_W78,MGM_W77,MGM_W76);
   and MGM_G96(MGM_W79,rb_delay,MGM_W78);
   and MGM_G97(MGM_W80,si_delay,MGM_W79);
   and MGM_G98(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W80);
   not MGM_G99(MGM_W81,clkb_delay);
   and MGM_G100(MGM_W82,d_delay,MGM_W81);
   and MGM_G101(MGM_W83,rb_delay,MGM_W82);
   not MGM_G102(MGM_W84,si_delay);
   and MGM_G103(MGM_W85,MGM_W84,MGM_W83);
   not MGM_G104(MGM_W86,ssb_delay);
   and MGM_G105(ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W86,MGM_W85);
   not MGM_G106(MGM_W87,clkb_delay);
   and MGM_G107(MGM_W88,d_delay,MGM_W87);
   and MGM_G108(MGM_W89,rb_delay,MGM_W88);
   not MGM_G109(MGM_W90,si_delay);
   and MGM_G110(MGM_W91,MGM_W90,MGM_W89);
   and MGM_G111(ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W91);
   not MGM_G112(MGM_W92,clkb_delay);
   and MGM_G113(MGM_W93,d_delay,MGM_W92);
   and MGM_G114(MGM_W94,rb_delay,MGM_W93);
   and MGM_G115(MGM_W95,si_delay,MGM_W94);
   not MGM_G116(MGM_W96,ssb_delay);
   and MGM_G117(ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W96,MGM_W95);
   not MGM_G118(MGM_W97,clkb_delay);
   and MGM_G119(MGM_W98,d_delay,MGM_W97);
   and MGM_G120(MGM_W99,rb_delay,MGM_W98);
   and MGM_G121(MGM_W100,si_delay,MGM_W99);
   and MGM_G122(ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W100);
   not MGM_G123(MGM_W101,d_delay);
   and MGM_G124(MGM_W102,MGM_W101,clkb_delay);
   and MGM_G125(MGM_W103,rb_delay,MGM_W102);
   not MGM_G126(MGM_W104,si_delay);
   and MGM_G127(MGM_W105,MGM_W104,MGM_W103);
   not MGM_G128(MGM_W106,ssb_delay);
   and MGM_G129(ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W106,MGM_W105);
   not MGM_G130(MGM_W107,d_delay);
   and MGM_G131(MGM_W108,MGM_W107,clkb_delay);
   and MGM_G132(MGM_W109,rb_delay,MGM_W108);
   not MGM_G133(MGM_W110,si_delay);
   and MGM_G134(MGM_W111,MGM_W110,MGM_W109);
   and MGM_G135(ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W111);
   not MGM_G136(MGM_W112,d_delay);
   and MGM_G137(MGM_W113,MGM_W112,clkb_delay);
   and MGM_G138(MGM_W114,rb_delay,MGM_W113);
   and MGM_G139(MGM_W115,si_delay,MGM_W114);
   not MGM_G140(MGM_W116,ssb_delay);
   and MGM_G141(ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W116,MGM_W115);
   not MGM_G142(MGM_W117,d_delay);
   and MGM_G143(MGM_W118,MGM_W117,clkb_delay);
   and MGM_G144(MGM_W119,rb_delay,MGM_W118);
   and MGM_G145(MGM_W120,si_delay,MGM_W119);
   and MGM_G146(ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W120);
   and MGM_G147(MGM_W121,d_delay,clkb_delay);
   and MGM_G148(MGM_W122,rb_delay,MGM_W121);
   not MGM_G149(MGM_W123,si_delay);
   and MGM_G150(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G151(MGM_W125,ssb_delay);
   and MGM_G152(ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W125,MGM_W124);
   and MGM_G153(MGM_W126,d_delay,clkb_delay);
   and MGM_G154(MGM_W127,rb_delay,MGM_W126);
   not MGM_G155(MGM_W128,si_delay);
   and MGM_G156(MGM_W129,MGM_W128,MGM_W127);
   and MGM_G157(ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W129);
   and MGM_G158(MGM_W130,d_delay,clkb_delay);
   and MGM_G159(MGM_W131,rb_delay,MGM_W130);
   and MGM_G160(MGM_W132,si_delay,MGM_W131);
   not MGM_G161(MGM_W133,ssb_delay);
   and MGM_G162(ENABLE_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W133,MGM_W132);
   and MGM_G163(MGM_W134,d_delay,clkb_delay);
   and MGM_G164(MGM_W135,rb_delay,MGM_W134);
   and MGM_G165(MGM_W136,si_delay,MGM_W135);
   and MGM_G166(ENABLE_clkb_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W136);
   not MGM_G167(MGM_W137,clkb_delay);
   not MGM_G168(MGM_W138,d_delay);
   and MGM_G169(MGM_W139,MGM_W138,MGM_W137);
   not MGM_G170(MGM_W140,si_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   not MGM_G172(MGM_W142,ssb_delay);
   and MGM_G173(ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W142,MGM_W141);
   not MGM_G174(MGM_W143,clkb_delay);
   not MGM_G175(MGM_W144,d_delay);
   and MGM_G176(MGM_W145,MGM_W144,MGM_W143);
   not MGM_G177(MGM_W146,si_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W147);
   not MGM_G180(MGM_W148,clkb_delay);
   not MGM_G181(MGM_W149,d_delay);
   and MGM_G182(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G183(MGM_W151,si_delay,MGM_W150);
   not MGM_G184(MGM_W152,ssb_delay);
   and MGM_G185(ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W153,clkb_delay);
   not MGM_G187(MGM_W154,d_delay);
   and MGM_G188(MGM_W155,MGM_W154,MGM_W153);
   and MGM_G189(MGM_W156,si_delay,MGM_W155);
   and MGM_G190(ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W156);
   not MGM_G191(MGM_W157,clkb_delay);
   and MGM_G192(MGM_W158,d_delay,MGM_W157);
   not MGM_G193(MGM_W159,si_delay);
   and MGM_G194(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G195(MGM_W161,ssb_delay);
   and MGM_G196(ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W161,MGM_W160);
   not MGM_G197(MGM_W162,clkb_delay);
   and MGM_G198(MGM_W163,d_delay,MGM_W162);
   not MGM_G199(MGM_W164,si_delay);
   and MGM_G200(MGM_W165,MGM_W164,MGM_W163);
   and MGM_G201(ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W165);
   not MGM_G202(MGM_W166,clkb_delay);
   and MGM_G203(MGM_W167,d_delay,MGM_W166);
   and MGM_G204(MGM_W168,si_delay,MGM_W167);
   not MGM_G205(MGM_W169,ssb_delay);
   and MGM_G206(ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb,MGM_W169,MGM_W168);
   not MGM_G207(MGM_W170,clkb_delay);
   and MGM_G208(MGM_W171,d_delay,MGM_W170);
   and MGM_G209(MGM_W172,si_delay,MGM_W171);
   and MGM_G210(ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W172);
   not MGM_G211(MGM_W173,d_delay);
   and MGM_G212(MGM_W174,MGM_W173,clkb_delay);
   not MGM_G213(MGM_W175,si_delay);
   and MGM_G214(MGM_W176,MGM_W175,MGM_W174);
   not MGM_G215(MGM_W177,ssb_delay);
   and MGM_G216(ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W177,MGM_W176);
   not MGM_G217(MGM_W178,d_delay);
   and MGM_G218(MGM_W179,MGM_W178,clkb_delay);
   not MGM_G219(MGM_W180,si_delay);
   and MGM_G220(MGM_W181,MGM_W180,MGM_W179);
   and MGM_G221(ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W181);
   not MGM_G222(MGM_W182,d_delay);
   and MGM_G223(MGM_W183,MGM_W182,clkb_delay);
   and MGM_G224(MGM_W184,si_delay,MGM_W183);
   not MGM_G225(MGM_W185,ssb_delay);
   and MGM_G226(ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W185,MGM_W184);
   not MGM_G227(MGM_W186,d_delay);
   and MGM_G228(MGM_W187,MGM_W186,clkb_delay);
   and MGM_G229(MGM_W188,si_delay,MGM_W187);
   and MGM_G230(ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W188);
   and MGM_G231(MGM_W189,d_delay,clkb_delay);
   not MGM_G232(MGM_W190,si_delay);
   and MGM_G233(MGM_W191,MGM_W190,MGM_W189);
   not MGM_G234(MGM_W192,ssb_delay);
   and MGM_G235(ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W192,MGM_W191);
   and MGM_G236(MGM_W193,d_delay,clkb_delay);
   not MGM_G237(MGM_W194,si_delay);
   and MGM_G238(MGM_W195,MGM_W194,MGM_W193);
   and MGM_G239(ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W195);
   and MGM_G240(MGM_W196,d_delay,clkb_delay);
   and MGM_G241(MGM_W197,si_delay,MGM_W196);
   not MGM_G242(MGM_W198,ssb_delay);
   and MGM_G243(ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb,MGM_W198,MGM_W197);
   and MGM_G244(MGM_W199,d_delay,clkb_delay);
   and MGM_G245(MGM_W200,si_delay,MGM_W199);
   and MGM_G246(ENABLE_clkb_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W200);
   not MGM_G247(MGM_W201,d_delay);
   and MGM_G248(MGM_W202,psb_delay,MGM_W201);
   and MGM_G249(MGM_W203,si_delay,MGM_W202);
   not MGM_G250(MGM_W204,ssb_delay);
   and MGM_G251(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W204,MGM_W203);
   and MGM_G252(MGM_W205,psb_delay,d_delay);
   not MGM_G253(MGM_W206,si_delay);
   and MGM_G254(MGM_W207,MGM_W206,MGM_W205);
   and MGM_G255(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W207);
   and MGM_G256(MGM_W208,psb_delay,d_delay);
   and MGM_G257(MGM_W209,si_delay,MGM_W208);
   not MGM_G258(MGM_W210,ssb_delay);
   and MGM_G259(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W210,MGM_W209);
   and MGM_G260(MGM_W211,psb_delay,d_delay);
   and MGM_G261(MGM_W212,si_delay,MGM_W211);
   and MGM_G262(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W212);
   not MGM_G263(MGM_W213,clkb_delay);
   not MGM_G264(MGM_W214,d_delay);
   and MGM_G265(MGM_W215,MGM_W214,MGM_W213);
   and MGM_G266(MGM_W216,psb_delay,MGM_W215);
   not MGM_G267(MGM_W217,si_delay);
   and MGM_G268(MGM_W218,MGM_W217,MGM_W216);
   not MGM_G269(MGM_W219,ssb_delay);
   and MGM_G270(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W219,MGM_W218);
   not MGM_G271(MGM_W220,clkb_delay);
   not MGM_G272(MGM_W221,d_delay);
   and MGM_G273(MGM_W222,MGM_W221,MGM_W220);
   and MGM_G274(MGM_W223,psb_delay,MGM_W222);
   not MGM_G275(MGM_W224,si_delay);
   and MGM_G276(MGM_W225,MGM_W224,MGM_W223);
   and MGM_G277(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W225);
   not MGM_G278(MGM_W226,clkb_delay);
   not MGM_G279(MGM_W227,d_delay);
   and MGM_G280(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G281(MGM_W229,psb_delay,MGM_W228);
   and MGM_G282(MGM_W230,si_delay,MGM_W229);
   not MGM_G283(MGM_W231,ssb_delay);
   and MGM_G284(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W231,MGM_W230);
   not MGM_G285(MGM_W232,clkb_delay);
   not MGM_G286(MGM_W233,d_delay);
   and MGM_G287(MGM_W234,MGM_W233,MGM_W232);
   and MGM_G288(MGM_W235,psb_delay,MGM_W234);
   and MGM_G289(MGM_W236,si_delay,MGM_W235);
   and MGM_G290(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W236);
   not MGM_G291(MGM_W237,clkb_delay);
   and MGM_G292(MGM_W238,d_delay,MGM_W237);
   and MGM_G293(MGM_W239,psb_delay,MGM_W238);
   not MGM_G294(MGM_W240,si_delay);
   and MGM_G295(MGM_W241,MGM_W240,MGM_W239);
   not MGM_G296(MGM_W242,ssb_delay);
   and MGM_G297(ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W242,MGM_W241);
   not MGM_G298(MGM_W243,clkb_delay);
   and MGM_G299(MGM_W244,d_delay,MGM_W243);
   and MGM_G300(MGM_W245,psb_delay,MGM_W244);
   not MGM_G301(MGM_W246,si_delay);
   and MGM_G302(MGM_W247,MGM_W246,MGM_W245);
   and MGM_G303(ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W247);
   not MGM_G304(MGM_W248,clkb_delay);
   and MGM_G305(MGM_W249,d_delay,MGM_W248);
   and MGM_G306(MGM_W250,psb_delay,MGM_W249);
   and MGM_G307(MGM_W251,si_delay,MGM_W250);
   not MGM_G308(MGM_W252,ssb_delay);
   and MGM_G309(ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W252,MGM_W251);
   not MGM_G310(MGM_W253,clkb_delay);
   and MGM_G311(MGM_W254,d_delay,MGM_W253);
   and MGM_G312(MGM_W255,psb_delay,MGM_W254);
   and MGM_G313(MGM_W256,si_delay,MGM_W255);
   and MGM_G314(ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W256);
   not MGM_G315(MGM_W257,d_delay);
   and MGM_G316(MGM_W258,MGM_W257,clkb_delay);
   and MGM_G317(MGM_W259,psb_delay,MGM_W258);
   not MGM_G318(MGM_W260,si_delay);
   and MGM_G319(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G320(MGM_W262,ssb_delay);
   and MGM_G321(ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   not MGM_G322(MGM_W263,d_delay);
   and MGM_G323(MGM_W264,MGM_W263,clkb_delay);
   and MGM_G324(MGM_W265,psb_delay,MGM_W264);
   not MGM_G325(MGM_W266,si_delay);
   and MGM_G326(MGM_W267,MGM_W266,MGM_W265);
   and MGM_G327(ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W267);
   not MGM_G328(MGM_W268,d_delay);
   and MGM_G329(MGM_W269,MGM_W268,clkb_delay);
   and MGM_G330(MGM_W270,psb_delay,MGM_W269);
   and MGM_G331(MGM_W271,si_delay,MGM_W270);
   not MGM_G332(MGM_W272,ssb_delay);
   and MGM_G333(ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W272,MGM_W271);
   not MGM_G334(MGM_W273,d_delay);
   and MGM_G335(MGM_W274,MGM_W273,clkb_delay);
   and MGM_G336(MGM_W275,psb_delay,MGM_W274);
   and MGM_G337(MGM_W276,si_delay,MGM_W275);
   and MGM_G338(ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W276);
   and MGM_G339(MGM_W277,d_delay,clkb_delay);
   and MGM_G340(MGM_W278,psb_delay,MGM_W277);
   not MGM_G341(MGM_W279,si_delay);
   and MGM_G342(MGM_W280,MGM_W279,MGM_W278);
   not MGM_G343(MGM_W281,ssb_delay);
   and MGM_G344(ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W281,MGM_W280);
   and MGM_G345(MGM_W282,d_delay,clkb_delay);
   and MGM_G346(MGM_W283,psb_delay,MGM_W282);
   not MGM_G347(MGM_W284,si_delay);
   and MGM_G348(MGM_W285,MGM_W284,MGM_W283);
   and MGM_G349(ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W285);
   and MGM_G350(MGM_W286,d_delay,clkb_delay);
   and MGM_G351(MGM_W287,psb_delay,MGM_W286);
   and MGM_G352(MGM_W288,si_delay,MGM_W287);
   not MGM_G353(MGM_W289,ssb_delay);
   and MGM_G354(ENABLE_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W289,MGM_W288);
   and MGM_G355(MGM_W290,d_delay,clkb_delay);
   and MGM_G356(MGM_W291,psb_delay,MGM_W290);
   and MGM_G357(MGM_W292,si_delay,MGM_W291);
   and MGM_G358(ENABLE_clkb_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W292);
   not MGM_G359(MGM_W293,d_delay);
   and MGM_G360(MGM_W294,psb_delay,MGM_W293);
   and MGM_G361(MGM_W295,rb_delay,MGM_W294);
   not MGM_G362(MGM_W296,ssb_delay);
   and MGM_G363(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W296,MGM_W295);
   and MGM_G364(MGM_W297,psb_delay,d_delay);
   and MGM_G365(MGM_W298,rb_delay,MGM_W297);
   not MGM_G366(MGM_W299,ssb_delay);
   and MGM_G367(ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W299,MGM_W298);
   not MGM_G368(MGM_W300,d_delay);
   and MGM_G369(MGM_W301,psb_delay,MGM_W300);
   and MGM_G370(MGM_W302,rb_delay,MGM_W301);
   and MGM_G371(ENABLE_NOT_d_AND_psb_AND_rb_AND_si,si_delay,MGM_W302);
   and MGM_G372(MGM_W303,psb_delay,d_delay);
   and MGM_G373(MGM_W304,rb_delay,MGM_W303);
   not MGM_G374(MGM_W305,si_delay);
   and MGM_G375(ENABLE_d_AND_psb_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy08fah1n16x5( clkb, d, o, psb, rb, si, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, psb, rb, si, ssb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy08fah_func b15fqy08fah1n16x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy08fah_func b15fqy08fah1n16x5_behav_inst(.clkb(clkb),.d(d),.o(o),.psb(psb),.rb(rb),.si(si),.ssb(ssb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   wire si_delay ;
   wire ssb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy08fah_func b15fqy08fah1n16x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy08fah_func b15fqy08fah1n16x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.si(si_delay),.ssb(ssb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(MGM_W2,rb_delay,MGM_W1);
   not MGM_G3(MGM_W3,si_delay);
   and MGM_G4(MGM_W4,MGM_W3,MGM_W2);
   not MGM_G5(MGM_W5,ssb_delay);
   and MGM_G6(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W5,MGM_W4);
   not MGM_G7(MGM_W6,d_delay);
   and MGM_G8(MGM_W7,psb_delay,MGM_W6);
   and MGM_G9(MGM_W8,rb_delay,MGM_W7);
   not MGM_G10(MGM_W9,si_delay);
   and MGM_G11(MGM_W10,MGM_W9,MGM_W8);
   and MGM_G12(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W10);
   not MGM_G13(MGM_W11,d_delay);
   and MGM_G14(MGM_W12,psb_delay,MGM_W11);
   and MGM_G15(MGM_W13,rb_delay,MGM_W12);
   and MGM_G16(MGM_W14,si_delay,MGM_W13);
   not MGM_G17(MGM_W15,ssb_delay);
   and MGM_G18(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W15,MGM_W14);
   not MGM_G19(MGM_W16,d_delay);
   and MGM_G20(MGM_W17,psb_delay,MGM_W16);
   and MGM_G21(MGM_W18,rb_delay,MGM_W17);
   and MGM_G22(MGM_W19,si_delay,MGM_W18);
   and MGM_G23(ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W19);
   and MGM_G24(MGM_W20,psb_delay,d_delay);
   and MGM_G25(MGM_W21,rb_delay,MGM_W20);
   not MGM_G26(MGM_W22,si_delay);
   and MGM_G27(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G28(MGM_W24,ssb_delay);
   and MGM_G29(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W24,MGM_W23);
   and MGM_G30(MGM_W25,psb_delay,d_delay);
   and MGM_G31(MGM_W26,rb_delay,MGM_W25);
   not MGM_G32(MGM_W27,si_delay);
   and MGM_G33(MGM_W28,MGM_W27,MGM_W26);
   and MGM_G34(ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W28);
   and MGM_G35(MGM_W29,psb_delay,d_delay);
   and MGM_G36(MGM_W30,rb_delay,MGM_W29);
   and MGM_G37(MGM_W31,si_delay,MGM_W30);
   not MGM_G38(MGM_W32,ssb_delay);
   and MGM_G39(ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb,MGM_W32,MGM_W31);
   and MGM_G40(MGM_W33,psb_delay,d_delay);
   and MGM_G41(MGM_W34,rb_delay,MGM_W33);
   and MGM_G42(MGM_W35,si_delay,MGM_W34);
   and MGM_G43(ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W35);
   and MGM_G44(MGM_W36,rb_delay,psb_delay);
   not MGM_G45(MGM_W37,si_delay);
   and MGM_G46(MGM_W38,MGM_W37,MGM_W36);
   and MGM_G47(ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W38);
   and MGM_G48(MGM_W39,rb_delay,psb_delay);
   and MGM_G49(MGM_W40,si_delay,MGM_W39);
   and MGM_G50(ENABLE_psb_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W40);
   not MGM_G51(MGM_W41,d_delay);
   and MGM_G52(MGM_W42,rb_delay,MGM_W41);
   not MGM_G53(MGM_W43,si_delay);
   and MGM_G54(MGM_W44,MGM_W43,MGM_W42);
   not MGM_G55(MGM_W45,ssb_delay);
   and MGM_G56(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W45,MGM_W44);
   not MGM_G57(MGM_W46,d_delay);
   and MGM_G58(MGM_W47,rb_delay,MGM_W46);
   not MGM_G59(MGM_W48,si_delay);
   and MGM_G60(MGM_W49,MGM_W48,MGM_W47);
   and MGM_G61(ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W49);
   not MGM_G62(MGM_W50,d_delay);
   and MGM_G63(MGM_W51,rb_delay,MGM_W50);
   and MGM_G64(MGM_W52,si_delay,MGM_W51);
   and MGM_G65(ENABLE_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W52);
   and MGM_G66(MGM_W53,rb_delay,d_delay);
   not MGM_G67(MGM_W54,si_delay);
   and MGM_G68(MGM_W55,MGM_W54,MGM_W53);
   not MGM_G69(MGM_W56,ssb_delay);
   and MGM_G70(ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W56,MGM_W55);
   not MGM_G71(MGM_W57,clkb_delay);
   not MGM_G72(MGM_W58,d_delay);
   and MGM_G73(MGM_W59,MGM_W58,MGM_W57);
   and MGM_G74(MGM_W60,rb_delay,MGM_W59);
   not MGM_G75(MGM_W61,si_delay);
   and MGM_G76(MGM_W62,MGM_W61,MGM_W60);
   not MGM_G77(MGM_W63,ssb_delay);
   and MGM_G78(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W63,MGM_W62);
   not MGM_G79(MGM_W64,clkb_delay);
   not MGM_G80(MGM_W65,d_delay);
   and MGM_G81(MGM_W66,MGM_W65,MGM_W64);
   and MGM_G82(MGM_W67,rb_delay,MGM_W66);
   not MGM_G83(MGM_W68,si_delay);
   and MGM_G84(MGM_W69,MGM_W68,MGM_W67);
   and MGM_G85(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W69);
   not MGM_G86(MGM_W70,clkb_delay);
   not MGM_G87(MGM_W71,d_delay);
   and MGM_G88(MGM_W72,MGM_W71,MGM_W70);
   and MGM_G89(MGM_W73,rb_delay,MGM_W72);
   and MGM_G90(MGM_W74,si_delay,MGM_W73);
   not MGM_G91(MGM_W75,ssb_delay);
   and MGM_G92(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W75,MGM_W74);
   not MGM_G93(MGM_W76,clkb_delay);
   not MGM_G94(MGM_W77,d_delay);
   and MGM_G95(MGM_W78,MGM_W77,MGM_W76);
   and MGM_G96(MGM_W79,rb_delay,MGM_W78);
   and MGM_G97(MGM_W80,si_delay,MGM_W79);
   and MGM_G98(ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W80);
   not MGM_G99(MGM_W81,clkb_delay);
   and MGM_G100(MGM_W82,d_delay,MGM_W81);
   and MGM_G101(MGM_W83,rb_delay,MGM_W82);
   not MGM_G102(MGM_W84,si_delay);
   and MGM_G103(MGM_W85,MGM_W84,MGM_W83);
   not MGM_G104(MGM_W86,ssb_delay);
   and MGM_G105(ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W86,MGM_W85);
   not MGM_G106(MGM_W87,clkb_delay);
   and MGM_G107(MGM_W88,d_delay,MGM_W87);
   and MGM_G108(MGM_W89,rb_delay,MGM_W88);
   not MGM_G109(MGM_W90,si_delay);
   and MGM_G110(MGM_W91,MGM_W90,MGM_W89);
   and MGM_G111(ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W91);
   not MGM_G112(MGM_W92,clkb_delay);
   and MGM_G113(MGM_W93,d_delay,MGM_W92);
   and MGM_G114(MGM_W94,rb_delay,MGM_W93);
   and MGM_G115(MGM_W95,si_delay,MGM_W94);
   not MGM_G116(MGM_W96,ssb_delay);
   and MGM_G117(ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W96,MGM_W95);
   not MGM_G118(MGM_W97,clkb_delay);
   and MGM_G119(MGM_W98,d_delay,MGM_W97);
   and MGM_G120(MGM_W99,rb_delay,MGM_W98);
   and MGM_G121(MGM_W100,si_delay,MGM_W99);
   and MGM_G122(ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W100);
   not MGM_G123(MGM_W101,d_delay);
   and MGM_G124(MGM_W102,MGM_W101,clkb_delay);
   and MGM_G125(MGM_W103,rb_delay,MGM_W102);
   not MGM_G126(MGM_W104,si_delay);
   and MGM_G127(MGM_W105,MGM_W104,MGM_W103);
   not MGM_G128(MGM_W106,ssb_delay);
   and MGM_G129(ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W106,MGM_W105);
   not MGM_G130(MGM_W107,d_delay);
   and MGM_G131(MGM_W108,MGM_W107,clkb_delay);
   and MGM_G132(MGM_W109,rb_delay,MGM_W108);
   not MGM_G133(MGM_W110,si_delay);
   and MGM_G134(MGM_W111,MGM_W110,MGM_W109);
   and MGM_G135(ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W111);
   not MGM_G136(MGM_W112,d_delay);
   and MGM_G137(MGM_W113,MGM_W112,clkb_delay);
   and MGM_G138(MGM_W114,rb_delay,MGM_W113);
   and MGM_G139(MGM_W115,si_delay,MGM_W114);
   not MGM_G140(MGM_W116,ssb_delay);
   and MGM_G141(ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W116,MGM_W115);
   not MGM_G142(MGM_W117,d_delay);
   and MGM_G143(MGM_W118,MGM_W117,clkb_delay);
   and MGM_G144(MGM_W119,rb_delay,MGM_W118);
   and MGM_G145(MGM_W120,si_delay,MGM_W119);
   and MGM_G146(ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W120);
   and MGM_G147(MGM_W121,d_delay,clkb_delay);
   and MGM_G148(MGM_W122,rb_delay,MGM_W121);
   not MGM_G149(MGM_W123,si_delay);
   and MGM_G150(MGM_W124,MGM_W123,MGM_W122);
   not MGM_G151(MGM_W125,ssb_delay);
   and MGM_G152(ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb,MGM_W125,MGM_W124);
   and MGM_G153(MGM_W126,d_delay,clkb_delay);
   and MGM_G154(MGM_W127,rb_delay,MGM_W126);
   not MGM_G155(MGM_W128,si_delay);
   and MGM_G156(MGM_W129,MGM_W128,MGM_W127);
   and MGM_G157(ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W129);
   and MGM_G158(MGM_W130,d_delay,clkb_delay);
   and MGM_G159(MGM_W131,rb_delay,MGM_W130);
   and MGM_G160(MGM_W132,si_delay,MGM_W131);
   not MGM_G161(MGM_W133,ssb_delay);
   and MGM_G162(ENABLE_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb,MGM_W133,MGM_W132);
   and MGM_G163(MGM_W134,d_delay,clkb_delay);
   and MGM_G164(MGM_W135,rb_delay,MGM_W134);
   and MGM_G165(MGM_W136,si_delay,MGM_W135);
   and MGM_G166(ENABLE_clkb_AND_d_AND_rb_AND_si_AND_ssb,ssb_delay,MGM_W136);
   not MGM_G167(MGM_W137,clkb_delay);
   not MGM_G168(MGM_W138,d_delay);
   and MGM_G169(MGM_W139,MGM_W138,MGM_W137);
   not MGM_G170(MGM_W140,si_delay);
   and MGM_G171(MGM_W141,MGM_W140,MGM_W139);
   not MGM_G172(MGM_W142,ssb_delay);
   and MGM_G173(ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W142,MGM_W141);
   not MGM_G174(MGM_W143,clkb_delay);
   not MGM_G175(MGM_W144,d_delay);
   and MGM_G176(MGM_W145,MGM_W144,MGM_W143);
   not MGM_G177(MGM_W146,si_delay);
   and MGM_G178(MGM_W147,MGM_W146,MGM_W145);
   and MGM_G179(ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W147);
   not MGM_G180(MGM_W148,clkb_delay);
   not MGM_G181(MGM_W149,d_delay);
   and MGM_G182(MGM_W150,MGM_W149,MGM_W148);
   and MGM_G183(MGM_W151,si_delay,MGM_W150);
   not MGM_G184(MGM_W152,ssb_delay);
   and MGM_G185(ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W152,MGM_W151);
   not MGM_G186(MGM_W153,clkb_delay);
   not MGM_G187(MGM_W154,d_delay);
   and MGM_G188(MGM_W155,MGM_W154,MGM_W153);
   and MGM_G189(MGM_W156,si_delay,MGM_W155);
   and MGM_G190(ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W156);
   not MGM_G191(MGM_W157,clkb_delay);
   and MGM_G192(MGM_W158,d_delay,MGM_W157);
   not MGM_G193(MGM_W159,si_delay);
   and MGM_G194(MGM_W160,MGM_W159,MGM_W158);
   not MGM_G195(MGM_W161,ssb_delay);
   and MGM_G196(ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W161,MGM_W160);
   not MGM_G197(MGM_W162,clkb_delay);
   and MGM_G198(MGM_W163,d_delay,MGM_W162);
   not MGM_G199(MGM_W164,si_delay);
   and MGM_G200(MGM_W165,MGM_W164,MGM_W163);
   and MGM_G201(ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W165);
   not MGM_G202(MGM_W166,clkb_delay);
   and MGM_G203(MGM_W167,d_delay,MGM_W166);
   and MGM_G204(MGM_W168,si_delay,MGM_W167);
   not MGM_G205(MGM_W169,ssb_delay);
   and MGM_G206(ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb,MGM_W169,MGM_W168);
   not MGM_G207(MGM_W170,clkb_delay);
   and MGM_G208(MGM_W171,d_delay,MGM_W170);
   and MGM_G209(MGM_W172,si_delay,MGM_W171);
   and MGM_G210(ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W172);
   not MGM_G211(MGM_W173,d_delay);
   and MGM_G212(MGM_W174,MGM_W173,clkb_delay);
   not MGM_G213(MGM_W175,si_delay);
   and MGM_G214(MGM_W176,MGM_W175,MGM_W174);
   not MGM_G215(MGM_W177,ssb_delay);
   and MGM_G216(ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb,MGM_W177,MGM_W176);
   not MGM_G217(MGM_W178,d_delay);
   and MGM_G218(MGM_W179,MGM_W178,clkb_delay);
   not MGM_G219(MGM_W180,si_delay);
   and MGM_G220(MGM_W181,MGM_W180,MGM_W179);
   and MGM_G221(ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W181);
   not MGM_G222(MGM_W182,d_delay);
   and MGM_G223(MGM_W183,MGM_W182,clkb_delay);
   and MGM_G224(MGM_W184,si_delay,MGM_W183);
   not MGM_G225(MGM_W185,ssb_delay);
   and MGM_G226(ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb,MGM_W185,MGM_W184);
   not MGM_G227(MGM_W186,d_delay);
   and MGM_G228(MGM_W187,MGM_W186,clkb_delay);
   and MGM_G229(MGM_W188,si_delay,MGM_W187);
   and MGM_G230(ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb,ssb_delay,MGM_W188);
   and MGM_G231(MGM_W189,d_delay,clkb_delay);
   not MGM_G232(MGM_W190,si_delay);
   and MGM_G233(MGM_W191,MGM_W190,MGM_W189);
   not MGM_G234(MGM_W192,ssb_delay);
   and MGM_G235(ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb,MGM_W192,MGM_W191);
   and MGM_G236(MGM_W193,d_delay,clkb_delay);
   not MGM_G237(MGM_W194,si_delay);
   and MGM_G238(MGM_W195,MGM_W194,MGM_W193);
   and MGM_G239(ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb,ssb_delay,MGM_W195);
   and MGM_G240(MGM_W196,d_delay,clkb_delay);
   and MGM_G241(MGM_W197,si_delay,MGM_W196);
   not MGM_G242(MGM_W198,ssb_delay);
   and MGM_G243(ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb,MGM_W198,MGM_W197);
   and MGM_G244(MGM_W199,d_delay,clkb_delay);
   and MGM_G245(MGM_W200,si_delay,MGM_W199);
   and MGM_G246(ENABLE_clkb_AND_d_AND_si_AND_ssb,ssb_delay,MGM_W200);
   not MGM_G247(MGM_W201,d_delay);
   and MGM_G248(MGM_W202,psb_delay,MGM_W201);
   and MGM_G249(MGM_W203,si_delay,MGM_W202);
   not MGM_G250(MGM_W204,ssb_delay);
   and MGM_G251(ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W204,MGM_W203);
   and MGM_G252(MGM_W205,psb_delay,d_delay);
   not MGM_G253(MGM_W206,si_delay);
   and MGM_G254(MGM_W207,MGM_W206,MGM_W205);
   and MGM_G255(ENABLE_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W207);
   and MGM_G256(MGM_W208,psb_delay,d_delay);
   and MGM_G257(MGM_W209,si_delay,MGM_W208);
   not MGM_G258(MGM_W210,ssb_delay);
   and MGM_G259(ENABLE_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W210,MGM_W209);
   and MGM_G260(MGM_W211,psb_delay,d_delay);
   and MGM_G261(MGM_W212,si_delay,MGM_W211);
   and MGM_G262(ENABLE_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W212);
   not MGM_G263(MGM_W213,clkb_delay);
   not MGM_G264(MGM_W214,d_delay);
   and MGM_G265(MGM_W215,MGM_W214,MGM_W213);
   and MGM_G266(MGM_W216,psb_delay,MGM_W215);
   not MGM_G267(MGM_W217,si_delay);
   and MGM_G268(MGM_W218,MGM_W217,MGM_W216);
   not MGM_G269(MGM_W219,ssb_delay);
   and MGM_G270(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W219,MGM_W218);
   not MGM_G271(MGM_W220,clkb_delay);
   not MGM_G272(MGM_W221,d_delay);
   and MGM_G273(MGM_W222,MGM_W221,MGM_W220);
   and MGM_G274(MGM_W223,psb_delay,MGM_W222);
   not MGM_G275(MGM_W224,si_delay);
   and MGM_G276(MGM_W225,MGM_W224,MGM_W223);
   and MGM_G277(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W225);
   not MGM_G278(MGM_W226,clkb_delay);
   not MGM_G279(MGM_W227,d_delay);
   and MGM_G280(MGM_W228,MGM_W227,MGM_W226);
   and MGM_G281(MGM_W229,psb_delay,MGM_W228);
   and MGM_G282(MGM_W230,si_delay,MGM_W229);
   not MGM_G283(MGM_W231,ssb_delay);
   and MGM_G284(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W231,MGM_W230);
   not MGM_G285(MGM_W232,clkb_delay);
   not MGM_G286(MGM_W233,d_delay);
   and MGM_G287(MGM_W234,MGM_W233,MGM_W232);
   and MGM_G288(MGM_W235,psb_delay,MGM_W234);
   and MGM_G289(MGM_W236,si_delay,MGM_W235);
   and MGM_G290(ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W236);
   not MGM_G291(MGM_W237,clkb_delay);
   and MGM_G292(MGM_W238,d_delay,MGM_W237);
   and MGM_G293(MGM_W239,psb_delay,MGM_W238);
   not MGM_G294(MGM_W240,si_delay);
   and MGM_G295(MGM_W241,MGM_W240,MGM_W239);
   not MGM_G296(MGM_W242,ssb_delay);
   and MGM_G297(ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W242,MGM_W241);
   not MGM_G298(MGM_W243,clkb_delay);
   and MGM_G299(MGM_W244,d_delay,MGM_W243);
   and MGM_G300(MGM_W245,psb_delay,MGM_W244);
   not MGM_G301(MGM_W246,si_delay);
   and MGM_G302(MGM_W247,MGM_W246,MGM_W245);
   and MGM_G303(ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W247);
   not MGM_G304(MGM_W248,clkb_delay);
   and MGM_G305(MGM_W249,d_delay,MGM_W248);
   and MGM_G306(MGM_W250,psb_delay,MGM_W249);
   and MGM_G307(MGM_W251,si_delay,MGM_W250);
   not MGM_G308(MGM_W252,ssb_delay);
   and MGM_G309(ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W252,MGM_W251);
   not MGM_G310(MGM_W253,clkb_delay);
   and MGM_G311(MGM_W254,d_delay,MGM_W253);
   and MGM_G312(MGM_W255,psb_delay,MGM_W254);
   and MGM_G313(MGM_W256,si_delay,MGM_W255);
   and MGM_G314(ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W256);
   not MGM_G315(MGM_W257,d_delay);
   and MGM_G316(MGM_W258,MGM_W257,clkb_delay);
   and MGM_G317(MGM_W259,psb_delay,MGM_W258);
   not MGM_G318(MGM_W260,si_delay);
   and MGM_G319(MGM_W261,MGM_W260,MGM_W259);
   not MGM_G320(MGM_W262,ssb_delay);
   and MGM_G321(ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W262,MGM_W261);
   not MGM_G322(MGM_W263,d_delay);
   and MGM_G323(MGM_W264,MGM_W263,clkb_delay);
   and MGM_G324(MGM_W265,psb_delay,MGM_W264);
   not MGM_G325(MGM_W266,si_delay);
   and MGM_G326(MGM_W267,MGM_W266,MGM_W265);
   and MGM_G327(ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W267);
   not MGM_G328(MGM_W268,d_delay);
   and MGM_G329(MGM_W269,MGM_W268,clkb_delay);
   and MGM_G330(MGM_W270,psb_delay,MGM_W269);
   and MGM_G331(MGM_W271,si_delay,MGM_W270);
   not MGM_G332(MGM_W272,ssb_delay);
   and MGM_G333(ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W272,MGM_W271);
   not MGM_G334(MGM_W273,d_delay);
   and MGM_G335(MGM_W274,MGM_W273,clkb_delay);
   and MGM_G336(MGM_W275,psb_delay,MGM_W274);
   and MGM_G337(MGM_W276,si_delay,MGM_W275);
   and MGM_G338(ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W276);
   and MGM_G339(MGM_W277,d_delay,clkb_delay);
   and MGM_G340(MGM_W278,psb_delay,MGM_W277);
   not MGM_G341(MGM_W279,si_delay);
   and MGM_G342(MGM_W280,MGM_W279,MGM_W278);
   not MGM_G343(MGM_W281,ssb_delay);
   and MGM_G344(ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb,MGM_W281,MGM_W280);
   and MGM_G345(MGM_W282,d_delay,clkb_delay);
   and MGM_G346(MGM_W283,psb_delay,MGM_W282);
   not MGM_G347(MGM_W284,si_delay);
   and MGM_G348(MGM_W285,MGM_W284,MGM_W283);
   and MGM_G349(ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb,ssb_delay,MGM_W285);
   and MGM_G350(MGM_W286,d_delay,clkb_delay);
   and MGM_G351(MGM_W287,psb_delay,MGM_W286);
   and MGM_G352(MGM_W288,si_delay,MGM_W287);
   not MGM_G353(MGM_W289,ssb_delay);
   and MGM_G354(ENABLE_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb,MGM_W289,MGM_W288);
   and MGM_G355(MGM_W290,d_delay,clkb_delay);
   and MGM_G356(MGM_W291,psb_delay,MGM_W290);
   and MGM_G357(MGM_W292,si_delay,MGM_W291);
   and MGM_G358(ENABLE_clkb_AND_d_AND_psb_AND_si_AND_ssb,ssb_delay,MGM_W292);
   not MGM_G359(MGM_W293,d_delay);
   and MGM_G360(MGM_W294,psb_delay,MGM_W293);
   and MGM_G361(MGM_W295,rb_delay,MGM_W294);
   not MGM_G362(MGM_W296,ssb_delay);
   and MGM_G363(ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W296,MGM_W295);
   and MGM_G364(MGM_W297,psb_delay,d_delay);
   and MGM_G365(MGM_W298,rb_delay,MGM_W297);
   not MGM_G366(MGM_W299,ssb_delay);
   and MGM_G367(ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb,MGM_W299,MGM_W298);
   not MGM_G368(MGM_W300,d_delay);
   and MGM_G369(MGM_W301,psb_delay,MGM_W300);
   and MGM_G370(MGM_W302,rb_delay,MGM_W301);
   and MGM_G371(ENABLE_NOT_d_AND_psb_AND_rb_AND_si,si_delay,MGM_W302);
   and MGM_G372(MGM_W303,psb_delay,d_delay);
   and MGM_G373(MGM_W304,rb_delay,MGM_W303);
   not MGM_G374(MGM_W305,si_delay);
   and MGM_G375(ENABLE_d_AND_psb_AND_rb_AND_NOT_si,MGM_W305,MGM_W304);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && psb==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && rb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b0 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b0 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1 && psb==1'b1 && si==1'b1 && ssb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      // recrem psb-clkb-negedge
      $recrem(posedge psb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clkb_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_clkb_AND_d_AND_rb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // recrem rb-clkb-negedge
      $recrem(posedge rb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      negedge clkb &&& (ENABLE_d_AND_psb_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_NOT_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      posedge rb &&& (ENABLE_clkb_AND_d_AND_si_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clkb_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_NOT_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_si_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d_AND_psb_AND_si_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      negedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold si- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      posedge si &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,si_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d_AND_psb_AND_rb_AND_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      negedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      // setuphold ssb- clkb-HL
      $setuphold(negedge clkb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      posedge ssb &&& (ENABLE_d_AND_psb_AND_rb_AND_NOT_si == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,ssb_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fqy203ah_func( clk, d1, d2, o1, o2, rb, si1, si2, ssb, notifier0, notifier1 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, rb, si1, si2, ssb, notifier0, notifier1;
   output o1, o2;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d2, si2, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier1 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C1, rb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D1, d1, si1, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, MGM_C1, 1'b0, MGM_CLK1, MGM_D1, vcc, vssx, notifier0 );
   INTCseq_cdiar2ah_0( o1, IQ1, vcc, vssx );
   INTCseq_cdiar2ah_0( o2, IQ2, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_fdw003ah_5( MGM_D0, d2, si2, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, notifier1 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk );
   INTCseq_cdiar2ah_1( MGM_C1, rb );
   INTCseq_fdw003ah_5( MGM_D1, d1, si1, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, MGM_C1, 1'b0, MGM_CLK1, MGM_D1, notifier0 );
   INTCseq_cdiar2ah_0( o1, IQ1 );
   INTCseq_cdiar2ah_0( o2, IQ2 );
`endif

endmodule
`endcelldefine



`celldefine
module b15fqy203ah1n02x5( clk, d1, d2, o1, o2, rb, si1, si2, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, rb, si1, si2, ssb;
   output o1, o2;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy203ah_func b15fqy203ah1n02x5_behav_inst(.clk(clk),.rb(rb),.ssb(ssb),.o1(o1),.o2(o2),.d1(d1),.d2(d2),.si1(si1),.si2(si2),.notifier0(1'b0),.notifier1(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy203ah_func b15fqy203ah1n02x5_behav_inst(.clk(clk),.rb(rb),.ssb(ssb),.o1(o1),.o2(o2),.d1(d1),.d2(d2),.si1(si1),.si2(si2),.notifier0(1'b0),.notifier1(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire rb_delay ;
   wire ssb_delay ;
   wire d1_delay ;
   wire d2_delay ;
   wire si1_delay ;
   wire si2_delay ;
   reg notifier;
   reg notifier0;
   reg notifier1;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
     notifier1 = (notifier1 !== notifier) ? notifier : ~notifier1;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy203ah_func b15fqy203ah1n02x5_inst(.clk(clk_delay),.rb(rb_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.d1(d1_delay),.d2(d2_delay),.si1(si1_delay),.si2(si2_delay),.notifier0(notifier0),.notifier1(notifier1),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy203ah_func b15fqy203ah1n02x5_inst(.clk(clk_delay),.rb(rb_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.d1(d1_delay),.d2(d2_delay),.si1(si1_delay),.si2(si2_delay),.notifier0(notifier0),.notifier1(notifier1));
   `endif
   
   // spec_gates_begin
   buf MGM_G0(ENABLE_rb,rb_delay);
   not MGM_G1(MGM_W0,d1_delay);
   not MGM_G2(MGM_W1,d2_delay);
   and MGM_G3(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G4(MGM_W3,si1_delay);
   and MGM_G5(MGM_W4,MGM_W3,MGM_W2);
   and MGM_G6(MGM_W5,si2_delay,MGM_W4);
   not MGM_G7(MGM_W6,ssb_delay);
   and MGM_G8(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W6,MGM_W5);
   not MGM_G9(MGM_W7,d1_delay);
   not MGM_G10(MGM_W8,d2_delay);
   and MGM_G11(MGM_W9,MGM_W8,MGM_W7);
   and MGM_G12(MGM_W10,si1_delay,MGM_W9);
   not MGM_G13(MGM_W11,si2_delay);
   and MGM_G14(MGM_W12,MGM_W11,MGM_W10);
   not MGM_G15(MGM_W13,ssb_delay);
   and MGM_G16(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W13,MGM_W12);
   not MGM_G17(MGM_W14,d1_delay);
   not MGM_G18(MGM_W15,d2_delay);
   and MGM_G19(MGM_W16,MGM_W15,MGM_W14);
   and MGM_G20(MGM_W17,si1_delay,MGM_W16);
   and MGM_G21(MGM_W18,si2_delay,MGM_W17);
   not MGM_G22(MGM_W19,ssb_delay);
   and MGM_G23(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W19,MGM_W18);
   not MGM_G24(MGM_W20,d1_delay);
   and MGM_G25(MGM_W21,d2_delay,MGM_W20);
   not MGM_G26(MGM_W22,si1_delay);
   and MGM_G27(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G28(MGM_W24,si2_delay);
   and MGM_G29(MGM_W25,MGM_W24,MGM_W23);
   and MGM_G30(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W25);
   not MGM_G31(MGM_W26,d1_delay);
   and MGM_G32(MGM_W27,d2_delay,MGM_W26);
   not MGM_G33(MGM_W28,si1_delay);
   and MGM_G34(MGM_W29,MGM_W28,MGM_W27);
   and MGM_G35(MGM_W30,si2_delay,MGM_W29);
   not MGM_G36(MGM_W31,ssb_delay);
   and MGM_G37(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W31,MGM_W30);
   not MGM_G38(MGM_W32,d1_delay);
   and MGM_G39(MGM_W33,d2_delay,MGM_W32);
   not MGM_G40(MGM_W34,si1_delay);
   and MGM_G41(MGM_W35,MGM_W34,MGM_W33);
   and MGM_G42(MGM_W36,si2_delay,MGM_W35);
   and MGM_G43(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W36);
   not MGM_G44(MGM_W37,d1_delay);
   and MGM_G45(MGM_W38,d2_delay,MGM_W37);
   and MGM_G46(MGM_W39,si1_delay,MGM_W38);
   not MGM_G47(MGM_W40,si2_delay);
   and MGM_G48(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G49(MGM_W42,ssb_delay);
   and MGM_G50(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W42,MGM_W41);
   not MGM_G51(MGM_W43,d1_delay);
   and MGM_G52(MGM_W44,d2_delay,MGM_W43);
   and MGM_G53(MGM_W45,si1_delay,MGM_W44);
   not MGM_G54(MGM_W46,si2_delay);
   and MGM_G55(MGM_W47,MGM_W46,MGM_W45);
   and MGM_G56(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W47);
   not MGM_G57(MGM_W48,d1_delay);
   and MGM_G58(MGM_W49,d2_delay,MGM_W48);
   and MGM_G59(MGM_W50,si1_delay,MGM_W49);
   and MGM_G60(MGM_W51,si2_delay,MGM_W50);
   not MGM_G61(MGM_W52,ssb_delay);
   and MGM_G62(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W52,MGM_W51);
   not MGM_G63(MGM_W53,d1_delay);
   and MGM_G64(MGM_W54,d2_delay,MGM_W53);
   and MGM_G65(MGM_W55,si1_delay,MGM_W54);
   and MGM_G66(MGM_W56,si2_delay,MGM_W55);
   and MGM_G67(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W56);
   not MGM_G68(MGM_W57,d2_delay);
   and MGM_G69(MGM_W58,MGM_W57,d1_delay);
   not MGM_G70(MGM_W59,si1_delay);
   and MGM_G71(MGM_W60,MGM_W59,MGM_W58);
   not MGM_G72(MGM_W61,si2_delay);
   and MGM_G73(MGM_W62,MGM_W61,MGM_W60);
   and MGM_G74(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W62);
   not MGM_G75(MGM_W63,d2_delay);
   and MGM_G76(MGM_W64,MGM_W63,d1_delay);
   not MGM_G77(MGM_W65,si1_delay);
   and MGM_G78(MGM_W66,MGM_W65,MGM_W64);
   and MGM_G79(MGM_W67,si2_delay,MGM_W66);
   not MGM_G80(MGM_W68,ssb_delay);
   and MGM_G81(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W68,MGM_W67);
   not MGM_G82(MGM_W69,d2_delay);
   and MGM_G83(MGM_W70,MGM_W69,d1_delay);
   not MGM_G84(MGM_W71,si1_delay);
   and MGM_G85(MGM_W72,MGM_W71,MGM_W70);
   and MGM_G86(MGM_W73,si2_delay,MGM_W72);
   and MGM_G87(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W73);
   not MGM_G88(MGM_W74,d2_delay);
   and MGM_G89(MGM_W75,MGM_W74,d1_delay);
   and MGM_G90(MGM_W76,si1_delay,MGM_W75);
   not MGM_G91(MGM_W77,si2_delay);
   and MGM_G92(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G93(MGM_W79,ssb_delay);
   and MGM_G94(ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G95(MGM_W80,d2_delay);
   and MGM_G96(MGM_W81,MGM_W80,d1_delay);
   and MGM_G97(MGM_W82,si1_delay,MGM_W81);
   not MGM_G98(MGM_W83,si2_delay);
   and MGM_G99(MGM_W84,MGM_W83,MGM_W82);
   and MGM_G100(ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W84);
   not MGM_G101(MGM_W85,d2_delay);
   and MGM_G102(MGM_W86,MGM_W85,d1_delay);
   and MGM_G103(MGM_W87,si1_delay,MGM_W86);
   and MGM_G104(MGM_W88,si2_delay,MGM_W87);
   not MGM_G105(MGM_W89,ssb_delay);
   and MGM_G106(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W89,MGM_W88);
   not MGM_G107(MGM_W90,d2_delay);
   and MGM_G108(MGM_W91,MGM_W90,d1_delay);
   and MGM_G109(MGM_W92,si1_delay,MGM_W91);
   and MGM_G110(MGM_W93,si2_delay,MGM_W92);
   and MGM_G111(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W93);
   and MGM_G112(MGM_W94,d2_delay,d1_delay);
   not MGM_G113(MGM_W95,si1_delay);
   and MGM_G114(MGM_W96,MGM_W95,MGM_W94);
   not MGM_G115(MGM_W97,si2_delay);
   and MGM_G116(MGM_W98,MGM_W97,MGM_W96);
   and MGM_G117(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W98);
   and MGM_G118(MGM_W99,d2_delay,d1_delay);
   not MGM_G119(MGM_W100,si1_delay);
   and MGM_G120(MGM_W101,MGM_W100,MGM_W99);
   and MGM_G121(MGM_W102,si2_delay,MGM_W101);
   not MGM_G122(MGM_W103,ssb_delay);
   and MGM_G123(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W103,MGM_W102);
   and MGM_G124(MGM_W104,d2_delay,d1_delay);
   not MGM_G125(MGM_W105,si1_delay);
   and MGM_G126(MGM_W106,MGM_W105,MGM_W104);
   and MGM_G127(MGM_W107,si2_delay,MGM_W106);
   and MGM_G128(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W107);
   and MGM_G129(MGM_W108,d2_delay,d1_delay);
   and MGM_G130(MGM_W109,si1_delay,MGM_W108);
   not MGM_G131(MGM_W110,si2_delay);
   and MGM_G132(MGM_W111,MGM_W110,MGM_W109);
   not MGM_G133(MGM_W112,ssb_delay);
   and MGM_G134(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W112,MGM_W111);
   and MGM_G135(MGM_W113,d2_delay,d1_delay);
   and MGM_G136(MGM_W114,si1_delay,MGM_W113);
   not MGM_G137(MGM_W115,si2_delay);
   and MGM_G138(MGM_W116,MGM_W115,MGM_W114);
   and MGM_G139(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W116);
   and MGM_G140(MGM_W117,d2_delay,d1_delay);
   and MGM_G141(MGM_W118,si1_delay,MGM_W117);
   and MGM_G142(MGM_W119,si2_delay,MGM_W118);
   not MGM_G143(MGM_W120,ssb_delay);
   and MGM_G144(ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W120,MGM_W119);
   and MGM_G145(MGM_W121,d2_delay,d1_delay);
   and MGM_G146(MGM_W122,si1_delay,MGM_W121);
   and MGM_G147(MGM_W123,si2_delay,MGM_W122);
   and MGM_G148(ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W123);
   not MGM_G149(MGM_W124,clk_delay);
   not MGM_G150(MGM_W125,d1_delay);
   and MGM_G151(MGM_W126,MGM_W125,MGM_W124);
   not MGM_G152(MGM_W127,d2_delay);
   and MGM_G153(MGM_W128,MGM_W127,MGM_W126);
   not MGM_G154(MGM_W129,si1_delay);
   and MGM_G155(MGM_W130,MGM_W129,MGM_W128);
   not MGM_G156(MGM_W131,si2_delay);
   and MGM_G157(MGM_W132,MGM_W131,MGM_W130);
   not MGM_G158(MGM_W133,ssb_delay);
   and MGM_G159(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W133,MGM_W132);
   not MGM_G160(MGM_W134,clk_delay);
   not MGM_G161(MGM_W135,d1_delay);
   and MGM_G162(MGM_W136,MGM_W135,MGM_W134);
   not MGM_G163(MGM_W137,d2_delay);
   and MGM_G164(MGM_W138,MGM_W137,MGM_W136);
   not MGM_G165(MGM_W139,si1_delay);
   and MGM_G166(MGM_W140,MGM_W139,MGM_W138);
   not MGM_G167(MGM_W141,si2_delay);
   and MGM_G168(MGM_W142,MGM_W141,MGM_W140);
   and MGM_G169(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W142);
   not MGM_G170(MGM_W143,clk_delay);
   not MGM_G171(MGM_W144,d1_delay);
   and MGM_G172(MGM_W145,MGM_W144,MGM_W143);
   not MGM_G173(MGM_W146,d2_delay);
   and MGM_G174(MGM_W147,MGM_W146,MGM_W145);
   not MGM_G175(MGM_W148,si1_delay);
   and MGM_G176(MGM_W149,MGM_W148,MGM_W147);
   and MGM_G177(MGM_W150,si2_delay,MGM_W149);
   not MGM_G178(MGM_W151,ssb_delay);
   and MGM_G179(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W151,MGM_W150);
   not MGM_G180(MGM_W152,clk_delay);
   not MGM_G181(MGM_W153,d1_delay);
   and MGM_G182(MGM_W154,MGM_W153,MGM_W152);
   not MGM_G183(MGM_W155,d2_delay);
   and MGM_G184(MGM_W156,MGM_W155,MGM_W154);
   not MGM_G185(MGM_W157,si1_delay);
   and MGM_G186(MGM_W158,MGM_W157,MGM_W156);
   and MGM_G187(MGM_W159,si2_delay,MGM_W158);
   and MGM_G188(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W159);
   not MGM_G189(MGM_W160,clk_delay);
   not MGM_G190(MGM_W161,d1_delay);
   and MGM_G191(MGM_W162,MGM_W161,MGM_W160);
   not MGM_G192(MGM_W163,d2_delay);
   and MGM_G193(MGM_W164,MGM_W163,MGM_W162);
   and MGM_G194(MGM_W165,si1_delay,MGM_W164);
   not MGM_G195(MGM_W166,si2_delay);
   and MGM_G196(MGM_W167,MGM_W166,MGM_W165);
   not MGM_G197(MGM_W168,ssb_delay);
   and MGM_G198(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W168,MGM_W167);
   not MGM_G199(MGM_W169,clk_delay);
   not MGM_G200(MGM_W170,d1_delay);
   and MGM_G201(MGM_W171,MGM_W170,MGM_W169);
   not MGM_G202(MGM_W172,d2_delay);
   and MGM_G203(MGM_W173,MGM_W172,MGM_W171);
   and MGM_G204(MGM_W174,si1_delay,MGM_W173);
   not MGM_G205(MGM_W175,si2_delay);
   and MGM_G206(MGM_W176,MGM_W175,MGM_W174);
   and MGM_G207(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W176);
   not MGM_G208(MGM_W177,clk_delay);
   not MGM_G209(MGM_W178,d1_delay);
   and MGM_G210(MGM_W179,MGM_W178,MGM_W177);
   not MGM_G211(MGM_W180,d2_delay);
   and MGM_G212(MGM_W181,MGM_W180,MGM_W179);
   and MGM_G213(MGM_W182,si1_delay,MGM_W181);
   and MGM_G214(MGM_W183,si2_delay,MGM_W182);
   not MGM_G215(MGM_W184,ssb_delay);
   and MGM_G216(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W184,MGM_W183);
   not MGM_G217(MGM_W185,clk_delay);
   not MGM_G218(MGM_W186,d1_delay);
   and MGM_G219(MGM_W187,MGM_W186,MGM_W185);
   not MGM_G220(MGM_W188,d2_delay);
   and MGM_G221(MGM_W189,MGM_W188,MGM_W187);
   and MGM_G222(MGM_W190,si1_delay,MGM_W189);
   and MGM_G223(MGM_W191,si2_delay,MGM_W190);
   and MGM_G224(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W191);
   not MGM_G225(MGM_W192,clk_delay);
   not MGM_G226(MGM_W193,d1_delay);
   and MGM_G227(MGM_W194,MGM_W193,MGM_W192);
   and MGM_G228(MGM_W195,d2_delay,MGM_W194);
   not MGM_G229(MGM_W196,si1_delay);
   and MGM_G230(MGM_W197,MGM_W196,MGM_W195);
   not MGM_G231(MGM_W198,si2_delay);
   and MGM_G232(MGM_W199,MGM_W198,MGM_W197);
   not MGM_G233(MGM_W200,ssb_delay);
   and MGM_G234(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W200,MGM_W199);
   not MGM_G235(MGM_W201,clk_delay);
   not MGM_G236(MGM_W202,d1_delay);
   and MGM_G237(MGM_W203,MGM_W202,MGM_W201);
   and MGM_G238(MGM_W204,d2_delay,MGM_W203);
   not MGM_G239(MGM_W205,si1_delay);
   and MGM_G240(MGM_W206,MGM_W205,MGM_W204);
   not MGM_G241(MGM_W207,si2_delay);
   and MGM_G242(MGM_W208,MGM_W207,MGM_W206);
   and MGM_G243(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W208);
   not MGM_G244(MGM_W209,clk_delay);
   not MGM_G245(MGM_W210,d1_delay);
   and MGM_G246(MGM_W211,MGM_W210,MGM_W209);
   and MGM_G247(MGM_W212,d2_delay,MGM_W211);
   not MGM_G248(MGM_W213,si1_delay);
   and MGM_G249(MGM_W214,MGM_W213,MGM_W212);
   and MGM_G250(MGM_W215,si2_delay,MGM_W214);
   not MGM_G251(MGM_W216,ssb_delay);
   and MGM_G252(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W216,MGM_W215);
   not MGM_G253(MGM_W217,clk_delay);
   not MGM_G254(MGM_W218,d1_delay);
   and MGM_G255(MGM_W219,MGM_W218,MGM_W217);
   and MGM_G256(MGM_W220,d2_delay,MGM_W219);
   not MGM_G257(MGM_W221,si1_delay);
   and MGM_G258(MGM_W222,MGM_W221,MGM_W220);
   and MGM_G259(MGM_W223,si2_delay,MGM_W222);
   and MGM_G260(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W223);
   not MGM_G261(MGM_W224,clk_delay);
   not MGM_G262(MGM_W225,d1_delay);
   and MGM_G263(MGM_W226,MGM_W225,MGM_W224);
   and MGM_G264(MGM_W227,d2_delay,MGM_W226);
   and MGM_G265(MGM_W228,si1_delay,MGM_W227);
   not MGM_G266(MGM_W229,si2_delay);
   and MGM_G267(MGM_W230,MGM_W229,MGM_W228);
   not MGM_G268(MGM_W231,ssb_delay);
   and MGM_G269(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W231,MGM_W230);
   not MGM_G270(MGM_W232,clk_delay);
   not MGM_G271(MGM_W233,d1_delay);
   and MGM_G272(MGM_W234,MGM_W233,MGM_W232);
   and MGM_G273(MGM_W235,d2_delay,MGM_W234);
   and MGM_G274(MGM_W236,si1_delay,MGM_W235);
   not MGM_G275(MGM_W237,si2_delay);
   and MGM_G276(MGM_W238,MGM_W237,MGM_W236);
   and MGM_G277(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W238);
   not MGM_G278(MGM_W239,clk_delay);
   not MGM_G279(MGM_W240,d1_delay);
   and MGM_G280(MGM_W241,MGM_W240,MGM_W239);
   and MGM_G281(MGM_W242,d2_delay,MGM_W241);
   and MGM_G282(MGM_W243,si1_delay,MGM_W242);
   and MGM_G283(MGM_W244,si2_delay,MGM_W243);
   not MGM_G284(MGM_W245,ssb_delay);
   and MGM_G285(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W245,MGM_W244);
   not MGM_G286(MGM_W246,clk_delay);
   not MGM_G287(MGM_W247,d1_delay);
   and MGM_G288(MGM_W248,MGM_W247,MGM_W246);
   and MGM_G289(MGM_W249,d2_delay,MGM_W248);
   and MGM_G290(MGM_W250,si1_delay,MGM_W249);
   and MGM_G291(MGM_W251,si2_delay,MGM_W250);
   and MGM_G292(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W251);
   not MGM_G293(MGM_W252,clk_delay);
   and MGM_G294(MGM_W253,d1_delay,MGM_W252);
   not MGM_G295(MGM_W254,d2_delay);
   and MGM_G296(MGM_W255,MGM_W254,MGM_W253);
   not MGM_G297(MGM_W256,si1_delay);
   and MGM_G298(MGM_W257,MGM_W256,MGM_W255);
   not MGM_G299(MGM_W258,si2_delay);
   and MGM_G300(MGM_W259,MGM_W258,MGM_W257);
   not MGM_G301(MGM_W260,ssb_delay);
   and MGM_G302(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W260,MGM_W259);
   not MGM_G303(MGM_W261,clk_delay);
   and MGM_G304(MGM_W262,d1_delay,MGM_W261);
   not MGM_G305(MGM_W263,d2_delay);
   and MGM_G306(MGM_W264,MGM_W263,MGM_W262);
   not MGM_G307(MGM_W265,si1_delay);
   and MGM_G308(MGM_W266,MGM_W265,MGM_W264);
   not MGM_G309(MGM_W267,si2_delay);
   and MGM_G310(MGM_W268,MGM_W267,MGM_W266);
   and MGM_G311(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W268);
   not MGM_G312(MGM_W269,clk_delay);
   and MGM_G313(MGM_W270,d1_delay,MGM_W269);
   not MGM_G314(MGM_W271,d2_delay);
   and MGM_G315(MGM_W272,MGM_W271,MGM_W270);
   not MGM_G316(MGM_W273,si1_delay);
   and MGM_G317(MGM_W274,MGM_W273,MGM_W272);
   and MGM_G318(MGM_W275,si2_delay,MGM_W274);
   not MGM_G319(MGM_W276,ssb_delay);
   and MGM_G320(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W276,MGM_W275);
   not MGM_G321(MGM_W277,clk_delay);
   and MGM_G322(MGM_W278,d1_delay,MGM_W277);
   not MGM_G323(MGM_W279,d2_delay);
   and MGM_G324(MGM_W280,MGM_W279,MGM_W278);
   not MGM_G325(MGM_W281,si1_delay);
   and MGM_G326(MGM_W282,MGM_W281,MGM_W280);
   and MGM_G327(MGM_W283,si2_delay,MGM_W282);
   and MGM_G328(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W283);
   not MGM_G329(MGM_W284,clk_delay);
   and MGM_G330(MGM_W285,d1_delay,MGM_W284);
   not MGM_G331(MGM_W286,d2_delay);
   and MGM_G332(MGM_W287,MGM_W286,MGM_W285);
   and MGM_G333(MGM_W288,si1_delay,MGM_W287);
   not MGM_G334(MGM_W289,si2_delay);
   and MGM_G335(MGM_W290,MGM_W289,MGM_W288);
   not MGM_G336(MGM_W291,ssb_delay);
   and MGM_G337(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W291,MGM_W290);
   not MGM_G338(MGM_W292,clk_delay);
   and MGM_G339(MGM_W293,d1_delay,MGM_W292);
   not MGM_G340(MGM_W294,d2_delay);
   and MGM_G341(MGM_W295,MGM_W294,MGM_W293);
   and MGM_G342(MGM_W296,si1_delay,MGM_W295);
   not MGM_G343(MGM_W297,si2_delay);
   and MGM_G344(MGM_W298,MGM_W297,MGM_W296);
   and MGM_G345(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W298);
   not MGM_G346(MGM_W299,clk_delay);
   and MGM_G347(MGM_W300,d1_delay,MGM_W299);
   not MGM_G348(MGM_W301,d2_delay);
   and MGM_G349(MGM_W302,MGM_W301,MGM_W300);
   and MGM_G350(MGM_W303,si1_delay,MGM_W302);
   and MGM_G351(MGM_W304,si2_delay,MGM_W303);
   not MGM_G352(MGM_W305,ssb_delay);
   and MGM_G353(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W305,MGM_W304);
   not MGM_G354(MGM_W306,clk_delay);
   and MGM_G355(MGM_W307,d1_delay,MGM_W306);
   not MGM_G356(MGM_W308,d2_delay);
   and MGM_G357(MGM_W309,MGM_W308,MGM_W307);
   and MGM_G358(MGM_W310,si1_delay,MGM_W309);
   and MGM_G359(MGM_W311,si2_delay,MGM_W310);
   and MGM_G360(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W311);
   not MGM_G361(MGM_W312,clk_delay);
   and MGM_G362(MGM_W313,d1_delay,MGM_W312);
   and MGM_G363(MGM_W314,d2_delay,MGM_W313);
   not MGM_G364(MGM_W315,si1_delay);
   and MGM_G365(MGM_W316,MGM_W315,MGM_W314);
   not MGM_G366(MGM_W317,si2_delay);
   and MGM_G367(MGM_W318,MGM_W317,MGM_W316);
   not MGM_G368(MGM_W319,ssb_delay);
   and MGM_G369(ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W319,MGM_W318);
   not MGM_G370(MGM_W320,clk_delay);
   and MGM_G371(MGM_W321,d1_delay,MGM_W320);
   and MGM_G372(MGM_W322,d2_delay,MGM_W321);
   not MGM_G373(MGM_W323,si1_delay);
   and MGM_G374(MGM_W324,MGM_W323,MGM_W322);
   not MGM_G375(MGM_W325,si2_delay);
   and MGM_G376(MGM_W326,MGM_W325,MGM_W324);
   and MGM_G377(ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W326);
   not MGM_G378(MGM_W327,clk_delay);
   and MGM_G379(MGM_W328,d1_delay,MGM_W327);
   and MGM_G380(MGM_W329,d2_delay,MGM_W328);
   not MGM_G381(MGM_W330,si1_delay);
   and MGM_G382(MGM_W331,MGM_W330,MGM_W329);
   and MGM_G383(MGM_W332,si2_delay,MGM_W331);
   not MGM_G384(MGM_W333,ssb_delay);
   and MGM_G385(ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W333,MGM_W332);
   not MGM_G386(MGM_W334,clk_delay);
   and MGM_G387(MGM_W335,d1_delay,MGM_W334);
   and MGM_G388(MGM_W336,d2_delay,MGM_W335);
   not MGM_G389(MGM_W337,si1_delay);
   and MGM_G390(MGM_W338,MGM_W337,MGM_W336);
   and MGM_G391(MGM_W339,si2_delay,MGM_W338);
   and MGM_G392(ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W339);
   not MGM_G393(MGM_W340,clk_delay);
   and MGM_G394(MGM_W341,d1_delay,MGM_W340);
   and MGM_G395(MGM_W342,d2_delay,MGM_W341);
   and MGM_G396(MGM_W343,si1_delay,MGM_W342);
   not MGM_G397(MGM_W344,si2_delay);
   and MGM_G398(MGM_W345,MGM_W344,MGM_W343);
   not MGM_G399(MGM_W346,ssb_delay);
   and MGM_G400(ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W346,MGM_W345);
   not MGM_G401(MGM_W347,clk_delay);
   and MGM_G402(MGM_W348,d1_delay,MGM_W347);
   and MGM_G403(MGM_W349,d2_delay,MGM_W348);
   and MGM_G404(MGM_W350,si1_delay,MGM_W349);
   not MGM_G405(MGM_W351,si2_delay);
   and MGM_G406(MGM_W352,MGM_W351,MGM_W350);
   and MGM_G407(ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W352);
   not MGM_G408(MGM_W353,clk_delay);
   and MGM_G409(MGM_W354,d1_delay,MGM_W353);
   and MGM_G410(MGM_W355,d2_delay,MGM_W354);
   and MGM_G411(MGM_W356,si1_delay,MGM_W355);
   and MGM_G412(MGM_W357,si2_delay,MGM_W356);
   not MGM_G413(MGM_W358,ssb_delay);
   and MGM_G414(ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W358,MGM_W357);
   not MGM_G415(MGM_W359,clk_delay);
   and MGM_G416(MGM_W360,d1_delay,MGM_W359);
   and MGM_G417(MGM_W361,d2_delay,MGM_W360);
   and MGM_G418(MGM_W362,si1_delay,MGM_W361);
   and MGM_G419(MGM_W363,si2_delay,MGM_W362);
   and MGM_G420(ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W363);
   not MGM_G421(MGM_W364,d1_delay);
   and MGM_G422(MGM_W365,MGM_W364,clk_delay);
   not MGM_G423(MGM_W366,d2_delay);
   and MGM_G424(MGM_W367,MGM_W366,MGM_W365);
   not MGM_G425(MGM_W368,si1_delay);
   and MGM_G426(MGM_W369,MGM_W368,MGM_W367);
   not MGM_G427(MGM_W370,si2_delay);
   and MGM_G428(MGM_W371,MGM_W370,MGM_W369);
   not MGM_G429(MGM_W372,ssb_delay);
   and MGM_G430(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W372,MGM_W371);
   not MGM_G431(MGM_W373,d1_delay);
   and MGM_G432(MGM_W374,MGM_W373,clk_delay);
   not MGM_G433(MGM_W375,d2_delay);
   and MGM_G434(MGM_W376,MGM_W375,MGM_W374);
   not MGM_G435(MGM_W377,si1_delay);
   and MGM_G436(MGM_W378,MGM_W377,MGM_W376);
   not MGM_G437(MGM_W379,si2_delay);
   and MGM_G438(MGM_W380,MGM_W379,MGM_W378);
   and MGM_G439(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W380);
   not MGM_G440(MGM_W381,d1_delay);
   and MGM_G441(MGM_W382,MGM_W381,clk_delay);
   not MGM_G442(MGM_W383,d2_delay);
   and MGM_G443(MGM_W384,MGM_W383,MGM_W382);
   not MGM_G444(MGM_W385,si1_delay);
   and MGM_G445(MGM_W386,MGM_W385,MGM_W384);
   and MGM_G446(MGM_W387,si2_delay,MGM_W386);
   not MGM_G447(MGM_W388,ssb_delay);
   and MGM_G448(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W388,MGM_W387);
   not MGM_G449(MGM_W389,d1_delay);
   and MGM_G450(MGM_W390,MGM_W389,clk_delay);
   not MGM_G451(MGM_W391,d2_delay);
   and MGM_G452(MGM_W392,MGM_W391,MGM_W390);
   not MGM_G453(MGM_W393,si1_delay);
   and MGM_G454(MGM_W394,MGM_W393,MGM_W392);
   and MGM_G455(MGM_W395,si2_delay,MGM_W394);
   and MGM_G456(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W395);
   not MGM_G457(MGM_W396,d1_delay);
   and MGM_G458(MGM_W397,MGM_W396,clk_delay);
   not MGM_G459(MGM_W398,d2_delay);
   and MGM_G460(MGM_W399,MGM_W398,MGM_W397);
   and MGM_G461(MGM_W400,si1_delay,MGM_W399);
   not MGM_G462(MGM_W401,si2_delay);
   and MGM_G463(MGM_W402,MGM_W401,MGM_W400);
   not MGM_G464(MGM_W403,ssb_delay);
   and MGM_G465(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W403,MGM_W402);
   not MGM_G466(MGM_W404,d1_delay);
   and MGM_G467(MGM_W405,MGM_W404,clk_delay);
   not MGM_G468(MGM_W406,d2_delay);
   and MGM_G469(MGM_W407,MGM_W406,MGM_W405);
   and MGM_G470(MGM_W408,si1_delay,MGM_W407);
   not MGM_G471(MGM_W409,si2_delay);
   and MGM_G472(MGM_W410,MGM_W409,MGM_W408);
   and MGM_G473(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W410);
   not MGM_G474(MGM_W411,d1_delay);
   and MGM_G475(MGM_W412,MGM_W411,clk_delay);
   not MGM_G476(MGM_W413,d2_delay);
   and MGM_G477(MGM_W414,MGM_W413,MGM_W412);
   and MGM_G478(MGM_W415,si1_delay,MGM_W414);
   and MGM_G479(MGM_W416,si2_delay,MGM_W415);
   not MGM_G480(MGM_W417,ssb_delay);
   and MGM_G481(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W417,MGM_W416);
   not MGM_G482(MGM_W418,d1_delay);
   and MGM_G483(MGM_W419,MGM_W418,clk_delay);
   not MGM_G484(MGM_W420,d2_delay);
   and MGM_G485(MGM_W421,MGM_W420,MGM_W419);
   and MGM_G486(MGM_W422,si1_delay,MGM_W421);
   and MGM_G487(MGM_W423,si2_delay,MGM_W422);
   and MGM_G488(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W423);
   not MGM_G489(MGM_W424,d1_delay);
   and MGM_G490(MGM_W425,MGM_W424,clk_delay);
   and MGM_G491(MGM_W426,d2_delay,MGM_W425);
   not MGM_G492(MGM_W427,si1_delay);
   and MGM_G493(MGM_W428,MGM_W427,MGM_W426);
   not MGM_G494(MGM_W429,si2_delay);
   and MGM_G495(MGM_W430,MGM_W429,MGM_W428);
   not MGM_G496(MGM_W431,ssb_delay);
   and MGM_G497(ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W431,MGM_W430);
   not MGM_G498(MGM_W432,d1_delay);
   and MGM_G499(MGM_W433,MGM_W432,clk_delay);
   and MGM_G500(MGM_W434,d2_delay,MGM_W433);
   not MGM_G501(MGM_W435,si1_delay);
   and MGM_G502(MGM_W436,MGM_W435,MGM_W434);
   not MGM_G503(MGM_W437,si2_delay);
   and MGM_G504(MGM_W438,MGM_W437,MGM_W436);
   and MGM_G505(ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W438);
   not MGM_G506(MGM_W439,d1_delay);
   and MGM_G507(MGM_W440,MGM_W439,clk_delay);
   and MGM_G508(MGM_W441,d2_delay,MGM_W440);
   not MGM_G509(MGM_W442,si1_delay);
   and MGM_G510(MGM_W443,MGM_W442,MGM_W441);
   and MGM_G511(MGM_W444,si2_delay,MGM_W443);
   not MGM_G512(MGM_W445,ssb_delay);
   and MGM_G513(ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W445,MGM_W444);
   not MGM_G514(MGM_W446,d1_delay);
   and MGM_G515(MGM_W447,MGM_W446,clk_delay);
   and MGM_G516(MGM_W448,d2_delay,MGM_W447);
   not MGM_G517(MGM_W449,si1_delay);
   and MGM_G518(MGM_W450,MGM_W449,MGM_W448);
   and MGM_G519(MGM_W451,si2_delay,MGM_W450);
   and MGM_G520(ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W451);
   not MGM_G521(MGM_W452,d1_delay);
   and MGM_G522(MGM_W453,MGM_W452,clk_delay);
   and MGM_G523(MGM_W454,d2_delay,MGM_W453);
   and MGM_G524(MGM_W455,si1_delay,MGM_W454);
   not MGM_G525(MGM_W456,si2_delay);
   and MGM_G526(MGM_W457,MGM_W456,MGM_W455);
   not MGM_G527(MGM_W458,ssb_delay);
   and MGM_G528(ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W458,MGM_W457);
   not MGM_G529(MGM_W459,d1_delay);
   and MGM_G530(MGM_W460,MGM_W459,clk_delay);
   and MGM_G531(MGM_W461,d2_delay,MGM_W460);
   and MGM_G532(MGM_W462,si1_delay,MGM_W461);
   not MGM_G533(MGM_W463,si2_delay);
   and MGM_G534(MGM_W464,MGM_W463,MGM_W462);
   and MGM_G535(ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W464);
   not MGM_G536(MGM_W465,d1_delay);
   and MGM_G537(MGM_W466,MGM_W465,clk_delay);
   and MGM_G538(MGM_W467,d2_delay,MGM_W466);
   and MGM_G539(MGM_W468,si1_delay,MGM_W467);
   and MGM_G540(MGM_W469,si2_delay,MGM_W468);
   not MGM_G541(MGM_W470,ssb_delay);
   and MGM_G542(ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W470,MGM_W469);
   not MGM_G543(MGM_W471,d1_delay);
   and MGM_G544(MGM_W472,MGM_W471,clk_delay);
   and MGM_G545(MGM_W473,d2_delay,MGM_W472);
   and MGM_G546(MGM_W474,si1_delay,MGM_W473);
   and MGM_G547(MGM_W475,si2_delay,MGM_W474);
   and MGM_G548(ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W475);
   and MGM_G549(MGM_W476,d1_delay,clk_delay);
   not MGM_G550(MGM_W477,d2_delay);
   and MGM_G551(MGM_W478,MGM_W477,MGM_W476);
   not MGM_G552(MGM_W479,si1_delay);
   and MGM_G553(MGM_W480,MGM_W479,MGM_W478);
   not MGM_G554(MGM_W481,si2_delay);
   and MGM_G555(MGM_W482,MGM_W481,MGM_W480);
   not MGM_G556(MGM_W483,ssb_delay);
   and MGM_G557(ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W483,MGM_W482);
   and MGM_G558(MGM_W484,d1_delay,clk_delay);
   not MGM_G559(MGM_W485,d2_delay);
   and MGM_G560(MGM_W486,MGM_W485,MGM_W484);
   not MGM_G561(MGM_W487,si1_delay);
   and MGM_G562(MGM_W488,MGM_W487,MGM_W486);
   not MGM_G563(MGM_W489,si2_delay);
   and MGM_G564(MGM_W490,MGM_W489,MGM_W488);
   and MGM_G565(ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W490);
   and MGM_G566(MGM_W491,d1_delay,clk_delay);
   not MGM_G567(MGM_W492,d2_delay);
   and MGM_G568(MGM_W493,MGM_W492,MGM_W491);
   not MGM_G569(MGM_W494,si1_delay);
   and MGM_G570(MGM_W495,MGM_W494,MGM_W493);
   and MGM_G571(MGM_W496,si2_delay,MGM_W495);
   not MGM_G572(MGM_W497,ssb_delay);
   and MGM_G573(ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W497,MGM_W496);
   and MGM_G574(MGM_W498,d1_delay,clk_delay);
   not MGM_G575(MGM_W499,d2_delay);
   and MGM_G576(MGM_W500,MGM_W499,MGM_W498);
   not MGM_G577(MGM_W501,si1_delay);
   and MGM_G578(MGM_W502,MGM_W501,MGM_W500);
   and MGM_G579(MGM_W503,si2_delay,MGM_W502);
   and MGM_G580(ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W503);
   and MGM_G581(MGM_W504,d1_delay,clk_delay);
   not MGM_G582(MGM_W505,d2_delay);
   and MGM_G583(MGM_W506,MGM_W505,MGM_W504);
   and MGM_G584(MGM_W507,si1_delay,MGM_W506);
   not MGM_G585(MGM_W508,si2_delay);
   and MGM_G586(MGM_W509,MGM_W508,MGM_W507);
   not MGM_G587(MGM_W510,ssb_delay);
   and MGM_G588(ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W510,MGM_W509);
   and MGM_G589(MGM_W511,d1_delay,clk_delay);
   not MGM_G590(MGM_W512,d2_delay);
   and MGM_G591(MGM_W513,MGM_W512,MGM_W511);
   and MGM_G592(MGM_W514,si1_delay,MGM_W513);
   not MGM_G593(MGM_W515,si2_delay);
   and MGM_G594(MGM_W516,MGM_W515,MGM_W514);
   and MGM_G595(ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W516);
   and MGM_G596(MGM_W517,d1_delay,clk_delay);
   not MGM_G597(MGM_W518,d2_delay);
   and MGM_G598(MGM_W519,MGM_W518,MGM_W517);
   and MGM_G599(MGM_W520,si1_delay,MGM_W519);
   and MGM_G600(MGM_W521,si2_delay,MGM_W520);
   not MGM_G601(MGM_W522,ssb_delay);
   and MGM_G602(ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W522,MGM_W521);
   and MGM_G603(MGM_W523,d1_delay,clk_delay);
   not MGM_G604(MGM_W524,d2_delay);
   and MGM_G605(MGM_W525,MGM_W524,MGM_W523);
   and MGM_G606(MGM_W526,si1_delay,MGM_W525);
   and MGM_G607(MGM_W527,si2_delay,MGM_W526);
   and MGM_G608(ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W527);
   and MGM_G609(MGM_W528,d1_delay,clk_delay);
   and MGM_G610(MGM_W529,d2_delay,MGM_W528);
   not MGM_G611(MGM_W530,si1_delay);
   and MGM_G612(MGM_W531,MGM_W530,MGM_W529);
   not MGM_G613(MGM_W532,si2_delay);
   and MGM_G614(MGM_W533,MGM_W532,MGM_W531);
   not MGM_G615(MGM_W534,ssb_delay);
   and MGM_G616(ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W534,MGM_W533);
   and MGM_G617(MGM_W535,d1_delay,clk_delay);
   and MGM_G618(MGM_W536,d2_delay,MGM_W535);
   not MGM_G619(MGM_W537,si1_delay);
   and MGM_G620(MGM_W538,MGM_W537,MGM_W536);
   not MGM_G621(MGM_W539,si2_delay);
   and MGM_G622(MGM_W540,MGM_W539,MGM_W538);
   and MGM_G623(ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W540);
   and MGM_G624(MGM_W541,d1_delay,clk_delay);
   and MGM_G625(MGM_W542,d2_delay,MGM_W541);
   not MGM_G626(MGM_W543,si1_delay);
   and MGM_G627(MGM_W544,MGM_W543,MGM_W542);
   and MGM_G628(MGM_W545,si2_delay,MGM_W544);
   not MGM_G629(MGM_W546,ssb_delay);
   and MGM_G630(ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W546,MGM_W545);
   and MGM_G631(MGM_W547,d1_delay,clk_delay);
   and MGM_G632(MGM_W548,d2_delay,MGM_W547);
   not MGM_G633(MGM_W549,si1_delay);
   and MGM_G634(MGM_W550,MGM_W549,MGM_W548);
   and MGM_G635(MGM_W551,si2_delay,MGM_W550);
   and MGM_G636(ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W551);
   and MGM_G637(MGM_W552,d1_delay,clk_delay);
   and MGM_G638(MGM_W553,d2_delay,MGM_W552);
   and MGM_G639(MGM_W554,si1_delay,MGM_W553);
   not MGM_G640(MGM_W555,si2_delay);
   and MGM_G641(MGM_W556,MGM_W555,MGM_W554);
   not MGM_G642(MGM_W557,ssb_delay);
   and MGM_G643(ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W557,MGM_W556);
   and MGM_G644(MGM_W558,d1_delay,clk_delay);
   and MGM_G645(MGM_W559,d2_delay,MGM_W558);
   and MGM_G646(MGM_W560,si1_delay,MGM_W559);
   not MGM_G647(MGM_W561,si2_delay);
   and MGM_G648(MGM_W562,MGM_W561,MGM_W560);
   and MGM_G649(ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W562);
   and MGM_G650(MGM_W563,d1_delay,clk_delay);
   and MGM_G651(MGM_W564,d2_delay,MGM_W563);
   and MGM_G652(MGM_W565,si1_delay,MGM_W564);
   and MGM_G653(MGM_W566,si2_delay,MGM_W565);
   not MGM_G654(MGM_W567,ssb_delay);
   and MGM_G655(ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W567,MGM_W566);
   and MGM_G656(MGM_W568,d1_delay,clk_delay);
   and MGM_G657(MGM_W569,d2_delay,MGM_W568);
   and MGM_G658(MGM_W570,si1_delay,MGM_W569);
   and MGM_G659(MGM_W571,si2_delay,MGM_W570);
   and MGM_G660(ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W571);
   not MGM_G661(MGM_W572,d1_delay);
   not MGM_G662(MGM_W573,d2_delay);
   and MGM_G663(MGM_W574,MGM_W573,MGM_W572);
   and MGM_G664(MGM_W575,rb_delay,MGM_W574);
   not MGM_G665(MGM_W576,si1_delay);
   and MGM_G666(MGM_W577,MGM_W576,MGM_W575);
   and MGM_G667(ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2,si2_delay,MGM_W577);
   not MGM_G668(MGM_W578,d1_delay);
   not MGM_G669(MGM_W579,d2_delay);
   and MGM_G670(MGM_W580,MGM_W579,MGM_W578);
   and MGM_G671(MGM_W581,rb_delay,MGM_W580);
   and MGM_G672(MGM_W582,si1_delay,MGM_W581);
   not MGM_G673(MGM_W583,si2_delay);
   and MGM_G674(ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2,MGM_W583,MGM_W582);
   not MGM_G675(MGM_W584,d1_delay);
   not MGM_G676(MGM_W585,d2_delay);
   and MGM_G677(MGM_W586,MGM_W585,MGM_W584);
   and MGM_G678(MGM_W587,rb_delay,MGM_W586);
   and MGM_G679(MGM_W588,si1_delay,MGM_W587);
   and MGM_G680(ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2,si2_delay,MGM_W588);
   not MGM_G681(MGM_W589,d1_delay);
   and MGM_G682(MGM_W590,d2_delay,MGM_W589);
   and MGM_G683(MGM_W591,rb_delay,MGM_W590);
   not MGM_G684(MGM_W592,si1_delay);
   and MGM_G685(MGM_W593,MGM_W592,MGM_W591);
   not MGM_G686(MGM_W594,si2_delay);
   and MGM_G687(ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2,MGM_W594,MGM_W593);
   not MGM_G688(MGM_W595,d1_delay);
   and MGM_G689(MGM_W596,d2_delay,MGM_W595);
   and MGM_G690(MGM_W597,rb_delay,MGM_W596);
   and MGM_G691(MGM_W598,si1_delay,MGM_W597);
   not MGM_G692(MGM_W599,si2_delay);
   and MGM_G693(ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2,MGM_W599,MGM_W598);
   not MGM_G694(MGM_W600,d1_delay);
   and MGM_G695(MGM_W601,d2_delay,MGM_W600);
   and MGM_G696(MGM_W602,rb_delay,MGM_W601);
   and MGM_G697(MGM_W603,si1_delay,MGM_W602);
   and MGM_G698(ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2,si2_delay,MGM_W603);
   not MGM_G699(MGM_W604,d2_delay);
   and MGM_G700(MGM_W605,MGM_W604,d1_delay);
   and MGM_G701(MGM_W606,rb_delay,MGM_W605);
   not MGM_G702(MGM_W607,si1_delay);
   and MGM_G703(MGM_W608,MGM_W607,MGM_W606);
   not MGM_G704(MGM_W609,si2_delay);
   and MGM_G705(ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2,MGM_W609,MGM_W608);
   not MGM_G706(MGM_W610,d2_delay);
   and MGM_G707(MGM_W611,MGM_W610,d1_delay);
   and MGM_G708(MGM_W612,rb_delay,MGM_W611);
   not MGM_G709(MGM_W613,si1_delay);
   and MGM_G710(MGM_W614,MGM_W613,MGM_W612);
   and MGM_G711(ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2,si2_delay,MGM_W614);
   not MGM_G712(MGM_W615,d2_delay);
   and MGM_G713(MGM_W616,MGM_W615,d1_delay);
   and MGM_G714(MGM_W617,rb_delay,MGM_W616);
   and MGM_G715(MGM_W618,si1_delay,MGM_W617);
   and MGM_G716(ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2,si2_delay,MGM_W618);
   and MGM_G717(MGM_W619,d2_delay,d1_delay);
   and MGM_G718(MGM_W620,rb_delay,MGM_W619);
   not MGM_G719(MGM_W621,si1_delay);
   and MGM_G720(MGM_W622,MGM_W621,MGM_W620);
   not MGM_G721(MGM_W623,si2_delay);
   and MGM_G722(ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2,MGM_W623,MGM_W622);
   and MGM_G723(MGM_W624,d2_delay,d1_delay);
   and MGM_G724(MGM_W625,rb_delay,MGM_W624);
   not MGM_G725(MGM_W626,si1_delay);
   and MGM_G726(MGM_W627,MGM_W626,MGM_W625);
   and MGM_G727(ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2,si2_delay,MGM_W627);
   and MGM_G728(MGM_W628,d2_delay,d1_delay);
   and MGM_G729(MGM_W629,rb_delay,MGM_W628);
   and MGM_G730(MGM_W630,si1_delay,MGM_W629);
   not MGM_G731(MGM_W631,si2_delay);
   and MGM_G732(ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2,MGM_W631,MGM_W630);
   and MGM_G733(ENABLE_ssb_AND_rb,rb_delay,ssb_delay);
   not MGM_G734(MGM_W632,ssb_delay);
   and MGM_G735(ENABLE_NOT_ssb_AND_rb,rb_delay,MGM_W632);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d1==1'b0 && rb==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_rb == 1'b1)
      ,0.0,0,notifier);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb,0.0,0,notifier);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,negedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,posedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d1 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d1 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d2 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d2 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si1 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si1 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si2 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si2 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy203ah1n03x5( clk, d1, d2, o1, o2, rb, si1, si2, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, rb, si1, si2, ssb;
   output o1, o2;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy203ah_func b15fqy203ah1n03x5_behav_inst(.clk(clk),.rb(rb),.ssb(ssb),.o1(o1),.o2(o2),.d1(d1),.d2(d2),.si1(si1),.si2(si2),.notifier0(1'b0),.notifier1(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy203ah_func b15fqy203ah1n03x5_behav_inst(.clk(clk),.rb(rb),.ssb(ssb),.o1(o1),.o2(o2),.d1(d1),.d2(d2),.si1(si1),.si2(si2),.notifier0(1'b0),.notifier1(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire rb_delay ;
   wire ssb_delay ;
   wire d1_delay ;
   wire d2_delay ;
   wire si1_delay ;
   wire si2_delay ;
   reg notifier;
   reg notifier0;
   reg notifier1;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
     notifier1 = (notifier1 !== notifier) ? notifier : ~notifier1;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy203ah_func b15fqy203ah1n03x5_inst(.clk(clk_delay),.rb(rb_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.d1(d1_delay),.d2(d2_delay),.si1(si1_delay),.si2(si2_delay),.notifier0(notifier0),.notifier1(notifier1),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy203ah_func b15fqy203ah1n03x5_inst(.clk(clk_delay),.rb(rb_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.d1(d1_delay),.d2(d2_delay),.si1(si1_delay),.si2(si2_delay),.notifier0(notifier0),.notifier1(notifier1));
   `endif
   
   // spec_gates_begin
   buf MGM_G0(ENABLE_rb,rb_delay);
   not MGM_G1(MGM_W0,d1_delay);
   not MGM_G2(MGM_W1,d2_delay);
   and MGM_G3(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G4(MGM_W3,si1_delay);
   and MGM_G5(MGM_W4,MGM_W3,MGM_W2);
   and MGM_G6(MGM_W5,si2_delay,MGM_W4);
   not MGM_G7(MGM_W6,ssb_delay);
   and MGM_G8(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W6,MGM_W5);
   not MGM_G9(MGM_W7,d1_delay);
   not MGM_G10(MGM_W8,d2_delay);
   and MGM_G11(MGM_W9,MGM_W8,MGM_W7);
   and MGM_G12(MGM_W10,si1_delay,MGM_W9);
   not MGM_G13(MGM_W11,si2_delay);
   and MGM_G14(MGM_W12,MGM_W11,MGM_W10);
   not MGM_G15(MGM_W13,ssb_delay);
   and MGM_G16(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W13,MGM_W12);
   not MGM_G17(MGM_W14,d1_delay);
   not MGM_G18(MGM_W15,d2_delay);
   and MGM_G19(MGM_W16,MGM_W15,MGM_W14);
   and MGM_G20(MGM_W17,si1_delay,MGM_W16);
   and MGM_G21(MGM_W18,si2_delay,MGM_W17);
   not MGM_G22(MGM_W19,ssb_delay);
   and MGM_G23(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W19,MGM_W18);
   not MGM_G24(MGM_W20,d1_delay);
   and MGM_G25(MGM_W21,d2_delay,MGM_W20);
   not MGM_G26(MGM_W22,si1_delay);
   and MGM_G27(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G28(MGM_W24,si2_delay);
   and MGM_G29(MGM_W25,MGM_W24,MGM_W23);
   and MGM_G30(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W25);
   not MGM_G31(MGM_W26,d1_delay);
   and MGM_G32(MGM_W27,d2_delay,MGM_W26);
   not MGM_G33(MGM_W28,si1_delay);
   and MGM_G34(MGM_W29,MGM_W28,MGM_W27);
   and MGM_G35(MGM_W30,si2_delay,MGM_W29);
   not MGM_G36(MGM_W31,ssb_delay);
   and MGM_G37(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W31,MGM_W30);
   not MGM_G38(MGM_W32,d1_delay);
   and MGM_G39(MGM_W33,d2_delay,MGM_W32);
   not MGM_G40(MGM_W34,si1_delay);
   and MGM_G41(MGM_W35,MGM_W34,MGM_W33);
   and MGM_G42(MGM_W36,si2_delay,MGM_W35);
   and MGM_G43(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W36);
   not MGM_G44(MGM_W37,d1_delay);
   and MGM_G45(MGM_W38,d2_delay,MGM_W37);
   and MGM_G46(MGM_W39,si1_delay,MGM_W38);
   not MGM_G47(MGM_W40,si2_delay);
   and MGM_G48(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G49(MGM_W42,ssb_delay);
   and MGM_G50(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W42,MGM_W41);
   not MGM_G51(MGM_W43,d1_delay);
   and MGM_G52(MGM_W44,d2_delay,MGM_W43);
   and MGM_G53(MGM_W45,si1_delay,MGM_W44);
   not MGM_G54(MGM_W46,si2_delay);
   and MGM_G55(MGM_W47,MGM_W46,MGM_W45);
   and MGM_G56(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W47);
   not MGM_G57(MGM_W48,d1_delay);
   and MGM_G58(MGM_W49,d2_delay,MGM_W48);
   and MGM_G59(MGM_W50,si1_delay,MGM_W49);
   and MGM_G60(MGM_W51,si2_delay,MGM_W50);
   not MGM_G61(MGM_W52,ssb_delay);
   and MGM_G62(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W52,MGM_W51);
   not MGM_G63(MGM_W53,d1_delay);
   and MGM_G64(MGM_W54,d2_delay,MGM_W53);
   and MGM_G65(MGM_W55,si1_delay,MGM_W54);
   and MGM_G66(MGM_W56,si2_delay,MGM_W55);
   and MGM_G67(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W56);
   not MGM_G68(MGM_W57,d2_delay);
   and MGM_G69(MGM_W58,MGM_W57,d1_delay);
   not MGM_G70(MGM_W59,si1_delay);
   and MGM_G71(MGM_W60,MGM_W59,MGM_W58);
   not MGM_G72(MGM_W61,si2_delay);
   and MGM_G73(MGM_W62,MGM_W61,MGM_W60);
   and MGM_G74(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W62);
   not MGM_G75(MGM_W63,d2_delay);
   and MGM_G76(MGM_W64,MGM_W63,d1_delay);
   not MGM_G77(MGM_W65,si1_delay);
   and MGM_G78(MGM_W66,MGM_W65,MGM_W64);
   and MGM_G79(MGM_W67,si2_delay,MGM_W66);
   not MGM_G80(MGM_W68,ssb_delay);
   and MGM_G81(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W68,MGM_W67);
   not MGM_G82(MGM_W69,d2_delay);
   and MGM_G83(MGM_W70,MGM_W69,d1_delay);
   not MGM_G84(MGM_W71,si1_delay);
   and MGM_G85(MGM_W72,MGM_W71,MGM_W70);
   and MGM_G86(MGM_W73,si2_delay,MGM_W72);
   and MGM_G87(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W73);
   not MGM_G88(MGM_W74,d2_delay);
   and MGM_G89(MGM_W75,MGM_W74,d1_delay);
   and MGM_G90(MGM_W76,si1_delay,MGM_W75);
   not MGM_G91(MGM_W77,si2_delay);
   and MGM_G92(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G93(MGM_W79,ssb_delay);
   and MGM_G94(ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G95(MGM_W80,d2_delay);
   and MGM_G96(MGM_W81,MGM_W80,d1_delay);
   and MGM_G97(MGM_W82,si1_delay,MGM_W81);
   not MGM_G98(MGM_W83,si2_delay);
   and MGM_G99(MGM_W84,MGM_W83,MGM_W82);
   and MGM_G100(ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W84);
   not MGM_G101(MGM_W85,d2_delay);
   and MGM_G102(MGM_W86,MGM_W85,d1_delay);
   and MGM_G103(MGM_W87,si1_delay,MGM_W86);
   and MGM_G104(MGM_W88,si2_delay,MGM_W87);
   not MGM_G105(MGM_W89,ssb_delay);
   and MGM_G106(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W89,MGM_W88);
   not MGM_G107(MGM_W90,d2_delay);
   and MGM_G108(MGM_W91,MGM_W90,d1_delay);
   and MGM_G109(MGM_W92,si1_delay,MGM_W91);
   and MGM_G110(MGM_W93,si2_delay,MGM_W92);
   and MGM_G111(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W93);
   and MGM_G112(MGM_W94,d2_delay,d1_delay);
   not MGM_G113(MGM_W95,si1_delay);
   and MGM_G114(MGM_W96,MGM_W95,MGM_W94);
   not MGM_G115(MGM_W97,si2_delay);
   and MGM_G116(MGM_W98,MGM_W97,MGM_W96);
   and MGM_G117(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W98);
   and MGM_G118(MGM_W99,d2_delay,d1_delay);
   not MGM_G119(MGM_W100,si1_delay);
   and MGM_G120(MGM_W101,MGM_W100,MGM_W99);
   and MGM_G121(MGM_W102,si2_delay,MGM_W101);
   not MGM_G122(MGM_W103,ssb_delay);
   and MGM_G123(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W103,MGM_W102);
   and MGM_G124(MGM_W104,d2_delay,d1_delay);
   not MGM_G125(MGM_W105,si1_delay);
   and MGM_G126(MGM_W106,MGM_W105,MGM_W104);
   and MGM_G127(MGM_W107,si2_delay,MGM_W106);
   and MGM_G128(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W107);
   and MGM_G129(MGM_W108,d2_delay,d1_delay);
   and MGM_G130(MGM_W109,si1_delay,MGM_W108);
   not MGM_G131(MGM_W110,si2_delay);
   and MGM_G132(MGM_W111,MGM_W110,MGM_W109);
   not MGM_G133(MGM_W112,ssb_delay);
   and MGM_G134(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W112,MGM_W111);
   and MGM_G135(MGM_W113,d2_delay,d1_delay);
   and MGM_G136(MGM_W114,si1_delay,MGM_W113);
   not MGM_G137(MGM_W115,si2_delay);
   and MGM_G138(MGM_W116,MGM_W115,MGM_W114);
   and MGM_G139(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W116);
   and MGM_G140(MGM_W117,d2_delay,d1_delay);
   and MGM_G141(MGM_W118,si1_delay,MGM_W117);
   and MGM_G142(MGM_W119,si2_delay,MGM_W118);
   not MGM_G143(MGM_W120,ssb_delay);
   and MGM_G144(ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W120,MGM_W119);
   and MGM_G145(MGM_W121,d2_delay,d1_delay);
   and MGM_G146(MGM_W122,si1_delay,MGM_W121);
   and MGM_G147(MGM_W123,si2_delay,MGM_W122);
   and MGM_G148(ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W123);
   not MGM_G149(MGM_W124,clk_delay);
   not MGM_G150(MGM_W125,d1_delay);
   and MGM_G151(MGM_W126,MGM_W125,MGM_W124);
   not MGM_G152(MGM_W127,d2_delay);
   and MGM_G153(MGM_W128,MGM_W127,MGM_W126);
   not MGM_G154(MGM_W129,si1_delay);
   and MGM_G155(MGM_W130,MGM_W129,MGM_W128);
   not MGM_G156(MGM_W131,si2_delay);
   and MGM_G157(MGM_W132,MGM_W131,MGM_W130);
   not MGM_G158(MGM_W133,ssb_delay);
   and MGM_G159(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W133,MGM_W132);
   not MGM_G160(MGM_W134,clk_delay);
   not MGM_G161(MGM_W135,d1_delay);
   and MGM_G162(MGM_W136,MGM_W135,MGM_W134);
   not MGM_G163(MGM_W137,d2_delay);
   and MGM_G164(MGM_W138,MGM_W137,MGM_W136);
   not MGM_G165(MGM_W139,si1_delay);
   and MGM_G166(MGM_W140,MGM_W139,MGM_W138);
   not MGM_G167(MGM_W141,si2_delay);
   and MGM_G168(MGM_W142,MGM_W141,MGM_W140);
   and MGM_G169(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W142);
   not MGM_G170(MGM_W143,clk_delay);
   not MGM_G171(MGM_W144,d1_delay);
   and MGM_G172(MGM_W145,MGM_W144,MGM_W143);
   not MGM_G173(MGM_W146,d2_delay);
   and MGM_G174(MGM_W147,MGM_W146,MGM_W145);
   not MGM_G175(MGM_W148,si1_delay);
   and MGM_G176(MGM_W149,MGM_W148,MGM_W147);
   and MGM_G177(MGM_W150,si2_delay,MGM_W149);
   not MGM_G178(MGM_W151,ssb_delay);
   and MGM_G179(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W151,MGM_W150);
   not MGM_G180(MGM_W152,clk_delay);
   not MGM_G181(MGM_W153,d1_delay);
   and MGM_G182(MGM_W154,MGM_W153,MGM_W152);
   not MGM_G183(MGM_W155,d2_delay);
   and MGM_G184(MGM_W156,MGM_W155,MGM_W154);
   not MGM_G185(MGM_W157,si1_delay);
   and MGM_G186(MGM_W158,MGM_W157,MGM_W156);
   and MGM_G187(MGM_W159,si2_delay,MGM_W158);
   and MGM_G188(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W159);
   not MGM_G189(MGM_W160,clk_delay);
   not MGM_G190(MGM_W161,d1_delay);
   and MGM_G191(MGM_W162,MGM_W161,MGM_W160);
   not MGM_G192(MGM_W163,d2_delay);
   and MGM_G193(MGM_W164,MGM_W163,MGM_W162);
   and MGM_G194(MGM_W165,si1_delay,MGM_W164);
   not MGM_G195(MGM_W166,si2_delay);
   and MGM_G196(MGM_W167,MGM_W166,MGM_W165);
   not MGM_G197(MGM_W168,ssb_delay);
   and MGM_G198(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W168,MGM_W167);
   not MGM_G199(MGM_W169,clk_delay);
   not MGM_G200(MGM_W170,d1_delay);
   and MGM_G201(MGM_W171,MGM_W170,MGM_W169);
   not MGM_G202(MGM_W172,d2_delay);
   and MGM_G203(MGM_W173,MGM_W172,MGM_W171);
   and MGM_G204(MGM_W174,si1_delay,MGM_W173);
   not MGM_G205(MGM_W175,si2_delay);
   and MGM_G206(MGM_W176,MGM_W175,MGM_W174);
   and MGM_G207(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W176);
   not MGM_G208(MGM_W177,clk_delay);
   not MGM_G209(MGM_W178,d1_delay);
   and MGM_G210(MGM_W179,MGM_W178,MGM_W177);
   not MGM_G211(MGM_W180,d2_delay);
   and MGM_G212(MGM_W181,MGM_W180,MGM_W179);
   and MGM_G213(MGM_W182,si1_delay,MGM_W181);
   and MGM_G214(MGM_W183,si2_delay,MGM_W182);
   not MGM_G215(MGM_W184,ssb_delay);
   and MGM_G216(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W184,MGM_W183);
   not MGM_G217(MGM_W185,clk_delay);
   not MGM_G218(MGM_W186,d1_delay);
   and MGM_G219(MGM_W187,MGM_W186,MGM_W185);
   not MGM_G220(MGM_W188,d2_delay);
   and MGM_G221(MGM_W189,MGM_W188,MGM_W187);
   and MGM_G222(MGM_W190,si1_delay,MGM_W189);
   and MGM_G223(MGM_W191,si2_delay,MGM_W190);
   and MGM_G224(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W191);
   not MGM_G225(MGM_W192,clk_delay);
   not MGM_G226(MGM_W193,d1_delay);
   and MGM_G227(MGM_W194,MGM_W193,MGM_W192);
   and MGM_G228(MGM_W195,d2_delay,MGM_W194);
   not MGM_G229(MGM_W196,si1_delay);
   and MGM_G230(MGM_W197,MGM_W196,MGM_W195);
   not MGM_G231(MGM_W198,si2_delay);
   and MGM_G232(MGM_W199,MGM_W198,MGM_W197);
   not MGM_G233(MGM_W200,ssb_delay);
   and MGM_G234(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W200,MGM_W199);
   not MGM_G235(MGM_W201,clk_delay);
   not MGM_G236(MGM_W202,d1_delay);
   and MGM_G237(MGM_W203,MGM_W202,MGM_W201);
   and MGM_G238(MGM_W204,d2_delay,MGM_W203);
   not MGM_G239(MGM_W205,si1_delay);
   and MGM_G240(MGM_W206,MGM_W205,MGM_W204);
   not MGM_G241(MGM_W207,si2_delay);
   and MGM_G242(MGM_W208,MGM_W207,MGM_W206);
   and MGM_G243(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W208);
   not MGM_G244(MGM_W209,clk_delay);
   not MGM_G245(MGM_W210,d1_delay);
   and MGM_G246(MGM_W211,MGM_W210,MGM_W209);
   and MGM_G247(MGM_W212,d2_delay,MGM_W211);
   not MGM_G248(MGM_W213,si1_delay);
   and MGM_G249(MGM_W214,MGM_W213,MGM_W212);
   and MGM_G250(MGM_W215,si2_delay,MGM_W214);
   not MGM_G251(MGM_W216,ssb_delay);
   and MGM_G252(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W216,MGM_W215);
   not MGM_G253(MGM_W217,clk_delay);
   not MGM_G254(MGM_W218,d1_delay);
   and MGM_G255(MGM_W219,MGM_W218,MGM_W217);
   and MGM_G256(MGM_W220,d2_delay,MGM_W219);
   not MGM_G257(MGM_W221,si1_delay);
   and MGM_G258(MGM_W222,MGM_W221,MGM_W220);
   and MGM_G259(MGM_W223,si2_delay,MGM_W222);
   and MGM_G260(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W223);
   not MGM_G261(MGM_W224,clk_delay);
   not MGM_G262(MGM_W225,d1_delay);
   and MGM_G263(MGM_W226,MGM_W225,MGM_W224);
   and MGM_G264(MGM_W227,d2_delay,MGM_W226);
   and MGM_G265(MGM_W228,si1_delay,MGM_W227);
   not MGM_G266(MGM_W229,si2_delay);
   and MGM_G267(MGM_W230,MGM_W229,MGM_W228);
   not MGM_G268(MGM_W231,ssb_delay);
   and MGM_G269(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W231,MGM_W230);
   not MGM_G270(MGM_W232,clk_delay);
   not MGM_G271(MGM_W233,d1_delay);
   and MGM_G272(MGM_W234,MGM_W233,MGM_W232);
   and MGM_G273(MGM_W235,d2_delay,MGM_W234);
   and MGM_G274(MGM_W236,si1_delay,MGM_W235);
   not MGM_G275(MGM_W237,si2_delay);
   and MGM_G276(MGM_W238,MGM_W237,MGM_W236);
   and MGM_G277(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W238);
   not MGM_G278(MGM_W239,clk_delay);
   not MGM_G279(MGM_W240,d1_delay);
   and MGM_G280(MGM_W241,MGM_W240,MGM_W239);
   and MGM_G281(MGM_W242,d2_delay,MGM_W241);
   and MGM_G282(MGM_W243,si1_delay,MGM_W242);
   and MGM_G283(MGM_W244,si2_delay,MGM_W243);
   not MGM_G284(MGM_W245,ssb_delay);
   and MGM_G285(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W245,MGM_W244);
   not MGM_G286(MGM_W246,clk_delay);
   not MGM_G287(MGM_W247,d1_delay);
   and MGM_G288(MGM_W248,MGM_W247,MGM_W246);
   and MGM_G289(MGM_W249,d2_delay,MGM_W248);
   and MGM_G290(MGM_W250,si1_delay,MGM_W249);
   and MGM_G291(MGM_W251,si2_delay,MGM_W250);
   and MGM_G292(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W251);
   not MGM_G293(MGM_W252,clk_delay);
   and MGM_G294(MGM_W253,d1_delay,MGM_W252);
   not MGM_G295(MGM_W254,d2_delay);
   and MGM_G296(MGM_W255,MGM_W254,MGM_W253);
   not MGM_G297(MGM_W256,si1_delay);
   and MGM_G298(MGM_W257,MGM_W256,MGM_W255);
   not MGM_G299(MGM_W258,si2_delay);
   and MGM_G300(MGM_W259,MGM_W258,MGM_W257);
   not MGM_G301(MGM_W260,ssb_delay);
   and MGM_G302(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W260,MGM_W259);
   not MGM_G303(MGM_W261,clk_delay);
   and MGM_G304(MGM_W262,d1_delay,MGM_W261);
   not MGM_G305(MGM_W263,d2_delay);
   and MGM_G306(MGM_W264,MGM_W263,MGM_W262);
   not MGM_G307(MGM_W265,si1_delay);
   and MGM_G308(MGM_W266,MGM_W265,MGM_W264);
   not MGM_G309(MGM_W267,si2_delay);
   and MGM_G310(MGM_W268,MGM_W267,MGM_W266);
   and MGM_G311(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W268);
   not MGM_G312(MGM_W269,clk_delay);
   and MGM_G313(MGM_W270,d1_delay,MGM_W269);
   not MGM_G314(MGM_W271,d2_delay);
   and MGM_G315(MGM_W272,MGM_W271,MGM_W270);
   not MGM_G316(MGM_W273,si1_delay);
   and MGM_G317(MGM_W274,MGM_W273,MGM_W272);
   and MGM_G318(MGM_W275,si2_delay,MGM_W274);
   not MGM_G319(MGM_W276,ssb_delay);
   and MGM_G320(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W276,MGM_W275);
   not MGM_G321(MGM_W277,clk_delay);
   and MGM_G322(MGM_W278,d1_delay,MGM_W277);
   not MGM_G323(MGM_W279,d2_delay);
   and MGM_G324(MGM_W280,MGM_W279,MGM_W278);
   not MGM_G325(MGM_W281,si1_delay);
   and MGM_G326(MGM_W282,MGM_W281,MGM_W280);
   and MGM_G327(MGM_W283,si2_delay,MGM_W282);
   and MGM_G328(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W283);
   not MGM_G329(MGM_W284,clk_delay);
   and MGM_G330(MGM_W285,d1_delay,MGM_W284);
   not MGM_G331(MGM_W286,d2_delay);
   and MGM_G332(MGM_W287,MGM_W286,MGM_W285);
   and MGM_G333(MGM_W288,si1_delay,MGM_W287);
   not MGM_G334(MGM_W289,si2_delay);
   and MGM_G335(MGM_W290,MGM_W289,MGM_W288);
   not MGM_G336(MGM_W291,ssb_delay);
   and MGM_G337(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W291,MGM_W290);
   not MGM_G338(MGM_W292,clk_delay);
   and MGM_G339(MGM_W293,d1_delay,MGM_W292);
   not MGM_G340(MGM_W294,d2_delay);
   and MGM_G341(MGM_W295,MGM_W294,MGM_W293);
   and MGM_G342(MGM_W296,si1_delay,MGM_W295);
   not MGM_G343(MGM_W297,si2_delay);
   and MGM_G344(MGM_W298,MGM_W297,MGM_W296);
   and MGM_G345(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W298);
   not MGM_G346(MGM_W299,clk_delay);
   and MGM_G347(MGM_W300,d1_delay,MGM_W299);
   not MGM_G348(MGM_W301,d2_delay);
   and MGM_G349(MGM_W302,MGM_W301,MGM_W300);
   and MGM_G350(MGM_W303,si1_delay,MGM_W302);
   and MGM_G351(MGM_W304,si2_delay,MGM_W303);
   not MGM_G352(MGM_W305,ssb_delay);
   and MGM_G353(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W305,MGM_W304);
   not MGM_G354(MGM_W306,clk_delay);
   and MGM_G355(MGM_W307,d1_delay,MGM_W306);
   not MGM_G356(MGM_W308,d2_delay);
   and MGM_G357(MGM_W309,MGM_W308,MGM_W307);
   and MGM_G358(MGM_W310,si1_delay,MGM_W309);
   and MGM_G359(MGM_W311,si2_delay,MGM_W310);
   and MGM_G360(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W311);
   not MGM_G361(MGM_W312,clk_delay);
   and MGM_G362(MGM_W313,d1_delay,MGM_W312);
   and MGM_G363(MGM_W314,d2_delay,MGM_W313);
   not MGM_G364(MGM_W315,si1_delay);
   and MGM_G365(MGM_W316,MGM_W315,MGM_W314);
   not MGM_G366(MGM_W317,si2_delay);
   and MGM_G367(MGM_W318,MGM_W317,MGM_W316);
   not MGM_G368(MGM_W319,ssb_delay);
   and MGM_G369(ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W319,MGM_W318);
   not MGM_G370(MGM_W320,clk_delay);
   and MGM_G371(MGM_W321,d1_delay,MGM_W320);
   and MGM_G372(MGM_W322,d2_delay,MGM_W321);
   not MGM_G373(MGM_W323,si1_delay);
   and MGM_G374(MGM_W324,MGM_W323,MGM_W322);
   not MGM_G375(MGM_W325,si2_delay);
   and MGM_G376(MGM_W326,MGM_W325,MGM_W324);
   and MGM_G377(ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W326);
   not MGM_G378(MGM_W327,clk_delay);
   and MGM_G379(MGM_W328,d1_delay,MGM_W327);
   and MGM_G380(MGM_W329,d2_delay,MGM_W328);
   not MGM_G381(MGM_W330,si1_delay);
   and MGM_G382(MGM_W331,MGM_W330,MGM_W329);
   and MGM_G383(MGM_W332,si2_delay,MGM_W331);
   not MGM_G384(MGM_W333,ssb_delay);
   and MGM_G385(ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W333,MGM_W332);
   not MGM_G386(MGM_W334,clk_delay);
   and MGM_G387(MGM_W335,d1_delay,MGM_W334);
   and MGM_G388(MGM_W336,d2_delay,MGM_W335);
   not MGM_G389(MGM_W337,si1_delay);
   and MGM_G390(MGM_W338,MGM_W337,MGM_W336);
   and MGM_G391(MGM_W339,si2_delay,MGM_W338);
   and MGM_G392(ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W339);
   not MGM_G393(MGM_W340,clk_delay);
   and MGM_G394(MGM_W341,d1_delay,MGM_W340);
   and MGM_G395(MGM_W342,d2_delay,MGM_W341);
   and MGM_G396(MGM_W343,si1_delay,MGM_W342);
   not MGM_G397(MGM_W344,si2_delay);
   and MGM_G398(MGM_W345,MGM_W344,MGM_W343);
   not MGM_G399(MGM_W346,ssb_delay);
   and MGM_G400(ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W346,MGM_W345);
   not MGM_G401(MGM_W347,clk_delay);
   and MGM_G402(MGM_W348,d1_delay,MGM_W347);
   and MGM_G403(MGM_W349,d2_delay,MGM_W348);
   and MGM_G404(MGM_W350,si1_delay,MGM_W349);
   not MGM_G405(MGM_W351,si2_delay);
   and MGM_G406(MGM_W352,MGM_W351,MGM_W350);
   and MGM_G407(ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W352);
   not MGM_G408(MGM_W353,clk_delay);
   and MGM_G409(MGM_W354,d1_delay,MGM_W353);
   and MGM_G410(MGM_W355,d2_delay,MGM_W354);
   and MGM_G411(MGM_W356,si1_delay,MGM_W355);
   and MGM_G412(MGM_W357,si2_delay,MGM_W356);
   not MGM_G413(MGM_W358,ssb_delay);
   and MGM_G414(ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W358,MGM_W357);
   not MGM_G415(MGM_W359,clk_delay);
   and MGM_G416(MGM_W360,d1_delay,MGM_W359);
   and MGM_G417(MGM_W361,d2_delay,MGM_W360);
   and MGM_G418(MGM_W362,si1_delay,MGM_W361);
   and MGM_G419(MGM_W363,si2_delay,MGM_W362);
   and MGM_G420(ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W363);
   not MGM_G421(MGM_W364,d1_delay);
   and MGM_G422(MGM_W365,MGM_W364,clk_delay);
   not MGM_G423(MGM_W366,d2_delay);
   and MGM_G424(MGM_W367,MGM_W366,MGM_W365);
   not MGM_G425(MGM_W368,si1_delay);
   and MGM_G426(MGM_W369,MGM_W368,MGM_W367);
   not MGM_G427(MGM_W370,si2_delay);
   and MGM_G428(MGM_W371,MGM_W370,MGM_W369);
   not MGM_G429(MGM_W372,ssb_delay);
   and MGM_G430(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W372,MGM_W371);
   not MGM_G431(MGM_W373,d1_delay);
   and MGM_G432(MGM_W374,MGM_W373,clk_delay);
   not MGM_G433(MGM_W375,d2_delay);
   and MGM_G434(MGM_W376,MGM_W375,MGM_W374);
   not MGM_G435(MGM_W377,si1_delay);
   and MGM_G436(MGM_W378,MGM_W377,MGM_W376);
   not MGM_G437(MGM_W379,si2_delay);
   and MGM_G438(MGM_W380,MGM_W379,MGM_W378);
   and MGM_G439(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W380);
   not MGM_G440(MGM_W381,d1_delay);
   and MGM_G441(MGM_W382,MGM_W381,clk_delay);
   not MGM_G442(MGM_W383,d2_delay);
   and MGM_G443(MGM_W384,MGM_W383,MGM_W382);
   not MGM_G444(MGM_W385,si1_delay);
   and MGM_G445(MGM_W386,MGM_W385,MGM_W384);
   and MGM_G446(MGM_W387,si2_delay,MGM_W386);
   not MGM_G447(MGM_W388,ssb_delay);
   and MGM_G448(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W388,MGM_W387);
   not MGM_G449(MGM_W389,d1_delay);
   and MGM_G450(MGM_W390,MGM_W389,clk_delay);
   not MGM_G451(MGM_W391,d2_delay);
   and MGM_G452(MGM_W392,MGM_W391,MGM_W390);
   not MGM_G453(MGM_W393,si1_delay);
   and MGM_G454(MGM_W394,MGM_W393,MGM_W392);
   and MGM_G455(MGM_W395,si2_delay,MGM_W394);
   and MGM_G456(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W395);
   not MGM_G457(MGM_W396,d1_delay);
   and MGM_G458(MGM_W397,MGM_W396,clk_delay);
   not MGM_G459(MGM_W398,d2_delay);
   and MGM_G460(MGM_W399,MGM_W398,MGM_W397);
   and MGM_G461(MGM_W400,si1_delay,MGM_W399);
   not MGM_G462(MGM_W401,si2_delay);
   and MGM_G463(MGM_W402,MGM_W401,MGM_W400);
   not MGM_G464(MGM_W403,ssb_delay);
   and MGM_G465(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W403,MGM_W402);
   not MGM_G466(MGM_W404,d1_delay);
   and MGM_G467(MGM_W405,MGM_W404,clk_delay);
   not MGM_G468(MGM_W406,d2_delay);
   and MGM_G469(MGM_W407,MGM_W406,MGM_W405);
   and MGM_G470(MGM_W408,si1_delay,MGM_W407);
   not MGM_G471(MGM_W409,si2_delay);
   and MGM_G472(MGM_W410,MGM_W409,MGM_W408);
   and MGM_G473(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W410);
   not MGM_G474(MGM_W411,d1_delay);
   and MGM_G475(MGM_W412,MGM_W411,clk_delay);
   not MGM_G476(MGM_W413,d2_delay);
   and MGM_G477(MGM_W414,MGM_W413,MGM_W412);
   and MGM_G478(MGM_W415,si1_delay,MGM_W414);
   and MGM_G479(MGM_W416,si2_delay,MGM_W415);
   not MGM_G480(MGM_W417,ssb_delay);
   and MGM_G481(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W417,MGM_W416);
   not MGM_G482(MGM_W418,d1_delay);
   and MGM_G483(MGM_W419,MGM_W418,clk_delay);
   not MGM_G484(MGM_W420,d2_delay);
   and MGM_G485(MGM_W421,MGM_W420,MGM_W419);
   and MGM_G486(MGM_W422,si1_delay,MGM_W421);
   and MGM_G487(MGM_W423,si2_delay,MGM_W422);
   and MGM_G488(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W423);
   not MGM_G489(MGM_W424,d1_delay);
   and MGM_G490(MGM_W425,MGM_W424,clk_delay);
   and MGM_G491(MGM_W426,d2_delay,MGM_W425);
   not MGM_G492(MGM_W427,si1_delay);
   and MGM_G493(MGM_W428,MGM_W427,MGM_W426);
   not MGM_G494(MGM_W429,si2_delay);
   and MGM_G495(MGM_W430,MGM_W429,MGM_W428);
   not MGM_G496(MGM_W431,ssb_delay);
   and MGM_G497(ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W431,MGM_W430);
   not MGM_G498(MGM_W432,d1_delay);
   and MGM_G499(MGM_W433,MGM_W432,clk_delay);
   and MGM_G500(MGM_W434,d2_delay,MGM_W433);
   not MGM_G501(MGM_W435,si1_delay);
   and MGM_G502(MGM_W436,MGM_W435,MGM_W434);
   not MGM_G503(MGM_W437,si2_delay);
   and MGM_G504(MGM_W438,MGM_W437,MGM_W436);
   and MGM_G505(ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W438);
   not MGM_G506(MGM_W439,d1_delay);
   and MGM_G507(MGM_W440,MGM_W439,clk_delay);
   and MGM_G508(MGM_W441,d2_delay,MGM_W440);
   not MGM_G509(MGM_W442,si1_delay);
   and MGM_G510(MGM_W443,MGM_W442,MGM_W441);
   and MGM_G511(MGM_W444,si2_delay,MGM_W443);
   not MGM_G512(MGM_W445,ssb_delay);
   and MGM_G513(ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W445,MGM_W444);
   not MGM_G514(MGM_W446,d1_delay);
   and MGM_G515(MGM_W447,MGM_W446,clk_delay);
   and MGM_G516(MGM_W448,d2_delay,MGM_W447);
   not MGM_G517(MGM_W449,si1_delay);
   and MGM_G518(MGM_W450,MGM_W449,MGM_W448);
   and MGM_G519(MGM_W451,si2_delay,MGM_W450);
   and MGM_G520(ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W451);
   not MGM_G521(MGM_W452,d1_delay);
   and MGM_G522(MGM_W453,MGM_W452,clk_delay);
   and MGM_G523(MGM_W454,d2_delay,MGM_W453);
   and MGM_G524(MGM_W455,si1_delay,MGM_W454);
   not MGM_G525(MGM_W456,si2_delay);
   and MGM_G526(MGM_W457,MGM_W456,MGM_W455);
   not MGM_G527(MGM_W458,ssb_delay);
   and MGM_G528(ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W458,MGM_W457);
   not MGM_G529(MGM_W459,d1_delay);
   and MGM_G530(MGM_W460,MGM_W459,clk_delay);
   and MGM_G531(MGM_W461,d2_delay,MGM_W460);
   and MGM_G532(MGM_W462,si1_delay,MGM_W461);
   not MGM_G533(MGM_W463,si2_delay);
   and MGM_G534(MGM_W464,MGM_W463,MGM_W462);
   and MGM_G535(ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W464);
   not MGM_G536(MGM_W465,d1_delay);
   and MGM_G537(MGM_W466,MGM_W465,clk_delay);
   and MGM_G538(MGM_W467,d2_delay,MGM_W466);
   and MGM_G539(MGM_W468,si1_delay,MGM_W467);
   and MGM_G540(MGM_W469,si2_delay,MGM_W468);
   not MGM_G541(MGM_W470,ssb_delay);
   and MGM_G542(ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W470,MGM_W469);
   not MGM_G543(MGM_W471,d1_delay);
   and MGM_G544(MGM_W472,MGM_W471,clk_delay);
   and MGM_G545(MGM_W473,d2_delay,MGM_W472);
   and MGM_G546(MGM_W474,si1_delay,MGM_W473);
   and MGM_G547(MGM_W475,si2_delay,MGM_W474);
   and MGM_G548(ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W475);
   and MGM_G549(MGM_W476,d1_delay,clk_delay);
   not MGM_G550(MGM_W477,d2_delay);
   and MGM_G551(MGM_W478,MGM_W477,MGM_W476);
   not MGM_G552(MGM_W479,si1_delay);
   and MGM_G553(MGM_W480,MGM_W479,MGM_W478);
   not MGM_G554(MGM_W481,si2_delay);
   and MGM_G555(MGM_W482,MGM_W481,MGM_W480);
   not MGM_G556(MGM_W483,ssb_delay);
   and MGM_G557(ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W483,MGM_W482);
   and MGM_G558(MGM_W484,d1_delay,clk_delay);
   not MGM_G559(MGM_W485,d2_delay);
   and MGM_G560(MGM_W486,MGM_W485,MGM_W484);
   not MGM_G561(MGM_W487,si1_delay);
   and MGM_G562(MGM_W488,MGM_W487,MGM_W486);
   not MGM_G563(MGM_W489,si2_delay);
   and MGM_G564(MGM_W490,MGM_W489,MGM_W488);
   and MGM_G565(ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W490);
   and MGM_G566(MGM_W491,d1_delay,clk_delay);
   not MGM_G567(MGM_W492,d2_delay);
   and MGM_G568(MGM_W493,MGM_W492,MGM_W491);
   not MGM_G569(MGM_W494,si1_delay);
   and MGM_G570(MGM_W495,MGM_W494,MGM_W493);
   and MGM_G571(MGM_W496,si2_delay,MGM_W495);
   not MGM_G572(MGM_W497,ssb_delay);
   and MGM_G573(ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W497,MGM_W496);
   and MGM_G574(MGM_W498,d1_delay,clk_delay);
   not MGM_G575(MGM_W499,d2_delay);
   and MGM_G576(MGM_W500,MGM_W499,MGM_W498);
   not MGM_G577(MGM_W501,si1_delay);
   and MGM_G578(MGM_W502,MGM_W501,MGM_W500);
   and MGM_G579(MGM_W503,si2_delay,MGM_W502);
   and MGM_G580(ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W503);
   and MGM_G581(MGM_W504,d1_delay,clk_delay);
   not MGM_G582(MGM_W505,d2_delay);
   and MGM_G583(MGM_W506,MGM_W505,MGM_W504);
   and MGM_G584(MGM_W507,si1_delay,MGM_W506);
   not MGM_G585(MGM_W508,si2_delay);
   and MGM_G586(MGM_W509,MGM_W508,MGM_W507);
   not MGM_G587(MGM_W510,ssb_delay);
   and MGM_G588(ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W510,MGM_W509);
   and MGM_G589(MGM_W511,d1_delay,clk_delay);
   not MGM_G590(MGM_W512,d2_delay);
   and MGM_G591(MGM_W513,MGM_W512,MGM_W511);
   and MGM_G592(MGM_W514,si1_delay,MGM_W513);
   not MGM_G593(MGM_W515,si2_delay);
   and MGM_G594(MGM_W516,MGM_W515,MGM_W514);
   and MGM_G595(ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W516);
   and MGM_G596(MGM_W517,d1_delay,clk_delay);
   not MGM_G597(MGM_W518,d2_delay);
   and MGM_G598(MGM_W519,MGM_W518,MGM_W517);
   and MGM_G599(MGM_W520,si1_delay,MGM_W519);
   and MGM_G600(MGM_W521,si2_delay,MGM_W520);
   not MGM_G601(MGM_W522,ssb_delay);
   and MGM_G602(ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W522,MGM_W521);
   and MGM_G603(MGM_W523,d1_delay,clk_delay);
   not MGM_G604(MGM_W524,d2_delay);
   and MGM_G605(MGM_W525,MGM_W524,MGM_W523);
   and MGM_G606(MGM_W526,si1_delay,MGM_W525);
   and MGM_G607(MGM_W527,si2_delay,MGM_W526);
   and MGM_G608(ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W527);
   and MGM_G609(MGM_W528,d1_delay,clk_delay);
   and MGM_G610(MGM_W529,d2_delay,MGM_W528);
   not MGM_G611(MGM_W530,si1_delay);
   and MGM_G612(MGM_W531,MGM_W530,MGM_W529);
   not MGM_G613(MGM_W532,si2_delay);
   and MGM_G614(MGM_W533,MGM_W532,MGM_W531);
   not MGM_G615(MGM_W534,ssb_delay);
   and MGM_G616(ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W534,MGM_W533);
   and MGM_G617(MGM_W535,d1_delay,clk_delay);
   and MGM_G618(MGM_W536,d2_delay,MGM_W535);
   not MGM_G619(MGM_W537,si1_delay);
   and MGM_G620(MGM_W538,MGM_W537,MGM_W536);
   not MGM_G621(MGM_W539,si2_delay);
   and MGM_G622(MGM_W540,MGM_W539,MGM_W538);
   and MGM_G623(ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W540);
   and MGM_G624(MGM_W541,d1_delay,clk_delay);
   and MGM_G625(MGM_W542,d2_delay,MGM_W541);
   not MGM_G626(MGM_W543,si1_delay);
   and MGM_G627(MGM_W544,MGM_W543,MGM_W542);
   and MGM_G628(MGM_W545,si2_delay,MGM_W544);
   not MGM_G629(MGM_W546,ssb_delay);
   and MGM_G630(ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W546,MGM_W545);
   and MGM_G631(MGM_W547,d1_delay,clk_delay);
   and MGM_G632(MGM_W548,d2_delay,MGM_W547);
   not MGM_G633(MGM_W549,si1_delay);
   and MGM_G634(MGM_W550,MGM_W549,MGM_W548);
   and MGM_G635(MGM_W551,si2_delay,MGM_W550);
   and MGM_G636(ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W551);
   and MGM_G637(MGM_W552,d1_delay,clk_delay);
   and MGM_G638(MGM_W553,d2_delay,MGM_W552);
   and MGM_G639(MGM_W554,si1_delay,MGM_W553);
   not MGM_G640(MGM_W555,si2_delay);
   and MGM_G641(MGM_W556,MGM_W555,MGM_W554);
   not MGM_G642(MGM_W557,ssb_delay);
   and MGM_G643(ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W557,MGM_W556);
   and MGM_G644(MGM_W558,d1_delay,clk_delay);
   and MGM_G645(MGM_W559,d2_delay,MGM_W558);
   and MGM_G646(MGM_W560,si1_delay,MGM_W559);
   not MGM_G647(MGM_W561,si2_delay);
   and MGM_G648(MGM_W562,MGM_W561,MGM_W560);
   and MGM_G649(ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W562);
   and MGM_G650(MGM_W563,d1_delay,clk_delay);
   and MGM_G651(MGM_W564,d2_delay,MGM_W563);
   and MGM_G652(MGM_W565,si1_delay,MGM_W564);
   and MGM_G653(MGM_W566,si2_delay,MGM_W565);
   not MGM_G654(MGM_W567,ssb_delay);
   and MGM_G655(ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W567,MGM_W566);
   and MGM_G656(MGM_W568,d1_delay,clk_delay);
   and MGM_G657(MGM_W569,d2_delay,MGM_W568);
   and MGM_G658(MGM_W570,si1_delay,MGM_W569);
   and MGM_G659(MGM_W571,si2_delay,MGM_W570);
   and MGM_G660(ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W571);
   not MGM_G661(MGM_W572,d1_delay);
   not MGM_G662(MGM_W573,d2_delay);
   and MGM_G663(MGM_W574,MGM_W573,MGM_W572);
   and MGM_G664(MGM_W575,rb_delay,MGM_W574);
   not MGM_G665(MGM_W576,si1_delay);
   and MGM_G666(MGM_W577,MGM_W576,MGM_W575);
   and MGM_G667(ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2,si2_delay,MGM_W577);
   not MGM_G668(MGM_W578,d1_delay);
   not MGM_G669(MGM_W579,d2_delay);
   and MGM_G670(MGM_W580,MGM_W579,MGM_W578);
   and MGM_G671(MGM_W581,rb_delay,MGM_W580);
   and MGM_G672(MGM_W582,si1_delay,MGM_W581);
   not MGM_G673(MGM_W583,si2_delay);
   and MGM_G674(ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2,MGM_W583,MGM_W582);
   not MGM_G675(MGM_W584,d1_delay);
   not MGM_G676(MGM_W585,d2_delay);
   and MGM_G677(MGM_W586,MGM_W585,MGM_W584);
   and MGM_G678(MGM_W587,rb_delay,MGM_W586);
   and MGM_G679(MGM_W588,si1_delay,MGM_W587);
   and MGM_G680(ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2,si2_delay,MGM_W588);
   not MGM_G681(MGM_W589,d1_delay);
   and MGM_G682(MGM_W590,d2_delay,MGM_W589);
   and MGM_G683(MGM_W591,rb_delay,MGM_W590);
   not MGM_G684(MGM_W592,si1_delay);
   and MGM_G685(MGM_W593,MGM_W592,MGM_W591);
   not MGM_G686(MGM_W594,si2_delay);
   and MGM_G687(ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2,MGM_W594,MGM_W593);
   not MGM_G688(MGM_W595,d1_delay);
   and MGM_G689(MGM_W596,d2_delay,MGM_W595);
   and MGM_G690(MGM_W597,rb_delay,MGM_W596);
   and MGM_G691(MGM_W598,si1_delay,MGM_W597);
   not MGM_G692(MGM_W599,si2_delay);
   and MGM_G693(ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2,MGM_W599,MGM_W598);
   not MGM_G694(MGM_W600,d1_delay);
   and MGM_G695(MGM_W601,d2_delay,MGM_W600);
   and MGM_G696(MGM_W602,rb_delay,MGM_W601);
   and MGM_G697(MGM_W603,si1_delay,MGM_W602);
   and MGM_G698(ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2,si2_delay,MGM_W603);
   not MGM_G699(MGM_W604,d2_delay);
   and MGM_G700(MGM_W605,MGM_W604,d1_delay);
   and MGM_G701(MGM_W606,rb_delay,MGM_W605);
   not MGM_G702(MGM_W607,si1_delay);
   and MGM_G703(MGM_W608,MGM_W607,MGM_W606);
   not MGM_G704(MGM_W609,si2_delay);
   and MGM_G705(ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2,MGM_W609,MGM_W608);
   not MGM_G706(MGM_W610,d2_delay);
   and MGM_G707(MGM_W611,MGM_W610,d1_delay);
   and MGM_G708(MGM_W612,rb_delay,MGM_W611);
   not MGM_G709(MGM_W613,si1_delay);
   and MGM_G710(MGM_W614,MGM_W613,MGM_W612);
   and MGM_G711(ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2,si2_delay,MGM_W614);
   not MGM_G712(MGM_W615,d2_delay);
   and MGM_G713(MGM_W616,MGM_W615,d1_delay);
   and MGM_G714(MGM_W617,rb_delay,MGM_W616);
   and MGM_G715(MGM_W618,si1_delay,MGM_W617);
   and MGM_G716(ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2,si2_delay,MGM_W618);
   and MGM_G717(MGM_W619,d2_delay,d1_delay);
   and MGM_G718(MGM_W620,rb_delay,MGM_W619);
   not MGM_G719(MGM_W621,si1_delay);
   and MGM_G720(MGM_W622,MGM_W621,MGM_W620);
   not MGM_G721(MGM_W623,si2_delay);
   and MGM_G722(ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2,MGM_W623,MGM_W622);
   and MGM_G723(MGM_W624,d2_delay,d1_delay);
   and MGM_G724(MGM_W625,rb_delay,MGM_W624);
   not MGM_G725(MGM_W626,si1_delay);
   and MGM_G726(MGM_W627,MGM_W626,MGM_W625);
   and MGM_G727(ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2,si2_delay,MGM_W627);
   and MGM_G728(MGM_W628,d2_delay,d1_delay);
   and MGM_G729(MGM_W629,rb_delay,MGM_W628);
   and MGM_G730(MGM_W630,si1_delay,MGM_W629);
   not MGM_G731(MGM_W631,si2_delay);
   and MGM_G732(ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2,MGM_W631,MGM_W630);
   and MGM_G733(ENABLE_ssb_AND_rb,rb_delay,ssb_delay);
   not MGM_G734(MGM_W632,ssb_delay);
   and MGM_G735(ENABLE_NOT_ssb_AND_rb,rb_delay,MGM_W632);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d1==1'b0 && rb==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_rb == 1'b1)
      ,0.0,0,notifier);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb,0.0,0,notifier);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,negedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,posedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d1 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d1 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d2 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d2 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si1 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si1 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si2 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si2 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy203ah1n04x5( clk, d1, d2, o1, o2, rb, si1, si2, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, rb, si1, si2, ssb;
   output o1, o2;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy203ah_func b15fqy203ah1n04x5_behav_inst(.clk(clk),.rb(rb),.ssb(ssb),.o1(o1),.o2(o2),.d1(d1),.d2(d2),.si1(si1),.si2(si2),.notifier0(1'b0),.notifier1(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy203ah_func b15fqy203ah1n04x5_behav_inst(.clk(clk),.rb(rb),.ssb(ssb),.o1(o1),.o2(o2),.d1(d1),.d2(d2),.si1(si1),.si2(si2),.notifier0(1'b0),.notifier1(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire rb_delay ;
   wire ssb_delay ;
   wire d1_delay ;
   wire d2_delay ;
   wire si1_delay ;
   wire si2_delay ;
   reg notifier;
   reg notifier0;
   reg notifier1;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
     notifier1 = (notifier1 !== notifier) ? notifier : ~notifier1;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy203ah_func b15fqy203ah1n04x5_inst(.clk(clk_delay),.rb(rb_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.d1(d1_delay),.d2(d2_delay),.si1(si1_delay),.si2(si2_delay),.notifier0(notifier0),.notifier1(notifier1),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy203ah_func b15fqy203ah1n04x5_inst(.clk(clk_delay),.rb(rb_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.d1(d1_delay),.d2(d2_delay),.si1(si1_delay),.si2(si2_delay),.notifier0(notifier0),.notifier1(notifier1));
   `endif
   
   // spec_gates_begin
   buf MGM_G0(ENABLE_rb,rb_delay);
   not MGM_G1(MGM_W0,d1_delay);
   not MGM_G2(MGM_W1,d2_delay);
   and MGM_G3(MGM_W2,MGM_W1,MGM_W0);
   not MGM_G4(MGM_W3,si1_delay);
   and MGM_G5(MGM_W4,MGM_W3,MGM_W2);
   and MGM_G6(MGM_W5,si2_delay,MGM_W4);
   not MGM_G7(MGM_W6,ssb_delay);
   and MGM_G8(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W6,MGM_W5);
   not MGM_G9(MGM_W7,d1_delay);
   not MGM_G10(MGM_W8,d2_delay);
   and MGM_G11(MGM_W9,MGM_W8,MGM_W7);
   and MGM_G12(MGM_W10,si1_delay,MGM_W9);
   not MGM_G13(MGM_W11,si2_delay);
   and MGM_G14(MGM_W12,MGM_W11,MGM_W10);
   not MGM_G15(MGM_W13,ssb_delay);
   and MGM_G16(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W13,MGM_W12);
   not MGM_G17(MGM_W14,d1_delay);
   not MGM_G18(MGM_W15,d2_delay);
   and MGM_G19(MGM_W16,MGM_W15,MGM_W14);
   and MGM_G20(MGM_W17,si1_delay,MGM_W16);
   and MGM_G21(MGM_W18,si2_delay,MGM_W17);
   not MGM_G22(MGM_W19,ssb_delay);
   and MGM_G23(ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W19,MGM_W18);
   not MGM_G24(MGM_W20,d1_delay);
   and MGM_G25(MGM_W21,d2_delay,MGM_W20);
   not MGM_G26(MGM_W22,si1_delay);
   and MGM_G27(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G28(MGM_W24,si2_delay);
   and MGM_G29(MGM_W25,MGM_W24,MGM_W23);
   and MGM_G30(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W25);
   not MGM_G31(MGM_W26,d1_delay);
   and MGM_G32(MGM_W27,d2_delay,MGM_W26);
   not MGM_G33(MGM_W28,si1_delay);
   and MGM_G34(MGM_W29,MGM_W28,MGM_W27);
   and MGM_G35(MGM_W30,si2_delay,MGM_W29);
   not MGM_G36(MGM_W31,ssb_delay);
   and MGM_G37(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W31,MGM_W30);
   not MGM_G38(MGM_W32,d1_delay);
   and MGM_G39(MGM_W33,d2_delay,MGM_W32);
   not MGM_G40(MGM_W34,si1_delay);
   and MGM_G41(MGM_W35,MGM_W34,MGM_W33);
   and MGM_G42(MGM_W36,si2_delay,MGM_W35);
   and MGM_G43(ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W36);
   not MGM_G44(MGM_W37,d1_delay);
   and MGM_G45(MGM_W38,d2_delay,MGM_W37);
   and MGM_G46(MGM_W39,si1_delay,MGM_W38);
   not MGM_G47(MGM_W40,si2_delay);
   and MGM_G48(MGM_W41,MGM_W40,MGM_W39);
   not MGM_G49(MGM_W42,ssb_delay);
   and MGM_G50(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W42,MGM_W41);
   not MGM_G51(MGM_W43,d1_delay);
   and MGM_G52(MGM_W44,d2_delay,MGM_W43);
   and MGM_G53(MGM_W45,si1_delay,MGM_W44);
   not MGM_G54(MGM_W46,si2_delay);
   and MGM_G55(MGM_W47,MGM_W46,MGM_W45);
   and MGM_G56(ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W47);
   not MGM_G57(MGM_W48,d1_delay);
   and MGM_G58(MGM_W49,d2_delay,MGM_W48);
   and MGM_G59(MGM_W50,si1_delay,MGM_W49);
   and MGM_G60(MGM_W51,si2_delay,MGM_W50);
   not MGM_G61(MGM_W52,ssb_delay);
   and MGM_G62(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W52,MGM_W51);
   not MGM_G63(MGM_W53,d1_delay);
   and MGM_G64(MGM_W54,d2_delay,MGM_W53);
   and MGM_G65(MGM_W55,si1_delay,MGM_W54);
   and MGM_G66(MGM_W56,si2_delay,MGM_W55);
   and MGM_G67(ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W56);
   not MGM_G68(MGM_W57,d2_delay);
   and MGM_G69(MGM_W58,MGM_W57,d1_delay);
   not MGM_G70(MGM_W59,si1_delay);
   and MGM_G71(MGM_W60,MGM_W59,MGM_W58);
   not MGM_G72(MGM_W61,si2_delay);
   and MGM_G73(MGM_W62,MGM_W61,MGM_W60);
   and MGM_G74(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W62);
   not MGM_G75(MGM_W63,d2_delay);
   and MGM_G76(MGM_W64,MGM_W63,d1_delay);
   not MGM_G77(MGM_W65,si1_delay);
   and MGM_G78(MGM_W66,MGM_W65,MGM_W64);
   and MGM_G79(MGM_W67,si2_delay,MGM_W66);
   not MGM_G80(MGM_W68,ssb_delay);
   and MGM_G81(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W68,MGM_W67);
   not MGM_G82(MGM_W69,d2_delay);
   and MGM_G83(MGM_W70,MGM_W69,d1_delay);
   not MGM_G84(MGM_W71,si1_delay);
   and MGM_G85(MGM_W72,MGM_W71,MGM_W70);
   and MGM_G86(MGM_W73,si2_delay,MGM_W72);
   and MGM_G87(ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W73);
   not MGM_G88(MGM_W74,d2_delay);
   and MGM_G89(MGM_W75,MGM_W74,d1_delay);
   and MGM_G90(MGM_W76,si1_delay,MGM_W75);
   not MGM_G91(MGM_W77,si2_delay);
   and MGM_G92(MGM_W78,MGM_W77,MGM_W76);
   not MGM_G93(MGM_W79,ssb_delay);
   and MGM_G94(ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W79,MGM_W78);
   not MGM_G95(MGM_W80,d2_delay);
   and MGM_G96(MGM_W81,MGM_W80,d1_delay);
   and MGM_G97(MGM_W82,si1_delay,MGM_W81);
   not MGM_G98(MGM_W83,si2_delay);
   and MGM_G99(MGM_W84,MGM_W83,MGM_W82);
   and MGM_G100(ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W84);
   not MGM_G101(MGM_W85,d2_delay);
   and MGM_G102(MGM_W86,MGM_W85,d1_delay);
   and MGM_G103(MGM_W87,si1_delay,MGM_W86);
   and MGM_G104(MGM_W88,si2_delay,MGM_W87);
   not MGM_G105(MGM_W89,ssb_delay);
   and MGM_G106(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W89,MGM_W88);
   not MGM_G107(MGM_W90,d2_delay);
   and MGM_G108(MGM_W91,MGM_W90,d1_delay);
   and MGM_G109(MGM_W92,si1_delay,MGM_W91);
   and MGM_G110(MGM_W93,si2_delay,MGM_W92);
   and MGM_G111(ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W93);
   and MGM_G112(MGM_W94,d2_delay,d1_delay);
   not MGM_G113(MGM_W95,si1_delay);
   and MGM_G114(MGM_W96,MGM_W95,MGM_W94);
   not MGM_G115(MGM_W97,si2_delay);
   and MGM_G116(MGM_W98,MGM_W97,MGM_W96);
   and MGM_G117(ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W98);
   and MGM_G118(MGM_W99,d2_delay,d1_delay);
   not MGM_G119(MGM_W100,si1_delay);
   and MGM_G120(MGM_W101,MGM_W100,MGM_W99);
   and MGM_G121(MGM_W102,si2_delay,MGM_W101);
   not MGM_G122(MGM_W103,ssb_delay);
   and MGM_G123(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W103,MGM_W102);
   and MGM_G124(MGM_W104,d2_delay,d1_delay);
   not MGM_G125(MGM_W105,si1_delay);
   and MGM_G126(MGM_W106,MGM_W105,MGM_W104);
   and MGM_G127(MGM_W107,si2_delay,MGM_W106);
   and MGM_G128(ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W107);
   and MGM_G129(MGM_W108,d2_delay,d1_delay);
   and MGM_G130(MGM_W109,si1_delay,MGM_W108);
   not MGM_G131(MGM_W110,si2_delay);
   and MGM_G132(MGM_W111,MGM_W110,MGM_W109);
   not MGM_G133(MGM_W112,ssb_delay);
   and MGM_G134(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W112,MGM_W111);
   and MGM_G135(MGM_W113,d2_delay,d1_delay);
   and MGM_G136(MGM_W114,si1_delay,MGM_W113);
   not MGM_G137(MGM_W115,si2_delay);
   and MGM_G138(MGM_W116,MGM_W115,MGM_W114);
   and MGM_G139(ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W116);
   and MGM_G140(MGM_W117,d2_delay,d1_delay);
   and MGM_G141(MGM_W118,si1_delay,MGM_W117);
   and MGM_G142(MGM_W119,si2_delay,MGM_W118);
   not MGM_G143(MGM_W120,ssb_delay);
   and MGM_G144(ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W120,MGM_W119);
   and MGM_G145(MGM_W121,d2_delay,d1_delay);
   and MGM_G146(MGM_W122,si1_delay,MGM_W121);
   and MGM_G147(MGM_W123,si2_delay,MGM_W122);
   and MGM_G148(ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W123);
   not MGM_G149(MGM_W124,clk_delay);
   not MGM_G150(MGM_W125,d1_delay);
   and MGM_G151(MGM_W126,MGM_W125,MGM_W124);
   not MGM_G152(MGM_W127,d2_delay);
   and MGM_G153(MGM_W128,MGM_W127,MGM_W126);
   not MGM_G154(MGM_W129,si1_delay);
   and MGM_G155(MGM_W130,MGM_W129,MGM_W128);
   not MGM_G156(MGM_W131,si2_delay);
   and MGM_G157(MGM_W132,MGM_W131,MGM_W130);
   not MGM_G158(MGM_W133,ssb_delay);
   and MGM_G159(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W133,MGM_W132);
   not MGM_G160(MGM_W134,clk_delay);
   not MGM_G161(MGM_W135,d1_delay);
   and MGM_G162(MGM_W136,MGM_W135,MGM_W134);
   not MGM_G163(MGM_W137,d2_delay);
   and MGM_G164(MGM_W138,MGM_W137,MGM_W136);
   not MGM_G165(MGM_W139,si1_delay);
   and MGM_G166(MGM_W140,MGM_W139,MGM_W138);
   not MGM_G167(MGM_W141,si2_delay);
   and MGM_G168(MGM_W142,MGM_W141,MGM_W140);
   and MGM_G169(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W142);
   not MGM_G170(MGM_W143,clk_delay);
   not MGM_G171(MGM_W144,d1_delay);
   and MGM_G172(MGM_W145,MGM_W144,MGM_W143);
   not MGM_G173(MGM_W146,d2_delay);
   and MGM_G174(MGM_W147,MGM_W146,MGM_W145);
   not MGM_G175(MGM_W148,si1_delay);
   and MGM_G176(MGM_W149,MGM_W148,MGM_W147);
   and MGM_G177(MGM_W150,si2_delay,MGM_W149);
   not MGM_G178(MGM_W151,ssb_delay);
   and MGM_G179(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W151,MGM_W150);
   not MGM_G180(MGM_W152,clk_delay);
   not MGM_G181(MGM_W153,d1_delay);
   and MGM_G182(MGM_W154,MGM_W153,MGM_W152);
   not MGM_G183(MGM_W155,d2_delay);
   and MGM_G184(MGM_W156,MGM_W155,MGM_W154);
   not MGM_G185(MGM_W157,si1_delay);
   and MGM_G186(MGM_W158,MGM_W157,MGM_W156);
   and MGM_G187(MGM_W159,si2_delay,MGM_W158);
   and MGM_G188(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W159);
   not MGM_G189(MGM_W160,clk_delay);
   not MGM_G190(MGM_W161,d1_delay);
   and MGM_G191(MGM_W162,MGM_W161,MGM_W160);
   not MGM_G192(MGM_W163,d2_delay);
   and MGM_G193(MGM_W164,MGM_W163,MGM_W162);
   and MGM_G194(MGM_W165,si1_delay,MGM_W164);
   not MGM_G195(MGM_W166,si2_delay);
   and MGM_G196(MGM_W167,MGM_W166,MGM_W165);
   not MGM_G197(MGM_W168,ssb_delay);
   and MGM_G198(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W168,MGM_W167);
   not MGM_G199(MGM_W169,clk_delay);
   not MGM_G200(MGM_W170,d1_delay);
   and MGM_G201(MGM_W171,MGM_W170,MGM_W169);
   not MGM_G202(MGM_W172,d2_delay);
   and MGM_G203(MGM_W173,MGM_W172,MGM_W171);
   and MGM_G204(MGM_W174,si1_delay,MGM_W173);
   not MGM_G205(MGM_W175,si2_delay);
   and MGM_G206(MGM_W176,MGM_W175,MGM_W174);
   and MGM_G207(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W176);
   not MGM_G208(MGM_W177,clk_delay);
   not MGM_G209(MGM_W178,d1_delay);
   and MGM_G210(MGM_W179,MGM_W178,MGM_W177);
   not MGM_G211(MGM_W180,d2_delay);
   and MGM_G212(MGM_W181,MGM_W180,MGM_W179);
   and MGM_G213(MGM_W182,si1_delay,MGM_W181);
   and MGM_G214(MGM_W183,si2_delay,MGM_W182);
   not MGM_G215(MGM_W184,ssb_delay);
   and MGM_G216(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W184,MGM_W183);
   not MGM_G217(MGM_W185,clk_delay);
   not MGM_G218(MGM_W186,d1_delay);
   and MGM_G219(MGM_W187,MGM_W186,MGM_W185);
   not MGM_G220(MGM_W188,d2_delay);
   and MGM_G221(MGM_W189,MGM_W188,MGM_W187);
   and MGM_G222(MGM_W190,si1_delay,MGM_W189);
   and MGM_G223(MGM_W191,si2_delay,MGM_W190);
   and MGM_G224(ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W191);
   not MGM_G225(MGM_W192,clk_delay);
   not MGM_G226(MGM_W193,d1_delay);
   and MGM_G227(MGM_W194,MGM_W193,MGM_W192);
   and MGM_G228(MGM_W195,d2_delay,MGM_W194);
   not MGM_G229(MGM_W196,si1_delay);
   and MGM_G230(MGM_W197,MGM_W196,MGM_W195);
   not MGM_G231(MGM_W198,si2_delay);
   and MGM_G232(MGM_W199,MGM_W198,MGM_W197);
   not MGM_G233(MGM_W200,ssb_delay);
   and MGM_G234(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W200,MGM_W199);
   not MGM_G235(MGM_W201,clk_delay);
   not MGM_G236(MGM_W202,d1_delay);
   and MGM_G237(MGM_W203,MGM_W202,MGM_W201);
   and MGM_G238(MGM_W204,d2_delay,MGM_W203);
   not MGM_G239(MGM_W205,si1_delay);
   and MGM_G240(MGM_W206,MGM_W205,MGM_W204);
   not MGM_G241(MGM_W207,si2_delay);
   and MGM_G242(MGM_W208,MGM_W207,MGM_W206);
   and MGM_G243(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W208);
   not MGM_G244(MGM_W209,clk_delay);
   not MGM_G245(MGM_W210,d1_delay);
   and MGM_G246(MGM_W211,MGM_W210,MGM_W209);
   and MGM_G247(MGM_W212,d2_delay,MGM_W211);
   not MGM_G248(MGM_W213,si1_delay);
   and MGM_G249(MGM_W214,MGM_W213,MGM_W212);
   and MGM_G250(MGM_W215,si2_delay,MGM_W214);
   not MGM_G251(MGM_W216,ssb_delay);
   and MGM_G252(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W216,MGM_W215);
   not MGM_G253(MGM_W217,clk_delay);
   not MGM_G254(MGM_W218,d1_delay);
   and MGM_G255(MGM_W219,MGM_W218,MGM_W217);
   and MGM_G256(MGM_W220,d2_delay,MGM_W219);
   not MGM_G257(MGM_W221,si1_delay);
   and MGM_G258(MGM_W222,MGM_W221,MGM_W220);
   and MGM_G259(MGM_W223,si2_delay,MGM_W222);
   and MGM_G260(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W223);
   not MGM_G261(MGM_W224,clk_delay);
   not MGM_G262(MGM_W225,d1_delay);
   and MGM_G263(MGM_W226,MGM_W225,MGM_W224);
   and MGM_G264(MGM_W227,d2_delay,MGM_W226);
   and MGM_G265(MGM_W228,si1_delay,MGM_W227);
   not MGM_G266(MGM_W229,si2_delay);
   and MGM_G267(MGM_W230,MGM_W229,MGM_W228);
   not MGM_G268(MGM_W231,ssb_delay);
   and MGM_G269(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W231,MGM_W230);
   not MGM_G270(MGM_W232,clk_delay);
   not MGM_G271(MGM_W233,d1_delay);
   and MGM_G272(MGM_W234,MGM_W233,MGM_W232);
   and MGM_G273(MGM_W235,d2_delay,MGM_W234);
   and MGM_G274(MGM_W236,si1_delay,MGM_W235);
   not MGM_G275(MGM_W237,si2_delay);
   and MGM_G276(MGM_W238,MGM_W237,MGM_W236);
   and MGM_G277(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W238);
   not MGM_G278(MGM_W239,clk_delay);
   not MGM_G279(MGM_W240,d1_delay);
   and MGM_G280(MGM_W241,MGM_W240,MGM_W239);
   and MGM_G281(MGM_W242,d2_delay,MGM_W241);
   and MGM_G282(MGM_W243,si1_delay,MGM_W242);
   and MGM_G283(MGM_W244,si2_delay,MGM_W243);
   not MGM_G284(MGM_W245,ssb_delay);
   and MGM_G285(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W245,MGM_W244);
   not MGM_G286(MGM_W246,clk_delay);
   not MGM_G287(MGM_W247,d1_delay);
   and MGM_G288(MGM_W248,MGM_W247,MGM_W246);
   and MGM_G289(MGM_W249,d2_delay,MGM_W248);
   and MGM_G290(MGM_W250,si1_delay,MGM_W249);
   and MGM_G291(MGM_W251,si2_delay,MGM_W250);
   and MGM_G292(ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W251);
   not MGM_G293(MGM_W252,clk_delay);
   and MGM_G294(MGM_W253,d1_delay,MGM_W252);
   not MGM_G295(MGM_W254,d2_delay);
   and MGM_G296(MGM_W255,MGM_W254,MGM_W253);
   not MGM_G297(MGM_W256,si1_delay);
   and MGM_G298(MGM_W257,MGM_W256,MGM_W255);
   not MGM_G299(MGM_W258,si2_delay);
   and MGM_G300(MGM_W259,MGM_W258,MGM_W257);
   not MGM_G301(MGM_W260,ssb_delay);
   and MGM_G302(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W260,MGM_W259);
   not MGM_G303(MGM_W261,clk_delay);
   and MGM_G304(MGM_W262,d1_delay,MGM_W261);
   not MGM_G305(MGM_W263,d2_delay);
   and MGM_G306(MGM_W264,MGM_W263,MGM_W262);
   not MGM_G307(MGM_W265,si1_delay);
   and MGM_G308(MGM_W266,MGM_W265,MGM_W264);
   not MGM_G309(MGM_W267,si2_delay);
   and MGM_G310(MGM_W268,MGM_W267,MGM_W266);
   and MGM_G311(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W268);
   not MGM_G312(MGM_W269,clk_delay);
   and MGM_G313(MGM_W270,d1_delay,MGM_W269);
   not MGM_G314(MGM_W271,d2_delay);
   and MGM_G315(MGM_W272,MGM_W271,MGM_W270);
   not MGM_G316(MGM_W273,si1_delay);
   and MGM_G317(MGM_W274,MGM_W273,MGM_W272);
   and MGM_G318(MGM_W275,si2_delay,MGM_W274);
   not MGM_G319(MGM_W276,ssb_delay);
   and MGM_G320(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W276,MGM_W275);
   not MGM_G321(MGM_W277,clk_delay);
   and MGM_G322(MGM_W278,d1_delay,MGM_W277);
   not MGM_G323(MGM_W279,d2_delay);
   and MGM_G324(MGM_W280,MGM_W279,MGM_W278);
   not MGM_G325(MGM_W281,si1_delay);
   and MGM_G326(MGM_W282,MGM_W281,MGM_W280);
   and MGM_G327(MGM_W283,si2_delay,MGM_W282);
   and MGM_G328(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W283);
   not MGM_G329(MGM_W284,clk_delay);
   and MGM_G330(MGM_W285,d1_delay,MGM_W284);
   not MGM_G331(MGM_W286,d2_delay);
   and MGM_G332(MGM_W287,MGM_W286,MGM_W285);
   and MGM_G333(MGM_W288,si1_delay,MGM_W287);
   not MGM_G334(MGM_W289,si2_delay);
   and MGM_G335(MGM_W290,MGM_W289,MGM_W288);
   not MGM_G336(MGM_W291,ssb_delay);
   and MGM_G337(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W291,MGM_W290);
   not MGM_G338(MGM_W292,clk_delay);
   and MGM_G339(MGM_W293,d1_delay,MGM_W292);
   not MGM_G340(MGM_W294,d2_delay);
   and MGM_G341(MGM_W295,MGM_W294,MGM_W293);
   and MGM_G342(MGM_W296,si1_delay,MGM_W295);
   not MGM_G343(MGM_W297,si2_delay);
   and MGM_G344(MGM_W298,MGM_W297,MGM_W296);
   and MGM_G345(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W298);
   not MGM_G346(MGM_W299,clk_delay);
   and MGM_G347(MGM_W300,d1_delay,MGM_W299);
   not MGM_G348(MGM_W301,d2_delay);
   and MGM_G349(MGM_W302,MGM_W301,MGM_W300);
   and MGM_G350(MGM_W303,si1_delay,MGM_W302);
   and MGM_G351(MGM_W304,si2_delay,MGM_W303);
   not MGM_G352(MGM_W305,ssb_delay);
   and MGM_G353(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W305,MGM_W304);
   not MGM_G354(MGM_W306,clk_delay);
   and MGM_G355(MGM_W307,d1_delay,MGM_W306);
   not MGM_G356(MGM_W308,d2_delay);
   and MGM_G357(MGM_W309,MGM_W308,MGM_W307);
   and MGM_G358(MGM_W310,si1_delay,MGM_W309);
   and MGM_G359(MGM_W311,si2_delay,MGM_W310);
   and MGM_G360(ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W311);
   not MGM_G361(MGM_W312,clk_delay);
   and MGM_G362(MGM_W313,d1_delay,MGM_W312);
   and MGM_G363(MGM_W314,d2_delay,MGM_W313);
   not MGM_G364(MGM_W315,si1_delay);
   and MGM_G365(MGM_W316,MGM_W315,MGM_W314);
   not MGM_G366(MGM_W317,si2_delay);
   and MGM_G367(MGM_W318,MGM_W317,MGM_W316);
   not MGM_G368(MGM_W319,ssb_delay);
   and MGM_G369(ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W319,MGM_W318);
   not MGM_G370(MGM_W320,clk_delay);
   and MGM_G371(MGM_W321,d1_delay,MGM_W320);
   and MGM_G372(MGM_W322,d2_delay,MGM_W321);
   not MGM_G373(MGM_W323,si1_delay);
   and MGM_G374(MGM_W324,MGM_W323,MGM_W322);
   not MGM_G375(MGM_W325,si2_delay);
   and MGM_G376(MGM_W326,MGM_W325,MGM_W324);
   and MGM_G377(ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W326);
   not MGM_G378(MGM_W327,clk_delay);
   and MGM_G379(MGM_W328,d1_delay,MGM_W327);
   and MGM_G380(MGM_W329,d2_delay,MGM_W328);
   not MGM_G381(MGM_W330,si1_delay);
   and MGM_G382(MGM_W331,MGM_W330,MGM_W329);
   and MGM_G383(MGM_W332,si2_delay,MGM_W331);
   not MGM_G384(MGM_W333,ssb_delay);
   and MGM_G385(ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W333,MGM_W332);
   not MGM_G386(MGM_W334,clk_delay);
   and MGM_G387(MGM_W335,d1_delay,MGM_W334);
   and MGM_G388(MGM_W336,d2_delay,MGM_W335);
   not MGM_G389(MGM_W337,si1_delay);
   and MGM_G390(MGM_W338,MGM_W337,MGM_W336);
   and MGM_G391(MGM_W339,si2_delay,MGM_W338);
   and MGM_G392(ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W339);
   not MGM_G393(MGM_W340,clk_delay);
   and MGM_G394(MGM_W341,d1_delay,MGM_W340);
   and MGM_G395(MGM_W342,d2_delay,MGM_W341);
   and MGM_G396(MGM_W343,si1_delay,MGM_W342);
   not MGM_G397(MGM_W344,si2_delay);
   and MGM_G398(MGM_W345,MGM_W344,MGM_W343);
   not MGM_G399(MGM_W346,ssb_delay);
   and MGM_G400(ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W346,MGM_W345);
   not MGM_G401(MGM_W347,clk_delay);
   and MGM_G402(MGM_W348,d1_delay,MGM_W347);
   and MGM_G403(MGM_W349,d2_delay,MGM_W348);
   and MGM_G404(MGM_W350,si1_delay,MGM_W349);
   not MGM_G405(MGM_W351,si2_delay);
   and MGM_G406(MGM_W352,MGM_W351,MGM_W350);
   and MGM_G407(ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W352);
   not MGM_G408(MGM_W353,clk_delay);
   and MGM_G409(MGM_W354,d1_delay,MGM_W353);
   and MGM_G410(MGM_W355,d2_delay,MGM_W354);
   and MGM_G411(MGM_W356,si1_delay,MGM_W355);
   and MGM_G412(MGM_W357,si2_delay,MGM_W356);
   not MGM_G413(MGM_W358,ssb_delay);
   and MGM_G414(ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W358,MGM_W357);
   not MGM_G415(MGM_W359,clk_delay);
   and MGM_G416(MGM_W360,d1_delay,MGM_W359);
   and MGM_G417(MGM_W361,d2_delay,MGM_W360);
   and MGM_G418(MGM_W362,si1_delay,MGM_W361);
   and MGM_G419(MGM_W363,si2_delay,MGM_W362);
   and MGM_G420(ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W363);
   not MGM_G421(MGM_W364,d1_delay);
   and MGM_G422(MGM_W365,MGM_W364,clk_delay);
   not MGM_G423(MGM_W366,d2_delay);
   and MGM_G424(MGM_W367,MGM_W366,MGM_W365);
   not MGM_G425(MGM_W368,si1_delay);
   and MGM_G426(MGM_W369,MGM_W368,MGM_W367);
   not MGM_G427(MGM_W370,si2_delay);
   and MGM_G428(MGM_W371,MGM_W370,MGM_W369);
   not MGM_G429(MGM_W372,ssb_delay);
   and MGM_G430(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W372,MGM_W371);
   not MGM_G431(MGM_W373,d1_delay);
   and MGM_G432(MGM_W374,MGM_W373,clk_delay);
   not MGM_G433(MGM_W375,d2_delay);
   and MGM_G434(MGM_W376,MGM_W375,MGM_W374);
   not MGM_G435(MGM_W377,si1_delay);
   and MGM_G436(MGM_W378,MGM_W377,MGM_W376);
   not MGM_G437(MGM_W379,si2_delay);
   and MGM_G438(MGM_W380,MGM_W379,MGM_W378);
   and MGM_G439(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W380);
   not MGM_G440(MGM_W381,d1_delay);
   and MGM_G441(MGM_W382,MGM_W381,clk_delay);
   not MGM_G442(MGM_W383,d2_delay);
   and MGM_G443(MGM_W384,MGM_W383,MGM_W382);
   not MGM_G444(MGM_W385,si1_delay);
   and MGM_G445(MGM_W386,MGM_W385,MGM_W384);
   and MGM_G446(MGM_W387,si2_delay,MGM_W386);
   not MGM_G447(MGM_W388,ssb_delay);
   and MGM_G448(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W388,MGM_W387);
   not MGM_G449(MGM_W389,d1_delay);
   and MGM_G450(MGM_W390,MGM_W389,clk_delay);
   not MGM_G451(MGM_W391,d2_delay);
   and MGM_G452(MGM_W392,MGM_W391,MGM_W390);
   not MGM_G453(MGM_W393,si1_delay);
   and MGM_G454(MGM_W394,MGM_W393,MGM_W392);
   and MGM_G455(MGM_W395,si2_delay,MGM_W394);
   and MGM_G456(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W395);
   not MGM_G457(MGM_W396,d1_delay);
   and MGM_G458(MGM_W397,MGM_W396,clk_delay);
   not MGM_G459(MGM_W398,d2_delay);
   and MGM_G460(MGM_W399,MGM_W398,MGM_W397);
   and MGM_G461(MGM_W400,si1_delay,MGM_W399);
   not MGM_G462(MGM_W401,si2_delay);
   and MGM_G463(MGM_W402,MGM_W401,MGM_W400);
   not MGM_G464(MGM_W403,ssb_delay);
   and MGM_G465(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W403,MGM_W402);
   not MGM_G466(MGM_W404,d1_delay);
   and MGM_G467(MGM_W405,MGM_W404,clk_delay);
   not MGM_G468(MGM_W406,d2_delay);
   and MGM_G469(MGM_W407,MGM_W406,MGM_W405);
   and MGM_G470(MGM_W408,si1_delay,MGM_W407);
   not MGM_G471(MGM_W409,si2_delay);
   and MGM_G472(MGM_W410,MGM_W409,MGM_W408);
   and MGM_G473(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W410);
   not MGM_G474(MGM_W411,d1_delay);
   and MGM_G475(MGM_W412,MGM_W411,clk_delay);
   not MGM_G476(MGM_W413,d2_delay);
   and MGM_G477(MGM_W414,MGM_W413,MGM_W412);
   and MGM_G478(MGM_W415,si1_delay,MGM_W414);
   and MGM_G479(MGM_W416,si2_delay,MGM_W415);
   not MGM_G480(MGM_W417,ssb_delay);
   and MGM_G481(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W417,MGM_W416);
   not MGM_G482(MGM_W418,d1_delay);
   and MGM_G483(MGM_W419,MGM_W418,clk_delay);
   not MGM_G484(MGM_W420,d2_delay);
   and MGM_G485(MGM_W421,MGM_W420,MGM_W419);
   and MGM_G486(MGM_W422,si1_delay,MGM_W421);
   and MGM_G487(MGM_W423,si2_delay,MGM_W422);
   and MGM_G488(ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W423);
   not MGM_G489(MGM_W424,d1_delay);
   and MGM_G490(MGM_W425,MGM_W424,clk_delay);
   and MGM_G491(MGM_W426,d2_delay,MGM_W425);
   not MGM_G492(MGM_W427,si1_delay);
   and MGM_G493(MGM_W428,MGM_W427,MGM_W426);
   not MGM_G494(MGM_W429,si2_delay);
   and MGM_G495(MGM_W430,MGM_W429,MGM_W428);
   not MGM_G496(MGM_W431,ssb_delay);
   and MGM_G497(ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W431,MGM_W430);
   not MGM_G498(MGM_W432,d1_delay);
   and MGM_G499(MGM_W433,MGM_W432,clk_delay);
   and MGM_G500(MGM_W434,d2_delay,MGM_W433);
   not MGM_G501(MGM_W435,si1_delay);
   and MGM_G502(MGM_W436,MGM_W435,MGM_W434);
   not MGM_G503(MGM_W437,si2_delay);
   and MGM_G504(MGM_W438,MGM_W437,MGM_W436);
   and MGM_G505(ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W438);
   not MGM_G506(MGM_W439,d1_delay);
   and MGM_G507(MGM_W440,MGM_W439,clk_delay);
   and MGM_G508(MGM_W441,d2_delay,MGM_W440);
   not MGM_G509(MGM_W442,si1_delay);
   and MGM_G510(MGM_W443,MGM_W442,MGM_W441);
   and MGM_G511(MGM_W444,si2_delay,MGM_W443);
   not MGM_G512(MGM_W445,ssb_delay);
   and MGM_G513(ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W445,MGM_W444);
   not MGM_G514(MGM_W446,d1_delay);
   and MGM_G515(MGM_W447,MGM_W446,clk_delay);
   and MGM_G516(MGM_W448,d2_delay,MGM_W447);
   not MGM_G517(MGM_W449,si1_delay);
   and MGM_G518(MGM_W450,MGM_W449,MGM_W448);
   and MGM_G519(MGM_W451,si2_delay,MGM_W450);
   and MGM_G520(ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W451);
   not MGM_G521(MGM_W452,d1_delay);
   and MGM_G522(MGM_W453,MGM_W452,clk_delay);
   and MGM_G523(MGM_W454,d2_delay,MGM_W453);
   and MGM_G524(MGM_W455,si1_delay,MGM_W454);
   not MGM_G525(MGM_W456,si2_delay);
   and MGM_G526(MGM_W457,MGM_W456,MGM_W455);
   not MGM_G527(MGM_W458,ssb_delay);
   and MGM_G528(ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W458,MGM_W457);
   not MGM_G529(MGM_W459,d1_delay);
   and MGM_G530(MGM_W460,MGM_W459,clk_delay);
   and MGM_G531(MGM_W461,d2_delay,MGM_W460);
   and MGM_G532(MGM_W462,si1_delay,MGM_W461);
   not MGM_G533(MGM_W463,si2_delay);
   and MGM_G534(MGM_W464,MGM_W463,MGM_W462);
   and MGM_G535(ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W464);
   not MGM_G536(MGM_W465,d1_delay);
   and MGM_G537(MGM_W466,MGM_W465,clk_delay);
   and MGM_G538(MGM_W467,d2_delay,MGM_W466);
   and MGM_G539(MGM_W468,si1_delay,MGM_W467);
   and MGM_G540(MGM_W469,si2_delay,MGM_W468);
   not MGM_G541(MGM_W470,ssb_delay);
   and MGM_G542(ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W470,MGM_W469);
   not MGM_G543(MGM_W471,d1_delay);
   and MGM_G544(MGM_W472,MGM_W471,clk_delay);
   and MGM_G545(MGM_W473,d2_delay,MGM_W472);
   and MGM_G546(MGM_W474,si1_delay,MGM_W473);
   and MGM_G547(MGM_W475,si2_delay,MGM_W474);
   and MGM_G548(ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W475);
   and MGM_G549(MGM_W476,d1_delay,clk_delay);
   not MGM_G550(MGM_W477,d2_delay);
   and MGM_G551(MGM_W478,MGM_W477,MGM_W476);
   not MGM_G552(MGM_W479,si1_delay);
   and MGM_G553(MGM_W480,MGM_W479,MGM_W478);
   not MGM_G554(MGM_W481,si2_delay);
   and MGM_G555(MGM_W482,MGM_W481,MGM_W480);
   not MGM_G556(MGM_W483,ssb_delay);
   and MGM_G557(ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W483,MGM_W482);
   and MGM_G558(MGM_W484,d1_delay,clk_delay);
   not MGM_G559(MGM_W485,d2_delay);
   and MGM_G560(MGM_W486,MGM_W485,MGM_W484);
   not MGM_G561(MGM_W487,si1_delay);
   and MGM_G562(MGM_W488,MGM_W487,MGM_W486);
   not MGM_G563(MGM_W489,si2_delay);
   and MGM_G564(MGM_W490,MGM_W489,MGM_W488);
   and MGM_G565(ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W490);
   and MGM_G566(MGM_W491,d1_delay,clk_delay);
   not MGM_G567(MGM_W492,d2_delay);
   and MGM_G568(MGM_W493,MGM_W492,MGM_W491);
   not MGM_G569(MGM_W494,si1_delay);
   and MGM_G570(MGM_W495,MGM_W494,MGM_W493);
   and MGM_G571(MGM_W496,si2_delay,MGM_W495);
   not MGM_G572(MGM_W497,ssb_delay);
   and MGM_G573(ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W497,MGM_W496);
   and MGM_G574(MGM_W498,d1_delay,clk_delay);
   not MGM_G575(MGM_W499,d2_delay);
   and MGM_G576(MGM_W500,MGM_W499,MGM_W498);
   not MGM_G577(MGM_W501,si1_delay);
   and MGM_G578(MGM_W502,MGM_W501,MGM_W500);
   and MGM_G579(MGM_W503,si2_delay,MGM_W502);
   and MGM_G580(ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W503);
   and MGM_G581(MGM_W504,d1_delay,clk_delay);
   not MGM_G582(MGM_W505,d2_delay);
   and MGM_G583(MGM_W506,MGM_W505,MGM_W504);
   and MGM_G584(MGM_W507,si1_delay,MGM_W506);
   not MGM_G585(MGM_W508,si2_delay);
   and MGM_G586(MGM_W509,MGM_W508,MGM_W507);
   not MGM_G587(MGM_W510,ssb_delay);
   and MGM_G588(ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W510,MGM_W509);
   and MGM_G589(MGM_W511,d1_delay,clk_delay);
   not MGM_G590(MGM_W512,d2_delay);
   and MGM_G591(MGM_W513,MGM_W512,MGM_W511);
   and MGM_G592(MGM_W514,si1_delay,MGM_W513);
   not MGM_G593(MGM_W515,si2_delay);
   and MGM_G594(MGM_W516,MGM_W515,MGM_W514);
   and MGM_G595(ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W516);
   and MGM_G596(MGM_W517,d1_delay,clk_delay);
   not MGM_G597(MGM_W518,d2_delay);
   and MGM_G598(MGM_W519,MGM_W518,MGM_W517);
   and MGM_G599(MGM_W520,si1_delay,MGM_W519);
   and MGM_G600(MGM_W521,si2_delay,MGM_W520);
   not MGM_G601(MGM_W522,ssb_delay);
   and MGM_G602(ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W522,MGM_W521);
   and MGM_G603(MGM_W523,d1_delay,clk_delay);
   not MGM_G604(MGM_W524,d2_delay);
   and MGM_G605(MGM_W525,MGM_W524,MGM_W523);
   and MGM_G606(MGM_W526,si1_delay,MGM_W525);
   and MGM_G607(MGM_W527,si2_delay,MGM_W526);
   and MGM_G608(ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W527);
   and MGM_G609(MGM_W528,d1_delay,clk_delay);
   and MGM_G610(MGM_W529,d2_delay,MGM_W528);
   not MGM_G611(MGM_W530,si1_delay);
   and MGM_G612(MGM_W531,MGM_W530,MGM_W529);
   not MGM_G613(MGM_W532,si2_delay);
   and MGM_G614(MGM_W533,MGM_W532,MGM_W531);
   not MGM_G615(MGM_W534,ssb_delay);
   and MGM_G616(ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W534,MGM_W533);
   and MGM_G617(MGM_W535,d1_delay,clk_delay);
   and MGM_G618(MGM_W536,d2_delay,MGM_W535);
   not MGM_G619(MGM_W537,si1_delay);
   and MGM_G620(MGM_W538,MGM_W537,MGM_W536);
   not MGM_G621(MGM_W539,si2_delay);
   and MGM_G622(MGM_W540,MGM_W539,MGM_W538);
   and MGM_G623(ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W540);
   and MGM_G624(MGM_W541,d1_delay,clk_delay);
   and MGM_G625(MGM_W542,d2_delay,MGM_W541);
   not MGM_G626(MGM_W543,si1_delay);
   and MGM_G627(MGM_W544,MGM_W543,MGM_W542);
   and MGM_G628(MGM_W545,si2_delay,MGM_W544);
   not MGM_G629(MGM_W546,ssb_delay);
   and MGM_G630(ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb,MGM_W546,MGM_W545);
   and MGM_G631(MGM_W547,d1_delay,clk_delay);
   and MGM_G632(MGM_W548,d2_delay,MGM_W547);
   not MGM_G633(MGM_W549,si1_delay);
   and MGM_G634(MGM_W550,MGM_W549,MGM_W548);
   and MGM_G635(MGM_W551,si2_delay,MGM_W550);
   and MGM_G636(ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb,ssb_delay,MGM_W551);
   and MGM_G637(MGM_W552,d1_delay,clk_delay);
   and MGM_G638(MGM_W553,d2_delay,MGM_W552);
   and MGM_G639(MGM_W554,si1_delay,MGM_W553);
   not MGM_G640(MGM_W555,si2_delay);
   and MGM_G641(MGM_W556,MGM_W555,MGM_W554);
   not MGM_G642(MGM_W557,ssb_delay);
   and MGM_G643(ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb,MGM_W557,MGM_W556);
   and MGM_G644(MGM_W558,d1_delay,clk_delay);
   and MGM_G645(MGM_W559,d2_delay,MGM_W558);
   and MGM_G646(MGM_W560,si1_delay,MGM_W559);
   not MGM_G647(MGM_W561,si2_delay);
   and MGM_G648(MGM_W562,MGM_W561,MGM_W560);
   and MGM_G649(ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb,ssb_delay,MGM_W562);
   and MGM_G650(MGM_W563,d1_delay,clk_delay);
   and MGM_G651(MGM_W564,d2_delay,MGM_W563);
   and MGM_G652(MGM_W565,si1_delay,MGM_W564);
   and MGM_G653(MGM_W566,si2_delay,MGM_W565);
   not MGM_G654(MGM_W567,ssb_delay);
   and MGM_G655(ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb,MGM_W567,MGM_W566);
   and MGM_G656(MGM_W568,d1_delay,clk_delay);
   and MGM_G657(MGM_W569,d2_delay,MGM_W568);
   and MGM_G658(MGM_W570,si1_delay,MGM_W569);
   and MGM_G659(MGM_W571,si2_delay,MGM_W570);
   and MGM_G660(ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_ssb,ssb_delay,MGM_W571);
   not MGM_G661(MGM_W572,d1_delay);
   not MGM_G662(MGM_W573,d2_delay);
   and MGM_G663(MGM_W574,MGM_W573,MGM_W572);
   and MGM_G664(MGM_W575,rb_delay,MGM_W574);
   not MGM_G665(MGM_W576,si1_delay);
   and MGM_G666(MGM_W577,MGM_W576,MGM_W575);
   and MGM_G667(ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2,si2_delay,MGM_W577);
   not MGM_G668(MGM_W578,d1_delay);
   not MGM_G669(MGM_W579,d2_delay);
   and MGM_G670(MGM_W580,MGM_W579,MGM_W578);
   and MGM_G671(MGM_W581,rb_delay,MGM_W580);
   and MGM_G672(MGM_W582,si1_delay,MGM_W581);
   not MGM_G673(MGM_W583,si2_delay);
   and MGM_G674(ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2,MGM_W583,MGM_W582);
   not MGM_G675(MGM_W584,d1_delay);
   not MGM_G676(MGM_W585,d2_delay);
   and MGM_G677(MGM_W586,MGM_W585,MGM_W584);
   and MGM_G678(MGM_W587,rb_delay,MGM_W586);
   and MGM_G679(MGM_W588,si1_delay,MGM_W587);
   and MGM_G680(ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2,si2_delay,MGM_W588);
   not MGM_G681(MGM_W589,d1_delay);
   and MGM_G682(MGM_W590,d2_delay,MGM_W589);
   and MGM_G683(MGM_W591,rb_delay,MGM_W590);
   not MGM_G684(MGM_W592,si1_delay);
   and MGM_G685(MGM_W593,MGM_W592,MGM_W591);
   not MGM_G686(MGM_W594,si2_delay);
   and MGM_G687(ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2,MGM_W594,MGM_W593);
   not MGM_G688(MGM_W595,d1_delay);
   and MGM_G689(MGM_W596,d2_delay,MGM_W595);
   and MGM_G690(MGM_W597,rb_delay,MGM_W596);
   and MGM_G691(MGM_W598,si1_delay,MGM_W597);
   not MGM_G692(MGM_W599,si2_delay);
   and MGM_G693(ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2,MGM_W599,MGM_W598);
   not MGM_G694(MGM_W600,d1_delay);
   and MGM_G695(MGM_W601,d2_delay,MGM_W600);
   and MGM_G696(MGM_W602,rb_delay,MGM_W601);
   and MGM_G697(MGM_W603,si1_delay,MGM_W602);
   and MGM_G698(ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2,si2_delay,MGM_W603);
   not MGM_G699(MGM_W604,d2_delay);
   and MGM_G700(MGM_W605,MGM_W604,d1_delay);
   and MGM_G701(MGM_W606,rb_delay,MGM_W605);
   not MGM_G702(MGM_W607,si1_delay);
   and MGM_G703(MGM_W608,MGM_W607,MGM_W606);
   not MGM_G704(MGM_W609,si2_delay);
   and MGM_G705(ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2,MGM_W609,MGM_W608);
   not MGM_G706(MGM_W610,d2_delay);
   and MGM_G707(MGM_W611,MGM_W610,d1_delay);
   and MGM_G708(MGM_W612,rb_delay,MGM_W611);
   not MGM_G709(MGM_W613,si1_delay);
   and MGM_G710(MGM_W614,MGM_W613,MGM_W612);
   and MGM_G711(ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2,si2_delay,MGM_W614);
   not MGM_G712(MGM_W615,d2_delay);
   and MGM_G713(MGM_W616,MGM_W615,d1_delay);
   and MGM_G714(MGM_W617,rb_delay,MGM_W616);
   and MGM_G715(MGM_W618,si1_delay,MGM_W617);
   and MGM_G716(ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2,si2_delay,MGM_W618);
   and MGM_G717(MGM_W619,d2_delay,d1_delay);
   and MGM_G718(MGM_W620,rb_delay,MGM_W619);
   not MGM_G719(MGM_W621,si1_delay);
   and MGM_G720(MGM_W622,MGM_W621,MGM_W620);
   not MGM_G721(MGM_W623,si2_delay);
   and MGM_G722(ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2,MGM_W623,MGM_W622);
   and MGM_G723(MGM_W624,d2_delay,d1_delay);
   and MGM_G724(MGM_W625,rb_delay,MGM_W624);
   not MGM_G725(MGM_W626,si1_delay);
   and MGM_G726(MGM_W627,MGM_W626,MGM_W625);
   and MGM_G727(ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2,si2_delay,MGM_W627);
   and MGM_G728(MGM_W628,d2_delay,d1_delay);
   and MGM_G729(MGM_W629,rb_delay,MGM_W628);
   and MGM_G730(MGM_W630,si1_delay,MGM_W629);
   not MGM_G731(MGM_W631,si2_delay);
   and MGM_G732(ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2,MGM_W631,MGM_W630);
   and MGM_G733(ENABLE_ssb_AND_rb,rb_delay,ssb_delay);
   not MGM_G734(MGM_W632,ssb_delay);
   and MGM_G735(ENABLE_NOT_ssb_AND_rb,rb_delay,MGM_W632);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d1==1'b0 && rb==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_rb == 1'b1)
      ,0.0,0,notifier);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_NOT_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_NOT_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_NOT_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_NOT_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_NOT_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clk_AND_d1_AND_d2_AND_si1_AND_si2_AND_ssb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb,0.0,0,notifier);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_NOT_d2_AND_rb_AND_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_NOT_si1_AND_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_rb_AND_si1_AND_NOT_si2 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,negedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,posedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d1 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d1 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d2 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d2 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si1 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si1 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si2 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si2 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_fqy403ah_func( clk, d1, d2, d3, d4, o1, o2, o3, o4, rb, si1, si2, si3, si4, ssb, notifier0, notifier1, notifier2, notifier3 `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, d3, d4, rb, si1, si2, si3, si4, ssb, notifier0, notifier1, notifier2, notifier3;
   output o1, o2, o3, o4;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_CLK0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D0, d4, si4, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ4, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, vcc, vssx, notifier3 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C1, rb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D1, d3, si3, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ3, MGM_C1, 1'b0, MGM_CLK1, MGM_D1, vcc, vssx, notifier2 );
   INTCseq_cdiar2ah_0( MGM_CLK2, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C2, rb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D2, d2, si2, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, MGM_C2, 1'b0, MGM_CLK2, MGM_D2, vcc, vssx, notifier1 );
   INTCseq_cdiar2ah_0( MGM_CLK3, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C3, rb, vcc, vssx );
   INTCseq_fdw003ah_5( MGM_D3, d1, si1, ssb, vcc, vssx );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, MGM_C3, 1'b0, MGM_CLK3, MGM_D3, vcc, vssx, notifier0 );
   INTCseq_cdiar2ah_0( o1, IQ1, vcc, vssx );
   INTCseq_cdiar2ah_0( o2, IQ2, vcc, vssx );
   INTCseq_cdiar2ah_0( o3, IQ3, vcc, vssx );
   INTCseq_cdiar2ah_0( o4, IQ4, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_CLK0, clk );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_fdw003ah_5( MGM_D0, d4, si4, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ4, MGM_C0, 1'b0, MGM_CLK0, MGM_D0, notifier3 );
   INTCseq_cdiar2ah_0( MGM_CLK1, clk );
   INTCseq_cdiar2ah_1( MGM_C1, rb );
   INTCseq_fdw003ah_5( MGM_D1, d3, si3, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ3, MGM_C1, 1'b0, MGM_CLK1, MGM_D1, notifier2 );
   INTCseq_cdiar2ah_0( MGM_CLK2, clk );
   INTCseq_cdiar2ah_1( MGM_C2, rb );
   INTCseq_fdw003ah_5( MGM_D2, d2, si2, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ2, MGM_C2, 1'b0, MGM_CLK2, MGM_D2, notifier1 );
   INTCseq_cdiar2ah_0( MGM_CLK3, clk );
   INTCseq_cdiar2ah_1( MGM_C3, rb );
   INTCseq_fdw003ah_5( MGM_D3, d1, si1, ssb );
   INTCseq_cdiar2ah_N_IQ_FF_UDP( IQ1, MGM_C3, 1'b0, MGM_CLK3, MGM_D3, notifier0 );
   INTCseq_cdiar2ah_0( o1, IQ1 );
   INTCseq_cdiar2ah_0( o2, IQ2 );
   INTCseq_cdiar2ah_0( o3, IQ3 );
   INTCseq_cdiar2ah_0( o4, IQ4 );
`endif

endmodule
`endcelldefine



`celldefine
module b15fqy403ah1d02x5( clk, d1, d2, d3, d4, o1, o2, o3, o4, rb, si1, si2, si3, si4, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, d3, d4, rb, si1, si2, si3, si4, ssb;
   output o1, o2, o3, o4;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy403ah_func b15fqy403ah1d02x5_behav_inst(.clk(clk),.rb(rb),.ssb(ssb),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.si1(si1),.si2(si2),.si3(si3),.si4(si4),.notifier0(1'b0),.notifier1(1'b0),.notifier2(1'b0),.notifier3(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy403ah_func b15fqy403ah1d02x5_behav_inst(.clk(clk),.rb(rb),.ssb(ssb),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.si1(si1),.si2(si2),.si3(si3),.si4(si4),.notifier0(1'b0),.notifier1(1'b0),.notifier2(1'b0),.notifier3(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire rb_delay ;
   wire ssb_delay ;
   wire d1_delay ;
   wire d2_delay ;
   wire d3_delay ;
   wire d4_delay ;
   wire si1_delay ;
   wire si2_delay ;
   wire si3_delay ;
   wire si4_delay ;
   reg notifier;
   reg notifier0;
   reg notifier1;
   reg notifier2;
   reg notifier3;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
     notifier1 = (notifier1 !== notifier) ? notifier : ~notifier1;
     notifier2 = (notifier2 !== notifier) ? notifier : ~notifier2;
     notifier3 = (notifier3 !== notifier) ? notifier : ~notifier3;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy403ah_func b15fqy403ah1d02x5_inst(.clk(clk_delay),.rb(rb_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1_delay),.d2(d2_delay),.d3(d3_delay),.d4(d4_delay),.si1(si1_delay),.si2(si2_delay),.si3(si3_delay),.si4(si4_delay),.notifier0(notifier0),.notifier1(notifier1),.notifier2(notifier2),.notifier3(notifier3),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy403ah_func b15fqy403ah1d02x5_inst(.clk(clk_delay),.rb(rb_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1_delay),.d2(d2_delay),.d3(d3_delay),.d4(d4_delay),.si1(si1_delay),.si2(si2_delay),.si3(si3_delay),.si4(si4_delay),.notifier0(notifier0),.notifier1(notifier1),.notifier2(notifier2),.notifier3(notifier3));
   `endif
   
   // spec_gates_begin
   buf MGM_G0(ENABLE_rb,rb_delay);
   and MGM_G1(MGM_W0,d2_delay,d1_delay);
   and MGM_G2(MGM_W1,d3_delay,MGM_W0);
   and MGM_G3(MGM_W2,d4_delay,MGM_W1);
   and MGM_G4(MGM_W3,si1_delay,MGM_W2);
   and MGM_G5(MGM_W4,si2_delay,MGM_W3);
   and MGM_G6(MGM_W5,si3_delay,MGM_W4);
   and MGM_G7(MGM_W6,si4_delay,MGM_W5);
   and MGM_G8(ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_si1_AND_si2_AND_si3_AND_si4_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d1_delay);
   not MGM_G10(MGM_W8,d2_delay);
   and MGM_G11(MGM_W9,MGM_W8,MGM_W7);
   not MGM_G12(MGM_W10,d3_delay);
   and MGM_G13(MGM_W11,MGM_W10,MGM_W9);
   not MGM_G14(MGM_W12,d4_delay);
   and MGM_G15(MGM_W13,MGM_W12,MGM_W11);
   and MGM_G16(MGM_W14,si1_delay,MGM_W13);
   and MGM_G17(MGM_W15,si2_delay,MGM_W14);
   and MGM_G18(MGM_W16,si3_delay,MGM_W15);
   and MGM_G19(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4,si4_delay,MGM_W16);
   and MGM_G20(MGM_W17,d2_delay,d1_delay);
   and MGM_G21(MGM_W18,d3_delay,MGM_W17);
   and MGM_G22(MGM_W19,d4_delay,MGM_W18);
   not MGM_G23(MGM_W20,si1_delay);
   and MGM_G24(MGM_W21,MGM_W20,MGM_W19);
   not MGM_G25(MGM_W22,si2_delay);
   and MGM_G26(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G27(MGM_W24,si3_delay);
   and MGM_G28(MGM_W25,MGM_W24,MGM_W23);
   not MGM_G29(MGM_W26,si4_delay);
   and MGM_G30(ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4,MGM_W26,MGM_W25);
   and MGM_G31(ENABLE_ssb_AND_rb,rb_delay,ssb_delay);
   not MGM_G32(MGM_W27,ssb_delay);
   and MGM_G33(ENABLE_NOT_ssb_AND_rb,rb_delay,MGM_W27);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d1==1'b0 && rb==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(d3==1'b0 && rb==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && rb==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && rb==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && rb==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && rb==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && rb==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && rb==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && rb==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b0 && si3==1'b0 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b0 && si3==1'b0 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b0 && si3==1'b1 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b0 && si3==1'b1 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b0 && si3==1'b0 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b0 && si3==1'b0 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b0 && si3==1'b1 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b0 && si3==1'b1 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(d4==1'b0 && rb==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && rb==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && rb==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && rb==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && rb==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && rb==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && rb==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && rb==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b0 && si4==1'b0 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b0 && si4==1'b0 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b0 && si4==1'b1 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b0 && si4==1'b1 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b0 && si4==1'b0 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b0 && si4==1'b0 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b0 && si4==1'b1 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b0 && si4==1'b1 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_rb == 1'b1)
      ,0.0,0,notifier);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_si1_AND_si2_AND_si3_AND_si4_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_si1_AND_si2_AND_si3_AND_si4_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb,0.0,0,notifier);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,negedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,posedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d1 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d1 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d2 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d2 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d3 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,d3_delay);
      
      // setuphold d3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d3 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,d3_delay);
      
      // setuphold d4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d4 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,d4_delay);
      
      // setuphold d4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d4 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,d4_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si1 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si1 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si2 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si2 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si3 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,si3_delay);
      
      // setuphold si3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si3 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,si3_delay);
      
      // setuphold si4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si4 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,si4_delay);
      
      // setuphold si4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si4 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,si4_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy403ah1d03x5( clk, d1, d2, d3, d4, o1, o2, o3, o4, rb, si1, si2, si3, si4, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, d3, d4, rb, si1, si2, si3, si4, ssb;
   output o1, o2, o3, o4;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy403ah_func b15fqy403ah1d03x5_behav_inst(.clk(clk),.rb(rb),.ssb(ssb),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.si1(si1),.si2(si2),.si3(si3),.si4(si4),.notifier0(1'b0),.notifier1(1'b0),.notifier2(1'b0),.notifier3(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy403ah_func b15fqy403ah1d03x5_behav_inst(.clk(clk),.rb(rb),.ssb(ssb),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.si1(si1),.si2(si2),.si3(si3),.si4(si4),.notifier0(1'b0),.notifier1(1'b0),.notifier2(1'b0),.notifier3(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire rb_delay ;
   wire ssb_delay ;
   wire d1_delay ;
   wire d2_delay ;
   wire d3_delay ;
   wire d4_delay ;
   wire si1_delay ;
   wire si2_delay ;
   wire si3_delay ;
   wire si4_delay ;
   reg notifier;
   reg notifier0;
   reg notifier1;
   reg notifier2;
   reg notifier3;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
     notifier1 = (notifier1 !== notifier) ? notifier : ~notifier1;
     notifier2 = (notifier2 !== notifier) ? notifier : ~notifier2;
     notifier3 = (notifier3 !== notifier) ? notifier : ~notifier3;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy403ah_func b15fqy403ah1d03x5_inst(.clk(clk_delay),.rb(rb_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1_delay),.d2(d2_delay),.d3(d3_delay),.d4(d4_delay),.si1(si1_delay),.si2(si2_delay),.si3(si3_delay),.si4(si4_delay),.notifier0(notifier0),.notifier1(notifier1),.notifier2(notifier2),.notifier3(notifier3),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy403ah_func b15fqy403ah1d03x5_inst(.clk(clk_delay),.rb(rb_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1_delay),.d2(d2_delay),.d3(d3_delay),.d4(d4_delay),.si1(si1_delay),.si2(si2_delay),.si3(si3_delay),.si4(si4_delay),.notifier0(notifier0),.notifier1(notifier1),.notifier2(notifier2),.notifier3(notifier3));
   `endif
   
   // spec_gates_begin
   buf MGM_G0(ENABLE_rb,rb_delay);
   and MGM_G1(MGM_W0,d2_delay,d1_delay);
   and MGM_G2(MGM_W1,d3_delay,MGM_W0);
   and MGM_G3(MGM_W2,d4_delay,MGM_W1);
   and MGM_G4(MGM_W3,si1_delay,MGM_W2);
   and MGM_G5(MGM_W4,si2_delay,MGM_W3);
   and MGM_G6(MGM_W5,si3_delay,MGM_W4);
   and MGM_G7(MGM_W6,si4_delay,MGM_W5);
   and MGM_G8(ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_si1_AND_si2_AND_si3_AND_si4_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d1_delay);
   not MGM_G10(MGM_W8,d2_delay);
   and MGM_G11(MGM_W9,MGM_W8,MGM_W7);
   not MGM_G12(MGM_W10,d3_delay);
   and MGM_G13(MGM_W11,MGM_W10,MGM_W9);
   not MGM_G14(MGM_W12,d4_delay);
   and MGM_G15(MGM_W13,MGM_W12,MGM_W11);
   and MGM_G16(MGM_W14,si1_delay,MGM_W13);
   and MGM_G17(MGM_W15,si2_delay,MGM_W14);
   and MGM_G18(MGM_W16,si3_delay,MGM_W15);
   and MGM_G19(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4,si4_delay,MGM_W16);
   and MGM_G20(MGM_W17,d2_delay,d1_delay);
   and MGM_G21(MGM_W18,d3_delay,MGM_W17);
   and MGM_G22(MGM_W19,d4_delay,MGM_W18);
   not MGM_G23(MGM_W20,si1_delay);
   and MGM_G24(MGM_W21,MGM_W20,MGM_W19);
   not MGM_G25(MGM_W22,si2_delay);
   and MGM_G26(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G27(MGM_W24,si3_delay);
   and MGM_G28(MGM_W25,MGM_W24,MGM_W23);
   not MGM_G29(MGM_W26,si4_delay);
   and MGM_G30(ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4,MGM_W26,MGM_W25);
   and MGM_G31(ENABLE_ssb_AND_rb,rb_delay,ssb_delay);
   not MGM_G32(MGM_W27,ssb_delay);
   and MGM_G33(ENABLE_NOT_ssb_AND_rb,rb_delay,MGM_W27);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d1==1'b0 && rb==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(d3==1'b0 && rb==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && rb==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && rb==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && rb==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && rb==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && rb==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && rb==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && rb==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b0 && si3==1'b0 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b0 && si3==1'b0 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b0 && si3==1'b1 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b0 && si3==1'b1 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b0 && si3==1'b0 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b0 && si3==1'b0 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b0 && si3==1'b1 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b0 && si3==1'b1 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(d4==1'b0 && rb==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && rb==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && rb==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && rb==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && rb==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && rb==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && rb==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && rb==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b0 && si4==1'b0 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b0 && si4==1'b0 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b0 && si4==1'b1 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b0 && si4==1'b1 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b0 && si4==1'b0 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b0 && si4==1'b0 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b0 && si4==1'b1 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b0 && si4==1'b1 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_rb == 1'b1)
      ,0.0,0,notifier);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_si1_AND_si2_AND_si3_AND_si4_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_si1_AND_si2_AND_si3_AND_si4_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb,0.0,0,notifier);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,negedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,posedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d1 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d1 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d2 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d2 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d3 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,d3_delay);
      
      // setuphold d3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d3 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,d3_delay);
      
      // setuphold d4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d4 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,d4_delay);
      
      // setuphold d4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d4 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,d4_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si1 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si1 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si2 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si2 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si3 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,si3_delay);
      
      // setuphold si3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si3 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,si3_delay);
      
      // setuphold si4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si4 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,si4_delay);
      
      // setuphold si4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si4 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,si4_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15fqy403ah1d04x5( clk, d1, d2, d3, d4, o1, o2, o3, o4, rb, si1, si2, si3, si4, ssb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d1, d2, d3, d4, rb, si1, si2, si3, si4, ssb;
   output o1, o2, o3, o4;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy403ah_func b15fqy403ah1d04x5_behav_inst(.clk(clk),.rb(rb),.ssb(ssb),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.si1(si1),.si2(si2),.si3(si3),.si4(si4),.notifier0(1'b0),.notifier1(1'b0),.notifier2(1'b0),.notifier3(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy403ah_func b15fqy403ah1d04x5_behav_inst(.clk(clk),.rb(rb),.ssb(ssb),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1),.d2(d2),.d3(d3),.d4(d4),.si1(si1),.si2(si2),.si3(si3),.si4(si4),.notifier0(1'b0),.notifier1(1'b0),.notifier2(1'b0),.notifier3(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire rb_delay ;
   wire ssb_delay ;
   wire d1_delay ;
   wire d2_delay ;
   wire d3_delay ;
   wire d4_delay ;
   wire si1_delay ;
   wire si2_delay ;
   wire si3_delay ;
   wire si4_delay ;
   reg notifier;
   reg notifier0;
   reg notifier1;
   reg notifier2;
   reg notifier3;
   
   always@(notifier) begin
     notifier0 = (notifier0 !== notifier) ? notifier : ~notifier0;
     notifier1 = (notifier1 !== notifier) ? notifier : ~notifier1;
     notifier2 = (notifier2 !== notifier) ? notifier : ~notifier2;
     notifier3 = (notifier3 !== notifier) ? notifier : ~notifier3;
   end
   
   
   `ifdef POWER_AWARE_MODE
      INTCseq_fqy403ah_func b15fqy403ah1d04x5_inst(.clk(clk_delay),.rb(rb_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1_delay),.d2(d2_delay),.d3(d3_delay),.d4(d4_delay),.si1(si1_delay),.si2(si2_delay),.si3(si3_delay),.si4(si4_delay),.notifier0(notifier0),.notifier1(notifier1),.notifier2(notifier2),.notifier3(notifier3),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_fqy403ah_func b15fqy403ah1d04x5_inst(.clk(clk_delay),.rb(rb_delay),.ssb(ssb_delay),.o1(o1),.o2(o2),.o3(o3),.o4(o4),.d1(d1_delay),.d2(d2_delay),.d3(d3_delay),.d4(d4_delay),.si1(si1_delay),.si2(si2_delay),.si3(si3_delay),.si4(si4_delay),.notifier0(notifier0),.notifier1(notifier1),.notifier2(notifier2),.notifier3(notifier3));
   `endif
   
   // spec_gates_begin
   buf MGM_G0(ENABLE_rb,rb_delay);
   and MGM_G1(MGM_W0,d2_delay,d1_delay);
   and MGM_G2(MGM_W1,d3_delay,MGM_W0);
   and MGM_G3(MGM_W2,d4_delay,MGM_W1);
   and MGM_G4(MGM_W3,si1_delay,MGM_W2);
   and MGM_G5(MGM_W4,si2_delay,MGM_W3);
   and MGM_G6(MGM_W5,si3_delay,MGM_W4);
   and MGM_G7(MGM_W6,si4_delay,MGM_W5);
   and MGM_G8(ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_si1_AND_si2_AND_si3_AND_si4_AND_ssb,ssb_delay,MGM_W6);
   not MGM_G9(MGM_W7,d1_delay);
   not MGM_G10(MGM_W8,d2_delay);
   and MGM_G11(MGM_W9,MGM_W8,MGM_W7);
   not MGM_G12(MGM_W10,d3_delay);
   and MGM_G13(MGM_W11,MGM_W10,MGM_W9);
   not MGM_G14(MGM_W12,d4_delay);
   and MGM_G15(MGM_W13,MGM_W12,MGM_W11);
   and MGM_G16(MGM_W14,si1_delay,MGM_W13);
   and MGM_G17(MGM_W15,si2_delay,MGM_W14);
   and MGM_G18(MGM_W16,si3_delay,MGM_W15);
   and MGM_G19(ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4,si4_delay,MGM_W16);
   and MGM_G20(MGM_W17,d2_delay,d1_delay);
   and MGM_G21(MGM_W18,d3_delay,MGM_W17);
   and MGM_G22(MGM_W19,d4_delay,MGM_W18);
   not MGM_G23(MGM_W20,si1_delay);
   and MGM_G24(MGM_W21,MGM_W20,MGM_W19);
   not MGM_G25(MGM_W22,si2_delay);
   and MGM_G26(MGM_W23,MGM_W22,MGM_W21);
   not MGM_G27(MGM_W24,si3_delay);
   and MGM_G28(MGM_W25,MGM_W24,MGM_W23);
   not MGM_G29(MGM_W26,si4_delay);
   and MGM_G30(ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4,MGM_W26,MGM_W25);
   and MGM_G31(ENABLE_ssb_AND_rb,rb_delay,ssb_delay);
   not MGM_G32(MGM_W27,ssb_delay);
   and MGM_G33(ENABLE_NOT_ssb_AND_rb,rb_delay,MGM_W27);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d1==1'b0 && rb==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b0 && rb==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(d1==1'b1 && rb==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc clk --> o1
      (posedge clk => (o1 : d1))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b0 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b0 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b0 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b1 && ssb==1'b0)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d1==1'b1 && si1==1'b1 && ssb==1'b1)
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o1
      (negedge rb => (o1 +: 1'b0))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b0 && rb==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(d2==1'b1 && rb==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc clk --> o2
      (posedge clk => (o2 : d2))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b0 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b0 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b0 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b1 && ssb==1'b0)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d2==1'b1 && si2==1'b1 && ssb==1'b1)
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o2
      (negedge rb => (o2 +: 1'b0))  = (0.0,0.0);
      
      if(d3==1'b0 && rb==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && rb==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && rb==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && rb==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b0 && rb==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && rb==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && rb==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(d3==1'b1 && rb==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc clk --> o3
      (posedge clk => (o3 : d3))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b0 && si3==1'b0 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b0 && si3==1'b0 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b0 && si3==1'b1 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b0 && si3==1'b1 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d3==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b0 && si3==1'b0 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b0 && si3==1'b0 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b0 && si3==1'b1 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b0 && si3==1'b1 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b1 && si3==1'b0 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b1 && si3==1'b0 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b1 && si3==1'b1 && ssb==1'b0)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d3==1'b1 && si3==1'b1 && ssb==1'b1)
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o3
      (negedge rb => (o3 +: 1'b0))  = (0.0,0.0);
      
      if(d4==1'b0 && rb==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && rb==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && rb==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && rb==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      ifnone
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b0 && rb==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && rb==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && rb==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(d4==1'b1 && rb==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc clk --> o4
      (posedge clk => (o4 : d4))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b0 && si4==1'b0 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b0 && si4==1'b0 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b0 && si4==1'b1 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b0 && si4==1'b1 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d4==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b0 && si4==1'b0 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b0 && si4==1'b0 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b0 && si4==1'b1 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b0 && si4==1'b1 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b1 && si4==1'b0 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b1 && si4==1'b0 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b1 && si4==1'b1 && ssb==1'b0)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d4==1'b1 && si4==1'b1 && ssb==1'b1)
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      ifnone
      // seq arc rb --> o4
      (negedge rb => (o4 +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clk &&& (ENABLE_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_rb == 1'b1)
      ,0.0,0,notifier);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_si1_AND_si2_AND_si3_AND_si4_AND_ssb == 1'b1),
      posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_si1_AND_si2_AND_si3_AND_si4_AND_ssb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // recrem rb-clk-posedge
      $recrem(posedge rb,posedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb,0.0,0,notifier);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      negedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      posedge ssb &&& (ENABLE_NOT_d1_AND_NOT_d2_AND_NOT_d3_AND_NOT_d4_AND_si1_AND_si2_AND_si3_AND_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      negedge ssb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      posedge ssb &&& (ENABLE_d1_AND_d2_AND_d3_AND_d4_AND_NOT_si1_AND_NOT_si2_AND_NOT_si3_AND_NOT_si4 == 1'b1),
      0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,negedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold ssb- clk-LH
      $setuphold(posedge clk,posedge ssb,0.0,0.0,notifier,,,clk_delay,ssb_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d1 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d1 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,d1_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d2 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d2 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,d2_delay);
      
      // setuphold d3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d3 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,d3_delay);
      
      // setuphold d3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d3 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,d3_delay);
      
      // setuphold d4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      negedge d4 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,d4_delay);
      
      // setuphold d4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_ssb_AND_rb == 1'b1),
      posedge d4 &&& (ENABLE_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,d4_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si1 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si1- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si1 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier0,,,clk_delay,si1_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si2 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si2- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si2 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier1,,,clk_delay,si2_delay);
      
      // setuphold si3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si3 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,si3_delay);
      
      // setuphold si3- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si3 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier2,,,clk_delay,si3_delay);
      
      // setuphold si4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      negedge si4 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,si4_delay);
      
      // setuphold si4- clk-LH
      $setuphold(posedge clk &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      posedge si4 &&& (ENABLE_NOT_ssb_AND_rb == 1'b1),
      0.0,0.0,notifier3,,,clk_delay,si4_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_lsn000ah_func( clk, d, o, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_EN0, clk, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, d, vcc, vssx );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, 1'b0, 1'b0, MGM_EN0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_EN0, clk );
   INTCseq_cdiar2ah_0( MGM_D0, d );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, 1'b0, 1'b0, MGM_EN0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15lsn000ah1n02x5( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn000ah_func b15lsn000ah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn000ah_func b15lsn000ah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn000ah_func b15lsn000ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn000ah_func b15lsn000ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lsn000ah1n03x5( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn000ah_func b15lsn000ah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn000ah_func b15lsn000ah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn000ah_func b15lsn000ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn000ah_func b15lsn000ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lsn000ah1n04x5( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn000ah_func b15lsn000ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn000ah_func b15lsn000ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn000ah_func b15lsn000ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn000ah_func b15lsn000ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lsn000ah1n06x5( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn000ah_func b15lsn000ah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn000ah_func b15lsn000ah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn000ah_func b15lsn000ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn000ah_func b15lsn000ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lsn000ah1n08x5( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn000ah_func b15lsn000ah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn000ah_func b15lsn000ah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn000ah_func b15lsn000ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn000ah_func b15lsn000ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lsn000ah1n12x5( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn000ah_func b15lsn000ah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn000ah_func b15lsn000ah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn000ah_func b15lsn000ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn000ah_func b15lsn000ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lsn000ah1n16x5( clk, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn000ah_func b15lsn000ah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn000ah_func b15lsn000ah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn000ah_func b15lsn000ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn000ah_func b15lsn000ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk,negedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk,posedge d,0.0,0.0,notifier,,,clk_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_lsn080ah_func( clkb, d, o, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_1( MGM_EN0, clkb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, d, vcc, vssx );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, 1'b0, 1'b0, MGM_EN0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_1( MGM_EN0, clkb );
   INTCseq_cdiar2ah_0( MGM_D0, d );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, 1'b0, 1'b0, MGM_EN0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15lsn080ah1n02x5( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn080ah_func b15lsn080ah1n02x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn080ah_func b15lsn080ah1n02x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn080ah_func b15lsn080ah1n02x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn080ah_func b15lsn080ah1n02x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lsn080ah1n03x5( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn080ah_func b15lsn080ah1n03x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn080ah_func b15lsn080ah1n03x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn080ah_func b15lsn080ah1n03x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn080ah_func b15lsn080ah1n03x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lsn080ah1n04x5( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn080ah_func b15lsn080ah1n04x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn080ah_func b15lsn080ah1n04x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn080ah_func b15lsn080ah1n04x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn080ah_func b15lsn080ah1n04x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lsn080ah1n06x5( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn080ah_func b15lsn080ah1n06x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn080ah_func b15lsn080ah1n06x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn080ah_func b15lsn080ah1n06x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn080ah_func b15lsn080ah1n06x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lsn080ah1n08x5( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn080ah_func b15lsn080ah1n08x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn080ah_func b15lsn080ah1n08x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn080ah_func b15lsn080ah1n08x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn080ah_func b15lsn080ah1n08x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lsn080ah1n12x5( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn080ah_func b15lsn080ah1n12x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn080ah_func b15lsn080ah1n12x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn080ah_func b15lsn080ah1n12x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn080ah_func b15lsn080ah1n12x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lsn080ah1n16x5( clkb, d, o `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn080ah_func b15lsn080ah1n16x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn080ah_func b15lsn080ah1n16x5_behav_inst(.clkb(clkb),.d(d),.o(o),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lsn080ah_func b15lsn080ah1n16x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lsn080ah_func b15lsn080ah1n16x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(ENABLE_NOT_d,d_delay);
   buf MGM_G1(ENABLE_d,d_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb,negedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb,posedge d,0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_lyn003ah_func( clk, d, o, rb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_EN0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, d, vcc, vssx );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, MGM_C0, 1'b0, MGM_EN0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_EN0, clk );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_cdiar2ah_0( MGM_D0, d );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, MGM_C0, 1'b0, MGM_EN0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15lyn003ah1n02x5( clk, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn003ah_func b15lyn003ah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn003ah_func b15lyn003ah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn003ah_func b15lyn003ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn003ah_func b15lyn003ah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-negedge
      $recrem(posedge rb,negedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn003ah1n03x5( clk, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn003ah_func b15lyn003ah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn003ah_func b15lyn003ah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn003ah_func b15lyn003ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn003ah_func b15lyn003ah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-negedge
      $recrem(posedge rb,negedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn003ah1n04x5( clk, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn003ah_func b15lyn003ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn003ah_func b15lyn003ah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn003ah_func b15lyn003ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn003ah_func b15lyn003ah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-negedge
      $recrem(posedge rb,negedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn003ah1n06x5( clk, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn003ah_func b15lyn003ah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn003ah_func b15lyn003ah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn003ah_func b15lyn003ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn003ah_func b15lyn003ah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-negedge
      $recrem(posedge rb,negedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn003ah1n08x5( clk, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn003ah_func b15lyn003ah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn003ah_func b15lyn003ah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn003ah_func b15lyn003ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn003ah_func b15lyn003ah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-negedge
      $recrem(posedge rb,negedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn003ah1n12x5( clk, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn003ah_func b15lyn003ah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn003ah_func b15lyn003ah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn003ah_func b15lyn003ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn003ah_func b15lyn003ah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-negedge
      $recrem(posedge rb,negedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn003ah1n16x5( clk, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn003ah_func b15lyn003ah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn003ah_func b15lyn003ah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn003ah_func b15lyn003ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn003ah_func b15lyn003ah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem rb-clk-negedge
      $recrem(posedge rb,negedge clk,0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_lyn00cah_func( clk, d, o, psb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_EN0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_P0, psb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, d, vcc, vssx );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, 1'b0, MGM_P0, MGM_EN0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_EN0, clk );
   INTCseq_cdiar2ah_1( MGM_P0, psb );
   INTCseq_cdiar2ah_0( MGM_D0, d );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, 1'b0, MGM_P0, MGM_EN0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15lyn00cah1n02x5( clk, d, o, psb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00cah_func b15lyn00cah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00cah_func b15lyn00cah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00cah_func b15lyn00cah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00cah_func b15lyn00cah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_psb,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_psb,psb_delay,d_delay);
   buf MGM_G3(ENABLE_psb,psb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (posedge psb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb == 1'b1),
      negedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb == 1'b1),
      posedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-negedge
      $recrem(posedge psb,negedge clk,0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn00cah1n03x5( clk, d, o, psb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00cah_func b15lyn00cah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00cah_func b15lyn00cah1n03x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00cah_func b15lyn00cah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00cah_func b15lyn00cah1n03x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_psb,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_psb,psb_delay,d_delay);
   buf MGM_G3(ENABLE_psb,psb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (posedge psb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb == 1'b1),
      negedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb == 1'b1),
      posedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-negedge
      $recrem(posedge psb,negedge clk,0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn00cah1n04x5( clk, d, o, psb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00cah_func b15lyn00cah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00cah_func b15lyn00cah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00cah_func b15lyn00cah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00cah_func b15lyn00cah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_psb,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_psb,psb_delay,d_delay);
   buf MGM_G3(ENABLE_psb,psb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (posedge psb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb == 1'b1),
      negedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb == 1'b1),
      posedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-negedge
      $recrem(posedge psb,negedge clk,0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn00cah1n06x5( clk, d, o, psb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00cah_func b15lyn00cah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00cah_func b15lyn00cah1n06x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00cah_func b15lyn00cah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00cah_func b15lyn00cah1n06x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_psb,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_psb,psb_delay,d_delay);
   buf MGM_G3(ENABLE_psb,psb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (posedge psb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb == 1'b1),
      negedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb == 1'b1),
      posedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-negedge
      $recrem(posedge psb,negedge clk,0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn00cah1n08x5( clk, d, o, psb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00cah_func b15lyn00cah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00cah_func b15lyn00cah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00cah_func b15lyn00cah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00cah_func b15lyn00cah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_psb,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_psb,psb_delay,d_delay);
   buf MGM_G3(ENABLE_psb,psb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (posedge psb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb == 1'b1),
      negedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb == 1'b1),
      posedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-negedge
      $recrem(posedge psb,negedge clk,0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn00cah1n12x5( clk, d, o, psb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00cah_func b15lyn00cah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00cah_func b15lyn00cah1n12x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00cah_func b15lyn00cah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00cah_func b15lyn00cah1n12x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_psb,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_psb,psb_delay,d_delay);
   buf MGM_G3(ENABLE_psb,psb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (posedge psb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb == 1'b1),
      negedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb == 1'b1),
      posedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-negedge
      $recrem(posedge psb,negedge clk,0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn00cah1n16x5( clk, d, o, psb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00cah_func b15lyn00cah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00cah_func b15lyn00cah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00cah_func b15lyn00cah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00cah_func b15lyn00cah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_psb,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_psb,psb_delay,d_delay);
   buf MGM_G3(ENABLE_psb,psb_delay);
   not MGM_G4(MGM_W1,clk_delay);
   not MGM_G5(MGM_W2,d_delay);
   and MGM_G6(ENABLE_NOT_clk_AND_NOT_d,MGM_W2,MGM_W1);
   not MGM_G7(MGM_W3,clk_delay);
   and MGM_G8(ENABLE_NOT_clk_AND_d,d_delay,MGM_W3);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (posedge psb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb == 1'b1),
      negedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb == 1'b1),
      posedge d &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-negedge
      $recrem(posedge psb,negedge clk,0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine


primitive INTCseq_lyn00fah_N_L_IQ_LATCH_UDP( Q, C, P, CK, D `ifdef POWER_AWARE_MODE , vcc, vssx `endif , N );
   output Q;
   reg Q;
   input C, P, CK, D, N; 
   `ifdef POWER_AWARE_MODE
   input vcc, vssx;
   `endif
   table 
  `ifdef POWER_AWARE_MODE
   //C  P  CK D  PW GN N  :  Q  :  Q 
     0  0  0  ?  1  0  ?  :  ?  :  -;
     ?  0  1  0  1  0  ?  :  ?  :  0;
     ?  0  ?  0  1  0  ?  :  0  :  0;
     ?  0  0  ?  1  0  ?  :  0  :  0;
     1  ?  ?  ?  1  0  ?  :  ?  :  0;
     0  ?  1  1  1  0  ?  :  ?  :  1;
     0  ?  ?  1  1  0  ?  :  1  :  1;
     0  ?  0  ?  1  0  ?  :  1  :  1;
     0  1  ?  ?  1  0  ?  :  ?  :  1;
     ?  ?  ?  ?  1  0  *  :  ?  :  x;
  `else
   //C  P  CK D  N  :  Q  :  Q 
     0  0  0  ?  ?  :  ?  :  -;
     ?  0  1  0  ?  :  ?  :  0;
     ?  0  ?  0  ?  :  0  :  0;
     ?  0  0  ?  ?  :  0  :  0;
     1  ?  ?  ?  ?  :  ?  :  0;
     0  ?  1  1  ?  :  ?  :  1;
     0  ?  ?  1  ?  :  1  :  1;
     0  ?  0  ?  ?  :  1  :  1;
     0  1  ?  ?  ?  :  ?  :  1;
     ?  ?  ?  ?  *  :  ?  :  x;
  `endif

endtable
endprimitive



`celldefine
module INTCseq_lyn00fah_func( clk, d, o, psb, rb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_0( MGM_EN0, clk, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_P0, psb, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, d, vcc, vssx );
   INTCseq_lyn00fah_N_L_IQ_LATCH_UDP( IQ, MGM_C0, MGM_P0, MGM_EN0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_0( MGM_EN0, clk );
   INTCseq_cdiar2ah_1( MGM_P0, psb );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_cdiar2ah_0( MGM_D0, d );
   INTCseq_lyn00fah_N_L_IQ_LATCH_UDP( IQ, MGM_C0, MGM_P0, MGM_EN0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15lyn00fah1n02x5( clk, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00fah_func b15lyn00fah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00fah_func b15lyn00fah1n02x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00fah_func b15lyn00fah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00fah_func b15lyn00fah1n02x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clk_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clk_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clk_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,clk_delay);
   not MGM_G15(MGM_W9,d_delay);
   and MGM_G16(ENABLE_NOT_clk_AND_NOT_d,MGM_W9,MGM_W8);
   not MGM_G17(MGM_W10,clk_delay);
   and MGM_G18(ENABLE_NOT_clk_AND_d,d_delay,MGM_W10);
   buf MGM_G19(ENABLE_psb,psb_delay);
   not MGM_G20(MGM_W11,clk_delay);
   not MGM_G21(MGM_W12,d_delay);
   and MGM_G22(MGM_W13,MGM_W12,MGM_W11);
   and MGM_G23(ENABLE_NOT_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W13);
   not MGM_G24(MGM_W14,clk_delay);
   and MGM_G25(MGM_W15,d_delay,MGM_W14);
   and MGM_G26(ENABLE_NOT_clk_AND_d_AND_psb,psb_delay,MGM_W15);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (posedge psb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-negedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      negedge clk &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-negedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      negedge clk &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn00fah1n04x5( clk, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00fah_func b15lyn00fah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00fah_func b15lyn00fah1n04x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00fah_func b15lyn00fah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00fah_func b15lyn00fah1n04x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clk_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clk_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clk_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,clk_delay);
   not MGM_G15(MGM_W9,d_delay);
   and MGM_G16(ENABLE_NOT_clk_AND_NOT_d,MGM_W9,MGM_W8);
   not MGM_G17(MGM_W10,clk_delay);
   and MGM_G18(ENABLE_NOT_clk_AND_d,d_delay,MGM_W10);
   buf MGM_G19(ENABLE_psb,psb_delay);
   not MGM_G20(MGM_W11,clk_delay);
   not MGM_G21(MGM_W12,d_delay);
   and MGM_G22(MGM_W13,MGM_W12,MGM_W11);
   and MGM_G23(ENABLE_NOT_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W13);
   not MGM_G24(MGM_W14,clk_delay);
   and MGM_G25(MGM_W15,d_delay,MGM_W14);
   and MGM_G26(ENABLE_NOT_clk_AND_d_AND_psb,psb_delay,MGM_W15);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (posedge psb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-negedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      negedge clk &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-negedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      negedge clk &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn00fah1n08x5( clk, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00fah_func b15lyn00fah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00fah_func b15lyn00fah1n08x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00fah_func b15lyn00fah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00fah_func b15lyn00fah1n08x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clk_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clk_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clk_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,clk_delay);
   not MGM_G15(MGM_W9,d_delay);
   and MGM_G16(ENABLE_NOT_clk_AND_NOT_d,MGM_W9,MGM_W8);
   not MGM_G17(MGM_W10,clk_delay);
   and MGM_G18(ENABLE_NOT_clk_AND_d,d_delay,MGM_W10);
   buf MGM_G19(ENABLE_psb,psb_delay);
   not MGM_G20(MGM_W11,clk_delay);
   not MGM_G21(MGM_W12,d_delay);
   and MGM_G22(MGM_W13,MGM_W12,MGM_W11);
   and MGM_G23(ENABLE_NOT_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W13);
   not MGM_G24(MGM_W14,clk_delay);
   and MGM_G25(MGM_W15,d_delay,MGM_W14);
   and MGM_G26(ENABLE_NOT_clk_AND_d_AND_psb,psb_delay,MGM_W15);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (posedge psb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-negedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      negedge clk &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-negedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      negedge clk &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn00fah1n16x5( clk, d, o, psb, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clk, d, psb, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00fah_func b15lyn00fah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00fah_func b15lyn00fah1n16x5_behav_inst(.clk(clk),.d(d),.o(o),.psb(psb),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clk_delay ;
   wire d_delay ;
   wire psb_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn00fah_func b15lyn00fah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn00fah_func b15lyn00fah1n16x5_inst(.clk(clk_delay),.d(d_delay),.o(o),.psb(psb_delay),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(MGM_W1,psb_delay,MGM_W0);
   and MGM_G2(ENABLE_NOT_d_AND_psb_AND_rb,rb_delay,MGM_W1);
   and MGM_G3(MGM_W2,psb_delay,d_delay);
   and MGM_G4(ENABLE_d_AND_psb_AND_rb,rb_delay,MGM_W2);
   and MGM_G5(ENABLE_psb_AND_rb,rb_delay,psb_delay);
   buf MGM_G6(ENABLE_rb,rb_delay);
   not MGM_G7(MGM_W3,clk_delay);
   not MGM_G8(MGM_W4,d_delay);
   and MGM_G9(MGM_W5,MGM_W4,MGM_W3);
   and MGM_G10(ENABLE_NOT_clk_AND_NOT_d_AND_rb,rb_delay,MGM_W5);
   not MGM_G11(MGM_W6,clk_delay);
   and MGM_G12(MGM_W7,d_delay,MGM_W6);
   and MGM_G13(ENABLE_NOT_clk_AND_d_AND_rb,rb_delay,MGM_W7);
   not MGM_G14(MGM_W8,clk_delay);
   not MGM_G15(MGM_W9,d_delay);
   and MGM_G16(ENABLE_NOT_clk_AND_NOT_d,MGM_W9,MGM_W8);
   not MGM_G17(MGM_W10,clk_delay);
   and MGM_G18(ENABLE_NOT_clk_AND_d,d_delay,MGM_W10);
   buf MGM_G19(ENABLE_psb,psb_delay);
   not MGM_G20(MGM_W11,clk_delay);
   not MGM_G21(MGM_W12,d_delay);
   and MGM_G22(MGM_W13,MGM_W12,MGM_W11);
   and MGM_G23(ENABLE_NOT_clk_AND_NOT_d_AND_psb,psb_delay,MGM_W13);
   not MGM_G24(MGM_W14,clk_delay);
   and MGM_G25(MGM_W15,d_delay,MGM_W14);
   and MGM_G26(ENABLE_NOT_clk_AND_d_AND_psb,psb_delay,MGM_W15);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b0 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(d==1'b1 && psb==1'b1 && rb==1'b1)
      // seq arc clk --> o
      (posedge clk => (o : d))  = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b1 && psb==1'b1 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (posedge psb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && rb==1'b1)
      // seq arc psb --> o
      (negedge psb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b0 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b0 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b0 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b0)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clk==1'b1 && d==1'b1 && psb==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      $width(posedge clk &&& (ENABLE_NOT_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(posedge clk &&& (ENABLE_d_AND_psb_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      negedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // setuphold d- clk-HL
      $setuphold(negedge clk &&& (ENABLE_psb_AND_rb == 1'b1),
      posedge d &&& (ENABLE_psb_AND_rb == 1'b1),
      0.0,0.0,notifier,,,clk_delay,d_delay);
      
      // recrem psb-clk-negedge
      $recrem(posedge psb &&& (ENABLE_rb == 1'b1),
      negedge clk &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,psb_delay,clk_delay);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge psb &&& (ENABLE_NOT_clk_AND_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // setuphold psb- rb-LH
      $setuphold(posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,rb_delay,psb_delay);
      
      // recrem rb-clk-negedge
      $recrem(posedge rb &&& (ENABLE_psb == 1'b1),
      negedge clk &&& (ENABLE_psb == 1'b1),
      0.0,0.0,notifier,,,rb_delay,clk_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_NOT_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      // setuphold rb- psb-LH
      $setuphold(posedge psb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      posedge rb &&& (ENABLE_NOT_clk_AND_d == 1'b1),
      0.0,0.0,notifier,,,psb_delay,rb_delay);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_NOT_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_NOT_clk_AND_d_AND_psb == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine



`celldefine
module INTCseq_lyn083ah_func( clkb, d, o, rb, notifier `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, rb, notifier;
   output o;
`ifdef POWER_AWARE_MODE
   inout  vcc;
   inout  vssx;
`endif

`ifdef POWER_AWARE_MODE
   INTCseq_cdiar2ah_1( MGM_EN0, clkb, vcc, vssx );
   INTCseq_cdiar2ah_1( MGM_C0, rb, vcc, vssx );
   INTCseq_cdiar2ah_0( MGM_D0, d, vcc, vssx );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, MGM_C0, 1'b0, MGM_EN0, MGM_D0, vcc, vssx, notifier );
   INTCseq_cdiar2ah_0( o, IQ, vcc, vssx );
`else
   INTCseq_cdiar2ah_1( MGM_EN0, clkb );
   INTCseq_cdiar2ah_1( MGM_C0, rb );
   INTCseq_cdiar2ah_0( MGM_D0, d );
   INTCseq_cilao5ah_N_IQ_LATCH_UDP( IQ, MGM_C0, 1'b0, MGM_EN0, MGM_D0, notifier );
   INTCseq_cdiar2ah_0( o, IQ );
`endif

endmodule
`endcelldefine



`celldefine
module b15lyn083ah1n02x5( clkb, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn083ah_func b15lyn083ah1n02x5_behav_inst(.clkb(clkb),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn083ah_func b15lyn083ah1n02x5_behav_inst(.clkb(clkb),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn083ah_func b15lyn083ah1n02x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn083ah_func b15lyn083ah1n02x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,d_delay);
   and MGM_G5(ENABLE_clkb_AND_NOT_d,MGM_W1,clkb_delay);
   and MGM_G6(ENABLE_clkb_AND_d,d_delay,clkb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem rb-clkb-posedge
      $recrem(posedge rb,posedge clkb,0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn083ah1n03x5( clkb, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn083ah_func b15lyn083ah1n03x5_behav_inst(.clkb(clkb),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn083ah_func b15lyn083ah1n03x5_behav_inst(.clkb(clkb),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn083ah_func b15lyn083ah1n03x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn083ah_func b15lyn083ah1n03x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,d_delay);
   and MGM_G5(ENABLE_clkb_AND_NOT_d,MGM_W1,clkb_delay);
   and MGM_G6(ENABLE_clkb_AND_d,d_delay,clkb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem rb-clkb-posedge
      $recrem(posedge rb,posedge clkb,0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn083ah1n04x5( clkb, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn083ah_func b15lyn083ah1n04x5_behav_inst(.clkb(clkb),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn083ah_func b15lyn083ah1n04x5_behav_inst(.clkb(clkb),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn083ah_func b15lyn083ah1n04x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn083ah_func b15lyn083ah1n04x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,d_delay);
   and MGM_G5(ENABLE_clkb_AND_NOT_d,MGM_W1,clkb_delay);
   and MGM_G6(ENABLE_clkb_AND_d,d_delay,clkb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem rb-clkb-posedge
      $recrem(posedge rb,posedge clkb,0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn083ah1n06x5( clkb, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn083ah_func b15lyn083ah1n06x5_behav_inst(.clkb(clkb),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn083ah_func b15lyn083ah1n06x5_behav_inst(.clkb(clkb),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn083ah_func b15lyn083ah1n06x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn083ah_func b15lyn083ah1n06x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,d_delay);
   and MGM_G5(ENABLE_clkb_AND_NOT_d,MGM_W1,clkb_delay);
   and MGM_G6(ENABLE_clkb_AND_d,d_delay,clkb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem rb-clkb-posedge
      $recrem(posedge rb,posedge clkb,0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn083ah1n08x5( clkb, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn083ah_func b15lyn083ah1n08x5_behav_inst(.clkb(clkb),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn083ah_func b15lyn083ah1n08x5_behav_inst(.clkb(clkb),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn083ah_func b15lyn083ah1n08x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn083ah_func b15lyn083ah1n08x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,d_delay);
   and MGM_G5(ENABLE_clkb_AND_NOT_d,MGM_W1,clkb_delay);
   and MGM_G6(ENABLE_clkb_AND_d,d_delay,clkb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem rb-clkb-posedge
      $recrem(posedge rb,posedge clkb,0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn083ah1n12x5( clkb, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn083ah_func b15lyn083ah1n12x5_behav_inst(.clkb(clkb),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn083ah_func b15lyn083ah1n12x5_behav_inst(.clkb(clkb),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn083ah_func b15lyn083ah1n12x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn083ah_func b15lyn083ah1n12x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,d_delay);
   and MGM_G5(ENABLE_clkb_AND_NOT_d,MGM_W1,clkb_delay);
   and MGM_G6(ENABLE_clkb_AND_d,d_delay,clkb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem rb-clkb-posedge
      $recrem(posedge rb,posedge clkb,0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine





`celldefine
module b15lyn083ah1n16x5( clkb, d, o, rb `ifdef POWER_AWARE_MODE , vcc, vssx `endif );
   input clkb, d, rb;
   output o;
`ifdef POWER_AWARE_MODE
   (* pg_type = "primary_power" *) inout vcc;
   (* pg_type = "primary_ground" *) inout vssx;
`endif

`ifdef FUNCTIONAL  //  functional //
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn083ah_func b15lyn083ah1n16x5_behav_inst(.clkb(clkb),.d(d),.o(o),.rb(rb),.notifier(1'b0),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn083ah_func b15lyn083ah1n16x5_behav_inst(.clkb(clkb),.d(d),.o(o),.rb(rb),.notifier(1'b0));
      
   `endif
   
`else
   wire clkb_delay ;
   wire d_delay ;
   wire rb_delay ;
   reg notifier;
   
   `ifdef POWER_AWARE_MODE
      INTCseq_lyn083ah_func b15lyn083ah1n16x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier),.vcc(vcc),.vssx(vssx));
   `else
      INTCseq_lyn083ah_func b15lyn083ah1n16x5_inst(.clkb(clkb_delay),.d(d_delay),.o(o),.rb(rb_delay),.notifier(notifier));
   `endif
   
   // spec_gates_begin
   not MGM_G0(MGM_W0,d_delay);
   and MGM_G1(ENABLE_NOT_d_AND_rb,rb_delay,MGM_W0);
   and MGM_G2(ENABLE_d_AND_rb,rb_delay,d_delay);
   buf MGM_G3(ENABLE_rb,rb_delay);
   not MGM_G4(MGM_W1,d_delay);
   and MGM_G5(ENABLE_clkb_AND_NOT_d,MGM_W1,clkb_delay);
   and MGM_G6(ENABLE_clkb_AND_d,d_delay,clkb_delay);
   // spec_gates_end
   specify


   // specify_block_begin
      if(d==1'b1 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(d==1'b0 && rb==1'b1)
      // seq arc clkb --> o
      (negedge clkb => (o : d))  = (0.0,0.0);
      
      if(clkb==1'b0 && rb==1'b1)
      // comb arc negedge d --> o
      (negedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0 && rb==1'b1)
      // comb arc posedge d --> o
      (posedge d => (o:d)) = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b0 && d==1'b1)
      // seq arc rb --> o
      (posedge rb => (o +: 1'b1))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b0)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      if(clkb==1'b1 && d==1'b1)
      // seq arc rb --> o
      (negedge rb => (o +: 1'b0))  = (0.0,0.0);
      
      $width(negedge clkb &&& (ENABLE_NOT_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge clkb &&& (ENABLE_d_AND_rb == 1'b1)
      ,0.0,0,notifier);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb &&& (ENABLE_rb == 1'b1),
      negedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // setuphold d- clkb-LH
      $setuphold(posedge clkb &&& (ENABLE_rb == 1'b1),
      posedge d &&& (ENABLE_rb == 1'b1),
      0.0,0.0,notifier,,,clkb_delay,d_delay);
      
      // recrem rb-clkb-posedge
      $recrem(posedge rb,posedge clkb,0.0,0.0,notifier,,,rb_delay,clkb_delay);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_NOT_d == 1'b1)
      ,0.0,0,notifier);
      
      $width(negedge rb &&& (ENABLE_clkb_AND_d == 1'b1)
      ,0.0,0,notifier);
      
      
   // specify_block_end 
   endspecify

`endif 


endmodule
`endcelldefine
