module pll (

);

ringpll u_ringpll (
    .clkpll, 
    .clkpll0, 
    .clkpll1, 
    .idvdisable_bo, 
    .idvfreqao, 
    .idvfreqbo, 
    .idvpulseo, 
    .idvtclko, 
    .idvtctrlo, 
    .idvtdo, 
    .idvtreso, 
    .lock, 
    .odfx_fscan_sdo, 
    .tdo, 
    .view_dig_out, 
    .viewanabus, 
    .bypass, 
    .clkpostdist, 
    .clkref, 
    .fraction, 
    .fz_cp1trim, 
    .fz_cp2trim, 
    .fz_cpnbias, 
    .fz_dca_cb, 
    .fz_dca_ctrl, 
    .fz_irefgen, 
    .fz_ldo_bypass, 
    .fz_ldo_extrefsel, 
    .fz_ldo_faststart, 
    .fz_ldo_fbtrim, 
    .fz_ldo_reftrim, 
    .fz_ldo_vinvoltsel, 
    .fz_lockcnt, 
    .fz_lockforce, 
    .fz_lockstickyb, 
    .fz_lockthresh, 
    .fz_lpfclksel, 
    .fz_nopfdpwrgate, 
    .fz_pfd_pw, 
    .fz_pfddly, 
    .fz_skadj, 
    .fz_spare, 
    .fz_startup, 
    .fz_tight_loopb, 
    .fz_vcosel, 
    .fz_vcotrim, 
    .idfx_fscan_byprstb, 
    .idfx_fscan_clkungate,
    .idfx_fscan_mode, 
    .idfx_fscan_rstbypen, 
    .idfx_fscan_sdi, 
    .idfx_fscan_shiften, 
    .idvdisable_bi, 
    .idvfreqai, 
    .idvfreqbi, 
    .idvpulsei, 
    .idvtclki, 
    .idvtctrli, 
    .idvtdi, 
    .idvtresi, 
    .ldo_enable, 
    .ldo_vref, 
    .mash_order_plus_one, 
    .mdiv_ratio, 
    .pllen, 
    .pllfwen_b, 
    .powergood_vnn, 
    .ratio, 
    .ssc_cyc_to_peak_m1, 
    .ssc_en, 
    .ssc_frac_step, 
    .tcapturedr, 
    .tck, 
    .tdi, 
    .treg_en, 
    .trst_n, 
    .tshiftdr, 
    .tupdatedr, 
    .vccdig_nom,
    .vccdist_nom, 
    .vccldo_hv, 
    .vcodiv_ratio, 
    .vnnaon_nom, 
    .vss, 
    .zdiv0_ratio, 
    .zdiv0_ratio_p5, 
    .zdiv1_ratio, 
    .zdiv1_ratio_p5
);

endmodule