module Noise_injection_block_Stuck (
    Random,
    S,
    VB,
    Iout
);

input Random;
input [15:0] S;
input [3:0] VB;
output Iout;

endmodule