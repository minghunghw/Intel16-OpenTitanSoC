module dummy_stub();

endmodule
