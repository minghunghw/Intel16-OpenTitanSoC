module sandbox (
   
)

endmodule