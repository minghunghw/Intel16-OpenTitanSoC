module peri_device (clk_i,
    rst_ni,
    gpio_o,
    tl_peri_device_i,
    tl_peri_device_o);
 input clk_i;
 input rst_ni;
 output [31:0] gpio_o;
 input [108:0] tl_peri_device_i;
 output [65:0] tl_peri_device_o;

 wire eq_x_101_n25;
 wire eq_x_106_n25;
 wire eq_x_111_n25;
 wire eq_x_116_n25;
 wire eq_x_121_n25;
 wire eq_x_126_n25;
 wire eq_x_131_n25;
 wire eq_x_136_n25;
 wire eq_x_141_n25;
 wire eq_x_146_n25;
 wire eq_x_151_n25;
 wire eq_x_156_n25;
 wire eq_x_161_n25;
 wire eq_x_166_n25;
 wire eq_x_171_n25;
 wire eq_x_176_n25;
 wire eq_x_181_n25;
 wire eq_x_186_n25;
 wire eq_x_191_n25;
 wire eq_x_196_n25;
 wire eq_x_201_n25;
 wire eq_x_206_n25;
 wire eq_x_211_n25;
 wire eq_x_216_n25;
 wire eq_x_221_n25;
 wire eq_x_226_n25;
 wire eq_x_231_n25;
 wire eq_x_76_n25;
 wire eq_x_81_n25;
 wire eq_x_86_n25;
 wire eq_x_91_n25;
 wire eq_x_96_n25;
 wire n1435;
 wire n1438;
 wire n1443;
 wire n1446;
 wire n1451;
 wire n1454;
 wire n1527;
 wire n1530;
 wire n2628;
 wire n2629;
 wire n2630;
 wire n2631;
 wire n2632;
 wire n2633;
 wire n2634;
 wire n2635;
 wire n2636;
 wire n2637;
 wire n2638;
 wire n2639;
 wire n2644;
 wire n2645;
 wire n2646;
 wire n2647;
 wire n2648;
 wire n2649;
 wire n2650;
 wire n2651;
 wire n2652;
 wire n2653;
 wire n2654;
 wire n2655;
 wire n2656;
 wire n2657;
 wire n2658;
 wire n2659;
 wire n2660;
 wire n2661;
 wire n2662;
 wire n2663;
 wire n2664;
 wire n2665;
 wire n2666;
 wire n2667;
 wire n2668;
 wire n2669;
 wire n2670;
 wire n2671;
 wire n2672;
 wire n2673;
 wire n2674;
 wire n2675;
 wire n2676;
 wire n2677;
 wire n2678;
 wire n2679;
 wire n2680;
 wire n2681;
 wire n2682;
 wire n2683;
 wire n2684;
 wire n2685;
 wire n2686;
 wire n2687;
 wire n2688;
 wire n2689;
 wire n2690;
 wire n2691;
 wire n2692;
 wire n2693;
 wire n2694;
 wire n2695;
 wire n2696;
 wire n2697;
 wire n2698;
 wire n2699;
 wire n2700;
 wire n2701;
 wire n2702;
 wire n2703;
 wire n2704;
 wire n2705;
 wire n2706;
 wire n2707;
 wire n2708;
 wire n2709;
 wire n2710;
 wire n2711;
 wire n2712;
 wire n2713;
 wire n2714;
 wire n2715;
 wire n2716;
 wire n2717;
 wire n2718;
 wire n2719;
 wire n2720;
 wire n2721;
 wire n2722;
 wire n2723;
 wire n2724;
 wire n2725;
 wire n2726;
 wire n2727;
 wire n2728;
 wire n2729;
 wire n2730;
 wire n2731;
 wire n2732;
 wire n2733;
 wire n2734;
 wire n2735;
 wire n2736;
 wire n2737;
 wire n2738;
 wire n2739;
 wire n2740;
 wire n2741;
 wire n2742;
 wire n2743;
 wire n2744;
 wire n2745;
 wire n2746;
 wire n2747;
 wire n2748;
 wire n2749;
 wire n2750;
 wire n2751;
 wire n2752;
 wire n2753;
 wire n2754;
 wire n2755;
 wire n2756;
 wire n2757;
 wire n2758;
 wire n2759;
 wire n2760;
 wire n2761;
 wire n2762;
 wire n2763;
 wire n2764;
 wire n2765;
 wire n2766;
 wire n2767;
 wire n2768;
 wire n2769;
 wire n2770;
 wire n2771;
 wire n2772;
 wire n2773;
 wire n2774;
 wire n2775;
 wire n2776;
 wire n2777;
 wire n2778;
 wire n2779;
 wire n2780;
 wire n2781;
 wire n2782;
 wire n2783;
 wire n2784;
 wire n2785;
 wire n2786;
 wire n2787;
 wire n2788;
 wire n2789;
 wire n2790;
 wire n2791;
 wire n2792;
 wire n2793;
 wire n2794;
 wire n2795;
 wire n2796;
 wire n2797;
 wire n2798;
 wire n2799;
 wire n2800;
 wire n2801;
 wire n2802;
 wire n2803;
 wire n2804;
 wire n2805;
 wire n2806;
 wire n2807;
 wire n2808;
 wire n2809;
 wire n2810;
 wire n2811;
 wire n2812;
 wire n2813;
 wire n2814;
 wire n2815;
 wire n2816;
 wire n2817;
 wire n2818;
 wire n2819;
 wire n2820;
 wire n2821;
 wire n2822;
 wire n2823;
 wire n2824;
 wire n2825;
 wire n2826;
 wire n2827;
 wire n2828;
 wire n2829;
 wire n2830;
 wire n2831;
 wire n2832;
 wire n2833;
 wire n2834;
 wire n2835;
 wire n2836;
 wire n2837;
 wire n2838;
 wire n2839;
 wire n2840;
 wire n2841;
 wire n2842;
 wire n2843;
 wire n2844;
 wire n2845;
 wire n2846;
 wire n2847;
 wire n2848;
 wire n2849;
 wire n2850;
 wire n2851;
 wire n2852;
 wire n2853;
 wire n2854;
 wire n2855;
 wire n2856;
 wire n2857;
 wire n2858;
 wire n2859;
 wire n2860;
 wire n2861;
 wire n2862;
 wire n2863;
 wire n2864;
 wire n2865;
 wire n2866;
 wire n2867;
 wire n2868;
 wire n2869;
 wire n2870;
 wire n2871;
 wire n2872;
 wire n2873;
 wire n2874;
 wire n2875;
 wire n2876;
 wire n2877;
 wire n2878;
 wire n2879;
 wire n2880;
 wire n2881;
 wire n2882;
 wire n2883;
 wire n2884;
 wire n2885;
 wire n2886;
 wire n2887;
 wire n2888;
 wire n2889;
 wire n2890;
 wire n2891;
 wire n2892;
 wire n2893;
 wire n2894;
 wire n2895;
 wire n2896;
 wire n2897;
 wire n2898;
 wire n2899;
 wire n2900;
 wire n2901;
 wire n2902;
 wire n2903;
 wire n2904;
 wire n2905;
 wire n2906;
 wire n2907;
 wire n2908;
 wire n2909;
 wire n2910;
 wire n2911;
 wire n2912;
 wire n2913;
 wire n2914;
 wire n2915;
 wire n2916;
 wire n2917;
 wire n2918;
 wire n2919;
 wire n2920;
 wire n2921;
 wire n2922;
 wire n2923;
 wire n2924;
 wire n2925;
 wire n2926;
 wire n2927;
 wire n2928;
 wire n2929;
 wire n2930;
 wire n2931;
 wire n2932;
 wire n2933;
 wire n2934;
 wire n2935;
 wire n2936;
 wire n2937;
 wire n2938;
 wire n2939;
 wire n2940;
 wire n2941;
 wire n2942;
 wire n2943;
 wire n2944;
 wire n2945;
 wire n2946;
 wire n2947;
 wire n2948;
 wire n2949;
 wire n2950;
 wire n2951;
 wire n2952;
 wire n2953;
 wire n2954;
 wire n2955;
 wire n2956;
 wire n2957;
 wire n2958;
 wire n2959;
 wire n2960;
 wire n2961;
 wire n2962;
 wire n2963;
 wire n2964;
 wire n2965;
 wire n2966;
 wire n2967;
 wire n2968;
 wire n2969;
 wire n2970;
 wire n2971;
 wire n2972;
 wire n2973;
 wire n2974;
 wire n2975;
 wire n2976;
 wire n2977;
 wire n2978;
 wire n2979;
 wire n2980;
 wire n2981;
 wire n2982;
 wire n2983;
 wire n2984;
 wire n2985;
 wire n2986;
 wire n2987;
 wire n2988;
 wire n2989;
 wire n2990;
 wire n2991;
 wire n2992;
 wire n2993;
 wire n2994;
 wire n2995;
 wire n2996;
 wire n2997;
 wire n2998;
 wire n2999;
 wire n3000;
 wire n3001;
 wire n3002;
 wire n3003;
 wire n3004;
 wire n3005;
 wire n3006;
 wire n3007;
 wire n3008;
 wire n3009;
 wire n3010;
 wire n3011;
 wire n3012;
 wire n3013;
 wire n3014;
 wire n3015;
 wire n3016;
 wire n3017;
 wire n3018;
 wire n3019;
 wire n3020;
 wire n3021;
 wire n3022;
 wire n3023;
 wire n3024;
 wire n3025;
 wire n3026;
 wire n3027;
 wire n3028;
 wire n3029;
 wire n3030;
 wire n3031;
 wire n3032;
 wire n3033;
 wire n3034;
 wire n3035;
 wire n3036;
 wire n3037;
 wire n3038;
 wire n3039;
 wire n3040;
 wire n3041;
 wire n3042;
 wire n3043;
 wire n3044;
 wire n3045;
 wire n3046;
 wire n3047;
 wire n3049;
 wire n3050;
 wire n3051;
 wire n3052;
 wire n3053;
 wire n3054;
 wire n3055;
 wire n3056;
 wire n3057;
 wire n3058;
 wire n3059;
 wire n3060;
 wire n3061;
 wire n3063;
 wire n3064;
 wire n3065;
 wire n3066;
 wire n3067;
 wire n3068;
 wire n3069;
 wire n3070;
 wire n3072;
 wire n3073;
 wire n3074;
 wire n3075;
 wire n3076;
 wire n3078;
 wire n3079;
 wire n3080;
 wire n3082;
 wire n3083;
 wire n3084;
 wire n3085;
 wire n3086;
 wire n3087;
 wire n3088;
 wire n3089;
 wire n3090;
 wire n3091;
 wire n3092;
 wire n3093;
 wire n3095;
 wire n3096;
 wire n3098;
 wire n3099;
 wire n3100;
 wire n3102;
 wire n3105;
 wire n3106;
 wire n3107;
 wire n3120;
 wire n3129;
 wire n3131;
 wire n3132;
 wire n3133;
 wire n3134;
 wire n3135;
 wire n3137;
 wire n3138;
 wire n3139;
 wire n3140;
 wire n3141;
 wire n3142;
 wire n3143;
 wire n3144;
 wire n3145;
 wire n3146;
 wire n3147;
 wire n3148;
 wire n3149;
 wire n3151;
 wire n3152;
 wire n3154;
 wire n3155;
 wire n3156;
 wire n3157;
 wire n3158;
 wire n3159;
 wire n3161;
 wire n3162;
 wire n3163;
 wire n3164;
 wire n3166;
 wire n3167;
 wire n3168;
 wire n3169;
 wire n3170;
 wire n3171;
 wire n3173;
 wire n3174;
 wire n3175;
 wire n3176;
 wire n3177;
 wire n3178;
 wire n3179;
 wire n3180;
 wire n3181;
 wire n3182;
 wire n3183;
 wire n3184;
 wire n3185;
 wire n3186;
 wire n3187;
 wire n3188;
 wire n3189;
 wire n3190;
 wire n3191;
 wire n3192;
 wire n3193;
 wire n3194;
 wire n3195;
 wire n3196;
 wire n3199;
 wire n3200;
 wire n3201;
 wire n3202;
 wire n3203;
 wire n3204;
 wire n3206;
 wire n3207;
 wire n3209;
 wire n3210;
 wire n3211;
 wire n3212;
 wire n3213;
 wire n3214;
 wire n3215;
 wire n3216;
 wire n3217;
 wire n3218;
 wire n3219;
 wire n3220;
 wire n3221;
 wire n3222;
 wire n3223;
 wire n3224;
 wire n3225;
 wire n3226;
 wire n3227;
 wire n3228;
 wire n3229;
 wire n3230;
 wire n3231;
 wire n3232;
 wire n3233;
 wire n3234;
 wire n3235;
 wire n3236;
 wire n3237;
 wire n3238;
 wire n3240;
 wire n3241;
 wire n3242;
 wire n3243;
 wire n3245;
 wire n3246;
 wire n3247;
 wire n3248;
 wire n3249;
 wire n3250;
 wire n3252;
 wire n3253;
 wire n3254;
 wire n3256;
 wire n3257;
 wire n3258;
 wire n3259;
 wire n3260;
 wire n3261;
 wire n3262;
 wire n3263;
 wire n3264;
 wire n3265;
 wire n3266;
 wire n3267;
 wire n3268;
 wire n3269;
 wire n3270;
 wire n3271;
 wire n3272;
 wire n3273;
 wire n3274;
 wire n3276;
 wire n3277;
 wire n3278;
 wire n3279;
 wire n3280;
 wire n3281;
 wire n3282;
 wire n3283;
 wire n3284;
 wire n3285;
 wire n3286;
 wire n3287;
 wire n3288;
 wire n3289;
 wire n3290;
 wire n3291;
 wire n3292;
 wire n3293;
 wire n3294;
 wire n3296;
 wire n3297;
 wire n3298;
 wire n3299;
 wire n3300;
 wire n3301;
 wire n3302;
 wire n3303;
 wire n3304;
 wire n3305;
 wire n3306;
 wire n3307;
 wire n3308;
 wire n3309;
 wire n3310;
 wire n3311;
 wire n3313;
 wire n3314;
 wire n3315;
 wire n3316;
 wire n3317;
 wire n3318;
 wire n3319;
 wire n3320;
 wire n3321;
 wire n3322;
 wire n3323;
 wire n3324;
 wire n3325;
 wire n3326;
 wire n3327;
 wire n3328;
 wire n3330;
 wire n3331;
 wire n3332;
 wire n3333;
 wire n3334;
 wire n3335;
 wire n3336;
 wire n3337;
 wire n3338;
 wire n3339;
 wire n3340;
 wire n3341;
 wire n3343;
 wire n3344;
 wire n3345;
 wire n3346;
 wire n3347;
 wire n3348;
 wire n3349;
 wire n3350;
 wire n3351;
 wire n3352;
 wire n3353;
 wire n3354;
 wire n3355;
 wire n3356;
 wire n3357;
 wire n3358;
 wire n3359;
 wire n3360;
 wire n3361;
 wire n3362;
 wire n3363;
 wire n3364;
 wire n3365;
 wire n3366;
 wire n3367;
 wire n3369;
 wire n3370;
 wire n3371;
 wire n3372;
 wire n3373;
 wire n3374;
 wire n3375;
 wire n3376;
 wire n3377;
 wire n3378;
 wire n3379;
 wire n3380;
 wire n3381;
 wire n3382;
 wire n3383;
 wire n3384;
 wire n3385;
 wire n3386;
 wire n3387;
 wire n3388;
 wire n3389;
 wire n3390;
 wire n3391;
 wire n3392;
 wire n3393;
 wire n3394;
 wire n3395;
 wire n3396;
 wire n3397;
 wire n3398;
 wire n3399;
 wire n3400;
 wire n3401;
 wire n3402;
 wire n3403;
 wire n3404;
 wire n3405;
 wire n3406;
 wire n3407;
 wire n3408;
 wire n3409;
 wire n3410;
 wire n3411;
 wire n3412;
 wire n3413;
 wire n3414;
 wire n3415;
 wire n3416;
 wire n3417;
 wire n3418;
 wire n3419;
 wire n3420;
 wire n3421;
 wire n3422;
 wire n3423;
 wire n3424;
 wire n3425;
 wire n3426;
 wire n3427;
 wire n3428;
 wire n3429;
 wire n3431;
 wire n3432;
 wire n3433;
 wire n3434;
 wire n3435;
 wire n3436;
 wire n3437;
 wire n3438;
 wire n3439;
 wire n3440;
 wire n3441;
 wire n3442;
 wire n3443;
 wire n3444;
 wire n3445;
 wire n3446;
 wire n3447;
 wire n3448;
 wire n3449;
 wire n3450;
 wire n3451;
 wire n3452;
 wire n3454;
 wire n3455;
 wire n3456;
 wire n3457;
 wire n3458;
 wire n3459;
 wire n3460;
 wire n3461;
 wire n3462;
 wire n3463;
 wire n3464;
 wire n3465;
 wire n3466;
 wire n3467;
 wire n3468;
 wire n3469;
 wire n3470;
 wire n3471;
 wire n3472;
 wire n3473;
 wire n3474;
 wire n3475;
 wire n3476;
 wire n3477;
 wire n3478;
 wire n3479;
 wire n3480;
 wire n3481;
 wire n3482;
 wire n3483;
 wire n3484;
 wire n3485;
 wire n3486;
 wire n3487;
 wire n3488;
 wire n3489;
 wire n3490;
 wire n3491;
 wire n3492;
 wire n3493;
 wire n3494;
 wire n3495;
 wire n3496;
 wire n3497;
 wire n3498;
 wire n3499;
 wire n3500;
 wire n3501;
 wire n3503;
 wire n3504;
 wire n3505;
 wire n3506;
 wire n3507;
 wire n3508;
 wire n3509;
 wire n3510;
 wire n3511;
 wire n3512;
 wire n3513;
 wire n3514;
 wire n3515;
 wire n3516;
 wire n3517;
 wire n3518;
 wire n3519;
 wire n3520;
 wire n3521;
 wire n3522;
 wire n3523;
 wire n3524;
 wire n3525;
 wire n3526;
 wire n3529;
 wire n3530;
 wire n3540;
 wire n3541;
 wire n3542;
 wire n3544;
 wire n3545;
 wire n3546;
 wire n3547;
 wire n3548;
 wire n3549;
 wire n3550;
 wire n3551;
 wire n3552;
 wire n3553;
 wire n3554;
 wire n3555;
 wire n3557;
 wire n3567;
 wire n3568;
 wire n3569;
 wire n3570;
 wire n3571;
 wire n3572;
 wire n3573;
 wire n3574;
 wire n3575;
 wire n3576;
 wire n3577;
 wire n3578;
 wire n3580;
 wire n3581;
 wire n3582;
 wire n3583;
 wire n3584;
 wire n3585;
 wire n3586;
 wire n3587;
 wire n3588;
 wire n3589;
 wire n3590;
 wire n3591;
 wire n3592;
 wire n3593;
 wire n3594;
 wire n3595;
 wire n3596;
 wire n3597;
 wire n3598;
 wire n3599;
 wire n3600;
 wire n3601;
 wire n3602;
 wire n3603;
 wire n3604;
 wire n3605;
 wire n3606;
 wire n3607;
 wire n3608;
 wire n3609;
 wire n3610;
 wire n3611;
 wire n3612;
 wire n3613;
 wire n3614;
 wire n3615;
 wire n3616;
 wire n3617;
 wire n3618;
 wire n3619;
 wire n3620;
 wire n3621;
 wire n3622;
 wire n3623;
 wire n3624;
 wire n3625;
 wire n3626;
 wire n3627;
 wire n3628;
 wire n3629;
 wire n3630;
 wire n3631;
 wire n3632;
 wire n3633;
 wire n3634;
 wire n3635;
 wire n3636;
 wire n3637;
 wire n3638;
 wire n3640;
 wire n3641;
 wire n3642;
 wire n3643;
 wire n3644;
 wire n3645;
 wire n3646;
 wire n3648;
 wire n3649;
 wire n3650;
 wire n3651;
 wire n3652;
 wire n3653;
 wire n3654;
 wire n3655;
 wire n3656;
 wire n3657;
 wire n3658;
 wire n3659;
 wire n3660;
 wire n3661;
 wire n3662;
 wire n3663;
 wire n3664;
 wire n3665;
 wire n3667;
 wire n3668;
 wire n3669;
 wire n3670;
 wire n3671;
 wire n3672;
 wire n3673;
 wire n3674;
 wire n3675;
 wire n3676;
 wire n3677;
 wire n3678;
 wire n3679;
 wire n3680;
 wire n3681;
 wire n3682;
 wire n3683;
 wire n3684;
 wire n3685;
 wire n3686;
 wire n3687;
 wire n3688;
 wire n3689;
 wire n3690;
 wire n3691;
 wire n3692;
 wire n3693;
 wire n3694;
 wire n3695;
 wire n3696;
 wire n3697;
 wire n3698;
 wire n3699;
 wire n3700;
 wire n3701;
 wire n3702;
 wire n3703;
 wire n3704;
 wire n3705;
 wire n3706;
 wire n3707;
 wire n3708;
 wire n3709;
 wire n3710;
 wire n3711;
 wire n3712;
 wire n3713;
 wire n3714;
 wire n3715;
 wire n3716;
 wire n3717;
 wire n3718;
 wire n3719;
 wire n3720;
 wire n3721;
 wire n3722;
 wire n3724;
 wire n3725;
 wire n3726;
 wire n3727;
 wire n3728;
 wire n3729;
 wire n3730;
 wire n3732;
 wire n3733;
 wire n3734;
 wire n3735;
 wire n3736;
 wire n3737;
 wire n3738;
 wire n3739;
 wire n3740;
 wire n3741;
 wire n3742;
 wire n3744;
 wire n3745;
 wire n3746;
 wire n3747;
 wire n3748;
 wire n3749;
 wire n3750;
 wire n3752;
 wire n3753;
 wire n3754;
 wire n3755;
 wire n3756;
 wire n3757;
 wire n3758;
 wire n3759;
 wire n3760;
 wire n3761;
 wire n3762;
 wire n3763;
 wire n3764;
 wire n3767;
 wire n3768;
 wire n3769;
 wire n3770;
 wire n3771;
 wire n3772;
 wire n3773;
 wire n3774;
 wire n3777;
 wire n3778;
 wire n3779;
 wire n3780;
 wire n3784;
 wire n3785;
 wire n3787;
 wire n3788;
 wire n3789;
 wire n3790;
 wire n3797;
 wire n3798;
 wire n3799;
 wire n3801;
 wire n3804;
 wire n3805;
 wire n3806;
 wire n3807;
 wire n3808;
 wire n3809;
 wire n3810;
 wire n3811;
 wire n3812;
 wire n3813;
 wire n3814;
 wire n3815;
 wire n3816;
 wire n3817;
 wire n3818;
 wire n3819;
 wire n3829;
 wire n3831;
 wire n3891;
 wire n3892;
 wire n3893;
 wire n3894;
 wire n3895;
 wire n3896;
 wire n3897;
 wire n3898;
 wire n3899;
 wire n3900;
 wire n3901;
 wire n3902;
 wire n3903;
 wire n3904;
 wire n3905;
 wire n3906;
 wire net93;
 wire net92;
 wire net91;
 wire net90;
 wire net89;
 wire net88;
 wire net87;
 wire net86;
 wire net85;
 wire net84;
 wire net83;
 wire net82;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire net75;
 wire net74;
 wire net73;
 wire net70;
 wire net69;
 wire net68;
 wire n3933;
 wire n3934;
 wire n3935;
 wire n3936;
 wire n3937;
 wire n3938;
 wire n3939;
 wire n3940;
 wire n3941;
 wire n3942;
 wire n3943;
 wire n3944;
 wire net67;
 wire net66;
 wire net65;
 wire net64;
 wire net63;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire net54;
 wire net53;
 wire net52;
 wire net51;
 wire net50;
 wire net49;
 wire net48;
 wire net47;
 wire net46;
 wire net45;
 wire net44;
 wire net43;
 wire net42;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire net36;
 wire net35;
 wire net34;
 wire net33;
 wire net32;
 wire net31;
 wire net30;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire net11;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire net71;
 wire net72;
 wire net81;
 wire clknet_leaf_0_clk_i;
 wire u_gpio_N113;
 wire u_gpio_N114;
 wire u_gpio_N115;
 wire u_gpio_N116;
 wire u_gpio_N117;
 wire u_gpio_N118;
 wire u_gpio_N119;
 wire u_gpio_N120;
 wire u_gpio_N121;
 wire u_gpio_N122;
 wire u_gpio_N123;
 wire u_gpio_N124;
 wire u_gpio_N125;
 wire u_gpio_N126;
 wire u_gpio_N127;
 wire u_gpio_N128;
 wire u_gpio_N129;
 wire u_gpio_N130;
 wire u_gpio_N131;
 wire u_gpio_N132;
 wire u_gpio_N133;
 wire u_gpio_N134;
 wire u_gpio_N135;
 wire u_gpio_N136;
 wire u_gpio_N137;
 wire u_gpio_N138;
 wire u_gpio_N139;
 wire u_gpio_N140;
 wire u_gpio_N141;
 wire u_gpio_N142;
 wire u_gpio_N143;
 wire u_gpio_N144;
 wire u_gpio_N145;
 wire u_gpio_N146;
 wire u_gpio_N38;
 wire u_gpio_N39;
 wire u_gpio_N40;
 wire u_gpio_N41;
 wire u_gpio_N42;
 wire u_gpio_N43;
 wire u_gpio_N44;
 wire u_gpio_N45;
 wire u_gpio_N46;
 wire u_gpio_N47;
 wire u_gpio_N48;
 wire u_gpio_N49;
 wire u_gpio_N50;
 wire u_gpio_N51;
 wire u_gpio_N52;
 wire u_gpio_N53;
 wire u_gpio_N54;
 wire u_gpio_N55;
 wire u_gpio_N56;
 wire u_gpio_N57;
 wire u_gpio_N58;
 wire u_gpio_N59;
 wire u_gpio_N60;
 wire u_gpio_N61;
 wire u_gpio_N62;
 wire u_gpio_N63;
 wire u_gpio_N64;
 wire u_gpio_N65;
 wire u_gpio_N66;
 wire u_gpio_N67;
 wire u_gpio_N68;
 wire u_gpio_N69;
 wire u_gpio_N70;
 wire u_gpio_N71;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_ack_level;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_nd;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_pd;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_req_trigger;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_test_set_d;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_n1;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_ping_set_d;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_ping_set_q;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nd;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_intq_0_;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_intq_0_;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_intq_0_;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_intq_0_;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q;
 wire u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_n5;
 wire u_gpio_gen_filter_0__u_filter_filter_q;
 wire u_gpio_gen_filter_0__u_filter_filter_synced;
 wire u_gpio_gen_filter_0__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_0__u_filter_stored_value_q;
 wire u_gpio_gen_filter_10__u_filter_filter_q;
 wire u_gpio_gen_filter_10__u_filter_filter_synced;
 wire u_gpio_gen_filter_10__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_10__u_filter_stored_value_q;
 wire u_gpio_gen_filter_11__u_filter_filter_q;
 wire u_gpio_gen_filter_11__u_filter_filter_synced;
 wire u_gpio_gen_filter_11__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_11__u_filter_stored_value_q;
 wire u_gpio_gen_filter_12__u_filter_filter_q;
 wire u_gpio_gen_filter_12__u_filter_filter_synced;
 wire u_gpio_gen_filter_12__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_12__u_filter_stored_value_q;
 wire u_gpio_gen_filter_13__u_filter_filter_q;
 wire u_gpio_gen_filter_13__u_filter_filter_synced;
 wire u_gpio_gen_filter_13__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_13__u_filter_stored_value_q;
 wire u_gpio_gen_filter_14__u_filter_filter_q;
 wire u_gpio_gen_filter_14__u_filter_filter_synced;
 wire u_gpio_gen_filter_14__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_14__u_filter_stored_value_q;
 wire u_gpio_gen_filter_15__u_filter_filter_q;
 wire u_gpio_gen_filter_15__u_filter_filter_synced;
 wire u_gpio_gen_filter_15__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_15__u_filter_stored_value_q;
 wire u_gpio_gen_filter_16__u_filter_filter_q;
 wire u_gpio_gen_filter_16__u_filter_filter_synced;
 wire u_gpio_gen_filter_16__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_16__u_filter_stored_value_q;
 wire u_gpio_gen_filter_17__u_filter_filter_q;
 wire u_gpio_gen_filter_17__u_filter_filter_synced;
 wire u_gpio_gen_filter_17__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_17__u_filter_stored_value_q;
 wire u_gpio_gen_filter_18__u_filter_filter_q;
 wire u_gpio_gen_filter_18__u_filter_filter_synced;
 wire u_gpio_gen_filter_18__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_18__u_filter_stored_value_q;
 wire u_gpio_gen_filter_19__u_filter_filter_q;
 wire u_gpio_gen_filter_19__u_filter_filter_synced;
 wire u_gpio_gen_filter_19__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_19__u_filter_stored_value_q;
 wire u_gpio_gen_filter_1__u_filter_filter_q;
 wire u_gpio_gen_filter_1__u_filter_filter_synced;
 wire u_gpio_gen_filter_1__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_1__u_filter_stored_value_q;
 wire u_gpio_gen_filter_20__u_filter_filter_q;
 wire u_gpio_gen_filter_20__u_filter_filter_synced;
 wire u_gpio_gen_filter_20__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_20__u_filter_stored_value_q;
 wire u_gpio_gen_filter_21__u_filter_filter_q;
 wire u_gpio_gen_filter_21__u_filter_filter_synced;
 wire u_gpio_gen_filter_21__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_21__u_filter_stored_value_q;
 wire u_gpio_gen_filter_22__u_filter_filter_q;
 wire u_gpio_gen_filter_22__u_filter_filter_synced;
 wire u_gpio_gen_filter_22__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_22__u_filter_stored_value_q;
 wire u_gpio_gen_filter_23__u_filter_filter_q;
 wire u_gpio_gen_filter_23__u_filter_filter_synced;
 wire u_gpio_gen_filter_23__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_23__u_filter_stored_value_q;
 wire u_gpio_gen_filter_24__u_filter_filter_q;
 wire u_gpio_gen_filter_24__u_filter_filter_synced;
 wire u_gpio_gen_filter_24__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_24__u_filter_stored_value_q;
 wire u_gpio_gen_filter_25__u_filter_filter_q;
 wire u_gpio_gen_filter_25__u_filter_filter_synced;
 wire u_gpio_gen_filter_25__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_25__u_filter_stored_value_q;
 wire u_gpio_gen_filter_26__u_filter_filter_q;
 wire u_gpio_gen_filter_26__u_filter_filter_synced;
 wire u_gpio_gen_filter_26__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_26__u_filter_stored_value_q;
 wire u_gpio_gen_filter_27__u_filter_filter_q;
 wire u_gpio_gen_filter_27__u_filter_filter_synced;
 wire u_gpio_gen_filter_27__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_27__u_filter_stored_value_q;
 wire u_gpio_gen_filter_28__u_filter_filter_q;
 wire u_gpio_gen_filter_28__u_filter_filter_synced;
 wire u_gpio_gen_filter_28__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_28__u_filter_stored_value_q;
 wire u_gpio_gen_filter_29__u_filter_filter_q;
 wire u_gpio_gen_filter_29__u_filter_filter_synced;
 wire u_gpio_gen_filter_29__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_29__u_filter_stored_value_q;
 wire u_gpio_gen_filter_2__u_filter_filter_q;
 wire u_gpio_gen_filter_2__u_filter_filter_synced;
 wire u_gpio_gen_filter_2__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_2__u_filter_stored_value_q;
 wire u_gpio_gen_filter_30__u_filter_filter_q;
 wire u_gpio_gen_filter_30__u_filter_filter_synced;
 wire u_gpio_gen_filter_30__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_30__u_filter_stored_value_q;
 wire u_gpio_gen_filter_31__u_filter_filter_q;
 wire u_gpio_gen_filter_31__u_filter_filter_synced;
 wire u_gpio_gen_filter_31__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_31__u_filter_stored_value_q;
 wire u_gpio_gen_filter_3__u_filter_filter_q;
 wire u_gpio_gen_filter_3__u_filter_filter_synced;
 wire u_gpio_gen_filter_3__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_3__u_filter_stored_value_q;
 wire u_gpio_gen_filter_4__u_filter_filter_q;
 wire u_gpio_gen_filter_4__u_filter_filter_synced;
 wire u_gpio_gen_filter_4__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_4__u_filter_stored_value_q;
 wire u_gpio_gen_filter_5__u_filter_filter_q;
 wire u_gpio_gen_filter_5__u_filter_filter_synced;
 wire u_gpio_gen_filter_5__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_5__u_filter_stored_value_q;
 wire u_gpio_gen_filter_6__u_filter_filter_q;
 wire u_gpio_gen_filter_6__u_filter_filter_synced;
 wire u_gpio_gen_filter_6__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_6__u_filter_stored_value_q;
 wire u_gpio_gen_filter_7__u_filter_filter_q;
 wire u_gpio_gen_filter_7__u_filter_filter_synced;
 wire u_gpio_gen_filter_7__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_7__u_filter_stored_value_q;
 wire u_gpio_gen_filter_8__u_filter_filter_q;
 wire u_gpio_gen_filter_8__u_filter_filter_synced;
 wire u_gpio_gen_filter_8__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_8__u_filter_stored_value_q;
 wire u_gpio_gen_filter_9__u_filter_filter_q;
 wire u_gpio_gen_filter_9__u_filter_filter_synced;
 wire u_gpio_gen_filter_9__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire u_gpio_gen_filter_9__u_filter_stored_value_q;
 wire u_gpio_intr_hw_N1;
 wire u_gpio_intr_hw_N10;
 wire u_gpio_intr_hw_N11;
 wire u_gpio_intr_hw_N12;
 wire u_gpio_intr_hw_N13;
 wire u_gpio_intr_hw_N14;
 wire u_gpio_intr_hw_N15;
 wire u_gpio_intr_hw_N16;
 wire u_gpio_intr_hw_N17;
 wire u_gpio_intr_hw_N18;
 wire u_gpio_intr_hw_N19;
 wire u_gpio_intr_hw_N2;
 wire u_gpio_intr_hw_N20;
 wire u_gpio_intr_hw_N21;
 wire u_gpio_intr_hw_N22;
 wire u_gpio_intr_hw_N23;
 wire u_gpio_intr_hw_N24;
 wire u_gpio_intr_hw_N25;
 wire u_gpio_intr_hw_N26;
 wire u_gpio_intr_hw_N27;
 wire u_gpio_intr_hw_N28;
 wire u_gpio_intr_hw_N29;
 wire u_gpio_intr_hw_N3;
 wire u_gpio_intr_hw_N30;
 wire u_gpio_intr_hw_N31;
 wire u_gpio_intr_hw_N32;
 wire u_gpio_intr_hw_N4;
 wire u_gpio_intr_hw_N5;
 wire u_gpio_intr_hw_N6;
 wire u_gpio_intr_hw_N7;
 wire u_gpio_intr_hw_N8;
 wire u_gpio_intr_hw_N9;
 wire u_gpio_net3588;
 wire u_gpio_net3594;
 wire u_gpio_net3599;
 wire u_gpio_net3604;
 wire u_gpio_u_reg_err_q;
 wire u_gpio_u_reg_reg_we_check_14_;
 wire u_gpio_u_reg_u_ctrl_en_input_filter_net3621;
 wire u_gpio_u_reg_u_ctrl_en_input_filter_net3627;
 wire u_gpio_u_reg_u_intr_ctrl_en_falling_net3621;
 wire u_gpio_u_reg_u_intr_ctrl_en_falling_net3627;
 wire u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621;
 wire u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627;
 wire u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621;
 wire u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627;
 wire u_gpio_u_reg_u_intr_ctrl_en_rising_net3621;
 wire u_gpio_u_reg_u_intr_ctrl_en_rising_net3627;
 wire u_gpio_u_reg_u_intr_enable_net3621;
 wire u_gpio_u_reg_u_intr_enable_net3627;
 wire u_gpio_u_reg_u_intr_state_n1;
 wire u_gpio_u_reg_u_intr_state_net3644;
 wire u_gpio_u_reg_u_intr_state_net3650;
 wire u_gpio_u_reg_u_reg_if_N14;
 wire u_gpio_u_reg_u_reg_if_N15;
 wire u_gpio_u_reg_u_reg_if_N16;
 wire u_gpio_u_reg_u_reg_if_N17;
 wire u_gpio_u_reg_u_reg_if_N18;
 wire u_gpio_u_reg_u_reg_if_N19;
 wire u_gpio_u_reg_u_reg_if_N20;
 wire u_gpio_u_reg_u_reg_if_N21;
 wire u_gpio_u_reg_u_reg_if_N22;
 wire u_gpio_u_reg_u_reg_if_N23;
 wire u_gpio_u_reg_u_reg_if_N24;
 wire u_gpio_u_reg_u_reg_if_N25;
 wire u_gpio_u_reg_u_reg_if_N26;
 wire u_gpio_u_reg_u_reg_if_N27;
 wire u_gpio_u_reg_u_reg_if_N28;
 wire u_gpio_u_reg_u_reg_if_N29;
 wire u_gpio_u_reg_u_reg_if_N30;
 wire u_gpio_u_reg_u_reg_if_N31;
 wire u_gpio_u_reg_u_reg_if_N32;
 wire u_gpio_u_reg_u_reg_if_N33;
 wire u_gpio_u_reg_u_reg_if_N34;
 wire u_gpio_u_reg_u_reg_if_N35;
 wire u_gpio_u_reg_u_reg_if_N36;
 wire u_gpio_u_reg_u_reg_if_N37;
 wire u_gpio_u_reg_u_reg_if_N38;
 wire u_gpio_u_reg_u_reg_if_N39;
 wire u_gpio_u_reg_u_reg_if_N40;
 wire u_gpio_u_reg_u_reg_if_N41;
 wire u_gpio_u_reg_u_reg_if_N42;
 wire u_gpio_u_reg_u_reg_if_N43;
 wire u_gpio_u_reg_u_reg_if_N44;
 wire u_gpio_u_reg_u_reg_if_N45;
 wire u_gpio_u_reg_u_reg_if_N46;
 wire u_gpio_u_reg_u_reg_if_N7;
 wire u_gpio_u_reg_u_reg_if_net3667;
 wire u_gpio_u_reg_u_reg_if_net3673;
 wire u_gpio_u_reg_u_reg_if_net3678;
 wire u_gpio_u_reg_u_reg_if_rd_req;
 wire u_xbar_periph_u_s1n_6_N59;
 wire u_xbar_periph_u_s1n_6_N60;
 wire u_xbar_periph_u_s1n_6_N61;
 wire u_xbar_periph_u_s1n_6_N62;
 wire u_xbar_periph_u_s1n_6_N63;
 wire u_xbar_periph_u_s1n_6_N64;
 wire u_xbar_periph_u_s1n_6_N65;
 wire u_xbar_periph_u_s1n_6_N66;
 wire u_xbar_periph_u_s1n_6_N67;
 wire u_xbar_periph_u_s1n_6_N68;
 wire u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_N12;
 wire u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_N8;
 wire u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_req_pending;
 wire u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_rsp_pending;
 wire u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713;
 wire u_xbar_periph_u_s1n_6_net3695;
 wire net1345;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_2_clk_i;
 wire clknet_leaf_3_clk_i;
 wire clknet_leaf_4_clk_i;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_6_clk_i;
 wire clknet_leaf_7_clk_i;
 wire clknet_leaf_8_clk_i;
 wire clknet_leaf_9_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_leaf_12_clk_i;
 wire clknet_0_clk_i;
 wire clknet_1_0__leaf_clk_i;
 wire clknet_1_1__leaf_clk_i;
 wire clknet_0_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713;
 wire clknet_1_0__leaf_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713;
 wire clknet_1_1__leaf_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713;
 wire clknet_0_u_xbar_periph_u_s1n_6_net3695;
 wire clknet_1_0__leaf_u_xbar_periph_u_s1n_6_net3695;
 wire clknet_1_1__leaf_u_xbar_periph_u_s1n_6_net3695;
 wire clknet_0_u_gpio_u_reg_u_reg_if_net3667;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3667;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3667;
 wire clknet_0_u_gpio_u_reg_u_reg_if_net3673;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3673;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3673;
 wire clknet_0_u_gpio_u_reg_u_reg_if_net3678;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3678;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3678;
 wire clknet_0_u_gpio_u_reg_u_intr_state_net3644;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_intr_state_net3644;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_intr_state_net3644;
 wire clknet_0_u_gpio_u_reg_u_intr_state_net3650;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_intr_state_net3650;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_intr_state_net3650;
 wire clknet_0_u_gpio_u_reg_u_intr_enable_net3621;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_intr_enable_net3621;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_intr_enable_net3621;
 wire clknet_0_u_gpio_u_reg_u_intr_enable_net3627;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_intr_enable_net3627;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_intr_enable_net3627;
 wire clknet_0_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621;
 wire clknet_0_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627;
 wire clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621;
 wire clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627;
 wire clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621;
 wire clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627;
 wire clknet_0_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621;
 wire clknet_0_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627;
 wire clknet_0_u_gpio_u_reg_u_ctrl_en_input_filter_net3621;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3621;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3621;
 wire clknet_0_u_gpio_u_reg_u_ctrl_en_input_filter_net3627;
 wire clknet_1_0__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3627;
 wire clknet_1_1__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3627;
 wire clknet_0_u_gpio_net3588;
 wire clknet_1_0__leaf_u_gpio_net3588;
 wire clknet_1_1__leaf_u_gpio_net3588;
 wire clknet_0_u_gpio_net3594;
 wire clknet_1_0__leaf_u_gpio_net3594;
 wire clknet_1_1__leaf_u_gpio_net3594;
 wire clknet_0_u_gpio_net3599;
 wire clknet_1_0__leaf_u_gpio_net3599;
 wire clknet_1_1__leaf_u_gpio_net3599;
 wire clknet_0_u_gpio_net3604;
 wire clknet_1_0__leaf_u_gpio_net3604;
 wire clknet_1_1__leaf_u_gpio_net3604;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire [31:0] gpio_2_xbar;
 wire [31:0] u_gpio_data_in_q;
 wire [2:0] u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_d;
 wire [2:0] u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q;
 wire [1:0] u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d;
 wire [1:0] u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q;
 wire [1:0] u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d;
 wire [1:0] u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q;
 wire [3:0] u_gpio_gen_filter_0__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_0__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_10__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_10__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_11__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_11__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_12__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_12__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_13__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_13__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_14__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_14__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_15__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_15__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_16__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_16__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_17__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_17__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_18__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_18__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_19__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_19__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_1__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_1__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_20__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_20__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_21__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_21__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_22__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_22__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_23__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_23__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_24__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_24__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_25__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_25__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_26__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_26__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_27__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_27__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_28__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_28__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_29__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_29__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_2__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_2__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_30__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_30__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_31__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_31__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_3__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_3__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_4__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_4__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_5__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_5__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_6__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_6__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_7__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_7__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_8__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_8__u_filter_diff_ctr_q;
 wire [3:0] u_gpio_gen_filter_9__u_filter_diff_ctr_d;
 wire [3:0] u_gpio_gen_filter_9__u_filter_diff_ctr_q;
 wire [223:0] u_gpio_reg2hw;
 wire [31:0] u_gpio_u_reg_data_in_qs;
 wire [15:0] u_gpio_u_reg_masked_oe_lower_data_qs;
 wire [15:0] u_gpio_u_reg_masked_oe_upper_data_qs;
 wire [31:0] u_gpio_u_reg_u_ctrl_en_input_filter_wr_data;
 wire [31:0] u_gpio_u_reg_u_data_in_wr_data;
 wire [31:0] u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data;
 wire [31:0] u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data;
 wire [31:0] u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data;
 wire [31:0] u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data;
 wire [31:0] u_gpio_u_reg_u_intr_enable_wr_data;
 wire [31:0] u_gpio_u_reg_u_intr_state_wr_data;
 wire [2:0] u_xbar_periph_u_s1n_6_dev_select_outstanding;
 wire [2:0] u_xbar_periph_u_s1n_6_dev_select_t;
 wire [2:0] u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type;
 wire [1:0] u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_opcode;
 wire [8:0] u_xbar_periph_u_s1n_6_num_req_outstanding;
 wire [24:0] u_xbar_periph_u_s1n_6_tl_u_i;

 b15inv000an1n03x5 U3215 (.a(net12),
    .o1(n1435));
 b15and002ar1n16x5 U3216 (.a(u_gpio_reg2hw[181]),
    .b(u_gpio_reg2hw[213]),
    .o(u_gpio_intr_hw_N11));
 b15and002an1n12x5 U3217 (.a(u_gpio_reg2hw[196]),
    .b(u_gpio_reg2hw[164]),
    .o(u_gpio_intr_hw_N28));
 b15and002ah1n08x5 U3218 (.a(u_gpio_reg2hw[205]),
    .b(u_gpio_reg2hw[173]),
    .o(u_gpio_intr_hw_N19));
 b15and002ar1n03x5 U3219 (.a(net281),
    .b(u_gpio_reg2hw[166]),
    .o(u_gpio_intr_hw_N26));
 b15and002al1n03x5 U3220 (.a(u_gpio_reg2hw[200]),
    .b(u_gpio_reg2hw[168]),
    .o(u_gpio_intr_hw_N24));
 b15and002al1n02x5 U3221 (.a(u_gpio_reg2hw[167]),
    .b(u_gpio_reg2hw[199]),
    .o(u_gpio_intr_hw_N25));
 b15and002ar1n03x5 U3222 (.a(u_gpio_reg2hw[192]),
    .b(u_gpio_reg2hw[160]),
    .o(u_gpio_intr_hw_N32));
 b15and002ah1n08x5 U3223 (.a(u_gpio_reg2hw[197]),
    .b(u_gpio_reg2hw[165]),
    .o(u_gpio_intr_hw_N27));
 b15and002as1n02x5 U3224 (.a(u_gpio_reg2hw[202]),
    .b(u_gpio_reg2hw[170]),
    .o(u_gpio_intr_hw_N22));
 b15and002as1n04x5 U3225 (.a(u_gpio_reg2hw[207]),
    .b(u_gpio_reg2hw[175]),
    .o(u_gpio_intr_hw_N17));
 b15and002as1n08x5 U3226 (.a(u_gpio_reg2hw[220]),
    .b(net286),
    .o(u_gpio_intr_hw_N4));
 b15and002al1n16x5 U3227 (.a(u_gpio_reg2hw[204]),
    .b(u_gpio_reg2hw[172]),
    .o(u_gpio_intr_hw_N20));
 b15and002al1n08x5 U3228 (.a(u_gpio_reg2hw[193]),
    .b(u_gpio_reg2hw[161]),
    .o(u_gpio_intr_hw_N31));
 b15and002al1n02x5 U3229 (.a(u_gpio_reg2hw[201]),
    .b(u_gpio_reg2hw[169]),
    .o(u_gpio_intr_hw_N23));
 b15and002al1n02x5 U3230 (.a(u_gpio_reg2hw[203]),
    .b(u_gpio_reg2hw[171]),
    .o(u_gpio_intr_hw_N21));
 b15and002al1n02x5 U3231 (.a(u_gpio_reg2hw[195]),
    .b(net284),
    .o(u_gpio_intr_hw_N29));
 b15and002ah1n02x5 U3232 (.a(u_gpio_reg2hw[206]),
    .b(u_gpio_reg2hw[174]),
    .o(u_gpio_intr_hw_N18));
 b15and002aq1n03x5 U3233 (.a(u_gpio_reg2hw[194]),
    .b(net285),
    .o(u_gpio_intr_hw_N30));
 b15and002ar1n08x5 U3234 (.a(u_gpio_reg2hw[187]),
    .b(u_gpio_reg2hw[219]),
    .o(u_gpio_intr_hw_N5));
 b15and002al1n02x5 U3235 (.a(u_gpio_reg2hw[185]),
    .b(u_gpio_reg2hw[217]),
    .o(u_gpio_intr_hw_N7));
 b15and002as1n08x5 U3236 (.a(u_gpio_reg2hw[189]),
    .b(u_gpio_reg2hw[221]),
    .o(u_gpio_intr_hw_N3));
 b15and002as1n02x5 U3237 (.a(u_gpio_reg2hw[190]),
    .b(net282),
    .o(u_gpio_intr_hw_N2));
 b15and002al1n08x5 U3238 (.a(u_gpio_reg2hw[191]),
    .b(u_gpio_reg2hw[223]),
    .o(u_gpio_intr_hw_N1));
 b15and002ah1n02x5 U3239 (.a(u_gpio_reg2hw[176]),
    .b(u_gpio_reg2hw[208]),
    .o(u_gpio_intr_hw_N16));
 b15and002ar1n02x5 U3240 (.a(u_gpio_reg2hw[180]),
    .b(u_gpio_reg2hw[212]),
    .o(u_gpio_intr_hw_N12));
 b15and002ar1n03x5 U3241 (.a(u_gpio_reg2hw[178]),
    .b(u_gpio_reg2hw[210]),
    .o(u_gpio_intr_hw_N14));
 b15and002ar1n08x5 U3242 (.a(u_gpio_reg2hw[184]),
    .b(u_gpio_reg2hw[216]),
    .o(u_gpio_intr_hw_N8));
 b15and002ar1n02x5 U3243 (.a(u_gpio_reg2hw[186]),
    .b(u_gpio_reg2hw[218]),
    .o(u_gpio_intr_hw_N6));
 b15and002ar1n02x5 U3244 (.a(u_gpio_reg2hw[177]),
    .b(u_gpio_reg2hw[209]),
    .o(u_gpio_intr_hw_N15));
 b15and002aq1n04x5 U3245 (.a(u_gpio_reg2hw[182]),
    .b(u_gpio_reg2hw[214]),
    .o(u_gpio_intr_hw_N10));
 b15and002al1n02x5 U3246 (.a(u_gpio_reg2hw[183]),
    .b(u_gpio_reg2hw[215]),
    .o(u_gpio_intr_hw_N9));
 b15and002ar1n08x5 U3247 (.a(u_gpio_reg2hw[179]),
    .b(u_gpio_reg2hw[211]),
    .o(u_gpio_intr_hw_N13));
 b15inv000as1n80x5 U3248 (.a(net505),
    .o1(n3891));
 b15inv000as1n80x5 U3249 (.a(net504),
    .o1(n3892));
 b15inv000as1n64x5 U3250 (.a(net31),
    .o1(n3893));
 b15inv000as1n48x5 U3251 (.a(net32),
    .o1(n3894));
 b15inv000ah1n48x5 U3252 (.a(net33),
    .o1(n3895));
 b15inv000as1n28x5 U3253 (.a(net34),
    .o1(n3896));
 b15inv040as1n40x5 U3254 (.a(net35),
    .o1(n3897));
 b15inv040as1n40x5 U3255 (.a(net36),
    .o1(n3898));
 b15inv040aq1n60x5 U3256 (.a(net503),
    .o1(n3899));
 b15inv000al1n04x5 U3257 (.a(u_xbar_periph_u_s1n_6_num_req_outstanding[0]),
    .o1(u_xbar_periph_u_s1n_6_N60));
 b15inv000al1n80x5 U3258 (.a(net502),
    .o1(n3900));
 b15inv000al1n80x5 U3259 (.a(net39),
    .o1(n3901));
 b15inv000aq1n80x5 U3260 (.a(net40),
    .o1(n3902));
 b15inv040as1n36x5 U3261 (.a(net41),
    .o1(n3903));
 b15inv040aq1n60x5 U3262 (.a(net42),
    .o1(n3904));
 b15inv000as1n80x5 U3263 (.a(net43),
    .o1(n3905));
 b15inv000as1n80x5 U3264 (.a(net44),
    .o1(n3906));
 b15ztpn00an1n08x5 PHY_94 ();
 b15ztpn00an1n08x5 PHY_93 ();
 b15ztpn00an1n08x5 PHY_92 ();
 b15ztpn00an1n08x5 PHY_91 ();
 b15ztpn00an1n08x5 PHY_90 ();
 b15ztpn00an1n08x5 PHY_89 ();
 b15ztpn00an1n08x5 PHY_88 ();
 b15ztpn00an1n08x5 PHY_87 ();
 b15ztpn00an1n08x5 PHY_86 ();
 b15ztpn00an1n08x5 PHY_85 ();
 b15ztpn00an1n08x5 PHY_84 ();
 b15ztpn00an1n08x5 PHY_83 ();
 b15ztpn00an1n08x5 PHY_82 ();
 b15ztpn00an1n08x5 PHY_81 ();
 b15ztpn00an1n08x5 PHY_80 ();
 b15ztpn00an1n08x5 PHY_79 ();
 b15ztpn00an1n08x5 PHY_78 ();
 b15ztpn00an1n08x5 PHY_77 ();
 b15ztpn00an1n08x5 PHY_76 ();
 b15ztpn00an1n08x5 PHY_75 ();
 b15ztpn00an1n08x5 PHY_74 ();
 b15ztpn00an1n08x5 PHY_73 ();
 b15ztpn00an1n08x5 PHY_72 ();
 b15ztpn00an1n08x5 PHY_71 ();
 b15ztpn00an1n08x5 PHY_70 ();
 b15ztpn00an1n08x5 PHY_69 ();
 b15inv000al1n02x5 U3291 (.a(net455),
    .o1(n3933));
 b15inv040as1n10x5 U3292 (.a(n3617),
    .o1(n3934));
 b15inv000aq1n28x5 U3293 (.a(net1860),
    .o1(n3935));
 b15inv040as1n20x5 U3294 (.a(n3134),
    .o1(n3936));
 b15inv040al1n12x5 U3295 (.a(net201),
    .o1(n3937));
 b15inv040as1n48x5 U3296 (.a(n3226),
    .o1(n3938));
 b15inv040as1n10x5 U3297 (.a(net210),
    .o1(n3939));
 b15inv000al1n24x5 U3298 (.a(net212),
    .o1(n3940));
 b15inv000an1n24x5 U3299 (.a(net214),
    .o1(n3941));
 b15qgbin1an1n15x5 U3300 (.a(net218),
    .o1(n3942));
 b15inv040as1n20x5 U3301 (.a(net219),
    .o1(n3943));
 b15inv020ar1n32x5 U3302 (.a(net179),
    .o1(n3944));
 b15inv000ar1n03x5 U3303 (.a(net1345),
    .o1(tl_peri_device_o[48]));
 b15inv000ar1n03x5 U3305 (.a(net1346),
    .o1(tl_peri_device_o[59]));
 b15inv000ar1n03x5 U3307 (.a(net1347),
    .o1(tl_peri_device_o[60]));
 b15inv000ar1n03x5 U3309 (.a(net1348),
    .o1(tl_peri_device_o[61]));
 b15ztpn00an1n08x5 PHY_68 ();
 b15ztpn00an1n08x5 PHY_67 ();
 b15ztpn00an1n08x5 PHY_66 ();
 b15ztpn00an1n08x5 PHY_65 ();
 b15ztpn00an1n08x5 PHY_64 ();
 b15ztpn00an1n08x5 PHY_63 ();
 b15ztpn00an1n08x5 PHY_62 ();
 b15ztpn00an1n08x5 PHY_61 ();
 b15ztpn00an1n08x5 PHY_60 ();
 b15ztpn00an1n08x5 PHY_59 ();
 b15ztpn00an1n08x5 PHY_58 ();
 b15ztpn00an1n08x5 PHY_57 ();
 b15ztpn00an1n08x5 PHY_56 ();
 b15inv020as1n08x5 U3325 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd),
    .o1(n2747));
 b15inv020as1n10x5 U3326 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd),
    .o1(n2746));
 b15oai013ar1n03x5 U3327 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd),
    .c(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .d(n2746),
    .o1(n2628));
 b15oai013as1n04x5 U3328 (.a(n2628),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd),
    .c(net2122),
    .d(n2747),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_n5));
 b15inv000al1n02x5 U3329 (.a(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_rsp_pending),
    .o1(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_N8));
 b15nandp3ah1n08x5 U3330 (.a(u_gpio_gen_filter_23__u_filter_diff_ctr_q[1]),
    .b(u_gpio_gen_filter_23__u_filter_diff_ctr_q[3]),
    .c(u_gpio_gen_filter_23__u_filter_diff_ctr_q[2]),
    .o1(n2731));
 b15xor002ah1n06x5 U3331 (.a(net444),
    .b(net1987),
    .out0(n2728));
 b15aoi012ah1n02x5 U3332 (.a(n2728),
    .b(net1971),
    .c(n2731),
    .o1(u_gpio_gen_filter_23__u_filter_diff_ctr_d[0]));
 b15and003aq1n04x5 U3333 (.a(u_gpio_gen_filter_15__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_15__u_filter_diff_ctr_q[0]),
    .c(net2117),
    .o(n2676));
 b15xor002ah1n08x5 U3334 (.a(net449),
    .b(net2071),
    .out0(n2736));
 b15oab012an1n03x5 U3335 (.a(n2736),
    .b(u_gpio_gen_filter_15__u_filter_diff_ctr_q[3]),
    .c(n2676),
    .out0(u_gpio_gen_filter_15__u_filter_diff_ctr_d[3]));
 b15ztpn00an1n08x5 PHY_55 ();
 b15ztpn00an1n08x5 PHY_54 ();
 b15xor002aq1n16x5 U3338 (.a(net451),
    .b(net2167),
    .out0(n2687));
 b15and002an1n03x5 U3339 (.a(net2036),
    .b(u_gpio_gen_filter_14__u_filter_diff_ctr_q[1]),
    .o(n2680));
 b15nandp3ar1n04x5 U3340 (.a(net2036),
    .b(u_gpio_gen_filter_14__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_14__u_filter_diff_ctr_q[2]),
    .o1(n2634));
 b15oai022an1n02x5 U3341 (.a(n2680),
    .b(u_gpio_gen_filter_14__u_filter_diff_ctr_q[2]),
    .c(net2182),
    .d(n2634),
    .o1(n2629));
 b15norp02an1n03x5 U3342 (.a(n2687),
    .b(net2183),
    .o1(u_gpio_gen_filter_14__u_filter_diff_ctr_d[2]));
 b15xor002aq1n16x5 U3343 (.a(u_gpio_gen_filter_2__u_filter_filter_synced),
    .b(u_gpio_gen_filter_2__u_filter_filter_q),
    .out0(n2685));
 b15and002ar1n03x5 U3344 (.a(net2184),
    .b(u_gpio_gen_filter_2__u_filter_diff_ctr_q[1]),
    .o(n2683));
 b15nand03an1n06x5 U3345 (.a(net1975),
    .b(u_gpio_gen_filter_2__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_2__u_filter_diff_ctr_q[2]),
    .o1(n2632));
 b15oai022ar1n02x5 U3346 (.a(n2683),
    .b(net2196),
    .c(net2169),
    .d(n2632),
    .o1(n2630));
 b15norp02ar1n02x5 U3347 (.a(n2685),
    .b(n2630),
    .o1(u_gpio_gen_filter_2__u_filter_diff_ctr_d[2]));
 b15and002ar1n02x5 U3348 (.a(u_gpio_gen_filter_23__u_filter_diff_ctr_q[1]),
    .b(u_gpio_gen_filter_23__u_filter_diff_ctr_q[0]),
    .o(n2675));
 b15nand03as1n06x5 U3349 (.a(u_gpio_gen_filter_23__u_filter_diff_ctr_q[1]),
    .b(u_gpio_gen_filter_23__u_filter_diff_ctr_q[2]),
    .c(net1971),
    .o1(n2729));
 b15oai022ar1n02x5 U3350 (.a(net2049),
    .b(n2675),
    .c(u_gpio_gen_filter_23__u_filter_diff_ctr_q[3]),
    .d(n2729),
    .o1(n2631));
 b15norp02ar1n02x5 U3351 (.a(n2728),
    .b(net2050),
    .o1(u_gpio_gen_filter_23__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3352 (.a(net2169),
    .o1(n2633));
 b15aoi012ar1n02x5 U3353 (.a(n2685),
    .b(n2633),
    .c(n2632),
    .o1(u_gpio_gen_filter_2__u_filter_diff_ctr_d[3]));
 b15inv000al1n02x5 U3354 (.a(u_gpio_gen_filter_14__u_filter_diff_ctr_q[3]),
    .o1(n2635));
 b15aoi012as1n02x5 U3355 (.a(n2687),
    .b(n2635),
    .c(n2634),
    .o1(u_gpio_gen_filter_14__u_filter_diff_ctr_d[3]));
 b15nand03as1n06x5 U3356 (.a(u_gpio_gen_filter_14__u_filter_diff_ctr_q[3]),
    .b(u_gpio_gen_filter_14__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_14__u_filter_diff_ctr_q[2]),
    .o1(n2686));
 b15aoi012ar1n02x5 U3357 (.a(n2687),
    .b(net2036),
    .c(n2686),
    .o1(u_gpio_gen_filter_14__u_filter_diff_ctr_d[0]));
 b15nand03as1n04x5 U3358 (.a(net2215),
    .b(u_gpio_gen_filter_2__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_2__u_filter_diff_ctr_q[2]),
    .o1(n2684));
 b15aoi012aq1n02x5 U3359 (.a(n2685),
    .b(net1975),
    .c(n2684),
    .o1(u_gpio_gen_filter_2__u_filter_diff_ctr_d[0]));
 b15and003ah1n03x5 U3360 (.a(u_gpio_gen_filter_25__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_25__u_filter_diff_ctr_q[1]),
    .c(net2032),
    .o(n2791));
 b15xor002ah1n16x5 U3361 (.a(net2030),
    .b(u_gpio_gen_filter_25__u_filter_filter_synced),
    .out0(n2792));
 b15oab012al1n02x5 U3362 (.a(n2792),
    .b(net2083),
    .c(n2791),
    .out0(u_gpio_gen_filter_25__u_filter_diff_ctr_d[3]));
 b15and003as1n03x5 U3363 (.a(net1977),
    .b(u_gpio_gen_filter_17__u_filter_diff_ctr_q[1]),
    .c(net2057),
    .o(n2799));
 b15xor002an1n16x5 U3364 (.a(u_gpio_gen_filter_17__u_filter_filter_q),
    .b(u_gpio_gen_filter_17__u_filter_filter_synced),
    .out0(n2800));
 b15oab012ar1n02x5 U3365 (.a(n2800),
    .b(net2090),
    .c(n2799),
    .out0(u_gpio_gen_filter_17__u_filter_diff_ctr_d[3]));
 b15and003ah1n03x5 U3366 (.a(u_gpio_gen_filter_0__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_0__u_filter_diff_ctr_q[1]),
    .c(net2004),
    .o(n2807));
 b15xor002as1n08x5 U3367 (.a(net1991),
    .b(u_gpio_gen_filter_0__u_filter_filter_synced),
    .out0(n2808));
 b15oab012ar1n02x5 U3368 (.a(n2808),
    .b(u_gpio_gen_filter_0__u_filter_diff_ctr_q[3]),
    .c(n2807),
    .out0(u_gpio_gen_filter_0__u_filter_diff_ctr_d[3]));
 b15and003aq1n03x5 U3369 (.a(u_gpio_gen_filter_11__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_11__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_11__u_filter_diff_ctr_q[2]),
    .o(n2689));
 b15xor002ah1n08x5 U3370 (.a(u_gpio_gen_filter_11__u_filter_filter_synced),
    .b(net2014),
    .out0(n2743));
 b15oab012as1n02x5 U3371 (.a(n2743),
    .b(net2019),
    .c(n2689),
    .out0(u_gpio_gen_filter_11__u_filter_diff_ctr_d[3]));
 b15and003as1n04x5 U3372 (.a(net2044),
    .b(u_gpio_gen_filter_19__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_19__u_filter_diff_ctr_q[1]),
    .o(n2712));
 b15xor002as1n12x5 U3373 (.a(net446),
    .b(net2067),
    .out0(n2707));
 b15oab012aq1n02x5 U3374 (.a(n2707),
    .b(net2078),
    .c(n2712),
    .out0(u_gpio_gen_filter_19__u_filter_diff_ctr_d[3]));
 b15and003al1n04x5 U3375 (.a(net2113),
    .b(u_gpio_gen_filter_24__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_24__u_filter_diff_ctr_q[1]),
    .o(n2718));
 b15xor002ar1n16x5 U3376 (.a(net443),
    .b(u_gpio_gen_filter_24__u_filter_filter_q),
    .out0(n2713));
 b15oab012al1n02x5 U3377 (.a(n2713),
    .b(net2198),
    .c(n2718),
    .out0(u_gpio_gen_filter_24__u_filter_diff_ctr_d[3]));
 b15and003ah1n04x5 U3378 (.a(u_gpio_gen_filter_6__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_6__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_6__u_filter_diff_ctr_q[2]),
    .o(n2688));
 b15xor002ah1n12x5 U3379 (.a(net440),
    .b(net2008),
    .out0(n2739));
 b15oab012ar1n02x5 U3380 (.a(n2739),
    .b(u_gpio_gen_filter_6__u_filter_diff_ctr_q[3]),
    .c(n2688),
    .out0(u_gpio_gen_filter_6__u_filter_diff_ctr_d[3]));
 b15inv040an1n08x5 U3381 (.a(u_gpio_gen_filter_27__u_filter_filter_synced),
    .o1(n3461));
 b15xor002an1n06x5 U3382 (.a(net2022),
    .b(n3461),
    .out0(n2726));
 b15inv040as1n03x5 U3383 (.a(n2726),
    .o1(n2697));
 b15inv000al1n02x5 U3384 (.a(u_gpio_gen_filter_27__u_filter_diff_ctr_q[0]),
    .o1(n2636));
 b15aoi013al1n02x5 U3385 (.a(n2636),
    .b(u_gpio_gen_filter_27__u_filter_diff_ctr_q[3]),
    .c(u_gpio_gen_filter_27__u_filter_diff_ctr_q[1]),
    .d(u_gpio_gen_filter_27__u_filter_diff_ctr_q[2]),
    .o1(n2637));
 b15nor002an1n02x5 U3386 (.a(n2697),
    .b(n2637),
    .o1(u_gpio_gen_filter_27__u_filter_diff_ctr_d[0]));
 b15inv040as1n10x5 U3387 (.a(u_gpio_gen_filter_7__u_filter_filter_synced),
    .o1(n3254));
 b15xor002an1n08x5 U3388 (.a(net2048),
    .b(n3254),
    .out0(n2724));
 b15inv000aq1n05x5 U3389 (.a(n2724),
    .o1(n2702));
 b15inv000al1n02x5 U3390 (.a(u_gpio_gen_filter_7__u_filter_diff_ctr_q[0]),
    .o1(n2638));
 b15aoi013al1n02x5 U3391 (.a(n2638),
    .b(u_gpio_gen_filter_7__u_filter_diff_ctr_q[3]),
    .c(u_gpio_gen_filter_7__u_filter_diff_ctr_q[1]),
    .d(u_gpio_gen_filter_7__u_filter_diff_ctr_q[2]),
    .o1(n2639));
 b15nor002ah1n02x5 U3392 (.a(n2702),
    .b(n2639),
    .o1(u_gpio_gen_filter_7__u_filter_diff_ctr_d[0]));
 b15and003aq1n03x5 U3393 (.a(net2098),
    .b(u_gpio_gen_filter_5__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_5__u_filter_diff_ctr_q[1]),
    .o(n2925));
 b15inv040ah1n10x5 U3394 (.a(u_gpio_gen_filter_5__u_filter_filter_synced),
    .o1(n3398));
 b15xor002as1n06x5 U3395 (.a(net2074),
    .b(n3398),
    .out0(n2924));
 b15inv040aq1n03x5 U3396 (.a(n2924),
    .o1(n2928));
 b15oab012al1n03x5 U3397 (.a(n2928),
    .b(net2114),
    .c(n2925),
    .out0(u_gpio_gen_filter_5__u_filter_diff_ctr_d[3]));
 b15ztpn00an1n08x5 PHY_53 ();
 b15ztpn00an1n08x5 PHY_52 ();
 b15ztpn00an1n08x5 PHY_51 ();
 b15ztpn00an1n08x5 PHY_50 ();
 b15ztpn00an1n08x5 PHY_49 ();
 b15ztpn00an1n08x5 PHY_48 ();
 b15ztpn00an1n08x5 PHY_47 ();
 b15ztpn00an1n08x5 PHY_46 ();
 b15inv040aq1n02x5 U3406 (.a(u_gpio_gen_filter_7__u_filter_diff_ctr_q[3]),
    .o1(n2698));
 b15nandp3al1n08x5 U3407 (.a(u_gpio_gen_filter_7__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_7__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_7__u_filter_diff_ctr_q[2]),
    .o1(n3813));
 b15aoi012aq1n06x5 U3408 (.a(n2702),
    .b(n2698),
    .c(n3813),
    .o1(u_gpio_gen_filter_7__u_filter_diff_ctr_d[3]));
 b15inv000al1n02x5 U3409 (.a(u_gpio_gen_filter_27__u_filter_diff_ctr_q[3]),
    .o1(n2693));
 b15nand03an1n06x5 U3410 (.a(u_gpio_gen_filter_27__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_27__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_27__u_filter_diff_ctr_q[2]),
    .o1(n3817));
 b15aoi012al1n02x5 U3411 (.a(n2697),
    .b(n2693),
    .c(n3817),
    .o1(u_gpio_gen_filter_27__u_filter_diff_ctr_d[3]));
 b15inv000al1n12x5 U3412 (.a(net2131),
    .o1(n2849));
 b15nandp3an1n12x5 U3413 (.o1(n2847),
    .a(u_gpio_gen_filter_20__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_20__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_20__u_filter_diff_ctr_q[2]));
 b15xor002ah1n12x5 U3414 (.a(u_gpio_gen_filter_20__u_filter_filter_synced),
    .b(net2100),
    .out0(n2846));
 b15aoi012al1n04x5 U3415 (.a(n2846),
    .b(n2849),
    .c(n2847),
    .o1(u_gpio_gen_filter_20__u_filter_diff_ctr_d[3]));
 b15inv040ah1n06x5 U3416 (.a(net1968),
    .o1(n2831));
 b15nand03al1n16x5 U3417 (.a(u_gpio_gen_filter_28__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_28__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_28__u_filter_diff_ctr_q[2]),
    .o1(n2829));
 b15xor002as1n08x5 U3418 (.a(u_gpio_gen_filter_28__u_filter_filter_synced),
    .b(net1956),
    .out0(n2828));
 b15aoi012ar1n02x5 U3419 (.a(n2828),
    .b(n2831),
    .c(n2829),
    .o1(u_gpio_gen_filter_28__u_filter_diff_ctr_d[3]));
 b15inv000an1n16x5 U3420 (.a(net2112),
    .o1(n2879));
 b15nand03ah1n12x5 U3421 (.a(u_gpio_gen_filter_31__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_31__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_31__u_filter_diff_ctr_q[2]),
    .o1(n2877));
 b15xor002as1n16x5 U3422 (.a(u_gpio_gen_filter_31__u_filter_filter_synced),
    .b(u_gpio_gen_filter_31__u_filter_filter_q),
    .out0(n2876));
 b15aoi012ar1n02x5 U3423 (.a(n2876),
    .b(n2879),
    .c(n2877),
    .o1(u_gpio_gen_filter_31__u_filter_diff_ctr_d[3]));
 b15inv020ah1n12x5 U3424 (.a(net2054),
    .o1(n2843));
 b15nand03an1n16x5 U3425 (.a(u_gpio_gen_filter_4__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_4__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_4__u_filter_diff_ctr_q[2]),
    .o1(n2841));
 b15xor002an1n16x5 U3426 (.a(net441),
    .b(net2129),
    .out0(n2840));
 b15aoi012an1n02x5 U3427 (.a(n2840),
    .b(n2843),
    .c(n2841),
    .o1(u_gpio_gen_filter_4__u_filter_diff_ctr_d[3]));
 b15inv040as1n06x5 U3428 (.a(net1996),
    .o1(n2885));
 b15nandp3an1n12x5 U3429 (.o1(n2883),
    .a(u_gpio_gen_filter_13__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_13__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_13__u_filter_diff_ctr_q[2]));
 b15xor002ah1n12x5 U3430 (.a(u_gpio_gen_filter_13__u_filter_filter_synced),
    .b(net2056),
    .out0(n2882));
 b15aoi012al1n02x5 U3431 (.a(n2882),
    .b(n2885),
    .c(n2883),
    .o1(u_gpio_gen_filter_13__u_filter_diff_ctr_d[3]));
 b15inv040ar1n03x5 U3432 (.a(u_gpio_gen_filter_6__u_filter_diff_ctr_q[3]),
    .o1(n2645));
 b15aoi012al1n02x5 U3433 (.a(u_gpio_gen_filter_6__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_6__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_6__u_filter_diff_ctr_q[0]),
    .o1(n2644));
 b15aoi112an1n03x5 U3434 (.a(net2009),
    .b(n2644),
    .c(n2688),
    .d(n2645),
    .o1(u_gpio_gen_filter_6__u_filter_diff_ctr_d[2]));
 b15inv000al1n10x5 U3435 (.a(u_gpio_gen_filter_29__u_filter_diff_ctr_q[3]),
    .o1(n2861));
 b15nand03aq1n12x5 U3436 (.a(u_gpio_gen_filter_29__u_filter_diff_ctr_q[0]),
    .b(net1952),
    .c(u_gpio_gen_filter_29__u_filter_diff_ctr_q[2]),
    .o1(n2859));
 b15xor002an1n12x5 U3437 (.a(u_gpio_gen_filter_29__u_filter_filter_synced),
    .b(net1949),
    .out0(n2858));
 b15aoi012an1n02x5 U3438 (.a(n2858),
    .b(n2861),
    .c(net1953),
    .o1(u_gpio_gen_filter_29__u_filter_diff_ctr_d[3]));
 b15inv000an1n08x5 U3439 (.a(net2025),
    .o1(n2837));
 b15nandp3ah1n08x5 U3440 (.a(net1973),
    .b(u_gpio_gen_filter_18__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_18__u_filter_diff_ctr_q[2]),
    .o1(n2835));
 b15xor002as1n12x5 U3441 (.a(u_gpio_gen_filter_18__u_filter_filter_synced),
    .b(net2000),
    .out0(n2834));
 b15aoi012an1n02x5 U3442 (.a(n2834),
    .b(n2837),
    .c(n2835),
    .o1(u_gpio_gen_filter_18__u_filter_diff_ctr_d[3]));
 b15qbfin1bn1n16x5 U3443 (.a(net2102),
    .o1(n2867));
 b15nand03aq1n16x5 U3444 (.a(u_gpio_gen_filter_1__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_1__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_1__u_filter_diff_ctr_q[2]),
    .o1(n2865));
 b15xor002as1n16x5 U3445 (.a(u_gpio_gen_filter_1__u_filter_filter_synced),
    .b(u_gpio_gen_filter_1__u_filter_filter_q),
    .out0(n2864));
 b15aoi012al1n02x5 U3446 (.a(n2864),
    .b(n2867),
    .c(n2865),
    .o1(u_gpio_gen_filter_1__u_filter_diff_ctr_d[3]));
 b15inv000al1n12x5 U3447 (.a(net2073),
    .o1(n2873));
 b15nand03as1n12x5 U3448 (.a(u_gpio_gen_filter_9__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_9__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_9__u_filter_diff_ctr_q[2]),
    .o1(n2871));
 b15xor002an1n12x5 U3449 (.a(net439),
    .b(net2040),
    .out0(n2870));
 b15aoi012an1n02x5 U3450 (.a(n2870),
    .b(n2873),
    .c(n2871),
    .o1(u_gpio_gen_filter_9__u_filter_diff_ctr_d[3]));
 b15inv020ah1n08x5 U3451 (.a(net2061),
    .o1(n2825));
 b15nand03ah1n12x5 U3452 (.a(u_gpio_gen_filter_12__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_12__u_filter_diff_ctr_q[1]),
    .c(net2065),
    .o1(n2823));
 b15xor002al1n16x5 U3453 (.a(u_gpio_gen_filter_12__u_filter_filter_synced),
    .b(u_gpio_gen_filter_12__u_filter_filter_q),
    .out0(n2822));
 b15aoi012ar1n02x5 U3454 (.a(n2822),
    .b(n2825),
    .c(n2823),
    .o1(u_gpio_gen_filter_12__u_filter_diff_ctr_d[3]));
 b15inv000as1n10x5 U3455 (.a(u_gpio_gen_filter_8__u_filter_diff_ctr_q[3]),
    .o1(n2819));
 b15nandp3ah1n12x5 U3456 (.o1(n2817),
    .a(u_gpio_gen_filter_8__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_8__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_8__u_filter_diff_ctr_q[2]));
 b15xor002as1n16x5 U3457 (.a(u_gpio_gen_filter_8__u_filter_filter_synced),
    .b(net2028),
    .out0(n2816));
 b15aoi012al1n12x5 U3458 (.a(n2816),
    .b(n2819),
    .c(n2817),
    .o1(u_gpio_gen_filter_8__u_filter_diff_ctr_d[3]));
 b15inv020as1n10x5 U3459 (.a(u_gpio_gen_filter_3__u_filter_diff_ctr_q[3]),
    .o1(n2855));
 b15nand03as1n12x5 U3460 (.a(u_gpio_gen_filter_3__u_filter_diff_ctr_q[0]),
    .b(net2171),
    .c(net1982),
    .o1(n2853));
 b15xor002as1n08x5 U3461 (.a(u_gpio_gen_filter_3__u_filter_filter_synced),
    .b(u_gpio_gen_filter_3__u_filter_filter_q),
    .out0(n2852));
 b15aoi012as1n02x5 U3462 (.a(n2852),
    .b(n2855),
    .c(net1983),
    .o1(u_gpio_gen_filter_3__u_filter_diff_ctr_d[3]));
 b15inv000al1n02x5 U3463 (.a(u_gpio_gen_filter_11__u_filter_diff_ctr_q[3]),
    .o1(n2647));
 b15aoi012ar1n02x5 U3464 (.a(u_gpio_gen_filter_11__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_11__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_11__u_filter_diff_ctr_q[0]),
    .o1(n2646));
 b15aoi112an1n02x5 U3465 (.a(n2743),
    .b(n2646),
    .c(n2689),
    .d(n2647),
    .o1(u_gpio_gen_filter_11__u_filter_diff_ctr_d[2]));
 b15inv020an1n04x5 U3466 (.a(u_gpio_gen_filter_15__u_filter_diff_ctr_q[3]),
    .o1(n3814));
 b15and002al1n02x5 U3467 (.a(u_gpio_gen_filter_15__u_filter_diff_ctr_q[0]),
    .b(net2117),
    .o(n2677));
 b15norp02ar1n02x5 U3468 (.a(u_gpio_gen_filter_15__u_filter_diff_ctr_q[2]),
    .b(n2677),
    .o1(n2648));
 b15aoi112ah1n02x5 U3469 (.a(n2648),
    .b(n2736),
    .c(net2118),
    .d(n3814),
    .o1(u_gpio_gen_filter_15__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3470 (.a(n2823),
    .o1(n2650));
 b15aoi012ar1n02x5 U3471 (.a(u_gpio_gen_filter_12__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_12__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_12__u_filter_diff_ctr_q[0]),
    .o1(n2649));
 b15aoi112ar1n02x5 U3472 (.a(n2649),
    .b(n2822),
    .c(n2650),
    .d(n2825),
    .o1(u_gpio_gen_filter_12__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3473 (.a(n2883),
    .o1(n2652));
 b15aoi012al1n02x5 U3474 (.a(net2051),
    .b(u_gpio_gen_filter_13__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_13__u_filter_diff_ctr_q[0]),
    .o1(n2651));
 b15aoi112ar1n03x5 U3475 (.a(n2651),
    .b(n2882),
    .c(n2652),
    .d(n2885),
    .o1(u_gpio_gen_filter_13__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3476 (.a(n2835),
    .o1(n2654));
 b15aoi012al1n02x5 U3477 (.a(u_gpio_gen_filter_18__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_18__u_filter_diff_ctr_q[1]),
    .c(net2035),
    .o1(n2653));
 b15aoi112aq1n03x5 U3478 (.a(n2653),
    .b(n2834),
    .c(n2654),
    .d(n2837),
    .o1(u_gpio_gen_filter_18__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3479 (.a(n2865),
    .o1(n2656));
 b15aoi012ah1n02x5 U3480 (.a(u_gpio_gen_filter_1__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_1__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_1__u_filter_diff_ctr_q[0]),
    .o1(n2655));
 b15aoi112as1n02x5 U3481 (.a(n2655),
    .b(n2864),
    .c(n2656),
    .d(n2867),
    .o1(u_gpio_gen_filter_1__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3482 (.a(n2829),
    .o1(n2658));
 b15aoi012al1n02x5 U3483 (.a(u_gpio_gen_filter_28__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_28__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_28__u_filter_diff_ctr_q[0]),
    .o1(n2657));
 b15aoi112ar1n03x5 U3484 (.a(n2657),
    .b(n2828),
    .c(n2658),
    .d(n2831),
    .o1(u_gpio_gen_filter_28__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3485 (.a(n2859),
    .o1(n2660));
 b15aoi012al1n02x5 U3486 (.a(u_gpio_gen_filter_29__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_29__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_29__u_filter_diff_ctr_q[0]),
    .o1(n2659));
 b15aoi112ah1n02x5 U3487 (.a(n2659),
    .b(n2858),
    .c(n2660),
    .d(n2861),
    .o1(u_gpio_gen_filter_29__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3488 (.a(n2877),
    .o1(n2662));
 b15aoi012ar1n02x5 U3489 (.a(u_gpio_gen_filter_31__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_31__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_31__u_filter_diff_ctr_q[0]),
    .o1(n2661));
 b15aoi112ar1n02x5 U3490 (.a(n2661),
    .b(n2876),
    .c(n2662),
    .d(n2879),
    .o1(u_gpio_gen_filter_31__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3491 (.a(n2841),
    .o1(n2664));
 b15aoi012al1n02x5 U3492 (.a(u_gpio_gen_filter_4__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_4__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_4__u_filter_diff_ctr_q[0]),
    .o1(n2663));
 b15aoi112as1n02x5 U3493 (.a(n2663),
    .b(n2840),
    .c(n2664),
    .d(n2843),
    .o1(u_gpio_gen_filter_4__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3494 (.a(n2871),
    .o1(n2666));
 b15aoi012ar1n02x5 U3495 (.a(u_gpio_gen_filter_9__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_9__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_9__u_filter_diff_ctr_q[0]),
    .o1(n2665));
 b15aoi112aq1n02x5 U3496 (.a(n2665),
    .b(n2870),
    .c(n2666),
    .d(n2873),
    .o1(u_gpio_gen_filter_9__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3497 (.a(n2847),
    .o1(n2668));
 b15aoi012al1n02x5 U3498 (.a(u_gpio_gen_filter_20__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_20__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_20__u_filter_diff_ctr_q[0]),
    .o1(n2667));
 b15aoi112al1n03x5 U3499 (.a(n2667),
    .b(n2846),
    .c(n2668),
    .d(n2849),
    .o1(u_gpio_gen_filter_20__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3500 (.a(n2853),
    .o1(n2670));
 b15aoi012ar1n02x5 U3501 (.a(net1982),
    .b(net2202),
    .c(u_gpio_gen_filter_3__u_filter_diff_ctr_q[0]),
    .o1(n2669));
 b15aoi112ar1n02x5 U3502 (.a(n2669),
    .b(n2852),
    .c(n2670),
    .d(n2855),
    .o1(u_gpio_gen_filter_3__u_filter_diff_ctr_d[2]));
 b15inv040al1n02x5 U3503 (.a(n2817),
    .o1(n2672));
 b15aoi012al1n02x5 U3504 (.a(u_gpio_gen_filter_8__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_8__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_8__u_filter_diff_ctr_q[0]),
    .o1(n2671));
 b15aoi112al1n04x5 U3505 (.a(n2671),
    .b(n2816),
    .c(n2672),
    .d(n2819),
    .o1(u_gpio_gen_filter_8__u_filter_diff_ctr_d[2]));
 b15nand02ar1n02x5 U3506 (.a(u_gpio_gen_filter_23__u_filter_diff_ctr_q[3]),
    .b(u_gpio_gen_filter_23__u_filter_diff_ctr_q[2]),
    .o1(n2674));
 b15norp02ar1n02x5 U3507 (.a(u_gpio_gen_filter_23__u_filter_diff_ctr_q[1]),
    .b(net2089),
    .o1(n2673));
 b15aoi112ar1n02x3 U3508 (.a(n2673),
    .b(n2728),
    .c(n2675),
    .d(n2674),
    .o1(u_gpio_gen_filter_23__u_filter_diff_ctr_d[1]));
 b15and003an1n03x5 U3509 (.a(u_gpio_gen_filter_22__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_22__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_22__u_filter_diff_ctr_q[1]),
    .o(n2887));
 b15inv020al1n28x5 U3510 (.a(u_gpio_gen_filter_22__u_filter_filter_synced),
    .o1(n3510));
 b15xor002as1n16x5 U3511 (.a(net2003),
    .b(n3510),
    .out0(n2889));
 b15inv000ah1n04x5 U3512 (.a(n2889),
    .o1(n2888));
 b15oab012ar1n02x5 U3513 (.a(n2888),
    .b(net1993),
    .c(n2887),
    .out0(u_gpio_gen_filter_22__u_filter_diff_ctr_d[3]));
 b15nor002as1n03x5 U3514 (.a(u_gpio_gen_filter_15__u_filter_diff_ctr_q[0]),
    .b(net2117),
    .o1(n3815));
 b15nand02ah1n04x5 U3515 (.a(u_gpio_gen_filter_15__u_filter_diff_ctr_q[3]),
    .b(n2676),
    .o1(n2737));
 b15oaoi13al1n03x5 U3516 (.a(n2736),
    .b(n2737),
    .c(n3815),
    .d(n2677),
    .o1(u_gpio_gen_filter_15__u_filter_diff_ctr_d[1]));
 b15nand02ah1n03x5 U3517 (.a(u_gpio_gen_filter_14__u_filter_diff_ctr_q[3]),
    .b(u_gpio_gen_filter_14__u_filter_diff_ctr_q[2]),
    .o1(n2679));
 b15nor002ar1n03x5 U3518 (.a(net2186),
    .b(u_gpio_gen_filter_14__u_filter_diff_ctr_q[1]),
    .o1(n2678));
 b15aoi112as1n06x5 U3519 (.a(n2687),
    .b(n2678),
    .c(n2680),
    .d(n2679),
    .o1(u_gpio_gen_filter_14__u_filter_diff_ctr_d[1]));
 b15nandp2al1n02x5 U3520 (.a(net2169),
    .b(u_gpio_gen_filter_2__u_filter_diff_ctr_q[2]),
    .o1(n2682));
 b15norp02ar1n02x5 U3521 (.a(net2184),
    .b(u_gpio_gen_filter_2__u_filter_diff_ctr_q[1]),
    .o1(n2681));
 b15aoi112ah1n02x5 U3522 (.a(n2685),
    .b(n2681),
    .c(n2683),
    .d(n2682),
    .o1(u_gpio_gen_filter_2__u_filter_diff_ctr_d[1]));
 b15nor002ah1n02x5 U3523 (.a(n2685),
    .b(n2684),
    .o1(eq_x_221_n25));
 b15nor002aq1n03x5 U3524 (.a(n2687),
    .b(n2686),
    .o1(eq_x_161_n25));
 b15nand02an1n12x5 U3525 (.a(u_gpio_gen_filter_6__u_filter_diff_ctr_q[3]),
    .b(n2688),
    .o1(n2741));
 b15aoi012ar1n06x5 U3526 (.a(net2009),
    .b(u_gpio_gen_filter_6__u_filter_diff_ctr_q[0]),
    .c(n2741),
    .o1(u_gpio_gen_filter_6__u_filter_diff_ctr_d[0]));
 b15inv020aq1n03x5 U3527 (.a(u_gpio_gen_filter_25__u_filter_diff_ctr_q[3]),
    .o1(n2790));
 b15aoi012ah1n02x5 U3528 (.a(net2032),
    .b(u_gpio_gen_filter_25__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_25__u_filter_diff_ctr_q[0]),
    .o1(n2797));
 b15aoi112an1n02x5 U3529 (.a(net2033),
    .b(n2792),
    .c(n2791),
    .d(n2790),
    .o1(u_gpio_gen_filter_25__u_filter_diff_ctr_d[2]));
 b15inv020an1n03x5 U3530 (.a(u_gpio_gen_filter_0__u_filter_diff_ctr_q[3]),
    .o1(n2806));
 b15aoi012al1n06x5 U3531 (.a(net2004),
    .b(u_gpio_gen_filter_0__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_0__u_filter_diff_ctr_q[0]),
    .o1(n2813));
 b15aoi112ar1n03x5 U3532 (.a(n2813),
    .b(n2808),
    .c(n2807),
    .d(n2806),
    .o1(u_gpio_gen_filter_0__u_filter_diff_ctr_d[2]));
 b15inv020as1n03x5 U3533 (.a(u_gpio_gen_filter_17__u_filter_diff_ctr_q[3]),
    .o1(n2798));
 b15aoi012ar1n06x5 U3534 (.a(net2057),
    .b(u_gpio_gen_filter_17__u_filter_diff_ctr_q[1]),
    .c(net1977),
    .o1(n2805));
 b15aoi112al1n02x5 U3535 (.a(net2058),
    .b(n2800),
    .c(n2799),
    .d(n2798),
    .o1(u_gpio_gen_filter_17__u_filter_diff_ctr_d[2]));
 b15nandp2aq1n08x5 U3536 (.a(u_gpio_gen_filter_19__u_filter_diff_ctr_q[3]),
    .b(n2712),
    .o1(n2752));
 b15aoi012al1n02x5 U3537 (.a(n2707),
    .b(u_gpio_gen_filter_19__u_filter_diff_ctr_q[0]),
    .c(n2752),
    .o1(u_gpio_gen_filter_19__u_filter_diff_ctr_d[0]));
 b15nandp2aq1n04x5 U3538 (.a(u_gpio_gen_filter_24__u_filter_diff_ctr_q[3]),
    .b(n2718),
    .o1(n2749));
 b15aoi012an1n02x5 U3539 (.a(n2713),
    .b(net2143),
    .c(n2749),
    .o1(u_gpio_gen_filter_24__u_filter_diff_ctr_d[0]));
 b15inv040al1n02x5 U3540 (.a(net2159),
    .o1(n2773));
 b15nand03aq1n04x5 U3541 (.a(u_gpio_gen_filter_30__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_30__u_filter_diff_ctr_q[1]),
    .c(net2138),
    .o1(n2719));
 b15inv040an1n08x5 U3542 (.a(u_gpio_gen_filter_30__u_filter_filter_synced),
    .o1(n3516));
 b15xor002an1n12x5 U3543 (.a(net2157),
    .b(n3516),
    .out0(n2768));
 b15inv000al1n04x5 U3544 (.a(n2768),
    .o1(n2771));
 b15aoi012aq1n02x5 U3545 (.a(n2771),
    .b(n2773),
    .c(n2719),
    .o1(u_gpio_gen_filter_30__u_filter_diff_ctr_d[3]));
 b15inv000aq1n02x5 U3546 (.a(u_gpio_gen_filter_10__u_filter_diff_ctr_q[3]),
    .o1(n2759));
 b15nandp3ah1n03x5 U3547 (.a(net2163),
    .b(u_gpio_gen_filter_10__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_10__u_filter_diff_ctr_q[2]),
    .o1(n2720));
 b15inv000ar1n16x5 U3548 (.a(u_gpio_gen_filter_10__u_filter_filter_synced),
    .o1(n3374));
 b15xor002an1n12x5 U3549 (.a(u_gpio_gen_filter_10__u_filter_filter_q),
    .b(n3374),
    .out0(n2754));
 b15inv000al1n03x5 U3550 (.a(n2754),
    .o1(n2757));
 b15aoi012al1n04x5 U3551 (.a(n2757),
    .b(n2759),
    .c(net2164),
    .o1(u_gpio_gen_filter_10__u_filter_diff_ctr_d[3]));
 b15inv000al1n02x5 U3552 (.a(net2133),
    .o1(n2787));
 b15nand03aq1n02x5 U3553 (.a(u_gpio_gen_filter_16__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_16__u_filter_diff_ctr_q[1]),
    .c(net2016),
    .o1(n2721));
 b15inv000an1n28x5 U3554 (.a(u_gpio_gen_filter_16__u_filter_filter_synced),
    .o1(n3404));
 b15xor002as1n08x5 U3555 (.a(net2063),
    .b(n3404),
    .out0(n2782));
 b15inv000ar1n04x5 U3556 (.a(n2782),
    .o1(n2785));
 b15aoi012ar1n02x5 U3557 (.a(n2785),
    .b(n2787),
    .c(n2721),
    .o1(u_gpio_gen_filter_16__u_filter_diff_ctr_d[3]));
 b15inv040al1n02x5 U3558 (.a(u_gpio_gen_filter_26__u_filter_diff_ctr_q[3]),
    .o1(n2766));
 b15nand03ah1n03x5 U3559 (.a(u_gpio_gen_filter_26__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_26__u_filter_diff_ctr_q[1]),
    .c(net2174),
    .o1(n2723));
 b15inv040al1n10x5 U3560 (.a(u_gpio_gen_filter_26__u_filter_filter_synced),
    .o1(n3491));
 b15xor002as1n06x5 U3561 (.a(u_gpio_gen_filter_26__u_filter_filter_q),
    .b(n3491),
    .out0(n2761));
 b15inv040as1n02x5 U3562 (.a(n2761),
    .o1(n2764));
 b15aoi012ah1n02x5 U3563 (.a(n2764),
    .b(n2766),
    .c(n2723),
    .o1(u_gpio_gen_filter_26__u_filter_diff_ctr_d[3]));
 b15inv040aq1n02x5 U3564 (.a(u_gpio_gen_filter_21__u_filter_diff_ctr_q[3]),
    .o1(n2780));
 b15nand03al1n08x5 U3565 (.a(u_gpio_gen_filter_21__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_21__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_21__u_filter_diff_ctr_q[2]),
    .o1(n2722));
 b15inv000al1n20x5 U3566 (.a(u_gpio_gen_filter_21__u_filter_filter_synced),
    .o1(n3335));
 b15xor002ah1n16x5 U3567 (.a(u_gpio_gen_filter_21__u_filter_filter_q),
    .b(n3335),
    .out0(n2775));
 b15inv040ar1n03x5 U3568 (.a(n2775),
    .o1(n2778));
 b15aoi012ar1n06x5 U3569 (.a(n2778),
    .b(n2780),
    .c(n2722),
    .o1(u_gpio_gen_filter_21__u_filter_diff_ctr_d[3]));
 b15nand02ar1n02x5 U3570 (.a(net2221),
    .b(u_gpio_gen_filter_11__u_filter_diff_ctr_q[1]),
    .o1(n2691));
 b15nand02an1n04x5 U3571 (.a(u_gpio_gen_filter_11__u_filter_diff_ctr_q[3]),
    .b(n2689),
    .o1(n2744));
 b15inv000al1n02x5 U3572 (.a(n2744),
    .o1(n2690));
 b15oaoi13ar1n02x3 U3573 (.a(n2690),
    .b(n2691),
    .c(u_gpio_gen_filter_11__u_filter_diff_ctr_q[0]),
    .d(u_gpio_gen_filter_11__u_filter_diff_ctr_q[1]),
    .o1(n2692));
 b15norp02ar1n02x5 U3574 (.a(n2692),
    .b(n2743),
    .o1(u_gpio_gen_filter_11__u_filter_diff_ctr_d[1]));
 b15nand02ar1n02x5 U3575 (.a(u_gpio_gen_filter_27__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_27__u_filter_diff_ctr_q[1]),
    .o1(n2695));
 b15nor002al1n02x5 U3576 (.a(n2693),
    .b(n3817),
    .o1(n2694));
 b15oaoi13an1n02x5 U3577 (.a(n2694),
    .b(n2695),
    .c(u_gpio_gen_filter_27__u_filter_diff_ctr_q[0]),
    .d(u_gpio_gen_filter_27__u_filter_diff_ctr_q[1]),
    .o1(n2696));
 b15nor002aq1n02x5 U3578 (.a(n2697),
    .b(n2696),
    .o1(u_gpio_gen_filter_27__u_filter_diff_ctr_d[1]));
 b15nand02ar1n02x5 U3579 (.a(u_gpio_gen_filter_7__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_7__u_filter_diff_ctr_q[1]),
    .o1(n2700));
 b15norp02al1n02x5 U3580 (.a(n2698),
    .b(n3813),
    .o1(n2699));
 b15oaoi13ar1n02x3 U3581 (.a(n2699),
    .b(n2700),
    .c(u_gpio_gen_filter_7__u_filter_diff_ctr_q[0]),
    .d(u_gpio_gen_filter_7__u_filter_diff_ctr_q[1]),
    .o1(n2701));
 b15norp02ar1n02x5 U3582 (.a(n2702),
    .b(n2701),
    .o1(u_gpio_gen_filter_7__u_filter_diff_ctr_d[1]));
 b15nandp2an1n04x5 U3583 (.a(u_gpio_gen_filter_19__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_19__u_filter_diff_ctr_q[1]),
    .o1(n2708));
 b15inv000al1n02x5 U3584 (.a(n2752),
    .o1(n2703));
 b15oaoi13ar1n02x3 U3585 (.a(n2703),
    .b(n2708),
    .c(u_gpio_gen_filter_19__u_filter_diff_ctr_q[0]),
    .d(u_gpio_gen_filter_19__u_filter_diff_ctr_q[1]),
    .o1(n2704));
 b15nor002al1n02x5 U3586 (.a(n2707),
    .b(n2704),
    .o1(u_gpio_gen_filter_19__u_filter_diff_ctr_d[1]));
 b15nand02an1n02x5 U3587 (.a(u_gpio_gen_filter_24__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_24__u_filter_diff_ctr_q[1]),
    .o1(n2714));
 b15inv000al1n02x5 U3588 (.a(n2749),
    .o1(n2705));
 b15oaoi13ar1n02x3 U3589 (.a(n2705),
    .b(n2714),
    .c(u_gpio_gen_filter_24__u_filter_diff_ctr_q[0]),
    .d(u_gpio_gen_filter_24__u_filter_diff_ctr_q[1]),
    .o1(n2706));
 b15norp02an1n02x5 U3590 (.a(n2713),
    .b(n2706),
    .o1(u_gpio_gen_filter_24__u_filter_diff_ctr_d[1]));
 b15inv000al1n02x5 U3591 (.a(u_gpio_gen_filter_19__u_filter_diff_ctr_q[2]),
    .o1(n2709));
 b15aoi012ar1n06x5 U3592 (.a(n2707),
    .b(n2709),
    .c(n2708),
    .o1(n2710));
 b15inv040ar1n02x5 U3593 (.a(n2710),
    .o1(n2711));
 b15nand02ah1n06x5 U3594 (.a(n2710),
    .b(u_gpio_gen_filter_19__u_filter_diff_ctr_q[3]),
    .o1(n2751));
 b15oai012ah1n06x5 U3595 (.a(n2751),
    .b(net2045),
    .c(n2711),
    .o1(u_gpio_gen_filter_19__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3596 (.a(net2113),
    .o1(n2715));
 b15aoi012ah1n02x5 U3597 (.a(n2713),
    .b(n2715),
    .c(n2714),
    .o1(n2716));
 b15inv000al1n02x5 U3598 (.a(n2716),
    .o1(n2717));
 b15nand02ah1n03x5 U3599 (.a(n2716),
    .b(u_gpio_gen_filter_24__u_filter_diff_ctr_q[3]),
    .o1(n2748));
 b15oai012al1n02x5 U3600 (.a(n2748),
    .b(n2718),
    .c(n2717),
    .o1(u_gpio_gen_filter_24__u_filter_diff_ctr_d[2]));
 b15nandp2as1n02x5 U3601 (.a(net1993),
    .b(n2889),
    .o1(n2886));
 b15aoi012an1n12x5 U3602 (.a(u_gpio_gen_filter_22__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_22__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_22__u_filter_diff_ctr_q[1]),
    .o1(n2894));
 b15oaoi13ah1n03x5 U3603 (.a(n2894),
    .b(net1994),
    .c(n2888),
    .d(n2887),
    .o1(u_gpio_gen_filter_22__u_filter_diff_ctr_d[2]));
 b15aoai13aq1n04x5 U3604 (.a(n2768),
    .b(net2138),
    .c(u_gpio_gen_filter_30__u_filter_diff_ctr_q[1]),
    .d(u_gpio_gen_filter_30__u_filter_diff_ctr_q[0]),
    .o1(n2772));
 b15oab012ar1n02x5 U3605 (.a(n2772),
    .b(u_gpio_gen_filter_30__u_filter_diff_ctr_q[3]),
    .c(n2719),
    .out0(u_gpio_gen_filter_30__u_filter_diff_ctr_d[2]));
 b15aoai13ar1n04x5 U3606 (.a(n2754),
    .b(net2220),
    .c(u_gpio_gen_filter_10__u_filter_diff_ctr_q[1]),
    .d(u_gpio_gen_filter_10__u_filter_diff_ctr_q[0]),
    .o1(n2758));
 b15oab012aq1n02x5 U3607 (.a(n2758),
    .b(u_gpio_gen_filter_10__u_filter_diff_ctr_q[3]),
    .c(net2164),
    .out0(u_gpio_gen_filter_10__u_filter_diff_ctr_d[2]));
 b15aoai13ah1n02x5 U3608 (.a(n2782),
    .b(net2016),
    .c(u_gpio_gen_filter_16__u_filter_diff_ctr_q[1]),
    .d(u_gpio_gen_filter_16__u_filter_diff_ctr_q[0]),
    .o1(n2786));
 b15oab012ar1n02x5 U3609 (.a(n2786),
    .b(u_gpio_gen_filter_16__u_filter_diff_ctr_q[3]),
    .c(n2721),
    .out0(u_gpio_gen_filter_16__u_filter_diff_ctr_d[2]));
 b15aoai13an1n06x5 U3610 (.a(n2775),
    .b(u_gpio_gen_filter_21__u_filter_diff_ctr_q[2]),
    .c(u_gpio_gen_filter_21__u_filter_diff_ctr_q[1]),
    .d(u_gpio_gen_filter_21__u_filter_diff_ctr_q[0]),
    .o1(n2779));
 b15oab012an1n02x5 U3611 (.a(n2779),
    .b(net2219),
    .c(n2722),
    .out0(u_gpio_gen_filter_21__u_filter_diff_ctr_d[2]));
 b15aoai13an1n03x5 U3612 (.a(n2761),
    .b(net2214),
    .c(u_gpio_gen_filter_26__u_filter_diff_ctr_q[1]),
    .d(u_gpio_gen_filter_26__u_filter_diff_ctr_q[0]),
    .o1(n2765));
 b15oab012ar1n02x5 U3613 (.a(n2765),
    .b(u_gpio_gen_filter_26__u_filter_diff_ctr_q[3]),
    .c(n2723),
    .out0(u_gpio_gen_filter_26__u_filter_diff_ctr_d[2]));
 b15aoai13aq1n06x5 U3614 (.a(n2724),
    .b(u_gpio_gen_filter_7__u_filter_diff_ctr_q[2]),
    .c(u_gpio_gen_filter_7__u_filter_diff_ctr_q[1]),
    .d(u_gpio_gen_filter_7__u_filter_diff_ctr_q[0]),
    .o1(n3812));
 b15nand03ah1n03x5 U3615 (.a(u_gpio_gen_filter_7__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_7__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_7__u_filter_diff_ctr_q[3]),
    .o1(n2725));
 b15nor002ar1n04x5 U3616 (.a(n3812),
    .b(n2725),
    .o1(eq_x_196_n25));
 b15aoai13aq1n04x5 U3617 (.a(n2726),
    .b(u_gpio_gen_filter_27__u_filter_diff_ctr_q[2]),
    .c(u_gpio_gen_filter_27__u_filter_diff_ctr_q[1]),
    .d(u_gpio_gen_filter_27__u_filter_diff_ctr_q[0]),
    .o1(n3816));
 b15nandp3ar1n03x5 U3618 (.a(u_gpio_gen_filter_27__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_27__u_filter_diff_ctr_q[1]),
    .c(u_gpio_gen_filter_27__u_filter_diff_ctr_q[3]),
    .o1(n2727));
 b15norp02aq1n04x5 U3619 (.a(n3816),
    .b(n2727),
    .o1(eq_x_96_n25));
 b15inv000al1n02x5 U3620 (.a(u_gpio_gen_filter_23__u_filter_diff_ctr_q[3]),
    .o1(n2730));
 b15aoi012as1n02x5 U3621 (.a(n2728),
    .b(n2730),
    .c(n2729),
    .o1(u_gpio_gen_filter_23__u_filter_diff_ctr_d[3]));
 b15nonb02ar1n12x5 U3622 (.a(u_gpio_gen_filter_23__u_filter_diff_ctr_d[3]),
    .b(n2731),
    .out0(eq_x_116_n25));
 b15norp02aq1n03x5 U3623 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nd),
    .o1(n2735));
 b15inv000al1n02x5 U3624 (.a(n2735),
    .o1(n2733));
 b15nand03al1n02x5 U3625 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq),
    .c(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq),
    .o1(n2732));
 b15oai013ah1n03x5 U3626 (.a(n2732),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq),
    .c(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq),
    .d(n2733),
    .o1(n2734));
 b15norp03al1n08x5 U3627 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[0]),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[1]),
    .c(n2734),
    .o1(n3038));
 b15aoi012aq1n08x5 U3628 (.a(n2735),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nd),
    .c(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .o1(n3039));
 b15nonb02ar1n03x5 U3629 (.a(n3038),
    .b(n3039),
    .out0(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[0]));
 b15aoi012ah1n04x5 U3630 (.a(n2736),
    .b(net2006),
    .c(n2737),
    .o1(u_gpio_gen_filter_15__u_filter_diff_ctr_d[0]));
 b15inv020ah1n12x5 U3631 (.a(net1784),
    .o1(n2906));
 b15orn003as1n24x5 U3632 (.a(n2906),
    .b(net1859),
    .c(net1915),
    .o(n3620));
 b15inv000an1n16x5 U3633 (.a(net1822),
    .o1(n3045));
 b15nor002an1n03x5 U3634 (.a(net1860),
    .b(net1823),
    .o1(net167));
 b15nand02ar1n02x5 U3635 (.a(u_gpio_gen_filter_6__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_6__u_filter_diff_ctr_q[1]),
    .o1(n2738));
 b15oai012an1n04x5 U3636 (.a(n2738),
    .b(u_gpio_gen_filter_6__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_6__u_filter_diff_ctr_q[1]),
    .o1(n2740));
 b15aoi012ah1n06x5 U3637 (.a(net2009),
    .b(n2741),
    .c(n2740),
    .o1(u_gpio_gen_filter_6__u_filter_diff_ctr_d[1]));
 b15nand03ar1n12x5 U3638 (.a(u_gpio_gen_filter_6__u_filter_diff_ctr_q[1]),
    .b(u_gpio_gen_filter_6__u_filter_diff_ctr_q[2]),
    .c(u_gpio_gen_filter_6__u_filter_diff_ctr_q[3]),
    .o1(n2742));
 b15nonb02an1n16x5 U3639 (.a(u_gpio_gen_filter_6__u_filter_diff_ctr_d[1]),
    .b(n2742),
    .out0(eq_x_201_n25));
 b15aoi012an1n04x5 U3640 (.a(n2743),
    .b(net2111),
    .c(n2744),
    .o1(u_gpio_gen_filter_11__u_filter_diff_ctr_d[0]));
 b15nand03as1n04x5 U3641 (.a(u_gpio_gen_filter_11__u_filter_diff_ctr_q[1]),
    .b(u_gpio_gen_filter_11__u_filter_diff_ctr_q[2]),
    .c(u_gpio_gen_filter_11__u_filter_diff_ctr_q[3]),
    .o1(n2745));
 b15nonb02al1n03x5 U3642 (.a(u_gpio_gen_filter_11__u_filter_diff_ctr_d[0]),
    .b(n2745),
    .out0(eq_x_176_n25));
 b15inv020as1n08x5 U3643 (.a(net1849),
    .o1(n2923));
 b15oai012aq1n32x5 U3644 (.a(net1915),
    .b(net1784),
    .c(net1859),
    .o1(n3617));
 b15oai012aq1n06x5 U3645 (.a(net1916),
    .b(net1860),
    .c(n2923),
    .o1(net122));
 b15xor002al1n16x5 U3646 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq),
    .b(n2746),
    .out0(n3215));
 b15xor002as1n08x5 U3647 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq),
    .b(n2747),
    .out0(n3216));
 b15aoi112ah1n06x5 U3648 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[0]),
    .c(n3215),
    .d(n3216),
    .o1(n3040));
 b15aoi022as1n16x5 U3649 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd),
    .c(n2747),
    .d(n2746),
    .o1(n3217));
 b15nonb02ar1n02x3 U3650 (.a(n3040),
    .b(n3217),
    .out0(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[0]));
 b15inv040ar1n02x5 U3651 (.a(u_gpio_gen_filter_24__u_filter_diff_ctr_q[1]),
    .o1(n2750));
 b15oaoi13an1n04x5 U3652 (.a(n2748),
    .b(n2749),
    .c(u_gpio_gen_filter_24__u_filter_diff_ctr_q[0]),
    .d(n2750),
    .o1(eq_x_111_n25));
 b15inv020ar1n05x5 U3653 (.a(u_gpio_gen_filter_19__u_filter_diff_ctr_q[1]),
    .o1(n2753));
 b15oaoi13as1n08x5 U3654 (.a(n2751),
    .b(n2752),
    .c(u_gpio_gen_filter_19__u_filter_diff_ctr_q[0]),
    .d(n2753),
    .o1(eq_x_136_n25));
 b15oai012an1n03x5 U3655 (.a(n2754),
    .b(net2163),
    .c(u_gpio_gen_filter_10__u_filter_diff_ctr_q[1]),
    .o1(n2755));
 b15nand04al1n08x5 U3656 (.a(u_gpio_gen_filter_10__u_filter_diff_ctr_q[1]),
    .b(u_gpio_gen_filter_10__u_filter_diff_ctr_q[3]),
    .c(net2190),
    .d(n2754),
    .o1(n2756));
 b15aoai13al1n06x5 U3657 (.a(n2756),
    .b(n2755),
    .c(u_gpio_gen_filter_10__u_filter_diff_ctr_q[1]),
    .d(net2079),
    .o1(u_gpio_gen_filter_10__u_filter_diff_ctr_d[1]));
 b15oai012ah1n04x5 U3658 (.a(n2756),
    .b(net2079),
    .c(n2757),
    .o1(u_gpio_gen_filter_10__u_filter_diff_ctr_d[0]));
 b15norp02an1n02x5 U3659 (.a(n2759),
    .b(n2758),
    .o1(n2760));
 b15and003as1n04x5 U3660 (.a(n2760),
    .b(u_gpio_gen_filter_10__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_10__u_filter_diff_ctr_d[0]),
    .o(eq_x_181_n25));
 b15oai012ah1n02x5 U3661 (.a(n2761),
    .b(u_gpio_gen_filter_26__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_26__u_filter_diff_ctr_q[1]),
    .o1(n2762));
 b15nand04ar1n12x5 U3662 (.a(u_gpio_gen_filter_26__u_filter_diff_ctr_q[1]),
    .b(u_gpio_gen_filter_26__u_filter_diff_ctr_q[3]),
    .c(net2207),
    .d(n2761),
    .o1(n2763));
 b15aoai13aq1n06x5 U3663 (.a(n2763),
    .b(n2762),
    .c(u_gpio_gen_filter_26__u_filter_diff_ctr_q[1]),
    .d(u_gpio_gen_filter_26__u_filter_diff_ctr_q[0]),
    .o1(u_gpio_gen_filter_26__u_filter_diff_ctr_d[1]));
 b15oai012aq1n06x5 U3664 (.a(n2763),
    .b(u_gpio_gen_filter_26__u_filter_diff_ctr_q[0]),
    .c(n2764),
    .o1(u_gpio_gen_filter_26__u_filter_diff_ctr_d[0]));
 b15norp02al1n02x5 U3665 (.a(n2766),
    .b(n2765),
    .o1(n2767));
 b15and003as1n02x5 U3666 (.a(n2767),
    .b(u_gpio_gen_filter_26__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_26__u_filter_diff_ctr_d[0]),
    .o(eq_x_101_n25));
 b15oai012ah1n02x5 U3667 (.a(n2768),
    .b(u_gpio_gen_filter_30__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_30__u_filter_diff_ctr_q[1]),
    .o1(n2769));
 b15nand04an1n08x5 U3668 (.a(u_gpio_gen_filter_30__u_filter_diff_ctr_q[1]),
    .b(u_gpio_gen_filter_30__u_filter_diff_ctr_q[3]),
    .c(net2138),
    .d(n2768),
    .o1(n2770));
 b15aoai13an1n06x5 U3669 (.a(net2139),
    .b(n2769),
    .c(u_gpio_gen_filter_30__u_filter_diff_ctr_q[1]),
    .d(u_gpio_gen_filter_30__u_filter_diff_ctr_q[0]),
    .o1(u_gpio_gen_filter_30__u_filter_diff_ctr_d[1]));
 b15oai012ar1n08x5 U3670 (.a(net2139),
    .b(u_gpio_gen_filter_30__u_filter_diff_ctr_q[0]),
    .c(n2771),
    .o1(u_gpio_gen_filter_30__u_filter_diff_ctr_d[0]));
 b15norp02al1n02x5 U3671 (.a(n2773),
    .b(n2772),
    .o1(n2774));
 b15and003ar1n03x5 U3672 (.a(n2774),
    .b(u_gpio_gen_filter_30__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_30__u_filter_diff_ctr_d[0]),
    .o(eq_x_81_n25));
 b15oai012ar1n02x5 U3673 (.a(n2775),
    .b(u_gpio_gen_filter_21__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_21__u_filter_diff_ctr_q[1]),
    .o1(n2776));
 b15nand04as1n03x5 U3674 (.a(u_gpio_gen_filter_21__u_filter_diff_ctr_q[1]),
    .b(net2187),
    .c(u_gpio_gen_filter_21__u_filter_diff_ctr_q[2]),
    .d(n2775),
    .o1(n2777));
 b15aoai13an1n03x5 U3675 (.a(net2188),
    .b(n2776),
    .c(u_gpio_gen_filter_21__u_filter_diff_ctr_q[1]),
    .d(u_gpio_gen_filter_21__u_filter_diff_ctr_q[0]),
    .o1(u_gpio_gen_filter_21__u_filter_diff_ctr_d[1]));
 b15oai012as1n03x5 U3676 (.a(n2777),
    .b(net2092),
    .c(n2778),
    .o1(u_gpio_gen_filter_21__u_filter_diff_ctr_d[0]));
 b15norp02an1n02x5 U3677 (.a(n2780),
    .b(n2779),
    .o1(n2781));
 b15and003ah1n03x5 U3678 (.a(n2781),
    .b(u_gpio_gen_filter_21__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_21__u_filter_diff_ctr_d[0]),
    .o(eq_x_126_n25));
 b15oai012ar1n02x5 U3679 (.a(n2782),
    .b(u_gpio_gen_filter_16__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_16__u_filter_diff_ctr_q[1]),
    .o1(n2783));
 b15nand04as1n06x5 U3680 (.a(u_gpio_gen_filter_16__u_filter_diff_ctr_q[1]),
    .b(u_gpio_gen_filter_16__u_filter_diff_ctr_q[3]),
    .c(net2016),
    .d(n2782),
    .o1(n2784));
 b15aoai13aq1n04x5 U3681 (.a(net2017),
    .b(n2783),
    .c(u_gpio_gen_filter_16__u_filter_diff_ctr_q[1]),
    .d(u_gpio_gen_filter_16__u_filter_diff_ctr_q[0]),
    .o1(u_gpio_gen_filter_16__u_filter_diff_ctr_d[1]));
 b15oai012an1n06x5 U3682 (.a(net2017),
    .b(net2038),
    .c(n2785),
    .o1(u_gpio_gen_filter_16__u_filter_diff_ctr_d[0]));
 b15nor002an1n03x5 U3683 (.a(n2787),
    .b(n2786),
    .o1(n2788));
 b15and003ah1n03x5 U3684 (.a(n2788),
    .b(u_gpio_gen_filter_16__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_16__u_filter_diff_ctr_d[0]),
    .o(eq_x_151_n25));
 b15aoai13al1n06x5 U3685 (.a(n2924),
    .b(net2098),
    .c(u_gpio_gen_filter_5__u_filter_diff_ctr_q[0]),
    .d(u_gpio_gen_filter_5__u_filter_diff_ctr_q[1]),
    .o1(n2789));
 b15nonb02al1n06x5 U3686 (.a(u_gpio_gen_filter_5__u_filter_diff_ctr_q[3]),
    .b(n2789),
    .out0(n2929));
 b15oabi12as1n02x5 U3687 (.a(n2929),
    .b(n2925),
    .c(n2789),
    .out0(u_gpio_gen_filter_5__u_filter_diff_ctr_d[2]));
 b15inv020as1n05x5 U3688 (.a(net1890),
    .o1(n2940));
 b15inv020ah1n05x5 U3689 (.a(net1795),
    .o1(n2918));
 b15oai022ah1n04x5 U3690 (.a(n3620),
    .b(n2940),
    .c(n3617),
    .d(net1796),
    .o1(net162));
 b15aoi022ah1n08x5 U3691 (.a(net1822),
    .b(n2940),
    .c(net1890),
    .d(net1823),
    .o1(n2922));
 b15oa0022ar1n03x5 U3692 (.a(n3617),
    .b(net1796),
    .c(net1891),
    .d(net1860),
    .o(net114));
 b15norp02ar1n03x5 U3693 (.a(n2790),
    .b(n2792),
    .o1(n2795));
 b15nandp2ar1n04x5 U3694 (.a(n2795),
    .b(n2791),
    .o1(n2793));
 b15oai012as1n04x5 U3695 (.a(n2793),
    .b(u_gpio_gen_filter_25__u_filter_diff_ctr_q[0]),
    .c(n2792),
    .o1(u_gpio_gen_filter_25__u_filter_diff_ctr_d[0]));
 b15oabi12al1n02x5 U3696 (.a(n2792),
    .b(u_gpio_gen_filter_25__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_25__u_filter_diff_ctr_q[1]),
    .out0(n2794));
 b15aoai13ar1n04x5 U3697 (.a(n2793),
    .b(n2794),
    .c(net2107),
    .d(u_gpio_gen_filter_25__u_filter_diff_ctr_q[0]),
    .o1(u_gpio_gen_filter_25__u_filter_diff_ctr_d[1]));
 b15nand03al1n02x5 U3698 (.a(n2795),
    .b(u_gpio_gen_filter_25__u_filter_diff_ctr_d[0]),
    .c(u_gpio_gen_filter_25__u_filter_diff_ctr_d[1]),
    .o1(n2796));
 b15norp02aq1n04x5 U3699 (.a(n2797),
    .b(n2796),
    .o1(eq_x_106_n25));
 b15norp02al1n04x5 U3700 (.a(n2798),
    .b(n2800),
    .o1(n2803));
 b15nand02aq1n04x5 U3701 (.a(n2803),
    .b(n2799),
    .o1(n2801));
 b15oai012ah1n06x5 U3702 (.a(n2801),
    .b(net1977),
    .c(n2800),
    .o1(u_gpio_gen_filter_17__u_filter_diff_ctr_d[0]));
 b15oabi12ar1n02x5 U3703 (.a(n2800),
    .b(u_gpio_gen_filter_17__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_17__u_filter_diff_ctr_q[1]),
    .out0(n2802));
 b15aoai13ah1n02x5 U3704 (.a(n2801),
    .b(n2802),
    .c(u_gpio_gen_filter_17__u_filter_diff_ctr_q[1]),
    .d(net1977),
    .o1(u_gpio_gen_filter_17__u_filter_diff_ctr_d[1]));
 b15nand03an1n03x5 U3705 (.a(n2803),
    .b(u_gpio_gen_filter_17__u_filter_diff_ctr_d[0]),
    .c(u_gpio_gen_filter_17__u_filter_diff_ctr_d[1]),
    .o1(n2804));
 b15nor002aq1n03x5 U3706 (.a(n2805),
    .b(n2804),
    .o1(eq_x_146_n25));
 b15nor002an1n03x5 U3707 (.a(n2806),
    .b(n2808),
    .o1(n2811));
 b15nand02al1n06x5 U3708 (.a(n2811),
    .b(n2807),
    .o1(n2809));
 b15oai012ah1n06x5 U3709 (.a(n2809),
    .b(u_gpio_gen_filter_0__u_filter_diff_ctr_q[0]),
    .c(n2808),
    .o1(u_gpio_gen_filter_0__u_filter_diff_ctr_d[0]));
 b15oabi12an1n04x5 U3710 (.a(n2808),
    .b(u_gpio_gen_filter_0__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_0__u_filter_diff_ctr_q[1]),
    .out0(n2810));
 b15aoai13as1n06x5 U3711 (.a(n2809),
    .b(n2810),
    .c(net2136),
    .d(u_gpio_gen_filter_0__u_filter_diff_ctr_q[0]),
    .o1(u_gpio_gen_filter_0__u_filter_diff_ctr_d[1]));
 b15nand03ah1n04x5 U3712 (.a(n2811),
    .b(u_gpio_gen_filter_0__u_filter_diff_ctr_d[0]),
    .c(u_gpio_gen_filter_0__u_filter_diff_ctr_d[1]),
    .o1(n2812));
 b15nor002ah1n04x5 U3713 (.a(n2813),
    .b(n2812),
    .o1(eq_x_231_n25));
 b15nand02ar1n02x5 U3714 (.a(u_gpio_gen_filter_8__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_8__u_filter_diff_ctr_q[1]),
    .o1(n2814));
 b15oai012an1n02x5 U3715 (.a(n2814),
    .b(u_gpio_gen_filter_8__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_8__u_filter_diff_ctr_q[1]),
    .o1(n2815));
 b15oaoi13an1n04x5 U3716 (.a(n2816),
    .b(n2815),
    .c(n2819),
    .d(n2817),
    .o1(u_gpio_gen_filter_8__u_filter_diff_ctr_d[1]));
 b15oaoi13as1n08x5 U3717 (.a(n2816),
    .b(u_gpio_gen_filter_8__u_filter_diff_ctr_q[0]),
    .c(n2819),
    .d(n2817),
    .o1(u_gpio_gen_filter_8__u_filter_diff_ctr_d[0]));
 b15nand03ar1n06x5 U3718 (.a(u_gpio_gen_filter_8__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_8__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_8__u_filter_diff_ctr_d[0]),
    .o1(n2818));
 b15nor002as1n06x5 U3719 (.a(n2819),
    .b(n2818),
    .o1(eq_x_191_n25));
 b15nand02ar1n02x5 U3720 (.a(u_gpio_gen_filter_12__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_12__u_filter_diff_ctr_q[1]),
    .o1(n2820));
 b15oai012ar1n04x5 U3721 (.a(n2820),
    .b(u_gpio_gen_filter_12__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_12__u_filter_diff_ctr_q[1]),
    .o1(n2821));
 b15oaoi13aq1n03x5 U3722 (.a(n2822),
    .b(n2821),
    .c(n2825),
    .d(n2823),
    .o1(u_gpio_gen_filter_12__u_filter_diff_ctr_d[1]));
 b15oaoi13as1n08x5 U3723 (.a(n2822),
    .b(u_gpio_gen_filter_12__u_filter_diff_ctr_q[0]),
    .c(n2825),
    .d(n2823),
    .o1(u_gpio_gen_filter_12__u_filter_diff_ctr_d[0]));
 b15nandp3aq1n02x5 U3724 (.a(net2065),
    .b(u_gpio_gen_filter_12__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_12__u_filter_diff_ctr_d[0]),
    .o1(n2824));
 b15norp02al1n03x5 U3725 (.a(n2825),
    .b(n2824),
    .o1(eq_x_171_n25));
 b15nand02ar1n02x5 U3726 (.a(u_gpio_gen_filter_28__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_28__u_filter_diff_ctr_q[1]),
    .o1(n2826));
 b15oai012ah1n03x5 U3727 (.a(n2826),
    .b(u_gpio_gen_filter_28__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_28__u_filter_diff_ctr_q[1]),
    .o1(n2827));
 b15oaoi13ar1n08x5 U3728 (.a(n2828),
    .b(n2827),
    .c(n2831),
    .d(n2829),
    .o1(u_gpio_gen_filter_28__u_filter_diff_ctr_d[1]));
 b15oaoi13ah1n04x5 U3729 (.a(n2828),
    .b(u_gpio_gen_filter_28__u_filter_diff_ctr_q[0]),
    .c(n2831),
    .d(n2829),
    .o1(u_gpio_gen_filter_28__u_filter_diff_ctr_d[0]));
 b15nand03an1n04x5 U3730 (.a(u_gpio_gen_filter_28__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_28__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_28__u_filter_diff_ctr_d[0]),
    .o1(n2830));
 b15norp02ah1n04x5 U3731 (.a(n2831),
    .b(n2830),
    .o1(eq_x_91_n25));
 b15nand02ar1n02x5 U3732 (.a(u_gpio_gen_filter_18__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_18__u_filter_diff_ctr_q[1]),
    .o1(n2832));
 b15oai012aq1n03x5 U3733 (.a(n2832),
    .b(net1973),
    .c(u_gpio_gen_filter_18__u_filter_diff_ctr_q[1]),
    .o1(n2833));
 b15oaoi13al1n04x5 U3734 (.a(n2834),
    .b(n2833),
    .c(n2837),
    .d(n2835),
    .o1(u_gpio_gen_filter_18__u_filter_diff_ctr_d[1]));
 b15oaoi13ah1n03x5 U3735 (.a(n2834),
    .b(net1973),
    .c(n2837),
    .d(n2835),
    .o1(u_gpio_gen_filter_18__u_filter_diff_ctr_d[0]));
 b15nand03al1n03x5 U3736 (.a(u_gpio_gen_filter_18__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_18__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_18__u_filter_diff_ctr_d[0]),
    .o1(n2836));
 b15norp02ar1n04x5 U3737 (.a(n2837),
    .b(n2836),
    .o1(eq_x_141_n25));
 b15nand02ar1n02x5 U3738 (.a(u_gpio_gen_filter_4__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_4__u_filter_diff_ctr_q[1]),
    .o1(n2838));
 b15oai012an1n03x5 U3739 (.a(n2838),
    .b(u_gpio_gen_filter_4__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_4__u_filter_diff_ctr_q[1]),
    .o1(n2839));
 b15oaoi13aq1n04x5 U3740 (.a(n2840),
    .b(n2839),
    .c(n2843),
    .d(n2841),
    .o1(u_gpio_gen_filter_4__u_filter_diff_ctr_d[1]));
 b15oaoi13an1n08x5 U3741 (.a(n2840),
    .b(u_gpio_gen_filter_4__u_filter_diff_ctr_q[0]),
    .c(n2843),
    .d(n2841),
    .o1(u_gpio_gen_filter_4__u_filter_diff_ctr_d[0]));
 b15nand03ar1n06x5 U3742 (.a(u_gpio_gen_filter_4__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_4__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_4__u_filter_diff_ctr_d[0]),
    .o1(n2842));
 b15norp02al1n02x5 U3743 (.a(n2843),
    .b(n2842),
    .o1(eq_x_211_n25));
 b15nand02ar1n02x5 U3744 (.a(u_gpio_gen_filter_20__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_20__u_filter_diff_ctr_q[1]),
    .o1(n2844));
 b15oai012al1n02x5 U3745 (.a(n2844),
    .b(u_gpio_gen_filter_20__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_20__u_filter_diff_ctr_q[1]),
    .o1(n2845));
 b15oaoi13ah1n03x5 U3746 (.a(n2846),
    .b(n2845),
    .c(n2849),
    .d(n2847),
    .o1(u_gpio_gen_filter_20__u_filter_diff_ctr_d[1]));
 b15oaoi13an1n04x5 U3747 (.a(n2846),
    .b(net2132),
    .c(n2849),
    .d(n2847),
    .o1(u_gpio_gen_filter_20__u_filter_diff_ctr_d[0]));
 b15nandp3ah1n04x5 U3748 (.a(u_gpio_gen_filter_20__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_20__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_20__u_filter_diff_ctr_d[0]),
    .o1(n2848));
 b15norp02ar1n08x5 U3749 (.a(n2849),
    .b(n2848),
    .o1(eq_x_131_n25));
 b15nand02ar1n02x5 U3750 (.a(u_gpio_gen_filter_3__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_3__u_filter_diff_ctr_q[1]),
    .o1(n2850));
 b15oai012ah1n02x5 U3751 (.a(n2850),
    .b(u_gpio_gen_filter_3__u_filter_diff_ctr_q[0]),
    .c(net2171),
    .o1(n2851));
 b15oaoi13as1n04x5 U3752 (.a(n2852),
    .b(net2172),
    .c(n2855),
    .d(net1983),
    .o1(u_gpio_gen_filter_3__u_filter_diff_ctr_d[1]));
 b15oaoi13as1n03x5 U3753 (.a(n2852),
    .b(net2109),
    .c(n2855),
    .d(net1983),
    .o1(u_gpio_gen_filter_3__u_filter_diff_ctr_d[0]));
 b15nand03ah1n04x5 U3754 (.a(net2218),
    .b(u_gpio_gen_filter_3__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_3__u_filter_diff_ctr_d[0]),
    .o1(n2854));
 b15nor002al1n04x5 U3755 (.a(n2855),
    .b(n2854),
    .o1(eq_x_216_n25));
 b15nand02ar1n02x5 U3756 (.a(u_gpio_gen_filter_29__u_filter_diff_ctr_q[0]),
    .b(net2096),
    .o1(n2856));
 b15oai012ah1n02x5 U3757 (.a(n2856),
    .b(u_gpio_gen_filter_29__u_filter_diff_ctr_q[0]),
    .c(net1952),
    .o1(n2857));
 b15oaoi13an1n04x5 U3758 (.a(n2858),
    .b(n2857),
    .c(n2861),
    .d(n2859),
    .o1(u_gpio_gen_filter_29__u_filter_diff_ctr_d[1]));
 b15oaoi13aq1n04x5 U3759 (.a(n2858),
    .b(net2088),
    .c(n2861),
    .d(n2859),
    .o1(u_gpio_gen_filter_29__u_filter_diff_ctr_d[0]));
 b15nand03ah1n06x5 U3760 (.a(u_gpio_gen_filter_29__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_29__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_29__u_filter_diff_ctr_d[0]),
    .o1(n2860));
 b15nor002an1n08x5 U3761 (.a(n2861),
    .b(n2860),
    .o1(eq_x_86_n25));
 b15nand02ar1n02x5 U3762 (.a(u_gpio_gen_filter_1__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_1__u_filter_diff_ctr_q[1]),
    .o1(n2862));
 b15oai012ar1n04x5 U3763 (.a(n2862),
    .b(u_gpio_gen_filter_1__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_1__u_filter_diff_ctr_q[1]),
    .o1(n2863));
 b15oaoi13al1n04x5 U3764 (.a(n2864),
    .b(n2863),
    .c(n2867),
    .d(n2865),
    .o1(u_gpio_gen_filter_1__u_filter_diff_ctr_d[1]));
 b15oaoi13al1n04x5 U3765 (.a(n2864),
    .b(net2180),
    .c(n2867),
    .d(n2865),
    .o1(u_gpio_gen_filter_1__u_filter_diff_ctr_d[0]));
 b15nandp3as1n08x5 U3766 (.a(u_gpio_gen_filter_1__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_1__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_1__u_filter_diff_ctr_d[0]),
    .o1(n2866));
 b15norp02ah1n24x5 U3767 (.a(n2867),
    .b(n2866),
    .o1(eq_x_226_n25));
 b15nand02ar1n02x5 U3768 (.a(u_gpio_gen_filter_9__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_9__u_filter_diff_ctr_q[1]),
    .o1(n2868));
 b15oai012aq1n02x5 U3769 (.a(n2868),
    .b(u_gpio_gen_filter_9__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_9__u_filter_diff_ctr_q[1]),
    .o1(n2869));
 b15oaoi13an1n04x5 U3770 (.a(n2870),
    .b(n2869),
    .c(n2873),
    .d(n2871),
    .o1(u_gpio_gen_filter_9__u_filter_diff_ctr_d[1]));
 b15oaoi13as1n08x5 U3771 (.a(n2870),
    .b(u_gpio_gen_filter_9__u_filter_diff_ctr_q[0]),
    .c(n2873),
    .d(n2871),
    .o1(u_gpio_gen_filter_9__u_filter_diff_ctr_d[0]));
 b15nand03aq1n06x5 U3772 (.a(u_gpio_gen_filter_9__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_9__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_9__u_filter_diff_ctr_d[0]),
    .o1(n2872));
 b15nor002ah1n08x5 U3773 (.a(n2873),
    .b(n2872),
    .o1(eq_x_186_n25));
 b15nand02ar1n02x5 U3774 (.a(u_gpio_gen_filter_31__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_31__u_filter_diff_ctr_q[1]),
    .o1(n2874));
 b15oai012aq1n03x5 U3775 (.a(n2874),
    .b(u_gpio_gen_filter_31__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_31__u_filter_diff_ctr_q[1]),
    .o1(n2875));
 b15oaoi13as1n08x5 U3776 (.a(n2876),
    .b(n2875),
    .c(n2879),
    .d(n2877),
    .o1(u_gpio_gen_filter_31__u_filter_diff_ctr_d[1]));
 b15oaoi13as1n08x5 U3777 (.a(n2876),
    .b(net2135),
    .c(n2879),
    .d(n2877),
    .o1(u_gpio_gen_filter_31__u_filter_diff_ctr_d[0]));
 b15nand03al1n24x5 U3778 (.a(u_gpio_gen_filter_31__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_31__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_31__u_filter_diff_ctr_d[0]),
    .o1(n2878));
 b15norp02ar1n48x5 U3779 (.a(n2879),
    .b(n2878),
    .o1(eq_x_76_n25));
 b15nand02ar1n02x5 U3780 (.a(u_gpio_gen_filter_13__u_filter_diff_ctr_q[0]),
    .b(u_gpio_gen_filter_13__u_filter_diff_ctr_q[1]),
    .o1(n2880));
 b15oai012aq1n03x5 U3781 (.a(n2880),
    .b(u_gpio_gen_filter_13__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_13__u_filter_diff_ctr_q[1]),
    .o1(n2881));
 b15oaoi13ar1n08x5 U3782 (.a(n2882),
    .b(n2881),
    .c(n2885),
    .d(n2883),
    .o1(u_gpio_gen_filter_13__u_filter_diff_ctr_d[1]));
 b15oaoi13ar1n08x5 U3783 (.a(n2882),
    .b(net2085),
    .c(n2885),
    .d(n2883),
    .o1(u_gpio_gen_filter_13__u_filter_diff_ctr_d[0]));
 b15nandp3ar1n04x5 U3784 (.a(u_gpio_gen_filter_13__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_13__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_13__u_filter_diff_ctr_d[0]),
    .o1(n2884));
 b15norp02as1n03x5 U3785 (.a(n2885),
    .b(n2884),
    .o1(eq_x_166_n25));
 b15inv020an1n04x5 U3786 (.a(n2886),
    .o1(n2892));
 b15nand02as1n04x5 U3787 (.a(n2892),
    .b(n2887),
    .o1(n2890));
 b15oai012al1n12x5 U3788 (.a(n2890),
    .b(u_gpio_gen_filter_22__u_filter_diff_ctr_q[0]),
    .c(n2888),
    .o1(u_gpio_gen_filter_22__u_filter_diff_ctr_d[0]));
 b15oai012an1n04x5 U3789 (.a(n2889),
    .b(u_gpio_gen_filter_22__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_22__u_filter_diff_ctr_q[1]),
    .o1(n2891));
 b15aoai13ah1n06x5 U3790 (.a(n2890),
    .b(n2891),
    .c(net2128),
    .d(u_gpio_gen_filter_22__u_filter_diff_ctr_q[0]),
    .o1(u_gpio_gen_filter_22__u_filter_diff_ctr_d[1]));
 b15nand03ah1n12x5 U3791 (.a(n2892),
    .b(u_gpio_gen_filter_22__u_filter_diff_ctr_d[0]),
    .c(u_gpio_gen_filter_22__u_filter_diff_ctr_d[1]),
    .o1(n2893));
 b15norp02al1n32x5 U3792 (.a(n2894),
    .b(n2893),
    .o1(eq_x_121_n25));
 b15inv000aq1n12x5 U3793 (.a(net1789),
    .o1(n3044));
 b15nor002aq1n04x5 U3794 (.a(n3620),
    .b(n3044),
    .o1(net166));
 b15inv000an1n08x5 U3795 (.a(net2222),
    .o1(n2897));
 b15inv000ar1n12x5 U3796 (.a(net1877),
    .o1(n2896));
 b15nandp2ah1n08x5 U3797 (.a(net1784),
    .b(n2896),
    .o1(n2895));
 b15oai012ah1n32x5 U3798 (.a(net1785),
    .b(n2897),
    .c(net1878),
    .o1(n3063));
 b15nanb02aq1n03x5 U3799 (.a(net1790),
    .b(net1786),
    .out0(net117));
 b15nor004an1n04x5 U3800 (.a(net62),
    .b(net59),
    .c(net69),
    .d(net70),
    .o1(n2901));
 b15nor004al1n02x5 U3801 (.a(net58),
    .b(net66),
    .c(net60),
    .d(net65),
    .o1(n2898));
 b15nona23as1n04x5 U3802 (.a(net63),
    .b(net64),
    .c(net67),
    .d(n2898),
    .out0(n2900));
 b15nanb02aq1n04x5 U3803 (.a(net61),
    .b(net68),
    .out0(n2899));
 b15nonb03as1n12x5 U3804 (.a(n2901),
    .b(n2900),
    .c(n2899),
    .out0(n2903));
 b15inv020aq1n10x5 U3805 (.a(net57),
    .o1(n2902));
 b15nand02aq1n48x5 U3806 (.a(n2903),
    .b(n2902),
    .o1(u_xbar_periph_u_s1n_6_dev_select_t[2]));
 b15inv000an1n06x5 U3807 (.a(net55),
    .o1(n2904));
 b15nonb02an1n08x5 U3808 (.a(net55),
    .b(net56),
    .out0(n3610));
 b15aob012an1n24x5 U3809 (.a(u_xbar_periph_u_s1n_6_dev_select_t[2]),
    .b(n2903),
    .c(n3610),
    .out0(n3613));
 b15oai012al1n24x5 U3810 (.a(n3613),
    .b(n2904),
    .c(u_xbar_periph_u_s1n_6_dev_select_t[2]),
    .o1(u_xbar_periph_u_s1n_6_dev_select_t[0]));
 b15inv020an1n04x5 U3811 (.a(net56),
    .o1(n2905));
 b15norp02ar1n08x5 U3812 (.a(u_xbar_periph_u_s1n_6_dev_select_t[2]),
    .b(n2905),
    .o1(u_xbar_periph_u_s1n_6_dev_select_t[1]));
 b15xor002ah1n16x5 U3813 (.a(u_xbar_periph_u_s1n_6_dev_select_t[0]),
    .b(n2906),
    .out0(n2913));
 b15xor002as1n03x5 U3814 (.a(u_xbar_periph_u_s1n_6_dev_select_t[1]),
    .b(net1859),
    .out0(n2908));
 b15qgbxo2an1n05x5 U3815 (.a(u_xbar_periph_u_s1n_6_dev_select_t[2]),
    .b(net2210),
    .out0(n2907));
 b15norp02aq1n16x5 U3816 (.a(n2908),
    .b(n2907),
    .o1(n2912));
 b15nor004as1n12x5 U3817 (.a(u_xbar_periph_u_s1n_6_num_req_outstanding[5]),
    .b(u_xbar_periph_u_s1n_6_num_req_outstanding[4]),
    .c(u_xbar_periph_u_s1n_6_num_req_outstanding[3]),
    .d(u_xbar_periph_u_s1n_6_num_req_outstanding[2]),
    .o1(n2911));
 b15orn003an1n08x5 U3818 (.a(u_xbar_periph_u_s1n_6_num_req_outstanding[8]),
    .b(u_xbar_periph_u_s1n_6_num_req_outstanding[7]),
    .c(u_xbar_periph_u_s1n_6_num_req_outstanding[6]),
    .o(n2909));
 b15norp03as1n24x5 U3819 (.a(n2909),
    .b(u_xbar_periph_u_s1n_6_num_req_outstanding[1]),
    .c(u_xbar_periph_u_s1n_6_num_req_outstanding[0]),
    .o1(n2910));
 b15aoi022as1n48x5 U3820 (.a(n2913),
    .b(n2912),
    .c(n2911),
    .d(n2910),
    .o1(n3616));
 b15nandp2al1n12x5 U3821 (.a(n3610),
    .b(net8),
    .o1(n2982));
 b15nor002aq1n04x5 U3822 (.a(n2982),
    .b(u_xbar_periph_u_s1n_6_tl_u_i[24]),
    .o1(n2914));
 b15nanb02ar1n24x5 U3823 (.a(u_xbar_periph_u_s1n_6_dev_select_t[2]),
    .b(n2914),
    .out0(n2915));
 b15norp02as1n48x5 U3824 (.a(n3616),
    .b(n2915),
    .o1(n3831));
 b15nor002an1n04x5 U3825 (.a(n3831),
    .b(n3045),
    .o1(n1530));
 b15nor002as1n03x5 U3826 (.a(n3831),
    .b(n3044),
    .o1(n1527));
 b15ztpn00an1n08x5 PHY_45 ();
 b15ztpn00an1n08x5 PHY_44 ();
 b15ao0022as1n04x5 U3829 (.a(n3935),
    .b(net2213),
    .c(n3934),
    .d(net1762),
    .o(net160));
 b15ao0022ar1n06x5 U3830 (.a(n3935),
    .b(u_xbar_periph_u_s1n_6_tl_u_i[12]),
    .c(n3934),
    .d(net1832),
    .o(net155));
 b15ao0022ar1n06x5 U3831 (.a(n3935),
    .b(u_xbar_periph_u_s1n_6_tl_u_i[14]),
    .c(n3934),
    .d(net1835),
    .o(net157));
 b15ao0022an1n06x5 U3832 (.a(n3935),
    .b(net1799),
    .c(n3934),
    .d(u_xbar_periph_u_s1n_6_tl_u_i[4]),
    .o(net158));
 b15ao0022an1n06x5 U3833 (.a(n3935),
    .b(u_xbar_periph_u_s1n_6_tl_u_i[18]),
    .c(n3934),
    .d(net1810),
    .o(net161));
 b15ao0022ar1n06x5 U3834 (.a(n3935),
    .b(u_xbar_periph_u_s1n_6_tl_u_i[11]),
    .c(n3934),
    .d(net1844),
    .o(net153));
 b15ao0022al1n06x5 U3835 (.a(n3935),
    .b(u_xbar_periph_u_s1n_6_tl_u_i[13]),
    .c(n3934),
    .d(net1816),
    .o(net156));
 b15ao0022aq1n06x5 U3836 (.a(n3935),
    .b(net1813),
    .c(n3934),
    .d(u_xbar_periph_u_s1n_6_tl_u_i[5]),
    .o(net159));
 b15aoi022as1n08x5 U3837 (.a(net1770),
    .b(u_xbar_periph_u_s1n_6_tl_u_i[10]),
    .c(n2923),
    .d(n3044),
    .o1(n2916));
 b15xor002an1n12x5 U3838 (.a(u_xbar_periph_u_s1n_6_tl_u_i[20]),
    .b(net1771),
    .out0(n2917));
 b15xor002al1n16x5 U3839 (.a(net1772),
    .b(net1766),
    .out0(n2941));
 b15aoi012an1n02x5 U3840 (.a(n3620),
    .b(net1773),
    .c(n2922),
    .o1(n2921));
 b15norp03as1n24x5 U3841 (.a(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_opcode[0]),
    .b(net1805),
    .c(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_opcode[1]),
    .o1(n3049));
 b15aboi22aq1n06x5 U3842 (.a(net1780),
    .b(net1795),
    .c(net1780),
    .d(net1796),
    .out0(n2919));
 b15xor002ah1n04x5 U3843 (.a(net1806),
    .b(n2919),
    .out0(n2943));
 b15norp02aq1n02x5 U3844 (.a(n3617),
    .b(n2943),
    .o1(n2920));
 b15oaoi13al1n04x5 U3845 (.a(n2920),
    .b(n2921),
    .c(net1773),
    .d(n2922),
    .o1(net172));
 b15oai122aq1n16x5 U3846 (.a(n3935),
    .b(net1822),
    .c(n2923),
    .d(net1823),
    .e(net1849),
    .o1(net113));
 b15inv000al1n06x5 U3847 (.a(n3831),
    .o1(n3638));
 b15aob012as1n03x5 U3848 (.a(n3638),
    .b(u_xbar_periph_u_s1n_6_tl_u_i[24]),
    .c(net2),
    .out0(u_gpio_u_reg_u_reg_if_N7));
 b15nor002as1n08x5 U3849 (.a(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_rsp_pending),
    .b(net1758),
    .o1(n3618));
 b15qgbno2an1n10x5 U3850 (.a(net1759),
    .b(net2),
    .o1(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_N12));
 b15nor002an1n08x5 U3851 (.a(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_N12),
    .b(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_rsp_pending),
    .o1(n3614));
 b15nano23as1n24x5 U3852 (.a(net8),
    .b(n3614),
    .c(n3616),
    .d(n3613),
    .out0(n3829));
 b15oai012an1n04x5 U3853 (.a(n2924),
    .b(u_gpio_gen_filter_5__u_filter_diff_ctr_q[0]),
    .c(u_gpio_gen_filter_5__u_filter_diff_ctr_q[1]),
    .o1(n2926));
 b15nandp2aq1n04x5 U3854 (.a(n2929),
    .b(n2925),
    .o1(n2927));
 b15aoai13al1n08x5 U3855 (.a(n2927),
    .b(n2926),
    .c(u_gpio_gen_filter_5__u_filter_diff_ctr_q[1]),
    .d(u_gpio_gen_filter_5__u_filter_diff_ctr_q[0]),
    .o1(u_gpio_gen_filter_5__u_filter_diff_ctr_d[1]));
 b15oai012aq1n06x5 U3856 (.a(n2927),
    .b(u_gpio_gen_filter_5__u_filter_diff_ctr_q[0]),
    .c(n2928),
    .o1(u_gpio_gen_filter_5__u_filter_diff_ctr_d[0]));
 b15and003ar1n03x5 U3857 (.a(n2929),
    .b(u_gpio_gen_filter_5__u_filter_diff_ctr_d[1]),
    .c(u_gpio_gen_filter_5__u_filter_diff_ctr_d[0]),
    .o(eq_x_206_n25));
 b15inv000ar1n06x5 U3858 (.a(net1880),
    .o1(n3051));
 b15inv000ah1n04x5 U3859 (.a(net1884),
    .o1(n3073));
 b15aoi022aq1n06x5 U3860 (.a(net1884),
    .b(net1880),
    .c(n3051),
    .d(n3073),
    .o1(n2931));
 b15inv040ah1n05x5 U3861 (.a(net1887),
    .o1(n3074));
 b15inv040as1n06x5 U3862 (.a(net1904),
    .o1(n3092));
 b15aoi022an1n16x5 U3863 (.a(gpio_2_xbar[26]),
    .b(n3074),
    .c(net1869),
    .d(n3092),
    .o1(n2930));
 b15xor002as1n06x5 U3864 (.a(n2931),
    .b(net1870),
    .out0(n2953));
 b15inv040as1n05x5 U3865 (.a(net1792),
    .o1(n3105));
 b15inv020as1n06x5 U3866 (.a(net1820),
    .o1(n3079));
 b15aoi022ar1n12x5 U3867 (.a(net1820),
    .b(net1793),
    .c(net1792),
    .d(n3079),
    .o1(n2936));
 b15qgbin1an1n05x5 U3868 (.a(net1828),
    .o1(n3089));
 b15inv020ah1n05x5 U3869 (.a(net1925),
    .o1(n3075));
 b15aoi022as1n12x5 U3870 (.a(gpio_2_xbar[21]),
    .b(net1828),
    .c(net1829),
    .d(n3075),
    .o1(n2958));
 b15inv020ah1n10x5 U3871 (.a(net1908),
    .o1(n3091));
 b15inv020as1n10x5 U3872 (.a(net1888),
    .o1(n3076));
 b15aoi022ar1n24x5 U3873 (.a(gpio_2_xbar[20]),
    .b(gpio_2_xbar[27]),
    .c(n3091),
    .d(n3076),
    .o1(n2932));
 b15xor002aq1n04x5 U3874 (.a(n2958),
    .b(n2932),
    .out0(n2934));
 b15inv040as1n05x5 U3875 (.a(net1842),
    .o1(n3067));
 b15inv000ar1n16x5 U3876 (.a(gpio_2_xbar[25]),
    .o1(n3093));
 b15aoi022aq1n16x5 U3877 (.a(gpio_2_xbar[25]),
    .b(net1842),
    .c(n3067),
    .d(n3093),
    .o1(n3055));
 b15inv000an1n05x5 U3878 (.a(net1840),
    .o1(n3082));
 b15inv000as1n06x5 U3879 (.a(net1847),
    .o1(n3085));
 b15aoi022an1n12x5 U3880 (.a(net1847),
    .b(net1840),
    .c(n3082),
    .d(net1848),
    .o1(n3053));
 b15xor002as1n02x5 U3881 (.a(n3055),
    .b(n3053),
    .out0(n2933));
 b15xor002as1n04x5 U3882 (.a(n2934),
    .b(n2933),
    .out0(n2935));
 b15xor002ah1n03x5 U3883 (.a(n2936),
    .b(n2935),
    .out0(n2938));
 b15aoi012ar1n02x5 U3884 (.a(net1860),
    .b(net1871),
    .c(n2938),
    .o1(n2937));
 b15oai012ah1n04x5 U3885 (.a(n2937),
    .b(net1871),
    .c(n2938),
    .o1(net144));
 b15inv000al1n02x5 U3886 (.a(net1773),
    .o1(n2939));
 b15aoi122ar1n04x5 U3887 (.a(n3620),
    .b(u_xbar_periph_u_s1n_6_tl_u_i[19]),
    .c(net1773),
    .d(n2940),
    .e(n2939),
    .o1(n2942));
 b15aoi012ah1n02x5 U3888 (.a(n2942),
    .b(n3934),
    .c(net1807),
    .o1(net112));
 b15nandp2ar1n02x5 U3889 (.a(n3935),
    .b(net1766),
    .o1(n2944));
 b15aob012al1n06x5 U3890 (.a(net1767),
    .b(net1806),
    .c(n3934),
    .out0(net165));
 b15inv040al1n02x5 U3891 (.a(net1768),
    .o1(net116));
 b15inv000al1n10x5 U3892 (.a(net1901),
    .o1(n3072));
 b15aoi022aq1n16x5 U3893 (.a(net1901),
    .b(net1908),
    .c(n3091),
    .d(n3072),
    .o1(n3014));
 b15inv040an1n08x5 U3894 (.a(net1857),
    .o1(n3083));
 b15inv040aq1n08x5 U3895 (.a(net1863),
    .o1(n3095));
 b15aoi022al1n04x5 U3896 (.a(net1863),
    .b(net1857),
    .c(n3083),
    .d(net1864),
    .o1(n2946));
 b15inv020as1n10x5 U3897 (.a(net1899),
    .o1(n3078));
 b15inv040as1n12x5 U3898 (.a(net1830),
    .o1(n3087));
 b15aoi022ar1n04x5 U3899 (.a(net1830),
    .b(n3078),
    .c(net1899),
    .d(n3087),
    .o1(n2945));
 b15xor002aq1n03x5 U3900 (.a(n2946),
    .b(n2945),
    .out0(n2948));
 b15inv040ah1n08x5 U3901 (.a(net1873),
    .o1(n3088));
 b15inv000aq1n12x5 U3902 (.a(net1911),
    .o1(n3084));
 b15aoi022as1n08x5 U3903 (.a(net1911),
    .b(net1873),
    .c(n3088),
    .d(net1912),
    .o1(n2947));
 b15xor002as1n03x5 U3904 (.a(n2948),
    .b(n2947),
    .out0(n2949));
 b15xor002as1n06x5 U3905 (.a(n3014),
    .b(net1929),
    .out0(n2950));
 b15inv000ah1n10x5 U3906 (.a(net1854),
    .o1(n3098));
 b15inv000aq1n12x5 U3907 (.a(net1893),
    .o1(n3068));
 b15aoi022al1n32x5 U3908 (.a(net1893),
    .b(net1854),
    .c(net1855),
    .d(net1894),
    .o1(n3060));
 b15xor002an1n08x5 U3909 (.a(n2950),
    .b(net1922),
    .out0(n2952));
 b15aoi012ar1n02x5 U3910 (.a(net1860),
    .b(net1871),
    .c(n2952),
    .o1(n2951));
 b15oai012ah1n04x5 U3911 (.a(n2951),
    .b(net1871),
    .c(n2952),
    .o1(net170));
 b15inv040aq1n04x5 U3912 (.a(net1802),
    .o1(n3086));
 b15aoi022as1n08x5 U3913 (.a(net1820),
    .b(net1802),
    .c(net1803),
    .d(n3079),
    .o1(n2955));
 b15inv040as1n05x5 U3914 (.a(net1826),
    .o1(n3096));
 b15aoi022an1n16x5 U3915 (.a(net1830),
    .b(net1826),
    .c(net1827),
    .d(net1831),
    .o1(n2954));
 b15xor002an1n16x5 U3916 (.a(n2955),
    .b(n2954),
    .out0(n3012));
 b15inv000aq1n12x5 U3917 (.a(net1902),
    .o1(n3090));
 b15aoi022ah1n24x5 U3918 (.a(net1902),
    .b(net1857),
    .c(n3083),
    .d(n3090),
    .o1(n3019));
 b15aoi022an1n12x5 U3919 (.a(net1863),
    .b(net1842),
    .c(n3067),
    .d(n3095),
    .o1(n2957));
 b15inv020ah1n12x5 U3920 (.a(net1913),
    .o1(n3100));
 b15aoi022an1n12x5 U3921 (.a(gpio_2_xbar[10]),
    .b(gpio_2_xbar[6]),
    .c(n3051),
    .d(n3100),
    .o1(n2956));
 b15qgbxo2an1n10x5 U3922 (.a(n2957),
    .b(n2956),
    .out0(n2959));
 b15xor002al1n08x5 U3923 (.a(n2959),
    .b(n2958),
    .out0(n2960));
 b15xor002al1n08x5 U3924 (.a(n3019),
    .b(n2960),
    .out0(n2961));
 b15inv040ar1n10x5 U3925 (.a(net1852),
    .o1(n3080));
 b15aoi022al1n24x5 U3926 (.a(net1852),
    .b(net1873),
    .c(n3088),
    .d(net1853),
    .o1(n3059));
 b15xor002as1n06x5 U3927 (.a(n2961),
    .b(net1874),
    .out0(n2963));
 b15aoi012ah1n02x5 U3928 (.a(net1860),
    .b(n3012),
    .c(net1875),
    .o1(n2962));
 b15oai012ar1n12x5 U3929 (.a(n2962),
    .b(n3012),
    .c(net1875),
    .o1(net164));
 b15inv040ah1n08x5 U3930 (.a(net7),
    .o1(n1451));
 b15inv000ar1n06x5 U3931 (.a(net9),
    .o1(n1443));
 b15nor002an1n24x5 U3932 (.a(net53),
    .b(net54),
    .o1(n3257));
 b15nandp3as1n24x5 U3933 (.a(n3257),
    .b(net52),
    .c(net51),
    .o1(n3042));
 b15inv000ar1n06x5 U3934 (.a(net45),
    .o1(n2964));
 b15norp02al1n03x5 U3935 (.a(n3042),
    .b(n2964),
    .o1(n2991));
 b15nand04aq1n08x5 U3936 (.a(net48),
    .b(net47),
    .c(net45),
    .d(net46),
    .o1(n2973));
 b15inv000aq1n04x5 U3937 (.a(n2973),
    .o1(n2990));
 b15inv000al1n02x5 U3938 (.a(net10),
    .o1(n2970));
 b15oai013ah1n03x5 U3939 (.a(net4),
    .b(net49),
    .c(net3),
    .d(net50),
    .o1(n2969));
 b15inv020aq1n03x5 U3940 (.a(net49),
    .o1(n2971));
 b15nonb03ah1n03x5 U3941 (.a(net50),
    .b(net45),
    .c(net46),
    .out0(n2979));
 b15aob012al1n02x5 U3942 (.a(n2979),
    .b(n2971),
    .c(net48),
    .out0(n2967));
 b15nor003as1n03x5 U3943 (.a(net48),
    .b(net47),
    .c(net50),
    .o1(n2978));
 b15aoi022al1n02x5 U3944 (.a(net49),
    .b(net45),
    .c(net46),
    .d(n2971),
    .o1(n2965));
 b15aoi112al1n02x5 U3945 (.a(net4),
    .b(net3),
    .c(n2978),
    .d(n2965),
    .o1(n2966));
 b15aoai13ah1n03x5 U3946 (.a(n2966),
    .b(n2967),
    .c(net49),
    .d(net47),
    .o1(n2968));
 b15oai112al1n08x5 U3947 (.a(n2969),
    .b(n2968),
    .c(net11),
    .d(n2970),
    .o1(n2989));
 b15inv000al1n02x5 U3948 (.a(net3),
    .o1(n2972));
 b15aoi112ah1n02x5 U3949 (.a(net48),
    .b(net46),
    .c(n2972),
    .d(n2971),
    .o1(n2975));
 b15nor003as1n02x5 U3950 (.a(net47),
    .b(net45),
    .c(net49),
    .o1(n2974));
 b15oai013an1n06x5 U3951 (.a(n2973),
    .b(net4),
    .c(n2975),
    .d(n2974),
    .o1(n2977));
 b15norp02ar1n02x5 U3952 (.a(net5),
    .b(n1451),
    .o1(n2976));
 b15oaoi13an1n03x5 U3953 (.a(n2976),
    .b(n1451),
    .c(net5),
    .d(n2977),
    .o1(n2988));
 b15norp02ar1n03x5 U3954 (.a(n2979),
    .b(n2978),
    .o1(n2980));
 b15oaoi13an1n02x5 U3955 (.a(net6),
    .b(net3),
    .c(net49),
    .d(n2980),
    .o1(n2986));
 b15aoi012ar1n02x5 U3956 (.a(net12),
    .b(net7),
    .c(net10),
    .o1(n2983));
 b15aoi022an1n02x5 U3957 (.a(net9),
    .b(net11),
    .c(net12),
    .d(n1443),
    .o1(n2981));
 b15nona22ar1n02x5 U3958 (.a(n2983),
    .b(n2982),
    .c(n2981),
    .out0(n2984));
 b15norp02ar1n02x5 U3959 (.a(u_xbar_periph_u_s1n_6_dev_select_t[2]),
    .b(n2984),
    .o1(n2985));
 b15nandp2ar1n03x5 U3960 (.a(n2986),
    .b(n2985),
    .o1(n2987));
 b15ornc04an1n16x5 U3961 (.a(n3616),
    .b(n2989),
    .c(n2988),
    .d(n2987),
    .o(n2992));
 b15oab012al1n04x5 U3962 (.a(n2992),
    .b(n2991),
    .c(n2990),
    .out0(n3026));
 b15nand02aq1n12x5 U3963 (.a(n3831),
    .b(n1451),
    .o1(n3025));
 b15nonb02ah1n08x5 U3964 (.a(n3025),
    .b(n2992),
    .out0(n3134));
 b15norp02ar1n03x5 U3965 (.a(n3026),
    .b(n3134),
    .o1(u_gpio_u_reg_u_reg_if_N46));
 b15aoi022ah1n08x5 U3966 (.a(net2210),
    .b(net1780),
    .c(n3935),
    .d(u_xbar_periph_u_s1n_6_tl_u_i[20]),
    .o1(n2993));
 b15nandp2ah1n02x5 U3967 (.a(net1781),
    .b(n3063),
    .o1(net115));
 b15nonb02aq1n02x5 U3968 (.a(net1786),
    .b(net1781),
    .out0(net163));
 b15inv000ah1n08x5 U3969 (.a(net1882),
    .o1(n3070));
 b15aoi022ah1n16x5 U3970 (.a(net1882),
    .b(net1888),
    .c(n3076),
    .d(n3070),
    .o1(n3016));
 b15aoi022aq1n12x5 U3971 (.a(net1852),
    .b(net1847),
    .c(n3085),
    .d(n3080),
    .o1(n2995));
 b15aoi022ah1n08x5 U3972 (.a(net1893),
    .b(net1863),
    .c(n3095),
    .d(n3068),
    .o1(n2994));
 b15qgbxo2an1n10x5 U3973 (.a(n2995),
    .b(n2994),
    .out0(n2999));
 b15aoi022ah1n06x5 U3974 (.a(net1902),
    .b(net1869),
    .c(n3074),
    .d(n3090),
    .o1(n2997));
 b15inv020ah1n12x5 U3975 (.a(net1897),
    .o1(n3102));
 b15aoi022an1n08x5 U3976 (.a(net1899),
    .b(net1897),
    .c(n3102),
    .d(n3078),
    .o1(n2996));
 b15xor002as1n06x5 U3977 (.a(n2997),
    .b(n2996),
    .out0(n2998));
 b15xor002an1n12x5 U3978 (.a(n2999),
    .b(n2998),
    .out0(n3000));
 b15xor002an1n16x5 U3979 (.a(n3016),
    .b(n3000),
    .out0(n3001));
 b15inv040as1n06x5 U3980 (.a(net1838),
    .o1(n3069));
 b15aoi022al1n16x5 U3981 (.a(net1838),
    .b(net1792),
    .c(net1793),
    .d(net1839),
    .o1(n3009));
 b15xor002an1n06x5 U3982 (.a(n3001),
    .b(n3009),
    .out0(n3004));
 b15aoi022ah1n04x5 U3983 (.a(net1802),
    .b(net1925),
    .c(n3075),
    .d(net1803),
    .o1(n3003));
 b15oai012ar1n03x5 U3984 (.a(n3935),
    .b(net1926),
    .c(n3004),
    .o1(n3002));
 b15aoai13aq1n04x5 U3985 (.a(net1786),
    .b(n3002),
    .c(n3004),
    .d(net1926),
    .o1(net154));
 b15aoi022al1n16x5 U3986 (.a(gpio_2_xbar[2]),
    .b(gpio_2_xbar[26]),
    .c(n3092),
    .d(n3072),
    .o1(n3008));
 b15aoi022ah1n16x5 U3987 (.a(net1897),
    .b(net1913),
    .c(n3100),
    .d(net1898),
    .o1(n3020));
 b15inv040an1n10x5 U3988 (.a(net1906),
    .o1(n3099));
 b15aoi022as1n16x5 U3989 (.a(net1906),
    .b(net1911),
    .c(net1912),
    .d(n3099),
    .o1(n3056));
 b15xor002as1n12x5 U3990 (.a(n3020),
    .b(n3056),
    .out0(n3006));
 b15aoi022al1n16x5 U3991 (.a(net2217),
    .b(gpio_2_xbar[25]),
    .c(n3093),
    .d(n3078),
    .o1(n3005));
 b15xor002ah1n12x5 U3992 (.a(n3006),
    .b(n3005),
    .out0(n3007));
 b15xor002ah1n16x5 U3993 (.a(n3008),
    .b(n3007),
    .out0(n3010));
 b15xor002ah1n04x5 U3994 (.a(n3010),
    .b(n3009),
    .out0(n3013));
 b15oai012ah1n03x5 U3995 (.a(n3935),
    .b(n3012),
    .c(n3013),
    .o1(n3011));
 b15aoai13al1n08x5 U3996 (.a(net1786),
    .b(n3011),
    .c(n3013),
    .d(n3012),
    .o1(net133));
 b15aoi022aq1n06x5 U3997 (.a(net1906),
    .b(net1854),
    .c(net1855),
    .d(n3099),
    .o1(n3015));
 b15xor002aq1n08x5 U3998 (.a(n3015),
    .b(n3014),
    .out0(n3017));
 b15xor002an1n12x5 U3999 (.a(n3017),
    .b(n3016),
    .out0(n3018));
 b15xor002ar1n08x5 U4000 (.a(n3019),
    .b(n3018),
    .out0(n3021));
 b15xor002aq1n08x5 U4001 (.a(n3021),
    .b(n3020),
    .out0(n3024));
 b15aoi022an1n06x5 U4002 (.a(net1840),
    .b(net1828),
    .c(net1829),
    .d(net1841),
    .o1(n3023));
 b15oai012al1n02x5 U4003 (.a(n3935),
    .b(net1919),
    .c(n3024),
    .o1(n3022));
 b15aoai13an1n04x5 U4004 (.a(net1786),
    .b(n3022),
    .c(n3024),
    .d(net1919),
    .o1(net171));
 b15nonb02as1n16x5 U4005 (.a(n3026),
    .b(n3025),
    .out0(n3256));
 b15inv000as1n48x5 U4006 (.a(net51),
    .o1(n3247));
 b15nandp2aq1n32x5 U4007 (.a(net53),
    .b(net54),
    .o1(n3529));
 b15norp03as1n24x5 U4008 (.a(n3247),
    .b(n3529),
    .c(net52),
    .o1(n3027));
 b15ztpn00an1n08x5 PHY_43 ();
 b15ztpn00an1n08x5 PHY_42 ();
 b15nand02ar1n24x5 U4011 (.a(n3256),
    .b(net433),
    .o1(n3028));
 b15ztpn00an1n08x5 PHY_41 ();
 b15ztpn00an1n08x5 PHY_40 ();
 b15inv000al1n20x5 U4014 (.a(net52),
    .o1(n3120));
 b15norp03an1n24x5 U4015 (.a(n3120),
    .b(n3247),
    .c(n3529),
    .o1(n3029));
 b15ztpn00an1n08x5 PHY_39 ();
 b15ztpn00an1n08x5 PHY_38 ();
 b15nandp2as1n24x5 U4018 (.a(net227),
    .b(net425),
    .o1(n3030));
 b15ztpn00an1n08x5 PHY_37 ();
 b15inv020as1n10x5 U4021 (.a(net54),
    .o1(n3131));
 b15nor002as1n16x5 U4022 (.a(net53),
    .b(n3131),
    .o1(n3246));
 b15inv020ah1n16x5 U4023 (.a(n3246),
    .o1(n3640));
 b15norp03aq1n24x5 U4024 (.a(n3120),
    .b(n3247),
    .c(n3640),
    .o1(n3031));
 b15ztpn00an1n08x5 PHY_36 ();
 b15ztpn00an1n08x5 PHY_35 ();
 b15nandp2aq1n32x5 U4027 (.a(net227),
    .b(net256),
    .o1(n3032));
 b15ztpn00an1n08x5 PHY_34 ();
 b15ztpn00an1n08x5 PHY_33 ();
 b15nandp2ah1n16x5 U4030 (.a(n3120),
    .b(n3247),
    .o1(n3137));
 b15norp02aq1n24x5 U4031 (.a(n3137),
    .b(n3529),
    .o1(n3033));
 b15ztpn00an1n08x5 PHY_32 ();
 b15ztpn00an1n08x5 PHY_31 ();
 b15nand02ah1n48x5 U4034 (.a(net227),
    .b(net278),
    .o1(n3034));
 b15ztpn00an1n08x5 PHY_30 ();
 b15ztpn00an1n08x5 PHY_29 ();
 b15nanb02an1n12x5 U4037 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[1]),
    .b(n3039),
    .out0(n3037));
 b15inv000ar1n06x5 U4038 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .o1(n3036));
 b15qgbna2an1n05x5 U4039 (.o1(n3035),
    .a(n3037),
    .b(net2084));
 b15oai012ar1n24x5 U4040 (.a(n3035),
    .b(n3037),
    .c(n3036),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_ack_level));
 b15nand02al1n12x5 U4041 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[0]),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[1]),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39));
 b15nonb03aq1n12x5 U4042 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39),
    .b(n3039),
    .c(n3038),
    .out0(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[1]));
 b15nand02an1n08x5 U4043 (.a(net2194),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39));
 b15nonb03al1n12x5 U4044 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39),
    .b(n3040),
    .c(n3217),
    .out0(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[1]));
 b15nor002ah1n06x5 U4045 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .o1(n3222));
 b15inv020aq1n08x5 U4046 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .o1(n3250));
 b15inv000al1n10x5 U4047 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .o1(n3808));
 b15nand02al1n02x5 U4048 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .b(n3808),
    .o1(n3225));
 b15nor002aq1n04x5 U4049 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[1]),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[1]),
    .o1(n3220));
 b15inv020as1n10x5 U4050 (.a(n3220),
    .o1(n3809));
 b15oaoi13ar1n03x5 U4051 (.a(n3809),
    .b(n3225),
    .c(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .d(n3808),
    .o1(n3041));
 b15oai012al1n06x5 U4052 (.a(n3041),
    .b(n3250),
    .c(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .o1(n3333));
 b15aoi012as1n04x5 U4053 (.a(n3333),
    .b(n3250),
    .c(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .o1(n3106));
 b15inv040as1n04x5 U4054 (.a(n3042),
    .o1(n3043));
 b15aoi013as1n08x5 U4055 (.a(net453),
    .b(net227),
    .c(n3043),
    .d(net13),
    .o1(n3213));
 b15aoi012ar1n02x5 U4056 (.a(n3213),
    .b(n3222),
    .c(n3106),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_test_set_d));
 b15nand04as1n16x5 U4057 (.a(n3935),
    .b(net1766),
    .c(net1823),
    .d(n3044),
    .o1(n3046));
 b15ztpn00an1n08x5 PHY_28 ();
 b15ztpn00an1n08x5 PHY_27 ();
 b15nand04as1n16x5 U4060 (.a(net1776),
    .b(n1438),
    .c(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type[1]),
    .d(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type[2]),
    .o1(n3047));
 b15nandp3aq1n24x5 U4061 (.a(net1806),
    .b(n3934),
    .c(net1777),
    .o1(n3050));
 b15ztpn00an1n08x5 PHY_26 ();
 b15ztpn00an1n08x5 PHY_25 ();
 b15oai012an1n04x5 U4064 (.a(net249),
    .b(net228),
    .c(net1881),
    .o1(net125));
 b15aoi022ah1n12x5 U4065 (.a(gpio_2_xbar[1]),
    .b(net1884),
    .c(n3073),
    .d(n3070),
    .o1(n3052));
 b15xor002as1n03x5 U4066 (.a(n3053),
    .b(n3052),
    .out0(n3054));
 b15xor002ar1n08x5 U4067 (.a(n3055),
    .b(n3054),
    .out0(n3057));
 b15qgbxo2an1n05x5 U4068 (.a(n3057),
    .b(n3056),
    .out0(n3058));
 b15xor002ar1n06x5 U4069 (.a(net1874),
    .b(n3058),
    .out0(n3061));
 b15xor002ah1n04x5 U4070 (.a(n3061),
    .b(net1922),
    .out0(n3066));
 b15aoi022ar1n12x5 U4071 (.a(net1826),
    .b(net1838),
    .c(net1839),
    .d(net1827),
    .o1(n3065));
 b15oai012an1n04x5 U4072 (.a(n3935),
    .b(n3065),
    .c(net1923),
    .o1(n3064));
 b15aoai13aq1n08x5 U4073 (.a(net1786),
    .b(n3064),
    .c(net1923),
    .d(n3065),
    .o1(net169));
 b15oai012as1n02x5 U4074 (.a(net250),
    .b(net1843),
    .c(net229),
    .o1(net123));
 b15oai012aq1n03x5 U4075 (.a(net249),
    .b(net1894),
    .c(net228),
    .o1(net121));
 b15oai012ar1n08x5 U4076 (.a(net250),
    .b(net1839),
    .c(net229),
    .o1(net124));
 b15oai012aq1n03x5 U4077 (.a(net249),
    .b(net1883),
    .c(net228),
    .o1(net119));
 b15oai012aq1n03x5 U4078 (.a(net249),
    .b(n3072),
    .c(net228),
    .o1(net120));
 b15ztpn00an1n08x5 PHY_24 ();
 b15ztpn00an1n08x5 PHY_23 ();
 b15oai012an1n03x5 U4081 (.a(net249),
    .b(net1885),
    .c(net228),
    .o1(net143));
 b15oai012as1n02x5 U4082 (.a(net249),
    .b(n3074),
    .c(net228),
    .o1(net139));
 b15oai012aq1n04x5 U4083 (.a(net250),
    .b(n3075),
    .c(net229),
    .o1(net141));
 b15oai012an1n04x5 U4084 (.a(net249),
    .b(net1889),
    .c(net228),
    .o1(net140));
 b15ztpn00an1n08x5 PHY_22 ();
 b15oai012aq1n03x5 U4086 (.a(net249),
    .b(net1900),
    .c(net228),
    .o1(net138));
 b15oai012al1n06x5 U4087 (.a(net250),
    .b(n3079),
    .c(net229),
    .o1(net137));
 b15oai012an1n04x5 U4088 (.a(net250),
    .b(net1853),
    .c(net229),
    .o1(net136));
 b15ztpn00an1n08x5 PHY_21 ();
 b15oai012aq1n03x5 U4090 (.a(net250),
    .b(net1841),
    .c(net229),
    .o1(net152));
 b15oai012an1n03x5 U4091 (.a(net250),
    .b(net1858),
    .c(net229),
    .o1(net134));
 b15oai012ar1n08x5 U4092 (.a(net249),
    .b(net1912),
    .c(net228),
    .o1(net132));
 b15oai012an1n04x5 U4093 (.a(net250),
    .b(net1848),
    .c(net229),
    .o1(net151));
 b15oai012ah1n03x5 U4094 (.a(net250),
    .b(net1803),
    .c(net229),
    .o1(net130));
 b15oai012as1n02x5 U4095 (.a(net250),
    .b(net1831),
    .c(net229),
    .o1(net150));
 b15oai012ar1n12x5 U4096 (.a(net249),
    .b(n3088),
    .c(net228),
    .o1(net128));
 b15oai012an1n04x5 U4097 (.a(net250),
    .b(net1829),
    .c(net229),
    .o1(net149));
 b15oai012al1n04x5 U4098 (.a(net249),
    .b(net1903),
    .c(net228),
    .o1(net126));
 b15oai012al1n04x5 U4099 (.a(net249),
    .b(net1909),
    .c(net228),
    .o1(net148));
 b15oai012al1n04x5 U4100 (.a(net249),
    .b(net1905),
    .c(net228),
    .o1(net147));
 b15oai012an1n03x5 U4101 (.a(net1778),
    .b(n3093),
    .c(n3046),
    .o1(net146));
 b15oai012al1n04x5 U4102 (.a(net250),
    .b(net1864),
    .c(net229),
    .o1(net145));
 b15oai012al1n06x5 U4103 (.a(net250),
    .b(net1827),
    .c(net229),
    .o1(net118));
 b15oai012aq1n03x5 U4104 (.a(net250),
    .b(net1855),
    .c(net229),
    .o1(net142));
 b15oai012al1n08x5 U4105 (.a(net249),
    .b(net1907),
    .c(net228),
    .o1(net131));
 b15oai012ar1n08x5 U4106 (.a(net249),
    .b(net1914),
    .c(net228),
    .o1(net129));
 b15oai012aq1n04x5 U4107 (.a(net249),
    .b(net1898),
    .c(net228),
    .o1(net127));
 b15oai012as1n04x5 U4108 (.a(net250),
    .b(net1793),
    .c(net229),
    .o1(net135));
 b15inv000al1n02x5 U4109 (.a(n3106),
    .o1(n3107));
 b15oai013al1n08x5 U4110 (.a(n3107),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .c(n3808),
    .d(n3809),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_d[2]));
 b15ztpn00an1n08x5 PHY_20 ();
 b15ztpn00an1n08x5 PHY_19 ();
 b15norp02an1n04x5 U4114 (.a(net485),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[28]));
 b15ztpn00an1n08x5 PHY_18 ();
 b15nor002aq1n03x5 U4116 (.a(n3901),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[26]));
 b15ztpn00an1n08x5 PHY_17 ();
 b15nor002al1n04x5 U4120 (.a(n3902),
    .b(n3030),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[27]));
 b15norp02as1n03x5 U4122 (.a(n3899),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[24]));
 b15nor002ah1n03x5 U4123 (.a(n3902),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[27]));
 b15ztpn00an1n08x5 PHY_16 ();
 b15norp02aq1n04x5 U4126 (.a(n3899),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[24]));
 b15norp02aq1n04x5 U4127 (.a(net485),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[28]));
 b15ztpn00an1n08x5 PHY_15 ();
 b15norp02al1n04x5 U4131 (.a(net478),
    .b(net221),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[31]));
 b15norp02an1n04x5 U4132 (.a(net485),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[28]));
 b15nor002ah1n04x5 U4133 (.a(n3902),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[27]));
 b15nor002as1n03x5 U4135 (.a(n3900),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[25]));
 b15norp02al1n04x5 U4137 (.a(net481),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[30]));
 b15nor002an1n03x5 U4138 (.a(n3902),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[27]));
 b15nor002al1n04x5 U4139 (.a(net478),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[31]));
 b15ztpn00an1n08x5 PHY_14 ();
 b15nor002al1n04x5 U4141 (.a(n3904),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[29]));
 b15norp02as1n03x5 U4142 (.a(net478),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[31]));
 b15nor002aq1n02x5 U4143 (.a(n3901),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[26]));
 b15norp02as1n03x5 U4144 (.a(n3904),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[29]));
 b15norp02aq1n04x5 U4145 (.a(n3900),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[25]));
 b15nor002an1n03x5 U4146 (.a(n3901),
    .b(net218),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[26]));
 b15norp02al1n03x5 U4147 (.a(net479),
    .b(n3030),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[31]));
 b15norp02an1n04x5 U4148 (.a(net481),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[30]));
 b15norp02as1n03x5 U4149 (.a(n3900),
    .b(net218),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[25]));
 b15nor002ar1n04x5 U4150 (.a(net481),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[30]));
 b15norp02an1n03x5 U4151 (.a(n3904),
    .b(net218),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[29]));
 b15nor002ar1n04x5 U4152 (.a(n3900),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[25]));
 b15nor002ar1n06x5 U4153 (.a(net484),
    .b(net218),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[28]));
 b15norp02as1n03x5 U4154 (.a(n3901),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[26]));
 b15norp02aq1n03x5 U4155 (.a(net483),
    .b(net218),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[30]));
 b15nor002ah1n03x5 U4156 (.a(n3904),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[29]));
 b15nor002aq1n06x5 U4157 (.a(n3899),
    .b(net218),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[24]));
 b15nor002as1n03x5 U4158 (.a(n3899),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[24]));
 b15inv020an1n64x5 U4159 (.a(net20),
    .o1(n3540));
 b15ztpn00an1n08x5 PHY_13 ();
 b15nor002aq1n03x5 U4161 (.a(n3540),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[7]));
 b15ztpn00an1n08x5 PHY_12 ();
 b15norp02as1n04x5 U4163 (.a(n3540),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[7]));
 b15ztpn00an1n08x5 PHY_11 ();
 b15nor002aq1n06x5 U4165 (.a(n3540),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[7]));
 b15ztpn00an1n08x5 PHY_10 ();
 b15nor002al1n06x5 U4167 (.a(n3540),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[7]));
 b15inv000as1n40x5 U4168 (.a(net16),
    .o1(n3550));
 b15norp02aq1n03x5 U4169 (.a(net476),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[3]));
 b15inv000as1n80x5 U4170 (.a(net507),
    .o1(n3542));
 b15norp02an1n04x5 U4171 (.a(net474),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[8]));
 b15inv000as1n24x5 U4172 (.a(net15),
    .o1(n3545));
 b15nor002ah1n02x5 U4173 (.a(net473),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[2]));
 b15inv000an1n80x5 U4174 (.a(net25),
    .o1(n3544));
 b15ztpn00an1n08x5 PHY_9 ();
 b15norp02an1n04x5 U4176 (.a(n3544),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[12]));
 b15inv040an1n60x5 U4177 (.a(net13),
    .o1(n3546));
 b15norp02aq1n04x5 U4178 (.a(n3546),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[0]));
 b15nor002ah1n04x5 U4179 (.a(n3546),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[0]));
 b15norp02al1n04x5 U4180 (.a(n3546),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[0]));
 b15inv040as1n40x5 U4181 (.a(net27),
    .o1(n3554));
 b15nor002an1n03x5 U4182 (.a(n3554),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[14]));
 b15inv000as1n40x5 U4183 (.a(net23),
    .o1(n3549));
 b15nor002ar1n04x5 U4184 (.a(net471),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[10]));
 b15inv000as1n80x5 U4185 (.a(net506),
    .o1(n3552));
 b15nor002ah1n02x5 U4186 (.a(net469),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[9]));
 b15ztpn00an1n08x5 PHY_8 ();
 b15nor002an1n06x5 U4188 (.a(n3544),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[12]));
 b15inv040as1n36x5 U4189 (.a(net26),
    .o1(n3547));
 b15nor002aq1n03x5 U4190 (.a(net466),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[13]));
 b15norp02as1n03x5 U4191 (.a(net468),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[9]));
 b15norp02an1n02x5 U4192 (.a(net473),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[2]));
 b15inv000as1n20x5 U4193 (.a(net18),
    .o1(n3553));
 b15norp02aq1n03x5 U4194 (.a(net465),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[5]));
 b15norp02ar1n04x5 U4195 (.a(net471),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[10]));
 b15nor002an1n03x5 U4196 (.a(net477),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[3]));
 b15norp02al1n04x5 U4197 (.a(net468),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[9]));
 b15inv000as1n24x5 U4198 (.a(net17),
    .o1(n3551));
 b15norp02aq1n04x5 U4199 (.a(net462),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[4]));
 b15inv040aq1n48x5 U4200 (.a(net28),
    .o1(n3555));
 b15nor002ar1n06x5 U4201 (.a(n3555),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[15]));
 b15inv020as1n56x5 U4202 (.a(net19),
    .o1(n3557));
 b15norp02al1n08x5 U4203 (.a(n3557),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[6]));
 b15nor002ah1n02x5 U4204 (.a(net474),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[8]));
 b15nor002aq1n03x5 U4205 (.a(net473),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[2]));
 b15inv020an1n80x5 U4206 (.a(net508),
    .o1(n3541));
 b15nor002as1n03x5 U4207 (.a(n3541),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[1]));
 b15nor002aq1n04x5 U4208 (.a(n3555),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[15]));
 b15nor002aq1n02x5 U4209 (.a(net476),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[3]));
 b15norp02as1n02x5 U4210 (.a(net463),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[4]));
 b15inv040as1n36x5 U4211 (.a(net24),
    .o1(n3548));
 b15norp02an1n04x5 U4212 (.a(net460),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[11]));
 b15norp02al1n04x5 U4213 (.a(net461),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[11]));
 b15ztpn00an1n08x5 PHY_7 ();
 b15norp02ar1n04x5 U4215 (.a(n3555),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[15]));
 b15norp02as1n02x5 U4216 (.a(net463),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[4]));
 b15nor002al1n02x5 U4217 (.a(net470),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[10]));
 b15nor002an1n03x5 U4218 (.a(net475),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[8]));
 b15norp02as1n03x5 U4219 (.a(net460),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[11]));
 b15norp02aq1n03x5 U4220 (.a(net467),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[13]));
 b15nor002ah1n02x5 U4221 (.a(net468),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[9]));
 b15ztpn00an1n08x5 PHY_6 ();
 b15norp02ar1n03x5 U4223 (.a(n3555),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[15]));
 b15nor002ar1n06x5 U4224 (.a(n3541),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[1]));
 b15nor002ah1n02x5 U4225 (.a(net470),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[10]));
 b15nor002ar1n04x5 U4226 (.a(n3541),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[1]));
 b15nor002al1n04x5 U4227 (.a(n3554),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[14]));
 b15nor002as1n02x5 U4228 (.a(n3554),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[14]));
 b15nor002ar1n04x5 U4229 (.a(net466),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[13]));
 b15nor002an1n02x5 U4230 (.a(n3551),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[4]));
 b15norp02ar1n03x5 U4231 (.a(net464),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[5]));
 b15nor002al1n03x5 U4232 (.a(n3544),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[12]));
 b15nor002an1n03x5 U4233 (.a(net460),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[11]));
 b15norp02an1n03x5 U4234 (.a(net464),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[5]));
 b15norp02an1n02x5 U4235 (.a(net476),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[3]));
 b15norp02as1n03x5 U4236 (.a(n3541),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[1]));
 b15nor002ar1n02x5 U4237 (.a(n3544),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[12]));
 b15nor002ar1n03x5 U4238 (.a(net474),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[8]));
 b15nor002aq1n06x5 U4239 (.a(net472),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[2]));
 b15nor002ah1n04x5 U4240 (.a(n3557),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[6]));
 b15nor002aq1n03x5 U4241 (.a(n3554),
    .b(net215),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[14]));
 b15nor002aq1n03x5 U4242 (.a(net466),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[13]));
 b15nor002an1n04x5 U4243 (.a(n3557),
    .b(net213),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[6]));
 b15nor002an1n03x5 U4244 (.a(net464),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[5]));
 b15nor002aq1n03x5 U4245 (.a(n3546),
    .b(net216),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[0]));
 b15nor002as1n02x5 U4246 (.a(n3557),
    .b(net220),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[6]));
 b15ztpn00an1n08x5 PHY_5 ();
 b15norp02as1n04x5 U4248 (.a(net490),
    .b(net218),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[21]));
 b15nor002ah1n02x5 U4249 (.a(net490),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[21]));
 b15nor002ah1n03x5 U4250 (.a(net491),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[21]));
 b15and003as1n24x5 U4251 (.a(n3257),
    .b(net51),
    .c(n3120),
    .o(n3665));
 b15ztpn00an1n08x5 PHY_4 ();
 b15nandp2ar1n48x5 U4253 (.a(n3256),
    .b(net421),
    .o1(n3129));
 b15ztpn00an1n08x5 PHY_3 ();
 b15ztpn00an1n08x5 PHY_2 ();
 b15norp02as1n03x5 U4256 (.a(n3540),
    .b(net211),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[7]));
 b15norp02as1n03x5 U4257 (.a(net491),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[21]));
 b15ztpn00an1n08x5 PHY_1 ();
 b15norp02al1n03x5 U4259 (.a(net496),
    .b(net218),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[17]));
 b15ztpn00an1n08x5 PHY_0 ();
 b15nor002an1n03x5 U4261 (.a(net501),
    .b(net218),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[16]));
 b15nor002aq1n03x5 U4263 (.a(net494),
    .b(net218),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[19]));
 b15nor002aq1n03x5 U4265 (.a(n3893),
    .b(net218),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[18]));
 b15norp02aq1n04x5 U4267 (.a(net489),
    .b(net218),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[22]));
 b15norp02an1n04x5 U4268 (.a(net488),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[22]));
 b15norp02as1n03x5 U4270 (.a(net487),
    .b(net218),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[23]));
 b15norp02al1n04x5 U4271 (.a(net486),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[23]));
 b15nor002an1n03x5 U4272 (.a(net497),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[17]));
 b15norp02as1n03x5 U4273 (.a(net495),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[19]));
 b15nor002al1n04x5 U4274 (.a(n3893),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[18]));
 b15nor002aq1n03x5 U4276 (.a(net492),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[20]));
 b15norp02ar1n08x5 U4277 (.a(net486),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[23]));
 b15norp02as1n04x5 U4278 (.a(net493),
    .b(net218),
    .o1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[20]));
 b15norp02an1n04x5 U4279 (.a(net492),
    .b(n3032),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[20]));
 b15nor002al1n06x5 U4280 (.a(net499),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[16]));
 b15norp02an1n04x5 U4281 (.a(net497),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[17]));
 b15nor002ar1n04x5 U4282 (.a(net499),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[16]));
 b15norp02an1n04x5 U4283 (.a(net495),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[19]));
 b15norp02ar1n08x5 U4284 (.a(net488),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[22]));
 b15nor002aq1n03x5 U4285 (.a(net492),
    .b(n3034),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[20]));
 b15norp02an1n04x5 U4286 (.a(net486),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[23]));
 b15norp02al1n04x5 U4287 (.a(net488),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[22]));
 b15nor002aq1n04x5 U4290 (.a(net466),
    .b(net211),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[13]));
 b15norp02ah1n04x5 U4291 (.a(net472),
    .b(net211),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[2]));
 b15nor002aq1n04x5 U4292 (.a(n3546),
    .b(net211),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[0]));
 b15nor002al1n06x5 U4293 (.a(net497),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[17]));
 b15nor002as1n03x5 U4294 (.a(net495),
    .b(net214),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[19]));
 b15nor002ah1n03x5 U4295 (.a(net469),
    .b(net211),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[9]));
 b15nor002an1n03x5 U4296 (.a(net465),
    .b(net211),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[5]));
 b15qgbno2an1n05x5 U4297 (.o1(u_gpio_u_reg_u_intr_enable_wr_data[3]),
    .a(net477),
    .b(net211));
 b15nor002ar1n04x5 U4298 (.a(n3554),
    .b(net211),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[14]));
 b15norp02an1n04x5 U4299 (.a(n3893),
    .b(net212),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[18]));
 b15nor002aq1n03x5 U4300 (.a(n3893),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[18]));
 b15nor002ah1n03x5 U4301 (.a(net463),
    .b(net211),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[4]));
 b15nor002an1n03x5 U4302 (.a(n3555),
    .b(net211),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[15]));
 b15norp02an1n04x5 U4303 (.a(net500),
    .b(net219),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[16]));
 b15norp02as1n03x5 U4304 (.a(n3557),
    .b(net211),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[6]));
 b15norp02as1n02x5 U4305 (.a(n3541),
    .b(net211),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[1]));
 b15qgbno2an1n05x5 U4306 (.o1(u_gpio_u_reg_u_intr_enable_wr_data[10]),
    .a(net471),
    .b(net211));
 b15nor002ar1n04x5 U4307 (.a(net475),
    .b(net211),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[8]));
 b15norp02ar1n04x5 U4308 (.a(n3544),
    .b(net211),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[12]));
 b15norp02al1n02x5 U4309 (.a(net461),
    .b(net211),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[11]));
 b15nor002aq1n03x5 U4310 (.a(net490),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[21]));
 b15norp02ar1n03x5 U4311 (.a(net501),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[16]));
 b15norp02al1n03x5 U4312 (.a(net494),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[19]));
 b15nor002ar1n03x5 U4313 (.a(n3893),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[18]));
 b15nor002aq1n03x5 U4314 (.a(net487),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[23]));
 b15nor002ar1n03x5 U4315 (.a(net493),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[20]));
 b15norp02aq1n03x5 U4316 (.a(net489),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[22]));
 b15norp02aq1n02x5 U4317 (.a(net496),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[17]));
 b15nor002an1n02x5 U4320 (.a(net483),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[30]));
 b15nor002an1n03x5 U4321 (.a(net484),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[28]));
 b15nor002ah1n02x5 U4322 (.a(n3901),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[26]));
 b15nor002an1n03x5 U4323 (.a(n3904),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[29]));
 b15norp02an1n04x5 U4324 (.a(net479),
    .b(n3129),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[31]));
 b15nor002aq1n03x5 U4325 (.a(n3899),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[24]));
 b15norp02aq1n04x5 U4326 (.a(n3902),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[27]));
 b15norp02ar1n04x5 U4327 (.a(n3900),
    .b(net210),
    .o1(u_gpio_u_reg_u_intr_enable_wr_data[25]));
 b15aoi022as1n04x5 U4330 (.a(u_gpio_reg2hw[31]),
    .b(net429),
    .c(net420),
    .d(u_gpio_reg2hw[191]),
    .o1(n3143));
 b15nand02ah1n32x5 U4331 (.a(net53),
    .b(n3131),
    .o1(n3642));
 b15norp03ah1n16x5 U4332 (.a(net52),
    .b(n3247),
    .c(n3642),
    .o1(n3797));
 b15aoi022as1n12x5 U4333 (.a(net301),
    .b(net433),
    .c(net269),
    .d(net103),
    .o1(n3142));
 b15nor002an1n24x5 U4334 (.a(n3137),
    .b(n3642),
    .o1(n3132));
 b15aoi022aq1n12x5 U4337 (.a(u_gpio_reg2hw[159]),
    .b(net253),
    .c(net263),
    .d(u_gpio_u_reg_data_in_qs[31]),
    .o1(n3141));
 b15nand02as1n48x5 U4338 (.a(net52),
    .b(n3247),
    .o1(n3641));
 b15norp02ar1n32x5 U4339 (.a(n3641),
    .b(n3529),
    .o1(n3133));
 b15nor004as1n12x5 U4344 (.a(net53),
    .b(net54),
    .c(net52),
    .d(net51),
    .o1(n3135));
 b15norp02al1n08x5 U4348 (.a(n3137),
    .b(n3640),
    .o1(n3798));
 b15aoi022al1n04x5 U4349 (.a(u_gpio_reg2hw[127]),
    .b(net278),
    .c(net390),
    .d(net246),
    .o1(n3138));
 b15aob012an1n04x5 U4350 (.a(n3138),
    .b(net455),
    .c(u_gpio_reg2hw[223]),
    .out0(n3139));
 b15aoi112as1n08x5 U4351 (.a(net225),
    .b(n3139),
    .c(u_gpio_reg2hw[63]),
    .d(net259),
    .o1(n3140));
 b15nand04as1n16x5 U4352 (.a(n3143),
    .b(net248),
    .c(n3141),
    .d(n3140),
    .o1(u_gpio_u_reg_u_reg_if_N45));
 b15aoi022ah1n12x5 U4353 (.a(u_gpio_reg2hw[91]),
    .b(net432),
    .c(net274),
    .d(net368),
    .o1(n3149));
 b15aoi022an1n12x5 U4354 (.a(net396),
    .b(net246),
    .c(net263),
    .d(u_gpio_u_reg_data_in_qs[27]),
    .o1(n3148));
 b15aoi022ar1n12x5 U4356 (.a(net292),
    .b(net259),
    .c(net420),
    .d(u_gpio_reg2hw[187]),
    .o1(n3147));
 b15aoi022as1n06x5 U4358 (.a(u_gpio_reg2hw[155]),
    .b(net253),
    .c(u_gpio_reg2hw[123]),
    .d(net276),
    .o1(n3144));
 b15aob012ah1n04x5 U4359 (.a(n3144),
    .b(net455),
    .c(u_gpio_reg2hw[219]),
    .out0(n3145));
 b15aoi112al1n08x5 U4360 (.a(net225),
    .b(n3145),
    .c(u_gpio_reg2hw[27]),
    .d(net427),
    .o1(n3146));
 b15nand04as1n16x5 U4361 (.a(n3149),
    .b(n3148),
    .c(n3147),
    .d(n3146),
    .o1(u_gpio_u_reg_u_reg_if_N41));
 b15aoi022ar1n04x5 U4363 (.a(u_gpio_reg2hw[25]),
    .b(net427),
    .c(u_gpio_reg2hw[153]),
    .d(net253),
    .o1(n3157));
 b15aoi022aq1n02x5 U4364 (.a(u_gpio_reg2hw[89]),
    .b(net432),
    .c(net270),
    .d(net370),
    .o1(n3156));
 b15aoi022aq1n02x5 U4365 (.a(u_gpio_reg2hw[57]),
    .b(net259),
    .c(net420),
    .d(u_gpio_reg2hw[185]),
    .o1(n3155));
 b15aoi022al1n02x5 U4368 (.a(net401),
    .b(net246),
    .c(net263),
    .d(u_gpio_u_reg_data_in_qs[25]),
    .o1(n3151));
 b15aob012aq1n04x5 U4369 (.a(n3151),
    .b(net455),
    .c(u_gpio_reg2hw[217]),
    .out0(n3152));
 b15aoi112as1n04x5 U4370 (.a(net225),
    .b(n3152),
    .c(u_gpio_reg2hw[121]),
    .d(net276),
    .o1(n3154));
 b15nand04an1n08x5 U4371 (.a(n3157),
    .b(n3156),
    .c(n3155),
    .d(n3154),
    .o1(u_gpio_u_reg_u_reg_if_N39));
 b15aoi022as1n12x5 U4372 (.a(net340),
    .b(net428),
    .c(u_gpio_reg2hw[150]),
    .d(net258),
    .o1(n3164));
 b15aoi022as1n04x5 U4373 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[6]),
    .b(net246),
    .c(net420),
    .d(u_gpio_reg2hw[182]),
    .o1(n3163));
 b15aoi022as1n08x5 U4374 (.a(net293),
    .b(net259),
    .c(net272),
    .d(net375),
    .o1(n3162));
 b15aoi022an1n12x5 U4377 (.a(u_gpio_reg2hw[118]),
    .b(net276),
    .c(net264),
    .d(u_gpio_u_reg_data_in_qs[22]),
    .o1(n3158));
 b15aob012an1n04x5 U4378 (.a(n3158),
    .b(net458),
    .c(u_gpio_reg2hw[214]),
    .out0(n3159));
 b15aoi112as1n08x5 U4379 (.a(net225),
    .b(n3159),
    .c(u_gpio_reg2hw[86]),
    .d(net431),
    .o1(n3161));
 b15nand04as1n16x5 U4380 (.a(n3164),
    .b(n3163),
    .c(n3162),
    .d(n3161),
    .o1(u_gpio_u_reg_u_reg_if_N36));
 b15aoi022an1n12x5 U4381 (.a(u_gpio_reg2hw[149]),
    .b(net252),
    .c(u_gpio_reg2hw[53]),
    .d(net259),
    .o1(n3171));
 b15aoi022al1n12x5 U4383 (.a(net341),
    .b(net428),
    .c(u_gpio_reg2hw[85]),
    .d(net431),
    .o1(n3170));
 b15aoi022aq1n16x5 U4384 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[5]),
    .b(net247),
    .c(net271),
    .d(net377),
    .o1(n3169));
 b15inv020aq1n08x5 U4385 (.a(u_gpio_reg2hw[213]),
    .o1(n3339));
 b15aoi022an1n02x5 U4386 (.a(net420),
    .b(u_gpio_reg2hw[181]),
    .c(net264),
    .d(u_gpio_u_reg_data_in_qs[21]),
    .o1(n3166));
 b15oai012ar1n06x5 U4387 (.a(n3166),
    .b(n3933),
    .c(n3339),
    .o1(n3167));
 b15aoi112as1n04x5 U4388 (.a(net225),
    .b(n3167),
    .c(u_gpio_reg2hw[117]),
    .d(net277),
    .o1(n3168));
 b15nand04aq1n12x5 U4389 (.a(n3171),
    .b(n3170),
    .c(n3169),
    .d(n3168),
    .o1(u_gpio_u_reg_u_reg_if_N35));
 b15aoi022ar1n32x5 U4391 (.a(u_gpio_reg2hw[146]),
    .b(net252),
    .c(u_gpio_reg2hw[50]),
    .d(net259),
    .o1(n3178));
 b15aoi022ar1n12x5 U4392 (.a(net306),
    .b(net430),
    .c(n3665),
    .d(u_gpio_reg2hw[178]),
    .o1(n3177));
 b15aoi022an1n48x5 U4393 (.a(net271),
    .b(net88),
    .c(net264),
    .d(u_gpio_u_reg_data_in_qs[18]),
    .o1(n3176));
 b15aoi022ar1n24x5 U4394 (.a(u_gpio_reg2hw[114]),
    .b(net277),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[2]),
    .d(net247),
    .o1(n3173));
 b15aob012as1n02x5 U4395 (.a(n3173),
    .b(net458),
    .c(u_gpio_reg2hw[210]),
    .out0(n3174));
 b15aoi112aq1n06x5 U4396 (.a(net225),
    .b(n3174),
    .c(net347),
    .d(net429),
    .o1(n3175));
 b15nand04as1n16x5 U4397 (.a(n3178),
    .b(n3177),
    .c(n3176),
    .d(n3175),
    .o1(u_gpio_u_reg_u_reg_if_N32));
 b15aoi022an1n12x5 U4398 (.a(u_gpio_reg2hw[144]),
    .b(net253),
    .c(net420),
    .d(u_gpio_reg2hw[176]),
    .o1(n3184));
 b15aoi022an1n32x5 U4399 (.a(net269),
    .b(net383),
    .c(net267),
    .d(u_gpio_u_reg_data_in_qs[16]),
    .o1(n3183));
 b15aoi022an1n16x5 U4400 (.a(u_gpio_reg2hw[16]),
    .b(net428),
    .c(net307),
    .d(n3027),
    .o1(n3182));
 b15aoi022an1n04x5 U4401 (.a(u_gpio_reg2hw[112]),
    .b(net277),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[0]),
    .d(net247),
    .o1(n3179));
 b15aob012an1n04x5 U4402 (.a(n3179),
    .b(net458),
    .c(u_gpio_reg2hw[208]),
    .out0(n3180));
 b15aoi112as1n08x5 U4403 (.a(net225),
    .b(n3180),
    .c(u_gpio_reg2hw[48]),
    .d(net259),
    .o1(n3181));
 b15nand04as1n16x5 U4404 (.a(n3184),
    .b(n3183),
    .c(n3182),
    .d(n3181),
    .o1(u_gpio_u_reg_u_reg_if_N30));
 b15aoi022ah1n12x5 U4405 (.a(net336),
    .b(net427),
    .c(net274),
    .d(net372),
    .o1(n3190));
 b15aoi022an1n06x5 U4406 (.a(u_gpio_reg2hw[152]),
    .b(net258),
    .c(net263),
    .d(u_gpio_u_reg_data_in_qs[24]),
    .o1(n3189));
 b15aoi022an1n12x5 U4407 (.a(net402),
    .b(net246),
    .c(net420),
    .d(u_gpio_reg2hw[184]),
    .o1(n3188));
 b15aoi022an1n04x5 U4408 (.a(u_gpio_reg2hw[56]),
    .b(net259),
    .c(u_gpio_reg2hw[120]),
    .d(net279),
    .o1(n3185));
 b15aob012ar1n06x5 U4409 (.a(n3185),
    .b(net459),
    .c(u_gpio_reg2hw[216]),
    .out0(n3186));
 b15aoi112ah1n06x5 U4410 (.a(net225),
    .b(n3186),
    .c(u_gpio_reg2hw[88]),
    .d(net432),
    .o1(n3187));
 b15nand04aq1n12x5 U4411 (.a(n3190),
    .b(n3189),
    .c(n3188),
    .d(n3187),
    .o1(u_gpio_u_reg_u_reg_if_N38));
 b15aoi022aq1n08x5 U4412 (.a(u_gpio_reg2hw[148]),
    .b(net252),
    .c(u_gpio_reg2hw[52]),
    .d(net259),
    .o1(n3196));
 b15aoi022as1n08x5 U4413 (.a(u_gpio_reg2hw[84]),
    .b(net431),
    .c(net272),
    .d(net378),
    .o1(n3195));
 b15aoi022aq1n12x5 U4414 (.a(net343),
    .b(net428),
    .c(u_gpio_reg2hw[116]),
    .d(net277),
    .o1(n3194));
 b15aoi022aq1n08x5 U4415 (.a(net420),
    .b(u_gpio_reg2hw[180]),
    .c(net264),
    .d(u_gpio_u_reg_data_in_qs[20]),
    .o1(n3191));
 b15aob012as1n02x5 U4416 (.a(n3191),
    .b(net455),
    .c(u_gpio_reg2hw[212]),
    .out0(n3192));
 b15aoi112aq1n08x5 U4417 (.a(net225),
    .b(n3192),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[4]),
    .d(net247),
    .o1(n3193));
 b15nand04as1n16x5 U4418 (.a(n3196),
    .b(n3195),
    .c(n3194),
    .d(n3193),
    .o1(u_gpio_u_reg_u_reg_if_N34));
 b15aoi022aq1n32x5 U4419 (.a(net409),
    .b(net247),
    .c(net273),
    .d(net381),
    .o1(n3204));
 b15aoi022ah1n32x5 U4420 (.a(u_gpio_reg2hw[49]),
    .b(net259),
    .c(u_gpio_reg2hw[113]),
    .d(net276),
    .o1(n3203));
 b15aoi022aq1n08x5 U4421 (.a(net420),
    .b(u_gpio_reg2hw[177]),
    .c(net262),
    .d(u_gpio_u_reg_data_in_qs[17]),
    .o1(n3202));
 b15aoi022an1n16x5 U4423 (.a(u_gpio_reg2hw[81]),
    .b(net431),
    .c(u_gpio_reg2hw[145]),
    .d(net252),
    .o1(n3199));
 b15aob012al1n06x5 U4424 (.a(n3199),
    .b(net455),
    .c(u_gpio_reg2hw[209]),
    .out0(n3200));
 b15aoi112as1n08x5 U4425 (.a(net225),
    .b(n3200),
    .c(u_gpio_reg2hw[17]),
    .d(net428),
    .o1(n3201));
 b15nand04as1n16x5 U4426 (.a(n3204),
    .b(n3203),
    .c(n3202),
    .d(n3201),
    .o1(u_gpio_u_reg_u_reg_if_N31));
 b15aoi022al1n32x5 U4427 (.a(net405),
    .b(net247),
    .c(net273),
    .d(net373),
    .o1(n3212));
 b15aoi022aq1n32x5 U4428 (.a(u_gpio_reg2hw[55]),
    .b(net259),
    .c(u_gpio_reg2hw[119]),
    .d(net276),
    .o1(n3211));
 b15aoi022aq1n08x5 U4429 (.a(net305),
    .b(net430),
    .c(net420),
    .d(u_gpio_reg2hw[183]),
    .o1(n3210));
 b15aoi022ar1n02x3 U4431 (.a(u_gpio_reg2hw[151]),
    .b(net252),
    .c(net262),
    .d(u_gpio_u_reg_data_in_qs[23]),
    .o1(n3206));
 b15aob012al1n04x5 U4432 (.a(n3206),
    .b(net455),
    .c(u_gpio_reg2hw[215]),
    .out0(n3207));
 b15aoi112ar1n08x5 U4433 (.a(net225),
    .b(n3207),
    .c(u_gpio_reg2hw[23]),
    .d(net428),
    .o1(n3209));
 b15nand04as1n16x5 U4434 (.a(n3212),
    .b(n3211),
    .c(n3210),
    .d(n3209),
    .o1(u_gpio_u_reg_u_reg_if_N37));
 b15nand02ah1n32x5 U4435 (.a(n3256),
    .b(net269),
    .o1(n3237));
 b15nano23as1n24x5 U4437 (.a(net53),
    .b(net52),
    .c(n3247),
    .d(net54),
    .out0(n3761));
 b15nandp2an1n16x5 U4438 (.a(n3256),
    .b(net417),
    .o1(n3226));
 b15nandp2ar1n02x5 U4439 (.a(net205),
    .b(n3226),
    .o1(u_gpio_N55));
 b15orn002aq1n32x5 U4440 (.a(u_gpio_u_reg_err_q),
    .b(net454),
    .o(u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_req_trigger));
 b15nonb02ah1n16x5 U4441 (.a(n3213),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_req_trigger),
    .out0(n3248));
 b15inv000al1n02x5 U4442 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[0]),
    .o1(n3214));
 b15oaoi13aq1n04x5 U4443 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .b(n3214),
    .c(n3216),
    .d(n3215),
    .o1(n3218));
 b15aoi012an1n06x5 U4444 (.a(net2029),
    .b(n3218),
    .c(n3217),
    .o1(n3811));
 b15nor003aq1n02x5 U4445 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .c(n3811),
    .o1(n3219));
 b15aoi012al1n04x5 U4446 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .b(n3248),
    .c(n3219),
    .o1(n3224));
 b15oai012ar1n02x5 U4447 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .c(n3222),
    .o1(n3221));
 b15aoai13ar1n02x3 U4448 (.a(n3220),
    .b(n3221),
    .c(n3222),
    .d(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .o1(n3223));
 b15oaoi13an1n02x5 U4449 (.a(n3223),
    .b(n3224),
    .c(n3250),
    .d(n3225),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_d[1]));
 b15nor002as1n06x5 U4451 (.a(net464),
    .b(n3896),
    .o1(n3288));
 b15aoai13al1n02x5 U4453 (.a(net199),
    .b(n3288),
    .c(net92),
    .d(n3896),
    .o1(n3227));
 b15oai012ar1n03x5 U4454 (.a(n3227),
    .b(net204),
    .c(n3896),
    .o1(u_gpio_N61));
 b15qgbno2an1n05x5 U4455 (.o1(n3271),
    .a(n3901),
    .b(n3549));
 b15aoai13ar1n06x5 U4456 (.a(net198),
    .b(n3271),
    .c(net97),
    .d(n3901),
    .o1(n3228));
 b15oai012aq1n03x5 U4457 (.a(n3228),
    .b(net207),
    .c(n3901),
    .o1(u_gpio_N66));
 b15norp02as1n12x5 U4458 (.a(n3554),
    .b(net482),
    .o1(n3267));
 b15aoai13as1n08x5 U4459 (.a(net200),
    .b(n3267),
    .c(net366),
    .d(net482),
    .o1(n3229));
 b15oai012al1n24x5 U4460 (.a(n3229),
    .b(net205),
    .c(net482),
    .o1(u_gpio_N70));
 b15norp02as1n04x5 U4461 (.a(n3902),
    .b(n3548),
    .o1(n3282));
 b15aoai13ar1n02x3 U4462 (.a(net198),
    .b(n3282),
    .c(net98),
    .d(n3902),
    .o1(n3230));
 b15oai012ah1n02x5 U4463 (.a(n3230),
    .b(net207),
    .c(n3902),
    .o1(u_gpio_N67));
 b15norp02al1n08x5 U4464 (.a(n3895),
    .b(n3551),
    .o1(n3263));
 b15aoai13as1n02x5 U4465 (.a(net199),
    .b(n3263),
    .c(net91),
    .d(n3895),
    .o1(n3231));
 b15oai012ar1n02x5 U4466 (.a(n3231),
    .b(net204),
    .c(n3895),
    .o1(u_gpio_N60));
 b15nor002ar1n06x5 U4467 (.a(n3545),
    .b(n3893),
    .o1(n3293));
 b15aoai13ar1n03x5 U4468 (.a(net199),
    .b(n3293),
    .c(net88),
    .d(n3893),
    .o1(n3232));
 b15oai012as1n03x5 U4469 (.a(n3232),
    .b(net208),
    .c(n3893),
    .o1(u_gpio_N58));
 b15nor002as1n08x5 U4470 (.a(n3899),
    .b(n3542),
    .o1(n3286));
 b15aoai13ar1n02x5 U4471 (.a(net198),
    .b(n3286),
    .c(net372),
    .d(n3899),
    .o1(n3233));
 b15oai012an1n02x5 U4472 (.a(n3233),
    .b(net207),
    .c(n3899),
    .o1(u_gpio_N64));
 b15norp02aq1n08x5 U4473 (.a(net495),
    .b(n3550),
    .o1(n3280));
 b15aoai13al1n02x5 U4474 (.a(net199),
    .b(n3280),
    .c(net89),
    .d(n3894),
    .o1(n3234));
 b15oai012aq1n04x5 U4475 (.a(n3234),
    .b(net208),
    .c(n3894),
    .o1(u_gpio_N59));
 b15norp02al1n12x5 U4476 (.a(n3541),
    .b(n3892),
    .o1(n3278));
 b15aoai13an1n02x5 U4477 (.a(net200),
    .b(n3278),
    .c(net87),
    .d(n3892),
    .o1(n3235));
 b15oai012aq1n04x5 U4478 (.a(n3235),
    .b(net206),
    .c(n3892),
    .o1(u_gpio_N57));
 b15nor002aq1n08x5 U4479 (.a(n3547),
    .b(n3904),
    .o1(n3261));
 b15aoai13ah1n02x5 U4480 (.a(net198),
    .b(n3261),
    .c(net100),
    .d(n3904),
    .o1(n3236));
 b15oai012ar1n04x5 U4481 (.a(n3236),
    .b(net207),
    .c(n3904),
    .o1(u_gpio_N69));
 b15nor002ar1n12x5 U4483 (.a(n3546),
    .b(n3891),
    .o1(n3273));
 b15aoai13ah1n03x5 U4484 (.a(net200),
    .b(n3273),
    .c(net384),
    .d(n3891),
    .o1(n3238));
 b15oai012al1n08x5 U4485 (.a(n3238),
    .b(net203),
    .c(n3891),
    .o1(u_gpio_N56));
 b15qgbno2an1n10x5 U4486 (.a(n3898),
    .b(n3540),
    .o1(n3265));
 b15aoai13an1n02x5 U4487 (.a(net200),
    .b(n3265),
    .c(net94),
    .d(n3898),
    .o1(n3240));
 b15oai012al1n02x5 U4488 (.a(n3240),
    .b(net205),
    .c(n3898),
    .o1(u_gpio_N63));
 b15nor002an1n12x5 U4489 (.a(n3900),
    .b(n3552),
    .o1(n3290));
 b15aoai13an1n02x5 U4490 (.a(net198),
    .b(n3290),
    .c(net96),
    .d(n3900),
    .o1(n3241));
 b15oai012al1n02x5 U4491 (.a(n3241),
    .b(net207),
    .c(n3900),
    .o1(u_gpio_N65));
 b15nor002aq1n16x5 U4492 (.a(n3555),
    .b(net480),
    .o1(n3269));
 b15aoai13as1n08x5 U4493 (.a(net200),
    .b(n3269),
    .c(net363),
    .d(n3906),
    .o1(n3242));
 b15oai012an1n16x5 U4494 (.a(n3242),
    .b(net205),
    .c(n3906),
    .o1(u_gpio_N71));
 b15norp02al1n16x5 U4495 (.a(net485),
    .b(n3544),
    .o1(n3284));
 b15aoai13al1n02x5 U4496 (.a(net198),
    .b(n3284),
    .c(net99),
    .d(n3903),
    .o1(n3243));
 b15oai012ar1n02x5 U4497 (.a(n3243),
    .b(net207),
    .c(n3903),
    .o1(u_gpio_N68));
 b15norp02as1n08x5 U4498 (.a(n3897),
    .b(n3557),
    .o1(n3276));
 b15aoai13aq1n03x5 U4499 (.a(net200),
    .b(n3276),
    .c(net376),
    .d(n3897),
    .o1(n3245));
 b15oai012al1n06x5 U4500 (.a(n3245),
    .b(net205),
    .c(n3897),
    .o1(u_gpio_N62));
 b15nor002aq1n16x5 U4501 (.a(n3640),
    .b(net52),
    .o1(n3760));
 b15inv020ah1n24x5 U4502 (.a(n3256),
    .o1(n3818));
 b15nonb02as1n16x5 U4503 (.a(net242),
    .b(n3818),
    .out0(u_gpio_N113));
 b15nor002al1n24x5 U4504 (.a(n3818),
    .b(n3641),
    .o1(n3530));
 b15nandp2al1n48x5 U4505 (.a(n3530),
    .b(n3246),
    .o1(n3330));
 b15nandp2aq1n32x5 U4506 (.a(u_gpio_N113),
    .b(n3247),
    .o1(n3296));
 b15nand02an1n04x5 U4508 (.a(net184),
    .b(net182),
    .o1(u_gpio_N130));
 b15aoi112ah1n04x5 U4509 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .c(n3811),
    .d(n3248),
    .o1(n3249));
 b15aoai13as1n08x5 U4510 (.a(n3808),
    .b(n3249),
    .c(n3250),
    .d(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .o1(n3332));
 b15nonb02al1n02x5 U4511 (.a(n3332),
    .b(n3809),
    .out0(u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_nd));
 b15norp02as1n08x5 U4512 (.a(n3809),
    .b(n3332),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_pd));
 b15aoi022as1n08x5 U4513 (.a(net505),
    .b(net509),
    .c(net411),
    .d(net499),
    .o1(n3252));
 b15oai022ah1n12x5 U4515 (.a(n3252),
    .b(net184),
    .c(net499),
    .d(net183),
    .o1(u_gpio_N131));
 b15nand02aq1n16x5 U4516 (.a(u_gpio_reg2hw[7]),
    .b(net2193),
    .o1(n3253));
 b15oai012ah1n48x5 U4517 (.a(n3253),
    .b(net320),
    .c(n3254),
    .o1(u_gpio_u_reg_u_data_in_wr_data[7]));
 b15nandp2ar1n32x5 U4519 (.a(net227),
    .b(net457),
    .o1(n3429));
 b15nonb02as1n03x5 U4521 (.a(u_gpio_reg2hw[135]),
    .b(u_gpio_data_in_q[7]),
    .out0(n3260));
 b15aoi012ah1n02x5 U4522 (.a(u_gpio_reg2hw[39]),
    .b(u_gpio_data_in_q[7]),
    .c(u_gpio_reg2hw[103]),
    .o1(n3258));
 b15nandp2as1n32x5 U4523 (.a(n3257),
    .b(n3530),
    .o1(n3343));
 b15oai022ar1n08x5 U4525 (.a(n3258),
    .b(u_gpio_u_reg_u_data_in_wr_data[7]),
    .c(net181),
    .d(n3540),
    .o1(n3259));
 b15oaoi13as1n08x5 U4526 (.a(n3259),
    .b(u_gpio_u_reg_u_data_in_wr_data[7]),
    .c(u_gpio_reg2hw[71]),
    .d(n3260),
    .o1(n3582));
 b15aboi22aq1n06x5 U4527 (.a(u_gpio_reg2hw[199]),
    .b(n3582),
    .c(net20),
    .d(n3937),
    .out0(u_gpio_u_reg_u_intr_state_wr_data[7]));
 b15norp03as1n24x5 U4528 (.a(n3818),
    .b(n3641),
    .c(n3642),
    .o1(n3292));
 b15aoai13as1n08x5 U4529 (.a(net194),
    .b(n3261),
    .c(net385),
    .d(n3904),
    .o1(n3262));
 b15oai012ah1n02x5 U4530 (.a(n3262),
    .b(net208),
    .c(n3547),
    .o1(u_gpio_N52));
 b15aoai13al1n03x5 U4531 (.a(net195),
    .b(n3263),
    .c(net105),
    .d(n3895),
    .o1(n3264));
 b15oai012ar1n02x5 U4532 (.a(n3264),
    .b(net204),
    .c(n3551),
    .o1(u_gpio_N43));
 b15aoai13al1n08x5 U4533 (.a(net196),
    .b(n3265),
    .c(net108),
    .d(n3898),
    .o1(n3266));
 b15oai012ah1n06x5 U4534 (.a(n3266),
    .b(net205),
    .c(n3540),
    .o1(u_gpio_N46));
 b15aoai13an1n02x5 U4535 (.a(net196),
    .b(n3267),
    .c(net84),
    .d(net482),
    .o1(n3268));
 b15oai012ar1n02x5 U4536 (.a(n3268),
    .b(net203),
    .c(n3554),
    .o1(u_gpio_N53));
 b15aoai13as1n08x5 U4537 (.a(net196),
    .b(n3269),
    .c(net85),
    .d(n3906),
    .o1(n3270));
 b15oai012aq1n12x5 U4538 (.a(n3270),
    .b(net203),
    .c(n3555),
    .o1(u_gpio_N54));
 b15aoai13aq1n08x5 U4539 (.a(net194),
    .b(n3271),
    .c(net389),
    .d(n3901),
    .o1(n3272));
 b15oai012ah1n24x5 U4540 (.a(n3272),
    .b(net207),
    .c(n3549),
    .o1(u_gpio_N49));
 b15aoai13al1n08x5 U4541 (.a(net196),
    .b(n3273),
    .c(net79),
    .d(n3891),
    .o1(n3274));
 b15oai012al1n08x5 U4542 (.a(n3274),
    .b(net203),
    .c(n3546),
    .o1(u_gpio_N39));
 b15aoai13al1n03x5 U4543 (.a(net196),
    .b(n3276),
    .c(net107),
    .d(n3897),
    .o1(n3277));
 b15oai012al1n02x5 U4544 (.a(n3277),
    .b(net205),
    .c(n3557),
    .o1(u_gpio_N45));
 b15aoai13as1n08x5 U4545 (.a(net196),
    .b(n3278),
    .c(net90),
    .d(n3892),
    .o1(n3279));
 b15oai012ar1n12x5 U4546 (.a(n3279),
    .b(net203),
    .c(n3541),
    .o1(u_gpio_N40));
 b15aoai13al1n08x5 U4547 (.a(net195),
    .b(n3280),
    .c(net104),
    .d(net495),
    .o1(n3281));
 b15oai012ar1n08x5 U4548 (.a(n3281),
    .b(net209),
    .c(n3550),
    .o1(u_gpio_N42));
 b15aoai13aq1n08x5 U4549 (.a(net194),
    .b(n3282),
    .c(net388),
    .d(n3902),
    .o1(n3283));
 b15oai012ah1n24x5 U4550 (.a(n3283),
    .b(net207),
    .c(n3548),
    .o1(u_gpio_N50));
 b15aoai13as1n08x5 U4551 (.a(net194),
    .b(n3284),
    .c(net386),
    .d(net484),
    .o1(n3285));
 b15oai012an1n24x5 U4552 (.a(n3285),
    .b(net207),
    .c(n3544),
    .o1(u_gpio_N51));
 b15aoai13as1n08x5 U4553 (.a(net194),
    .b(n3286),
    .c(net362),
    .d(n3899),
    .o1(n3287));
 b15oai012as1n24x5 U4554 (.a(n3287),
    .b(net207),
    .c(n3542),
    .o1(u_gpio_N47));
 b15aoai13ar1n02x5 U4555 (.a(net195),
    .b(n3288),
    .c(net106),
    .d(n3896),
    .o1(n3289));
 b15oai012al1n04x5 U4556 (.a(n3289),
    .b(net204),
    .c(n3553),
    .o1(u_gpio_N44));
 b15aoai13ah1n08x5 U4557 (.a(net194),
    .b(n3290),
    .c(net359),
    .d(n3900),
    .o1(n3291));
 b15oai012an1n32x5 U4558 (.a(n3291),
    .b(net207),
    .c(n3552),
    .o1(u_gpio_N48));
 b15aoai13ah1n03x5 U4559 (.a(net195),
    .b(n3293),
    .c(net101),
    .d(n3893),
    .o1(n3294));
 b15oai012ah1n02x5 U4560 (.a(n3294),
    .b(net209),
    .c(n3545),
    .o1(u_gpio_N41));
 b15aoi022an1n02x5 U4561 (.a(net505),
    .b(net509),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[0]),
    .d(net499),
    .o1(n3297));
 b15nandp2as1n48x5 U4562 (.a(net51),
    .b(u_gpio_N113),
    .o1(n3313));
 b15oai022ah1n02x5 U4564 (.a(n3297),
    .b(n3313),
    .c(n3546),
    .d(net183),
    .o1(u_gpio_N114));
 b15aoi022aq1n48x5 U4565 (.a(net40),
    .b(net24),
    .c(net412),
    .d(n3902),
    .o1(n3298));
 b15oai022an1n12x5 U4566 (.a(n3298),
    .b(n3313),
    .c(net461),
    .d(net182),
    .o1(u_gpio_N125));
 b15aoi022ah1n12x5 U4567 (.a(net31),
    .b(net15),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[2]),
    .d(n3893),
    .o1(n3299));
 b15oai022ar1n12x5 U4568 (.a(n3299),
    .b(n3313),
    .c(net472),
    .d(net183),
    .o1(u_gpio_N116));
 b15aoi022ah1n12x5 U4569 (.a(net42),
    .b(net26),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[13]),
    .d(n3904),
    .o1(n3300));
 b15oai022aq1n06x5 U4570 (.a(n3300),
    .b(n3313),
    .c(net467),
    .d(net182),
    .o1(u_gpio_N127));
 b15aoi022ah1n12x5 U4571 (.a(net32),
    .b(net16),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[3]),
    .d(n3894),
    .o1(n3301));
 b15oai022an1n06x5 U4572 (.a(n3301),
    .b(n3313),
    .c(n3550),
    .d(net183),
    .o1(u_gpio_N117));
 b15aoi022as1n08x5 U4573 (.a(net34),
    .b(net18),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[5]),
    .d(n3896),
    .o1(n3302));
 b15oai022as1n06x5 U4574 (.a(n3302),
    .b(n3313),
    .c(net465),
    .d(net183),
    .o1(u_gpio_N119));
 b15aoi022aq1n08x5 U4575 (.a(net33),
    .b(net17),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[4]),
    .d(n3895),
    .o1(n3303));
 b15oai022ah1n04x5 U4576 (.a(n3303),
    .b(n3313),
    .c(net462),
    .d(net183),
    .o1(u_gpio_N118));
 b15aoi022as1n08x5 U4577 (.a(net41),
    .b(net25),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[12]),
    .d(net484),
    .o1(n3304));
 b15oai022al1n08x5 U4578 (.a(n3304),
    .b(n3313),
    .c(n3544),
    .d(net182),
    .o1(u_gpio_N126));
 b15aoi022al1n04x5 U4579 (.a(net43),
    .b(net27),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[14]),
    .d(n3905),
    .o1(n3305));
 b15oai022ah1n02x5 U4580 (.a(n3305),
    .b(n3313),
    .c(n3554),
    .d(net183),
    .o1(u_gpio_N128));
 b15aoi022an1n06x5 U4581 (.a(net504),
    .b(net508),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[1]),
    .d(net498),
    .o1(n3306));
 b15oai022al1n08x5 U4582 (.a(n3306),
    .b(n3313),
    .c(n3541),
    .d(net183),
    .o1(u_gpio_N115));
 b15aoi022aq1n04x5 U4583 (.a(net35),
    .b(net19),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[6]),
    .d(net489),
    .o1(n3307));
 b15oai022ah1n06x5 U4584 (.a(n3307),
    .b(n3313),
    .c(n3557),
    .d(net183),
    .o1(u_gpio_N120));
 b15aoi022an1n04x5 U4585 (.a(net44),
    .b(net28),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[15]),
    .d(net480),
    .o1(n3308));
 b15oai022an1n06x5 U4586 (.a(n3308),
    .b(n3313),
    .c(n3555),
    .d(net183),
    .o1(u_gpio_N129));
 b15aoi022ar1n04x5 U4587 (.a(net36),
    .b(net20),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[7]),
    .d(net487),
    .o1(n3309));
 b15oai022aq1n06x5 U4588 (.a(n3309),
    .b(n3313),
    .c(n3540),
    .d(net183),
    .o1(u_gpio_N121));
 b15aoi022aq1n12x5 U4589 (.a(net502),
    .b(net506),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[9]),
    .d(n3900),
    .o1(n3310));
 b15oai022al1n12x5 U4590 (.a(n3310),
    .b(n3313),
    .c(net469),
    .d(net182),
    .o1(u_gpio_N123));
 b15aoi022ah1n06x5 U4591 (.a(net39),
    .b(net23),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[10]),
    .d(n3901),
    .o1(n3311));
 b15oai022aq1n12x5 U4592 (.a(n3311),
    .b(n3313),
    .c(net470),
    .d(net182),
    .o1(u_gpio_N124));
 b15aoi022ar1n12x5 U4593 (.a(net503),
    .b(net507),
    .c(u_gpio_u_reg_masked_oe_lower_data_qs[8]),
    .d(n3899),
    .o1(n3314));
 b15oai022as1n08x5 U4594 (.a(n3314),
    .b(n3313),
    .c(net475),
    .d(n3296),
    .o1(u_gpio_N122));
 b15aoi022aq1n02x5 U4595 (.a(net34),
    .b(net18),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[5]),
    .d(n3896),
    .o1(n3315));
 b15oai022ah1n04x5 U4596 (.a(n3315),
    .b(net184),
    .c(n3896),
    .d(net182),
    .o1(u_gpio_N136));
 b15aoi022al1n06x5 U4597 (.a(net41),
    .b(net25),
    .c(net395),
    .d(net484),
    .o1(n3316));
 b15oai022al1n08x5 U4598 (.a(n3316),
    .b(net184),
    .c(net484),
    .d(n3296),
    .o1(u_gpio_N143));
 b15aoi022an1n16x5 U4599 (.a(net35),
    .b(net19),
    .c(net406),
    .d(net489),
    .o1(n3317));
 b15oai022ah1n06x5 U4600 (.a(n3317),
    .b(net184),
    .c(net489),
    .d(net182),
    .o1(u_gpio_N137));
 b15aoi022an1n06x5 U4601 (.a(net39),
    .b(net23),
    .c(net399),
    .d(n3901),
    .o1(n3318));
 b15oai022ah1n08x5 U4602 (.a(n3318),
    .b(net184),
    .c(n3901),
    .d(net182),
    .o1(u_gpio_N141));
 b15aoi022aq1n16x5 U4603 (.a(net504),
    .b(net508),
    .c(net410),
    .d(net498),
    .o1(n3319));
 b15oai022aq1n08x5 U4604 (.a(n3319),
    .b(net184),
    .c(net498),
    .d(net183),
    .o1(u_gpio_N132));
 b15aoi022aq1n02x5 U4605 (.a(net32),
    .b(net16),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[3]),
    .d(n3894),
    .o1(n3320));
 b15oai022aq1n06x5 U4606 (.a(n3320),
    .b(net184),
    .c(n3894),
    .d(net182),
    .o1(u_gpio_N134));
 b15aoi022ar1n04x5 U4607 (.a(net31),
    .b(net15),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[2]),
    .d(n3893),
    .o1(n3321));
 b15oai022as1n02x5 U4608 (.a(n3321),
    .b(net184),
    .c(n3893),
    .d(net182),
    .o1(u_gpio_N133));
 b15aoi022an1n16x5 U4609 (.a(net44),
    .b(net28),
    .c(net391),
    .d(net480),
    .o1(n3322));
 b15oai022al1n08x5 U4610 (.a(n3322),
    .b(net184),
    .c(net480),
    .d(net182),
    .o1(u_gpio_N146));
 b15aoi022ar1n24x5 U4611 (.a(net36),
    .b(net20),
    .c(net404),
    .d(net487),
    .o1(n3323));
 b15oai022al1n06x5 U4612 (.a(n3323),
    .b(net184),
    .c(net487),
    .d(net183),
    .o1(u_gpio_N138));
 b15aoi022ar1n24x5 U4613 (.a(net43),
    .b(net27),
    .c(net392),
    .d(n3905),
    .o1(n3324));
 b15oai022as1n06x5 U4614 (.a(n3324),
    .b(net184),
    .c(n3905),
    .d(net183),
    .o1(u_gpio_N145));
 b15aoi022ah1n04x5 U4615 (.a(net42),
    .b(net26),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[13]),
    .d(n3904),
    .o1(n3325));
 b15oai022as1n06x5 U4616 (.a(n3325),
    .b(net184),
    .c(n3904),
    .d(net182),
    .o1(u_gpio_N144));
 b15aoi022an1n06x5 U4617 (.a(net502),
    .b(net506),
    .c(net401),
    .d(n3900),
    .o1(n3326));
 b15oai022aq1n06x5 U4618 (.a(n3326),
    .b(net184),
    .c(n3900),
    .d(net182),
    .o1(u_gpio_N140));
 b15aoi022an1n04x5 U4619 (.a(net33),
    .b(net17),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[4]),
    .d(n3895),
    .o1(n3327));
 b15oai022an1n06x5 U4620 (.a(n3327),
    .b(n3330),
    .c(n3895),
    .d(net182),
    .o1(u_gpio_N135));
 b15aoi022as1n32x5 U4621 (.a(net40),
    .b(net24),
    .c(net396),
    .d(n3902),
    .o1(n3328));
 b15oai022aq1n08x5 U4622 (.a(n3328),
    .b(net184),
    .c(n3902),
    .d(net183),
    .o1(u_gpio_N142));
 b15aoi022ar1n12x5 U4623 (.a(net503),
    .b(net507),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[8]),
    .d(n3899),
    .o1(n3331));
 b15oai022ar1n08x5 U4624 (.a(n3331),
    .b(net184),
    .c(n3899),
    .d(net182),
    .o1(u_gpio_N139));
 b15oai022an1n02x5 U4625 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .b(n3333),
    .c(n3809),
    .d(n3332),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_d[0]));
 b15qbfna2bn1n16x5 U4626 (.a(net342),
    .b(u_gpio_gen_filter_21__u_filter_stored_value_q),
    .o1(n3334));
 b15oai012as1n48x5 U4627 (.a(n3334),
    .b(net342),
    .c(n3335),
    .o1(u_gpio_u_reg_u_data_in_wr_data[21]));
 b15nonb02al1n06x5 U4628 (.a(u_gpio_reg2hw[149]),
    .b(u_gpio_data_in_q[21]),
    .out0(n3338));
 b15aoi012al1n04x5 U4629 (.a(u_gpio_reg2hw[53]),
    .b(u_gpio_data_in_q[21]),
    .c(u_gpio_reg2hw[117]),
    .o1(n3336));
 b15oai022an1n06x5 U4630 (.a(n3336),
    .b(u_gpio_u_reg_u_data_in_wr_data[21]),
    .c(net180),
    .d(net490),
    .o1(n3337));
 b15oaoi13as1n08x5 U4631 (.a(n3337),
    .b(u_gpio_u_reg_u_data_in_wr_data[21]),
    .c(u_gpio_reg2hw[85]),
    .d(n3338),
    .o1(n3581));
 b15aoi022ah1n08x5 U4632 (.a(n3937),
    .b(net34),
    .c(n3581),
    .d(n3339),
    .o1(u_gpio_u_reg_u_intr_state_wr_data[21]));
 b15inv040al1n10x5 U4633 (.a(u_gpio_gen_filter_3__u_filter_filter_synced),
    .o1(n3341));
 b15nand02aq1n16x5 U4634 (.a(u_gpio_reg2hw[3]),
    .b(u_gpio_gen_filter_3__u_filter_stored_value_q),
    .o1(n3340));
 b15oai012ah1n48x5 U4635 (.a(n3340),
    .b(net328),
    .c(n3341),
    .o1(u_gpio_u_reg_u_data_in_wr_data[3]));
 b15inv000an1n02x5 U4638 (.a(u_gpio_u_reg_u_data_in_wr_data[3]),
    .o1(n3344));
 b15aoai13ah1n08x5 U4639 (.a(n3344),
    .b(u_gpio_reg2hw[35]),
    .c(u_gpio_reg2hw[99]),
    .d(u_gpio_data_in_q[3]),
    .o1(n3347));
 b15inv040aq1n02x5 U4640 (.a(u_gpio_data_in_q[3]),
    .o1(n3345));
 b15aoai13as1n06x5 U4641 (.a(u_gpio_u_reg_u_data_in_wr_data[3]),
    .b(u_gpio_reg2hw[67]),
    .c(u_gpio_reg2hw[131]),
    .d(n3345),
    .o1(n3346));
 b15oai112as1n16x5 U4642 (.a(n3347),
    .b(n3346),
    .c(net181),
    .d(n3550),
    .o1(n3583));
 b15oa0022ar1n04x5 U4643 (.a(net477),
    .b(net201),
    .c(n3583),
    .d(u_gpio_reg2hw[195]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[3]));
 b15inv000ah1n08x5 U4644 (.a(u_gpio_gen_filter_1__u_filter_filter_synced),
    .o1(n3349));
 b15nandp2ah1n08x5 U4645 (.a(net357),
    .b(net2002),
    .o1(n3348));
 b15oai012aq1n48x5 U4646 (.a(n3348),
    .b(net357),
    .c(n3349),
    .o1(u_gpio_u_reg_u_data_in_wr_data[1]));
 b15inv000al1n02x5 U4647 (.a(u_gpio_u_reg_u_data_in_wr_data[1]),
    .o1(n3350));
 b15aoai13as1n06x5 U4648 (.a(n3350),
    .b(u_gpio_reg2hw[33]),
    .c(u_gpio_reg2hw[97]),
    .d(net2134),
    .o1(n3353));
 b15inv000aq1n02x5 U4649 (.a(u_gpio_data_in_q[1]),
    .o1(n3351));
 b15aoai13as1n06x5 U4650 (.a(u_gpio_u_reg_u_data_in_wr_data[1]),
    .b(u_gpio_reg2hw[65]),
    .c(u_gpio_reg2hw[129]),
    .d(n3351),
    .o1(n3352));
 b15oai112as1n16x5 U4651 (.a(n3353),
    .b(n3352),
    .c(net181),
    .d(n3541),
    .o1(n3571));
 b15oa0022as1n02x5 U4652 (.a(n3541),
    .b(net201),
    .c(n3571),
    .d(u_gpio_reg2hw[193]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[1]));
 b15inv000as1n08x5 U4653 (.a(u_gpio_gen_filter_13__u_filter_filter_synced),
    .o1(n3355));
 b15nandp2al1n12x5 U4654 (.a(net354),
    .b(u_gpio_gen_filter_13__u_filter_stored_value_q),
    .o1(n3354));
 b15oai012an1n48x5 U4655 (.a(n3354),
    .b(net354),
    .c(n3355),
    .o1(u_gpio_u_reg_u_data_in_wr_data[13]));
 b15inv000al1n02x5 U4656 (.a(u_gpio_u_reg_u_data_in_wr_data[13]),
    .o1(n3356));
 b15aoai13ar1n08x5 U4657 (.a(n3356),
    .b(net294),
    .c(u_gpio_reg2hw[109]),
    .d(u_gpio_data_in_q[13]),
    .o1(n3359));
 b15inv040ar1n02x5 U4658 (.a(u_gpio_data_in_q[13]),
    .o1(n3357));
 b15aoai13ah1n04x5 U4659 (.a(u_gpio_u_reg_u_data_in_wr_data[13]),
    .b(u_gpio_reg2hw[77]),
    .c(u_gpio_reg2hw[141]),
    .d(n3357),
    .o1(n3358));
 b15oai112as1n16x5 U4660 (.a(n3359),
    .b(n3358),
    .c(net181),
    .d(net466),
    .o1(n3587));
 b15oa0022an1n03x5 U4661 (.a(net467),
    .b(net201),
    .c(n3587),
    .d(u_gpio_reg2hw[205]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[13]));
 b15inv040aq1n06x5 U4662 (.a(net452),
    .o1(n3361));
 b15nand02ar1n16x5 U4663 (.a(net356),
    .b(u_gpio_gen_filter_12__u_filter_stored_value_q),
    .o1(n3360));
 b15oai012ah1n32x5 U4664 (.a(n3360),
    .b(net356),
    .c(n3361),
    .o1(u_gpio_u_reg_u_data_in_wr_data[12]));
 b15inv000al1n02x5 U4665 (.a(u_gpio_u_reg_u_data_in_wr_data[12]),
    .o1(n3362));
 b15aoai13ar1n08x5 U4666 (.a(n3362),
    .b(net296),
    .c(u_gpio_reg2hw[108]),
    .d(u_gpio_data_in_q[12]),
    .o1(n3365));
 b15inv000ah1n02x5 U4667 (.a(u_gpio_data_in_q[12]),
    .o1(n3363));
 b15aoai13ar1n08x5 U4668 (.a(u_gpio_u_reg_u_data_in_wr_data[12]),
    .b(u_gpio_reg2hw[76]),
    .c(u_gpio_reg2hw[140]),
    .d(n3363),
    .o1(n3364));
 b15oai112as1n16x5 U4669 (.a(n3365),
    .b(n3364),
    .c(net181),
    .d(n3544),
    .o1(n3591));
 b15oa0022aq1n03x5 U4670 (.a(n3544),
    .b(net202),
    .c(n3591),
    .d(u_gpio_reg2hw[204]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[12]));
 b15inv040ah1n05x5 U4671 (.a(net451),
    .o1(n3367));
 b15nandp2al1n12x5 U4672 (.a(net351),
    .b(net2189),
    .o1(n3366));
 b15oai012aq1n48x5 U4673 (.a(n3366),
    .b(net351),
    .c(n3367),
    .o1(u_gpio_u_reg_u_data_in_wr_data[14]));
 b15inv000al1n02x5 U4676 (.a(u_gpio_u_reg_u_data_in_wr_data[14]),
    .o1(n3369));
 b15aoai13aq1n06x5 U4677 (.a(n3369),
    .b(u_gpio_reg2hw[46]),
    .c(u_gpio_reg2hw[110]),
    .d(net2076),
    .o1(n3372));
 b15inv000al1n02x5 U4678 (.a(u_gpio_data_in_q[14]),
    .o1(n3370));
 b15aoai13aq1n06x5 U4679 (.a(u_gpio_u_reg_u_data_in_wr_data[14]),
    .b(u_gpio_reg2hw[78]),
    .c(u_gpio_reg2hw[142]),
    .d(n3370),
    .o1(n3371));
 b15oai112as1n16x5 U4680 (.a(n3372),
    .b(n3371),
    .c(net181),
    .d(n3554),
    .o1(n3568));
 b15oa0022ah1n02x5 U4681 (.a(n3554),
    .b(net201),
    .c(n3568),
    .d(u_gpio_reg2hw[206]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[14]));
 b15nandp2al1n05x5 U4682 (.a(u_gpio_reg2hw[10]),
    .b(net1963),
    .o1(n3373));
 b15oai012ah1n16x5 U4683 (.a(n3373),
    .b(u_gpio_reg2hw[10]),
    .c(n3374),
    .o1(u_gpio_u_reg_u_data_in_wr_data[10]));
 b15inv040al1n02x5 U4684 (.a(u_gpio_u_reg_u_data_in_wr_data[10]),
    .o1(n3375));
 b15aoai13aq1n08x5 U4685 (.a(n3375),
    .b(net298),
    .c(net315),
    .d(u_gpio_data_in_q[10]),
    .o1(n3378));
 b15inv040ar1n03x5 U4686 (.a(u_gpio_data_in_q[10]),
    .o1(n3376));
 b15aoai13an1n08x5 U4687 (.a(u_gpio_u_reg_u_data_in_wr_data[10]),
    .b(net311),
    .c(net291),
    .d(n3376),
    .o1(n3377));
 b15oai112as1n16x5 U4688 (.a(n3378),
    .b(n3377),
    .c(n3343),
    .d(net471),
    .o1(n3576));
 b15oa0022aq1n03x5 U4689 (.a(net471),
    .b(net201),
    .c(n3576),
    .d(u_gpio_reg2hw[202]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[10]));
 b15inv000as1n10x5 U4690 (.a(u_gpio_gen_filter_8__u_filter_filter_synced),
    .o1(n3380));
 b15nandp2ah1n08x5 U4691 (.a(net319),
    .b(u_gpio_gen_filter_8__u_filter_stored_value_q),
    .o1(n3379));
 b15oai012an1n48x5 U4692 (.a(n3379),
    .b(net319),
    .c(n3380),
    .o1(u_gpio_u_reg_u_data_in_wr_data[8]));
 b15inv000al1n02x5 U4693 (.a(u_gpio_u_reg_u_data_in_wr_data[8]),
    .o1(n3381));
 b15aoai13as1n06x5 U4694 (.a(n3381),
    .b(u_gpio_reg2hw[40]),
    .c(u_gpio_reg2hw[104]),
    .d(net2104),
    .o1(n3384));
 b15inv020an1n03x5 U4695 (.a(u_gpio_data_in_q[8]),
    .o1(n3382));
 b15aoai13ah1n06x5 U4696 (.a(u_gpio_u_reg_u_data_in_wr_data[8]),
    .b(net300),
    .c(u_gpio_reg2hw[136]),
    .d(n3382),
    .o1(n3383));
 b15oai112as1n16x5 U4697 (.a(n3384),
    .b(n3383),
    .c(net181),
    .d(net474),
    .o1(n3592));
 b15oa0022al1n04x5 U4698 (.a(net475),
    .b(net201),
    .c(n3592),
    .d(u_gpio_reg2hw[200]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[8]));
 b15inv000as1n08x5 U4699 (.a(u_gpio_gen_filter_2__u_filter_filter_synced),
    .o1(n3386));
 b15nand02an1n24x5 U4700 (.a(u_gpio_reg2hw[2]),
    .b(u_gpio_gen_filter_2__u_filter_stored_value_q),
    .o1(n3385));
 b15oai012as1n48x5 U4701 (.a(n3385),
    .b(net330),
    .c(n3386),
    .o1(u_gpio_u_reg_u_data_in_wr_data[2]));
 b15inv040al1n02x5 U4702 (.a(u_gpio_u_reg_u_data_in_wr_data[2]),
    .o1(n3387));
 b15aoai13ah1n08x5 U4703 (.a(n3387),
    .b(u_gpio_reg2hw[34]),
    .c(u_gpio_reg2hw[98]),
    .d(net2081),
    .o1(n3390));
 b15inv020ah1n03x5 U4704 (.a(u_gpio_data_in_q[2]),
    .o1(n3388));
 b15aoai13aq1n08x5 U4705 (.a(u_gpio_u_reg_u_data_in_wr_data[2]),
    .b(net304),
    .c(u_gpio_reg2hw[130]),
    .d(n3388),
    .o1(n3389));
 b15oai112as1n16x5 U4706 (.a(n3390),
    .b(n3389),
    .c(net181),
    .d(net472),
    .o1(n3588));
 b15oa0022ah1n03x5 U4707 (.a(net472),
    .b(net201),
    .c(net2082),
    .d(u_gpio_reg2hw[194]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[2]));
 b15inv040ar1n06x5 U4708 (.a(u_gpio_gen_filter_11__u_filter_filter_synced),
    .o1(n3392));
 b15nandp2as1n04x5 U4709 (.a(u_gpio_reg2hw[11]),
    .b(net2124),
    .o1(n3391));
 b15oai012an1n24x5 U4710 (.a(n3391),
    .b(u_gpio_reg2hw[11]),
    .c(n3392),
    .o1(u_gpio_u_reg_u_data_in_wr_data[11]));
 b15inv000aq1n02x5 U4711 (.a(u_gpio_u_reg_u_data_in_wr_data[11]),
    .o1(n3393));
 b15aoai13ar1n08x5 U4712 (.a(n3393),
    .b(net297),
    .c(net314),
    .d(u_gpio_data_in_q[11]),
    .o1(n3396));
 b15inv000ar1n03x5 U4713 (.a(u_gpio_data_in_q[11]),
    .o1(n3394));
 b15aoai13as1n06x5 U4714 (.a(u_gpio_u_reg_u_data_in_wr_data[11]),
    .b(net310),
    .c(net290),
    .d(n3394),
    .o1(n3395));
 b15oai112as1n16x5 U4715 (.a(n3396),
    .b(n3395),
    .c(net181),
    .d(net461),
    .o1(n3569));
 b15oa0022an1n02x5 U4716 (.a(net461),
    .b(net201),
    .c(n3569),
    .d(u_gpio_reg2hw[203]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[11]));
 b15nandp2ah1n08x5 U4717 (.a(net324),
    .b(u_gpio_gen_filter_5__u_filter_stored_value_q),
    .o1(n3397));
 b15oai012an1n48x5 U4718 (.a(n3397),
    .b(net324),
    .c(n3398),
    .o1(u_gpio_u_reg_u_data_in_wr_data[5]));
 b15inv000al1n02x5 U4719 (.a(u_gpio_u_reg_u_data_in_wr_data[5]),
    .o1(n3399));
 b15aoai13aq1n08x5 U4720 (.a(n3399),
    .b(u_gpio_reg2hw[37]),
    .c(u_gpio_reg2hw[101]),
    .d(u_gpio_data_in_q[5]),
    .o1(n3402));
 b15inv020ah1n03x5 U4721 (.a(u_gpio_data_in_q[5]),
    .o1(n3400));
 b15aoai13ar1n08x5 U4722 (.a(u_gpio_u_reg_u_data_in_wr_data[5]),
    .b(u_gpio_reg2hw[69]),
    .c(u_gpio_reg2hw[133]),
    .d(n3400),
    .o1(n3401));
 b15oai112as1n16x5 U4723 (.a(n3402),
    .b(n3401),
    .c(net181),
    .d(net465),
    .o1(n3573));
 b15oa0022al1n03x5 U4724 (.a(net465),
    .b(net201),
    .c(n3573),
    .d(u_gpio_reg2hw[197]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[5]));
 b15nandp2an1n12x5 U4725 (.a(net348),
    .b(u_gpio_gen_filter_16__u_filter_stored_value_q),
    .o1(n3403));
 b15oai012as1n48x5 U4726 (.a(n3403),
    .b(net348),
    .c(n3404),
    .o1(u_gpio_u_reg_u_data_in_wr_data[16]));
 b15inv000al1n02x5 U4727 (.a(u_gpio_u_reg_u_data_in_wr_data[16]),
    .o1(n3405));
 b15aoai13aq1n08x5 U4728 (.a(n3405),
    .b(u_gpio_reg2hw[48]),
    .c(u_gpio_reg2hw[112]),
    .d(net2177),
    .o1(n3408));
 b15inv020ar1n04x5 U4729 (.a(u_gpio_data_in_q[16]),
    .o1(n3406));
 b15aoai13an1n06x5 U4730 (.a(u_gpio_u_reg_u_data_in_wr_data[16]),
    .b(net308),
    .c(u_gpio_reg2hw[144]),
    .d(n3406),
    .o1(n3407));
 b15oai112as1n16x5 U4731 (.a(n3408),
    .b(n3407),
    .c(net180),
    .d(net500),
    .o1(n3575));
 b15oa0022an1n03x5 U4732 (.a(net500),
    .b(net202),
    .c(n3575),
    .d(u_gpio_reg2hw[208]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[16]));
 b15inv040as1n04x5 U4733 (.a(u_gpio_gen_filter_6__u_filter_filter_synced),
    .o1(n3410));
 b15nand02an1n02x5 U4734 (.a(u_gpio_reg2hw[6]),
    .b(u_gpio_gen_filter_6__u_filter_stored_value_q),
    .o1(n3409));
 b15oai012ar1n08x5 U4735 (.a(n3409),
    .b(u_gpio_reg2hw[6]),
    .c(n3410),
    .o1(u_gpio_u_reg_u_data_in_wr_data[6]));
 b15inv000al1n02x5 U4736 (.a(net241),
    .o1(n3411));
 b15aoai13as1n04x5 U4737 (.a(n3411),
    .b(u_gpio_reg2hw[38]),
    .c(u_gpio_reg2hw[102]),
    .d(u_gpio_data_in_q[6]),
    .o1(n3414));
 b15inv000al1n02x5 U4738 (.a(u_gpio_data_in_q[6]),
    .o1(n3412));
 b15aoai13an1n06x5 U4739 (.a(net241),
    .b(u_gpio_reg2hw[70]),
    .c(u_gpio_reg2hw[134]),
    .d(n3412),
    .o1(n3413));
 b15oai112as1n16x5 U4740 (.a(n3414),
    .b(n3413),
    .c(net181),
    .d(n3557),
    .o1(n3605));
 b15oa0022ah1n03x5 U4741 (.a(n3557),
    .b(net201),
    .c(n3605),
    .d(net2153),
    .o(u_gpio_u_reg_u_intr_state_wr_data[6]));
 b15inv040al1n02x5 U4742 (.a(u_gpio_gen_filter_20__u_filter_filter_synced),
    .o1(n3416));
 b15nandp2an1n02x5 U4743 (.a(u_gpio_reg2hw[20]),
    .b(u_gpio_gen_filter_20__u_filter_stored_value_q),
    .o1(n3415));
 b15oai012ar1n08x5 U4744 (.a(n3415),
    .b(u_gpio_reg2hw[20]),
    .c(n3416),
    .o1(u_gpio_u_reg_u_data_in_wr_data[20]));
 b15inv000al1n02x5 U4745 (.a(net240),
    .o1(n3417));
 b15aoai13aq1n08x5 U4746 (.a(n3417),
    .b(u_gpio_reg2hw[52]),
    .c(u_gpio_reg2hw[116]),
    .d(net2115),
    .o1(n3420));
 b15inv020as1n04x5 U4747 (.a(u_gpio_data_in_q[20]),
    .o1(n3418));
 b15aoai13aq1n06x5 U4748 (.a(net240),
    .b(u_gpio_reg2hw[84]),
    .c(u_gpio_reg2hw[148]),
    .d(n3418),
    .o1(n3419));
 b15oai112as1n16x5 U4749 (.a(n3420),
    .b(n3419),
    .c(net180),
    .d(n3895),
    .o1(n3567));
 b15oa0022ah1n02x5 U4750 (.a(n3895),
    .b(net202),
    .c(net2116),
    .d(u_gpio_reg2hw[212]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[20]));
 b15inv020as1n06x5 U4751 (.a(u_gpio_gen_filter_0__u_filter_filter_synced),
    .o1(n3422));
 b15nandp2al1n08x5 U4752 (.a(u_gpio_reg2hw[0]),
    .b(net2142),
    .o1(n3421));
 b15oai012an1n32x5 U4753 (.a(n3421),
    .b(u_gpio_reg2hw[0]),
    .c(n3422),
    .o1(u_gpio_u_reg_u_data_in_wr_data[0]));
 b15inv000al1n02x5 U4754 (.a(u_gpio_u_reg_u_data_in_wr_data[0]),
    .o1(n3423));
 b15aoai13al1n08x5 U4755 (.a(n3423),
    .b(u_gpio_reg2hw[32]),
    .c(u_gpio_reg2hw[96]),
    .d(u_gpio_data_in_q[0]),
    .o1(n3426));
 b15inv000an1n02x5 U4756 (.a(u_gpio_data_in_q[0]),
    .o1(n3424));
 b15aoai13as1n06x5 U4757 (.a(u_gpio_u_reg_u_data_in_wr_data[0]),
    .b(u_gpio_reg2hw[64]),
    .c(u_gpio_reg2hw[128]),
    .d(n3424),
    .o1(n3425));
 b15oai112as1n16x5 U4758 (.a(n3426),
    .b(n3425),
    .c(net181),
    .d(n3546),
    .o1(n3577));
 b15oa0022as1n03x5 U4759 (.a(n3546),
    .b(net201),
    .c(n3577),
    .d(u_gpio_reg2hw[192]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[0]));
 b15inv020as1n10x5 U4760 (.a(u_gpio_gen_filter_28__u_filter_filter_synced),
    .o1(n3428));
 b15nand02ar1n24x5 U4761 (.a(net333),
    .b(u_gpio_gen_filter_28__u_filter_stored_value_q),
    .o1(n3427));
 b15oai012ah1n48x5 U4762 (.a(n3427),
    .b(net332),
    .c(n3428),
    .o1(u_gpio_u_reg_u_data_in_wr_data[28]));
 b15inv000al1n02x5 U4765 (.a(u_gpio_u_reg_u_data_in_wr_data[28]),
    .o1(n3431));
 b15aoai13ah1n03x5 U4766 (.a(n3431),
    .b(u_gpio_reg2hw[60]),
    .c(u_gpio_reg2hw[124]),
    .d(net1946),
    .o1(n3434));
 b15inv000al1n02x5 U4767 (.a(net1946),
    .o1(n3432));
 b15aoai13ah1n03x5 U4768 (.a(u_gpio_u_reg_u_data_in_wr_data[28]),
    .b(u_gpio_reg2hw[92]),
    .c(u_gpio_reg2hw[156]),
    .d(n3432),
    .o1(n3433));
 b15oai112aq1n16x5 U4769 (.a(n3434),
    .b(n3433),
    .c(net180),
    .d(net485),
    .o1(n3595));
 b15oa0022as1n02x5 U4770 (.a(net485),
    .b(net202),
    .c(n3595),
    .d(u_gpio_reg2hw[220]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[28]));
 b15inv020ar1n08x5 U4771 (.a(net441),
    .o1(n3436));
 b15nand02as1n06x5 U4772 (.a(net325),
    .b(net2042),
    .o1(n3435));
 b15oai012as1n24x5 U4773 (.a(n3435),
    .b(net325),
    .c(n3436),
    .o1(u_gpio_u_reg_u_data_in_wr_data[4]));
 b15inv000al1n02x5 U4774 (.a(u_gpio_u_reg_u_data_in_wr_data[4]),
    .o1(n3437));
 b15aoai13al1n08x5 U4775 (.a(n3437),
    .b(u_gpio_reg2hw[36]),
    .c(u_gpio_reg2hw[100]),
    .d(u_gpio_data_in_q[4]),
    .o1(n3440));
 b15inv000al1n02x5 U4776 (.a(u_gpio_data_in_q[4]),
    .o1(n3438));
 b15aoai13aq1n06x5 U4777 (.a(u_gpio_u_reg_u_data_in_wr_data[4]),
    .b(u_gpio_reg2hw[68]),
    .c(u_gpio_reg2hw[132]),
    .d(n3438),
    .o1(n3439));
 b15oai112as1n16x5 U4778 (.a(n3440),
    .b(n3439),
    .c(net181),
    .d(net463),
    .o1(n3606));
 b15oa0022as1n02x5 U4779 (.a(net462),
    .b(net201),
    .c(n3606),
    .d(u_gpio_reg2hw[196]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[4]));
 b15inv000as1n08x5 U4780 (.a(net450),
    .o1(n3442));
 b15nand02an1n16x5 U4781 (.a(net350),
    .b(u_gpio_gen_filter_15__u_filter_stored_value_q),
    .o1(n3441));
 b15oai012as1n48x5 U4782 (.a(n3441),
    .b(net349),
    .c(n3442),
    .o1(u_gpio_u_reg_u_data_in_wr_data[15]));
 b15inv000al1n02x5 U4783 (.a(u_gpio_u_reg_u_data_in_wr_data[15]),
    .o1(n3443));
 b15aoai13as1n04x5 U4784 (.a(n3443),
    .b(u_gpio_reg2hw[47]),
    .c(net313),
    .d(net2024),
    .o1(n3446));
 b15inv000al1n02x5 U4785 (.a(u_gpio_data_in_q[15]),
    .o1(n3444));
 b15aoai13aq1n06x5 U4786 (.a(u_gpio_u_reg_u_data_in_wr_data[15]),
    .b(net309),
    .c(net289),
    .d(n3444),
    .o1(n3445));
 b15oai112as1n16x5 U4787 (.a(n3446),
    .b(n3445),
    .c(net181),
    .d(n3555),
    .o1(n3570));
 b15oa0022ah1n02x5 U4788 (.a(n3555),
    .b(net201),
    .c(n3570),
    .d(u_gpio_reg2hw[207]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[15]));
 b15inv000al1n02x5 U4789 (.a(u_gpio_gen_filter_9__u_filter_filter_synced),
    .o1(n3448));
 b15nand02al1n02x5 U4790 (.a(net318),
    .b(u_gpio_gen_filter_9__u_filter_stored_value_q),
    .o1(n3447));
 b15oai012al1n06x5 U4791 (.a(n3447),
    .b(net318),
    .c(n3448),
    .o1(u_gpio_u_reg_u_data_in_wr_data[9]));
 b15inv040al1n02x5 U4792 (.a(net239),
    .o1(n3449));
 b15aoai13as1n08x5 U4793 (.a(n3449),
    .b(u_gpio_reg2hw[41]),
    .c(u_gpio_reg2hw[105]),
    .d(net2155),
    .o1(n3452));
 b15inv040ar1n03x5 U4794 (.a(u_gpio_data_in_q[9]),
    .o1(n3450));
 b15aoai13as1n06x5 U4795 (.a(net239),
    .b(net299),
    .c(u_gpio_reg2hw[137]),
    .d(n3450),
    .o1(n3451));
 b15oai112as1n16x5 U4796 (.a(n3452),
    .b(n3451),
    .c(net181),
    .d(net468),
    .o1(n3586));
 b15oa0022al1n04x5 U4797 (.a(net469),
    .b(net201),
    .c(n3586),
    .d(u_gpio_reg2hw[201]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[9]));
 b15inv040an1n05x5 U4798 (.a(net442),
    .o1(n3455));
 b15nandp2al1n08x5 U4799 (.a(net336),
    .b(u_gpio_gen_filter_24__u_filter_stored_value_q),
    .o1(n3454));
 b15oai012al1n32x5 U4800 (.a(n3454),
    .b(net337),
    .c(n3455),
    .o1(u_gpio_u_reg_u_data_in_wr_data[24]));
 b15inv040al1n02x5 U4801 (.a(u_gpio_u_reg_u_data_in_wr_data[24]),
    .o1(n3456));
 b15aoai13as1n08x5 U4802 (.a(n3456),
    .b(u_gpio_reg2hw[56]),
    .c(u_gpio_reg2hw[120]),
    .d(net1951),
    .o1(n3459));
 b15inv020as1n03x5 U4803 (.a(net1951),
    .o1(n3457));
 b15aoai13as1n08x5 U4804 (.a(u_gpio_u_reg_u_data_in_wr_data[24]),
    .b(u_gpio_reg2hw[88]),
    .c(u_gpio_reg2hw[152]),
    .d(n3457),
    .o1(n3458));
 b15oai112ah1n16x5 U4805 (.a(n3459),
    .b(n3458),
    .c(net180),
    .d(n3899),
    .o1(n3596));
 b15oa0022aq1n02x5 U4806 (.a(n3899),
    .b(net202),
    .c(n3596),
    .d(u_gpio_reg2hw[216]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[24]));
 b15nand02al1n12x5 U4807 (.a(net334),
    .b(net2149),
    .o1(n3460));
 b15oai012an1n32x5 U4808 (.a(n3460),
    .b(net334),
    .c(n3461),
    .o1(u_gpio_u_reg_u_data_in_wr_data[27]));
 b15inv040al1n02x5 U4809 (.a(u_gpio_u_reg_u_data_in_wr_data[27]),
    .o1(n3462));
 b15aoai13al1n08x5 U4810 (.a(n3462),
    .b(net292),
    .c(u_gpio_reg2hw[123]),
    .d(net2176),
    .o1(n3465));
 b15inv020ah1n03x5 U4811 (.a(u_gpio_data_in_q[27]),
    .o1(n3463));
 b15aoai13ar1n08x5 U4812 (.a(u_gpio_u_reg_u_data_in_wr_data[27]),
    .b(u_gpio_reg2hw[91]),
    .c(u_gpio_reg2hw[155]),
    .d(n3463),
    .o1(n3464));
 b15oai112as1n16x5 U4813 (.a(n3465),
    .b(n3464),
    .c(net180),
    .d(n3902),
    .o1(n3572));
 b15oa0022ah1n02x5 U4814 (.a(n3902),
    .b(net202),
    .c(n3572),
    .d(u_gpio_reg2hw[219]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[27]));
 b15inv000ah1n05x5 U4815 (.a(net448),
    .o1(n3467));
 b15nandp2al1n08x5 U4816 (.a(net346),
    .b(u_gpio_gen_filter_18__u_filter_stored_value_q),
    .o1(n3466));
 b15oai012an1n32x5 U4817 (.a(n3466),
    .b(net346),
    .c(n3467),
    .o1(u_gpio_u_reg_u_data_in_wr_data[18]));
 b15inv040al1n02x5 U4818 (.a(u_gpio_u_reg_u_data_in_wr_data[18]),
    .o1(n3468));
 b15aoai13as1n06x5 U4819 (.a(n3468),
    .b(u_gpio_reg2hw[50]),
    .c(u_gpio_reg2hw[114]),
    .d(net2060),
    .o1(n3471));
 b15inv040al1n02x5 U4820 (.a(u_gpio_data_in_q[18]),
    .o1(n3469));
 b15aoai13as1n04x5 U4821 (.a(u_gpio_u_reg_u_data_in_wr_data[18]),
    .b(net306),
    .c(u_gpio_reg2hw[146]),
    .d(n3469),
    .o1(n3470));
 b15oai112as1n16x5 U4822 (.a(n3471),
    .b(n3470),
    .c(net180),
    .d(n3893),
    .o1(n3584));
 b15oa0022ar1n03x5 U4823 (.a(n3893),
    .b(net202),
    .c(n3584),
    .d(u_gpio_reg2hw[210]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[18]));
 b15inv040aq1n05x5 U4824 (.a(u_gpio_gen_filter_25__u_filter_filter_synced),
    .o1(n3473));
 b15qgbna2an1n10x5 U4825 (.a(net335),
    .b(u_gpio_gen_filter_25__u_filter_stored_value_q),
    .o1(n3472));
 b15oai012as1n32x5 U4826 (.a(n3472),
    .b(net335),
    .c(n3473),
    .o1(u_gpio_u_reg_u_data_in_wr_data[25]));
 b15inv000al1n02x5 U4827 (.a(u_gpio_u_reg_u_data_in_wr_data[25]),
    .o1(n3474));
 b15aoai13as1n06x5 U4828 (.a(n3474),
    .b(u_gpio_reg2hw[57]),
    .c(u_gpio_reg2hw[121]),
    .d(net1980),
    .o1(n3477));
 b15inv000as1n02x5 U4829 (.a(u_gpio_data_in_q[25]),
    .o1(n3475));
 b15aoai13ah1n06x5 U4830 (.a(u_gpio_u_reg_u_data_in_wr_data[25]),
    .b(u_gpio_reg2hw[89]),
    .c(u_gpio_reg2hw[153]),
    .d(n3475),
    .o1(n3476));
 b15oai112as1n16x5 U4831 (.a(n3477),
    .b(n3476),
    .c(net180),
    .d(n3900),
    .o1(n3589));
 b15oa0022aq1n02x5 U4832 (.a(n3900),
    .b(net202),
    .c(net1981),
    .d(u_gpio_reg2hw[217]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[25]));
 b15inv040as1n10x5 U4833 (.a(net447),
    .o1(n3479));
 b15nand02ah1n12x5 U4834 (.a(net345),
    .b(u_gpio_gen_filter_19__u_filter_stored_value_q),
    .o1(n3478));
 b15oai012aq1n48x5 U4835 (.a(n3478),
    .b(net345),
    .c(n3479),
    .o1(u_gpio_u_reg_u_data_in_wr_data[19]));
 b15inv040al1n02x5 U4836 (.a(u_gpio_u_reg_u_data_in_wr_data[19]),
    .o1(n3480));
 b15aoai13as1n08x5 U4837 (.a(n3480),
    .b(u_gpio_reg2hw[51]),
    .c(u_gpio_reg2hw[115]),
    .d(net2137),
    .o1(n3483));
 b15inv040al1n04x5 U4838 (.a(u_gpio_data_in_q[19]),
    .o1(n3481));
 b15aoai13an1n06x5 U4839 (.a(u_gpio_u_reg_u_data_in_wr_data[19]),
    .b(u_gpio_reg2hw[83]),
    .c(u_gpio_reg2hw[147]),
    .d(n3481),
    .o1(n3482));
 b15oai112as1n16x5 U4840 (.a(n3483),
    .b(n3482),
    .c(net180),
    .d(n3894),
    .o1(n3585));
 b15oa0022ar1n03x5 U4841 (.a(n3894),
    .b(net202),
    .c(n3585),
    .d(u_gpio_reg2hw[211]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[19]));
 b15inv020an1n06x5 U4842 (.a(u_gpio_gen_filter_29__u_filter_filter_synced),
    .o1(n3485));
 b15nand02an1n08x5 U4843 (.a(u_gpio_reg2hw[29]),
    .b(u_gpio_gen_filter_29__u_filter_stored_value_q),
    .o1(n3484));
 b15oai012as1n24x5 U4844 (.a(n3484),
    .b(u_gpio_reg2hw[29]),
    .c(n3485),
    .o1(u_gpio_u_reg_u_data_in_wr_data[29]));
 b15inv000al1n02x5 U4845 (.a(u_gpio_u_reg_u_data_in_wr_data[29]),
    .o1(n3486));
 b15aoai13an1n08x5 U4846 (.a(n3486),
    .b(u_gpio_reg2hw[61]),
    .c(u_gpio_reg2hw[125]),
    .d(net1965),
    .o1(n3489));
 b15inv000al1n03x5 U4847 (.a(u_gpio_data_in_q[29]),
    .o1(n3487));
 b15aoai13an1n08x5 U4848 (.a(u_gpio_u_reg_u_data_in_wr_data[29]),
    .b(u_gpio_reg2hw[93]),
    .c(u_gpio_reg2hw[157]),
    .d(n3487),
    .o1(n3488));
 b15oai112as1n16x5 U4849 (.a(n3489),
    .b(n3488),
    .c(net180),
    .d(n3904),
    .o1(n3593));
 b15oa0022ah1n02x5 U4850 (.a(n3904),
    .b(net202),
    .c(net1966),
    .d(u_gpio_reg2hw[221]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[29]));
 b15nand02al1n12x5 U4851 (.a(u_gpio_reg2hw[26]),
    .b(net2145),
    .o1(n3490));
 b15oai012aq1n32x5 U4852 (.a(n3490),
    .b(u_gpio_reg2hw[26]),
    .c(n3491),
    .o1(u_gpio_u_reg_u_data_in_wr_data[26]));
 b15inv000aq1n03x5 U4853 (.a(u_gpio_u_reg_u_data_in_wr_data[26]),
    .o1(n3492));
 b15aoai13an1n08x5 U4854 (.a(n3492),
    .b(u_gpio_reg2hw[58]),
    .c(net312),
    .d(net2205),
    .o1(n3495));
 b15inv000as1n02x5 U4855 (.a(u_gpio_data_in_q[26]),
    .o1(n3493));
 b15aoai13an1n08x5 U4856 (.a(u_gpio_u_reg_u_data_in_wr_data[26]),
    .b(u_gpio_reg2hw[90]),
    .c(u_gpio_reg2hw[154]),
    .d(n3493),
    .o1(n3494));
 b15oai112ah1n16x5 U4857 (.a(n3495),
    .b(n3494),
    .c(net180),
    .d(n3901),
    .o1(n3597));
 b15oa0022ar1n03x5 U4858 (.a(n3901),
    .b(net202),
    .c(n3597),
    .d(u_gpio_reg2hw[218]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[26]));
 b15inv000al1n06x5 U4859 (.a(u_gpio_gen_filter_31__u_filter_filter_synced),
    .o1(n3497));
 b15nand02al1n12x5 U4860 (.a(u_gpio_reg2hw[31]),
    .b(net2199),
    .o1(n3496));
 b15oai012aq1n32x5 U4861 (.a(n3496),
    .b(u_gpio_reg2hw[31]),
    .c(n3497),
    .o1(u_gpio_u_reg_u_data_in_wr_data[31]));
 b15inv000al1n02x5 U4862 (.a(u_gpio_u_reg_u_data_in_wr_data[31]),
    .o1(n3498));
 b15aoai13al1n08x5 U4863 (.a(n3498),
    .b(u_gpio_reg2hw[63]),
    .c(u_gpio_reg2hw[127]),
    .d(u_gpio_data_in_q[31]),
    .o1(n3501));
 b15inv040al1n02x5 U4864 (.a(u_gpio_data_in_q[31]),
    .o1(n3499));
 b15aoai13as1n06x5 U4865 (.a(u_gpio_u_reg_u_data_in_wr_data[31]),
    .b(net303),
    .c(u_gpio_reg2hw[159]),
    .d(n3499),
    .o1(n3500));
 b15oai112as1n16x5 U4866 (.a(n3501),
    .b(n3500),
    .c(net180),
    .d(net479),
    .o1(n3578));
 b15oa0022al1n06x5 U4867 (.a(net479),
    .b(n3429),
    .c(n3578),
    .d(u_gpio_reg2hw[223]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[31]));
 b15inv040ar1n02x5 U4868 (.a(u_gpio_gen_filter_17__u_filter_filter_synced),
    .o1(n3504));
 b15nandp2al1n02x5 U4869 (.a(u_gpio_reg2hw[17]),
    .b(u_gpio_gen_filter_17__u_filter_stored_value_q),
    .o1(n3503));
 b15oai012ar1n08x5 U4870 (.a(n3503),
    .b(u_gpio_reg2hw[17]),
    .c(n3504),
    .o1(u_gpio_u_reg_u_data_in_wr_data[17]));
 b15inv000al1n03x5 U4871 (.a(net238),
    .o1(n3505));
 b15aoai13ah1n08x5 U4872 (.a(n3505),
    .b(u_gpio_reg2hw[49]),
    .c(u_gpio_reg2hw[113]),
    .d(net2012),
    .o1(n3508));
 b15inv000al1n05x5 U4873 (.a(u_gpio_data_in_q[17]),
    .o1(n3506));
 b15aoai13as1n04x5 U4874 (.a(net238),
    .b(u_gpio_reg2hw[81]),
    .c(u_gpio_reg2hw[145]),
    .d(n3506),
    .o1(n3507));
 b15oai112as1n16x5 U4875 (.a(n3508),
    .b(n3507),
    .c(net180),
    .d(net497),
    .o1(n3590));
 b15oa0022an1n03x5 U4876 (.a(net497),
    .b(net202),
    .c(net2013),
    .d(u_gpio_reg2hw[209]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[17]));
 b15nand02an1n16x5 U4877 (.a(u_gpio_reg2hw[22]),
    .b(u_gpio_gen_filter_22__u_filter_stored_value_q),
    .o1(n3509));
 b15oai012ah1n48x5 U4878 (.a(n3509),
    .b(net339),
    .c(n3510),
    .o1(u_gpio_u_reg_u_data_in_wr_data[22]));
 b15inv000an1n02x5 U4879 (.a(u_gpio_u_reg_u_data_in_wr_data[22]),
    .o1(n3511));
 b15aoai13as1n08x5 U4880 (.a(n3511),
    .b(u_gpio_reg2hw[54]),
    .c(u_gpio_reg2hw[118]),
    .d(net1969),
    .o1(n3514));
 b15inv040ah1n03x5 U4881 (.a(u_gpio_data_in_q[22]),
    .o1(n3512));
 b15aoai13aq1n04x5 U4882 (.a(u_gpio_u_reg_u_data_in_wr_data[22]),
    .b(u_gpio_reg2hw[86]),
    .c(u_gpio_reg2hw[150]),
    .d(n3512),
    .o1(n3513));
 b15oai112as1n16x5 U4883 (.a(n3514),
    .b(n3513),
    .c(net180),
    .d(net488),
    .o1(n3594));
 b15oa0022as1n02x5 U4884 (.a(net489),
    .b(net202),
    .c(net1970),
    .d(u_gpio_reg2hw[214]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[22]));
 b15nand02ah1n06x5 U4885 (.a(u_gpio_reg2hw[30]),
    .b(net2077),
    .o1(n3515));
 b15oai012aq1n24x5 U4886 (.a(n3515),
    .b(u_gpio_reg2hw[30]),
    .c(n3516),
    .o1(u_gpio_u_reg_u_data_in_wr_data[30]));
 b15inv000al1n02x5 U4887 (.a(u_gpio_u_reg_u_data_in_wr_data[30]),
    .o1(n3517));
 b15aoai13an1n08x5 U4888 (.a(n3517),
    .b(u_gpio_reg2hw[62]),
    .c(u_gpio_reg2hw[126]),
    .d(u_gpio_data_in_q[30]),
    .o1(n3520));
 b15inv020ah1n03x5 U4889 (.a(u_gpio_data_in_q[30]),
    .o1(n3518));
 b15aoai13al1n08x5 U4890 (.a(u_gpio_u_reg_u_data_in_wr_data[30]),
    .b(u_gpio_reg2hw[94]),
    .c(u_gpio_reg2hw[158]),
    .d(n3518),
    .o1(n3519));
 b15oai112as1n16x5 U4891 (.a(n3520),
    .b(n3519),
    .c(net180),
    .d(net481),
    .o1(n3598));
 b15oa0022al1n03x5 U4892 (.a(net481),
    .b(net202),
    .c(n3598),
    .d(net2120),
    .o(u_gpio_u_reg_u_intr_state_wr_data[30]));
 b15inv000aq1n02x5 U4893 (.a(net445),
    .o1(n3522));
 b15nandp2al1n02x5 U4894 (.a(net338),
    .b(u_gpio_gen_filter_23__u_filter_stored_value_q),
    .o1(n3521));
 b15oai012al1n06x5 U4895 (.a(n3521),
    .b(net338),
    .c(n3522),
    .o1(u_gpio_u_reg_u_data_in_wr_data[23]));
 b15inv040as1n02x5 U4896 (.a(u_gpio_data_in_q[23]),
    .o1(n3523));
 b15aoai13ah1n04x5 U4897 (.a(net237),
    .b(net305),
    .c(u_gpio_reg2hw[151]),
    .d(n3523),
    .o1(n3526));
 b15inv040al1n02x5 U4898 (.a(net237),
    .o1(n3524));
 b15aoai13ah1n08x5 U4899 (.a(n3524),
    .b(u_gpio_reg2hw[55]),
    .c(u_gpio_reg2hw[119]),
    .d(net2150),
    .o1(n3525));
 b15oai112as1n16x5 U4900 (.a(n3526),
    .b(n3525),
    .c(net486),
    .d(net180),
    .o1(n3574));
 b15oa0022ar1n03x5 U4901 (.a(net487),
    .b(net202),
    .c(net2151),
    .d(u_gpio_reg2hw[215]),
    .o(u_gpio_u_reg_u_intr_state_wr_data[23]));
 b15nonb02ah1n03x5 U4902 (.a(n3530),
    .b(n3529),
    .out0(u_gpio_u_reg_reg_we_check_14_));
 b15norp02ar1n03x5 U4905 (.a(net481),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[30]));
 b15nor002ah1n02x5 U4906 (.a(n3899),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[24]));
 b15nor002ar1n03x5 U4907 (.a(n3901),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[26]));
 b15nor002aq1n02x5 U4908 (.a(net478),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[31]));
 b15nor002ar1n03x5 U4909 (.a(n3903),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[28]));
 b15norp02aq1n02x5 U4910 (.a(n3900),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[25]));
 b15nor002ar1n03x5 U4911 (.a(n3904),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[29]));
 b15norp02al1n03x5 U4912 (.a(n3902),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[27]));
 b15norp02ar1n04x5 U4914 (.a(n3540),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[7]));
 b15norp02as1n03x5 U4915 (.a(n3541),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[1]));
 b15nor002as1n02x5 U4916 (.a(net474),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[8]));
 b15norp02al1n04x5 U4918 (.a(n3544),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[12]));
 b15norp02al1n04x5 U4919 (.a(net473),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[2]));
 b15norp02an1n04x5 U4920 (.a(n3546),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[0]));
 b15nor002ar1n04x5 U4921 (.a(net467),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[13]));
 b15nor002an1n03x5 U4922 (.a(net460),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[11]));
 b15nor002an1n03x5 U4923 (.a(net470),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[10]));
 b15nor002aq1n03x5 U4924 (.a(net476),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[3]));
 b15nor002ar1n03x5 U4925 (.a(n3551),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[4]));
 b15norp02aq1n03x5 U4926 (.a(net468),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[9]));
 b15nor002ah1n02x5 U4927 (.a(net464),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[5]));
 b15nor002an1n03x5 U4928 (.a(n3554),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[14]));
 b15norp02as1n03x5 U4929 (.a(n3555),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[15]));
 b15norp02al1n04x5 U4930 (.a(n3557),
    .b(net173),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[6]));
 b15nor002ah1n02x5 U4931 (.a(net491),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[21]));
 b15nor002ar1n03x5 U4932 (.a(n3893),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[18]));
 b15nor002ar1n04x5 U4933 (.a(net486),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[23]));
 b15nor002ah1n02x5 U4934 (.a(net492),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[20]));
 b15nor002ah1n02x5 U4935 (.a(net495),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[19]));
 b15norp02al1n03x5 U4936 (.a(net497),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[17]));
 b15nor002an1n03x5 U4937 (.a(net488),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[22]));
 b15nor002an1n02x5 U4938 (.a(net500),
    .b(net174),
    .o1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[16]));
 b15nor004as1n08x5 U4939 (.a(n3570),
    .b(n3569),
    .c(n3568),
    .d(n3567),
    .o1(n3609));
 b15nor004ah1n06x5 U4940 (.a(n3574),
    .b(n3573),
    .c(n3572),
    .d(n3571),
    .o1(n3608));
 b15nor004al1n04x5 U4941 (.a(n3578),
    .b(n3577),
    .c(n3576),
    .d(n3575),
    .o1(n3580));
 b15nand04aq1n06x5 U4942 (.a(n3582),
    .b(n3581),
    .c(n3580),
    .d(net201),
    .o1(n3604));
 b15nor004ah1n03x5 U4943 (.a(n3586),
    .b(n3585),
    .c(n3584),
    .d(n3583),
    .o1(n3602));
 b15nor004an1n02x5 U4944 (.a(n3590),
    .b(n3589),
    .c(n3588),
    .d(n3587),
    .o1(n3601));
 b15nor004al1n03x5 U4945 (.a(n3594),
    .b(n3593),
    .c(n3592),
    .d(n3591),
    .o1(n3600));
 b15nor004as1n12x5 U4946 (.a(n3598),
    .b(n3597),
    .c(n3596),
    .d(n3595),
    .o1(n3599));
 b15nand04as1n06x5 U4947 (.a(n3602),
    .b(n3601),
    .c(n3600),
    .d(n3599),
    .o1(n3603));
 b15nor004aq1n08x5 U4948 (.a(n3606),
    .b(n3605),
    .c(n3604),
    .d(n3603),
    .o1(n3607));
 b15nandp3ah1n16x5 U4949 (.a(n3609),
    .b(n3608),
    .c(n3607),
    .o1(u_gpio_u_reg_u_intr_state_n1));
 b15inv000al1n02x5 U4950 (.a(u_xbar_periph_u_s1n_6_dev_select_t[2]),
    .o1(n3611));
 b15nand03ah1n06x5 U4951 (.a(n3611),
    .b(n3610),
    .c(net1865),
    .o1(n3612));
 b15oai112as1n16x5 U4952 (.a(net1866),
    .b(net8),
    .c(n3614),
    .d(n3613),
    .o1(n3615));
 b15norp02ah1n48x5 U4953 (.a(n3616),
    .b(net1867),
    .o1(net111));
 b15inv040ar1n06x5 U4954 (.a(u_xbar_periph_u_s1n_6_tl_u_i[24]),
    .o1(n3619));
 b15oai022ah1n24x5 U4955 (.a(n3620),
    .b(n3619),
    .c(net1759),
    .d(n3617),
    .o1(net168));
 b15nandp2aq1n24x5 U4956 (.a(net168),
    .b(net2),
    .o1(n3631));
 b15norp02ah1n48x5 U4957 (.a(net111),
    .b(n3631),
    .o1(n3629));
 b15xor002ah1n03x5 U4958 (.a(net2147),
    .b(n3629),
    .out0(n3622));
 b15xor002al1n08x5 U4959 (.a(n3622),
    .b(n3621),
    .out0(u_xbar_periph_u_s1n_6_N68));
 b15rm0023an1n04x5 U4960 (.c(n3623),
    .a(n3629),
    .b(u_xbar_periph_u_s1n_6_num_req_outstanding[7]),
    .carry(n3621),
    .sum(u_xbar_periph_u_s1n_6_N67));
 b15ru0023aq1n08x5 U4961 (.a(n3629),
    .b(u_xbar_periph_u_s1n_6_num_req_outstanding[6]),
    .c(n3624),
    .carry(n3623),
    .sum(u_xbar_periph_u_s1n_6_N66));
 b15ru0023aq1n08x5 U4962 (.a(n3629),
    .b(u_xbar_periph_u_s1n_6_num_req_outstanding[5]),
    .c(n3625),
    .carry(n3624),
    .sum(u_xbar_periph_u_s1n_6_N65));
 b15ru0023as1n06x5 U4963 (.a(n3629),
    .b(net2148),
    .c(n3626),
    .carry(n3625),
    .sum(u_xbar_periph_u_s1n_6_N64));
 b15rm0023al1n06x5 U4964 (.c(n3627),
    .a(n3629),
    .b(u_xbar_periph_u_s1n_6_num_req_outstanding[3]),
    .carry(n3626),
    .sum(u_xbar_periph_u_s1n_6_N63));
 b15ru0023as1n06x5 U4965 (.a(n3629),
    .b(net2160),
    .c(n3628),
    .carry(n3627),
    .sum(u_xbar_periph_u_s1n_6_N62));
 b15ru0023as1n06x5 U4966 (.a(n3629),
    .b(u_xbar_periph_u_s1n_6_num_req_outstanding[1]),
    .c(u_xbar_periph_u_s1n_6_num_req_outstanding[0]),
    .carry(n3628),
    .sum(u_xbar_periph_u_s1n_6_N61));
 b15inv000al1n05x5 U4967 (.a(n3629),
    .o1(n3630));
 b15aob012ah1n24x5 U4968 (.a(n3630),
    .b(net111),
    .c(n3631),
    .out0(u_xbar_periph_u_s1n_6_N59));
 b15aoi022aq1n16x5 U4969 (.a(u_gpio_reg2hw[94]),
    .b(net432),
    .c(u_gpio_reg2hw[158]),
    .d(net253),
    .o1(n3637));
 b15aoi022ar1n16x5 U4970 (.a(u_gpio_reg2hw[30]),
    .b(net427),
    .c(net268),
    .d(u_gpio_u_reg_data_in_qs[30]),
    .o1(n3636));
 b15aoi022ar1n32x5 U4971 (.a(u_gpio_reg2hw[62]),
    .b(net259),
    .c(u_gpio_reg2hw[126]),
    .d(net276),
    .o1(n3635));
 b15aoi022as1n16x5 U4972 (.a(net269),
    .b(net365),
    .c(net421),
    .d(u_gpio_reg2hw[190]),
    .o1(n3632));
 b15aob012aq1n04x5 U4973 (.a(n3632),
    .b(net455),
    .c(net282),
    .out0(n3633));
 b15aoi112as1n08x5 U4974 (.a(net225),
    .b(n3633),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[14]),
    .d(net246),
    .o1(n3634));
 b15nand04as1n16x5 U4975 (.a(n3637),
    .b(n3636),
    .c(n3635),
    .d(n3634),
    .o1(u_gpio_u_reg_u_reg_if_N44));
 b15nor004ar1n08x5 U4976 (.a(n3638),
    .b(net6),
    .c(n1451),
    .d(net5),
    .o1(u_gpio_u_reg_u_reg_if_rd_req));
 b15aoi022ah1n12x5 U4978 (.a(u_gpio_reg2hw[128]),
    .b(net256),
    .c(net242),
    .d(u_gpio_u_reg_masked_oe_lower_data_qs[0]),
    .o1(n3646));
 b15nor002ah1n24x5 U4979 (.a(n3641),
    .b(n3640),
    .o1(n3755));
 b15aoi022as1n06x5 U4980 (.a(net456),
    .b(u_gpio_reg2hw[192]),
    .c(net411),
    .d(net236),
    .o1(n3645));
 b15aoi022an1n12x5 U4981 (.a(u_gpio_reg2hw[64]),
    .b(net433),
    .c(u_gpio_reg2hw[32]),
    .d(net260),
    .o1(n3644));
 b15oabi12as1n24x5 U4982 (.a(net269),
    .b(n3642),
    .c(n3641),
    .out0(n3819));
 b15aoi022as1n48x5 U4983 (.a(net316),
    .b(net278),
    .c(net79),
    .d(net231),
    .o1(n3643));
 b15nand04as1n16x5 U4984 (.a(n3646),
    .b(n3645),
    .c(n3644),
    .d(n3643),
    .o1(n3650));
 b15aoi022ar1n24x5 U4986 (.a(net421),
    .b(u_gpio_reg2hw[160]),
    .c(net265),
    .d(net2203),
    .o1(n3649));
 b15aoi022al1n24x5 U4987 (.a(u_gpio_reg2hw[0]),
    .b(net423),
    .c(net418),
    .d(net383),
    .o1(n3648));
 b15nona23ah1n32x5 U4988 (.a(net222),
    .b(n3650),
    .c(n3649),
    .d(n3648),
    .out0(u_gpio_u_reg_u_reg_if_N14));
 b15aoi022al1n24x5 U4989 (.a(u_gpio_reg2hw[65]),
    .b(net433),
    .c(net417),
    .d(net382),
    .o1(n3654));
 b15aoi022aq1n08x5 U4990 (.a(net421),
    .b(u_gpio_reg2hw[161]),
    .c(net265),
    .d(u_gpio_u_reg_data_in_qs[1]),
    .o1(n3653));
 b15aoi022ah1n32x5 U4991 (.a(u_gpio_reg2hw[33]),
    .b(net260),
    .c(net245),
    .d(u_gpio_u_reg_masked_oe_lower_data_qs[1]),
    .o1(n3652));
 b15aoi022ah1n32x5 U4992 (.a(net407),
    .b(n3755),
    .c(net90),
    .d(net231),
    .o1(n3651));
 b15nand04as1n16x5 U4993 (.a(n3654),
    .b(n3653),
    .c(n3652),
    .d(n3651),
    .o1(n3657));
 b15aoi022as1n32x5 U4994 (.a(u_gpio_reg2hw[129]),
    .b(net256),
    .c(u_gpio_reg2hw[97]),
    .d(net278),
    .o1(n3656));
 b15aoi022ar1n16x5 U4995 (.a(net2141),
    .b(net423),
    .c(net457),
    .d(u_gpio_reg2hw[193]),
    .o1(n3655));
 b15nona23an1n32x5 U4996 (.a(net224),
    .b(n3657),
    .c(n3656),
    .d(n3655),
    .out0(u_gpio_u_reg_u_reg_if_N15));
 b15aoi022ah1n24x5 U4997 (.a(net329),
    .b(net425),
    .c(net455),
    .d(u_gpio_reg2hw[194]),
    .o1(n3661));
 b15aoi022an1n06x5 U4998 (.a(u_gpio_reg2hw[130]),
    .b(net252),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[2]),
    .d(net236),
    .o1(n3660));
 b15aoi022an1n12x5 U4999 (.a(net304),
    .b(net431),
    .c(net415),
    .d(net88),
    .o1(n3659));
 b15aoi022ar1n32x5 U5000 (.a(net243),
    .b(net393),
    .c(net101),
    .d(net232),
    .o1(n3658));
 b15nand04as1n06x5 U5001 (.a(n3661),
    .b(n3660),
    .c(n3659),
    .d(n3658),
    .o1(n3664));
 b15aoi022ah1n04x5 U5002 (.a(u_gpio_reg2hw[98]),
    .b(net277),
    .c(net266),
    .d(net2179),
    .o1(n3663));
 b15aoi022aq1n06x5 U5003 (.a(u_gpio_reg2hw[34]),
    .b(net260),
    .c(net422),
    .d(net285),
    .o1(n3662));
 b15nona23aq1n16x5 U5004 (.a(net223),
    .b(n3664),
    .c(n3663),
    .d(n3662),
    .out0(u_gpio_u_reg_u_reg_if_N16));
 b15aoi022an1n06x5 U5005 (.a(u_gpio_reg2hw[35]),
    .b(net260),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[3]),
    .d(net236),
    .o1(n3670));
 b15aoi022ar1n04x5 U5006 (.a(net243),
    .b(u_gpio_u_reg_masked_oe_lower_data_qs[3]),
    .c(net266),
    .d(net2110),
    .o1(n3669));
 b15aoi022as1n08x5 U5007 (.a(net327),
    .b(net424),
    .c(u_gpio_reg2hw[67]),
    .d(net433),
    .o1(n3668));
 b15aoi022aq1n32x5 U5009 (.a(net104),
    .b(net233),
    .c(net420),
    .d(net283),
    .o1(n3667));
 b15nand04as1n04x5 U5010 (.a(n3670),
    .b(n3669),
    .c(n3668),
    .d(n3667),
    .o1(n3673));
 b15aoi022ah1n06x5 U5011 (.a(u_gpio_reg2hw[99]),
    .b(net277),
    .c(net415),
    .d(net379),
    .o1(n3672));
 b15aoi022as1n04x5 U5012 (.a(u_gpio_reg2hw[131]),
    .b(net252),
    .c(net455),
    .d(u_gpio_reg2hw[195]),
    .o1(n3671));
 b15nona23an1n12x5 U5013 (.a(net223),
    .b(n3673),
    .c(n3672),
    .d(n3671),
    .out0(u_gpio_u_reg_u_reg_if_N17));
 b15aoi022ar1n12x5 U5014 (.a(net457),
    .b(u_gpio_reg2hw[196]),
    .c(net422),
    .d(u_gpio_reg2hw[164]),
    .o1(n3677));
 b15aoi022ar1n04x5 U5015 (.a(u_gpio_reg2hw[36]),
    .b(net260),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[4]),
    .d(net236),
    .o1(n3676));
 b15aoi022ar1n02x5 U5016 (.a(u_gpio_reg2hw[132]),
    .b(net256),
    .c(net266),
    .d(u_gpio_u_reg_data_in_qs[4]),
    .o1(n3675));
 b15aoi022aq1n16x5 U5017 (.a(net415),
    .b(net91),
    .c(net105),
    .d(net232),
    .o1(n3674));
 b15nand04ah1n04x5 U5018 (.a(n3677),
    .b(n3676),
    .c(n3675),
    .d(n3674),
    .o1(n3680));
 b15aoi022ar1n08x5 U5019 (.a(u_gpio_reg2hw[68]),
    .b(net433),
    .c(net243),
    .d(u_gpio_u_reg_masked_oe_lower_data_qs[4]),
    .o1(n3679));
 b15aoi022al1n12x5 U5020 (.a(net326),
    .b(net424),
    .c(u_gpio_reg2hw[100]),
    .d(net278),
    .o1(n3678));
 b15nona23al1n12x5 U5021 (.a(net223),
    .b(n3680),
    .c(n3679),
    .d(n3678),
    .out0(u_gpio_u_reg_u_reg_if_N18));
 b15aoi022al1n02x5 U5022 (.a(u_gpio_reg2hw[69]),
    .b(net433),
    .c(net266),
    .d(u_gpio_u_reg_data_in_qs[5]),
    .o1(n3684));
 b15aoi022an1n24x5 U5023 (.a(net323),
    .b(net425),
    .c(net415),
    .d(net377),
    .o1(n3683));
 b15aoi022al1n04x5 U5024 (.a(u_gpio_reg2hw[37]),
    .b(net260),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[5]),
    .d(net236),
    .o1(n3682));
 b15aoi022al1n32x5 U5025 (.a(net243),
    .b(u_gpio_u_reg_masked_oe_lower_data_qs[5]),
    .c(net106),
    .d(net232),
    .o1(n3681));
 b15nand04aq1n04x5 U5026 (.a(n3684),
    .b(n3683),
    .c(n3682),
    .d(n3681),
    .o1(n3687));
 b15aoi022ah1n08x5 U5027 (.a(net457),
    .b(u_gpio_reg2hw[197]),
    .c(net422),
    .d(u_gpio_reg2hw[165]),
    .o1(n3686));
 b15aoi022aq1n08x5 U5028 (.a(u_gpio_reg2hw[133]),
    .b(net256),
    .c(u_gpio_reg2hw[101]),
    .d(net278),
    .o1(n3685));
 b15nona23al1n16x5 U5029 (.a(net223),
    .b(n3687),
    .c(n3686),
    .d(n3685),
    .out0(u_gpio_u_reg_u_reg_if_N19));
 b15aoi022ar1n02x3 U5030 (.a(u_gpio_reg2hw[134]),
    .b(net257),
    .c(net417),
    .d(net376),
    .o1(n3691));
 b15aoi022ar1n02x3 U5031 (.a(u_gpio_reg2hw[38]),
    .b(net260),
    .c(net421),
    .d(u_gpio_reg2hw[166]),
    .o1(n3690));
 b15aoi022ar1n02x5 U5032 (.a(u_gpio_reg2hw[102]),
    .b(net278),
    .c(net406),
    .d(net236),
    .o1(n3689));
 b15aoi022ah1n16x5 U5033 (.a(net456),
    .b(net281),
    .c(net107),
    .d(net231),
    .o1(n3688));
 b15nand04as1n04x5 U5034 (.a(n3691),
    .b(n3690),
    .c(n3689),
    .d(n3688),
    .o1(n3694));
 b15aoi022ar1n02x5 U5035 (.a(n3760),
    .b(u_gpio_u_reg_masked_oe_lower_data_qs[6]),
    .c(net266),
    .d(u_gpio_u_reg_data_in_qs[6]),
    .o1(n3693));
 b15aoi022an1n02x5 U5036 (.a(net322),
    .b(net424),
    .c(u_gpio_reg2hw[70]),
    .d(net433),
    .o1(n3692));
 b15nona23aq1n05x5 U5037 (.a(net222),
    .b(n3694),
    .c(n3693),
    .d(n3692),
    .out0(u_gpio_u_reg_u_reg_if_N20));
 b15aoi022al1n08x5 U5038 (.a(u_gpio_reg2hw[71]),
    .b(net433),
    .c(net404),
    .d(net236),
    .o1(n3698));
 b15aoi022aq1n08x5 U5039 (.a(u_gpio_reg2hw[135]),
    .b(net257),
    .c(net421),
    .d(u_gpio_reg2hw[167]),
    .o1(n3697));
 b15aoi022an1n04x5 U5040 (.a(net321),
    .b(net424),
    .c(u_gpio_reg2hw[103]),
    .d(net278),
    .o1(n3696));
 b15aoi022al1n48x5 U5041 (.a(net108),
    .b(net231),
    .c(net265),
    .d(net435),
    .o1(n3695));
 b15nand04ah1n08x5 U5042 (.a(n3698),
    .b(n3697),
    .c(n3696),
    .d(n3695),
    .o1(n3701));
 b15aoi022ah1n16x5 U5043 (.a(u_gpio_reg2hw[39]),
    .b(net260),
    .c(net245),
    .d(u_gpio_u_reg_masked_oe_lower_data_qs[7]),
    .o1(n3700));
 b15aoi022an1n16x5 U5044 (.a(net458),
    .b(u_gpio_reg2hw[199]),
    .c(net417),
    .d(net373),
    .o1(n3699));
 b15nona23as1n32x5 U5045 (.a(net223),
    .b(n3701),
    .c(n3700),
    .d(n3699),
    .out0(u_gpio_u_reg_u_reg_if_N21));
 b15aoi022as1n16x5 U5046 (.a(net244),
    .b(u_gpio_u_reg_masked_oe_lower_data_qs[8]),
    .c(net416),
    .d(net371),
    .o1(n3705));
 b15aoi022an1n12x5 U5047 (.a(u_gpio_reg2hw[8]),
    .b(net426),
    .c(net421),
    .d(u_gpio_reg2hw[168]),
    .o1(n3704));
 b15aoi022ah1n24x5 U5048 (.a(u_gpio_reg2hw[136]),
    .b(net256),
    .c(u_gpio_reg2hw[104]),
    .d(net278),
    .o1(n3703));
 b15aoi022al1n48x5 U5049 (.a(net403),
    .b(net234),
    .c(net360),
    .d(net232),
    .o1(n3702));
 b15nand04as1n08x5 U5050 (.a(n3705),
    .b(n3704),
    .c(n3703),
    .d(n3702),
    .o1(n3708));
 b15aoi022as1n32x5 U5051 (.a(net300),
    .b(net433),
    .c(u_gpio_reg2hw[40]),
    .d(net260),
    .o1(n3707));
 b15aoi022as1n12x5 U5052 (.a(net455),
    .b(u_gpio_reg2hw[200]),
    .c(net267),
    .d(net1999),
    .o1(n3706));
 b15nona23aq1n32x5 U5053 (.a(net224),
    .b(n3708),
    .c(n3707),
    .d(n3706),
    .out0(u_gpio_u_reg_u_reg_if_N22));
 b15aoi022al1n04x5 U5054 (.a(u_gpio_reg2hw[137]),
    .b(net255),
    .c(net422),
    .d(u_gpio_reg2hw[169]),
    .o1(n3712));
 b15aoi022aq1n24x5 U5055 (.a(u_gpio_reg2hw[41]),
    .b(net260),
    .c(u_gpio_reg2hw[105]),
    .d(net278),
    .o1(n3711));
 b15aoi022ar1n32x5 U5056 (.a(u_gpio_reg2hw[9]),
    .b(net425),
    .c(net267),
    .d(u_gpio_u_reg_data_in_qs[9]),
    .o1(n3710));
 b15aoi022al1n24x5 U5057 (.a(net244),
    .b(u_gpio_u_reg_masked_oe_lower_data_qs[9]),
    .c(net110),
    .d(net232),
    .o1(n3709));
 b15nand04an1n08x5 U5058 (.a(n3712),
    .b(n3711),
    .c(n3710),
    .d(n3709),
    .o1(n3715));
 b15aoi022ah1n12x5 U5059 (.a(net299),
    .b(n3027),
    .c(net455),
    .d(u_gpio_reg2hw[201]),
    .o1(n3714));
 b15aoi022ah1n48x5 U5060 (.a(net400),
    .b(net234),
    .c(net419),
    .d(net370),
    .o1(n3713));
 b15nona23as1n32x5 U5061 (.a(net223),
    .b(n3715),
    .c(n3714),
    .d(n3713),
    .out0(u_gpio_u_reg_u_reg_if_N23));
 b15aoi022ah1n06x5 U5062 (.a(net291),
    .b(net251),
    .c(net315),
    .d(net275),
    .o1(n3719));
 b15aoi022aq1n06x5 U5063 (.a(net298),
    .b(net260),
    .c(net418),
    .d(net369),
    .o1(n3718));
 b15aoi022aq1n02x5 U5064 (.a(net311),
    .b(net430),
    .c(net399),
    .d(net235),
    .o1(n3717));
 b15aoi022ah1n08x5 U5065 (.a(net80),
    .b(net230),
    .c(net262),
    .d(u_gpio_u_reg_data_in_qs[10]),
    .o1(n3716));
 b15nand04ah1n08x5 U5066 (.a(n3719),
    .b(n3718),
    .c(n3717),
    .d(n3716),
    .o1(n3722));
 b15aoi022aq1n12x5 U5067 (.a(u_gpio_reg2hw[10]),
    .b(net425),
    .c(net421),
    .d(u_gpio_reg2hw[170]),
    .o1(n3721));
 b15aoi022ar1n24x5 U5068 (.a(net455),
    .b(u_gpio_reg2hw[202]),
    .c(net244),
    .d(u_gpio_u_reg_masked_oe_lower_data_qs[10]),
    .o1(n3720));
 b15nona23an1n32x5 U5069 (.a(net224),
    .b(n3722),
    .c(n3721),
    .d(n3720),
    .out0(u_gpio_u_reg_u_reg_if_N24));
 b15aoi022al1n06x5 U5070 (.a(net290),
    .b(net257),
    .c(net314),
    .d(net278),
    .o1(n3727));
 b15aoi022ah1n24x5 U5071 (.a(net397),
    .b(net234),
    .c(net416),
    .d(net368),
    .o1(n3726));
 b15aoi022an1n04x5 U5072 (.a(net421),
    .b(u_gpio_reg2hw[171]),
    .c(net267),
    .d(u_gpio_u_reg_data_in_qs[11]),
    .o1(n3725));
 b15aoi022al1n16x5 U5073 (.a(net244),
    .b(net413),
    .c(net81),
    .d(net230),
    .o1(n3724));
 b15nand04an1n08x5 U5074 (.a(n3727),
    .b(n3726),
    .c(n3725),
    .d(n3724),
    .o1(n3730));
 b15aoi022aq1n12x5 U5075 (.a(u_gpio_reg2hw[11]),
    .b(net426),
    .c(net310),
    .d(net433),
    .o1(n3729));
 b15aoi022ar1n16x5 U5076 (.a(net297),
    .b(net260),
    .c(net455),
    .d(u_gpio_reg2hw[203]),
    .o1(n3728));
 b15nona23aq1n32x5 U5077 (.a(net224),
    .b(n3730),
    .c(n3729),
    .d(n3728),
    .out0(u_gpio_u_reg_u_reg_if_N25));
 b15aoi022an1n16x5 U5078 (.a(net355),
    .b(net424),
    .c(u_gpio_reg2hw[76]),
    .d(net433),
    .o1(n3735));
 b15aoi022as1n48x5 U5079 (.a(net416),
    .b(net99),
    .c(net263),
    .d(net436),
    .o1(n3734));
 b15aoi022aq1n04x5 U5080 (.a(net244),
    .b(u_gpio_u_reg_masked_oe_lower_data_qs[12]),
    .c(net422),
    .d(u_gpio_reg2hw[172]),
    .o1(n3733));
 b15aoi022al1n24x5 U5081 (.a(net395),
    .b(net235),
    .c(net387),
    .d(net230),
    .o1(n3732));
 b15nand04al1n12x5 U5082 (.a(n3735),
    .b(n3734),
    .c(n3733),
    .d(n3732),
    .o1(n3738));
 b15aoi022ah1n24x5 U5083 (.a(u_gpio_reg2hw[140]),
    .b(net256),
    .c(u_gpio_reg2hw[108]),
    .d(net278),
    .o1(n3737));
 b15aoi022as1n12x5 U5084 (.a(net296),
    .b(net260),
    .c(net457),
    .d(u_gpio_reg2hw[204]),
    .o1(n3736));
 b15nona23as1n32x5 U5085 (.a(net223),
    .b(n3738),
    .c(n3737),
    .d(n3736),
    .out0(u_gpio_u_reg_u_reg_if_N26));
 b15aoi022al1n12x5 U5086 (.a(net295),
    .b(net259),
    .c(net415),
    .d(net367),
    .o1(n3742));
 b15aoi022as1n32x5 U5087 (.a(u_gpio_reg2hw[109]),
    .b(net278),
    .c(net266),
    .d(u_gpio_u_reg_data_in_qs[13]),
    .o1(n3741));
 b15aoi022ar1n12x5 U5088 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[13]),
    .b(net234),
    .c(net420),
    .d(u_gpio_reg2hw[173]),
    .o1(n3740));
 b15aoi022ah1n12x5 U5089 (.a(net458),
    .b(u_gpio_reg2hw[205]),
    .c(net83),
    .d(net230),
    .o1(n3739));
 b15nand04as1n16x5 U5090 (.a(n3742),
    .b(n3741),
    .c(n3740),
    .d(n3739),
    .o1(n3746));
 b15aoi022al1n32x5 U5091 (.a(net353),
    .b(net424),
    .c(u_gpio_reg2hw[77]),
    .d(net433),
    .o1(n3745));
 b15aoi022al1n24x5 U5092 (.a(u_gpio_reg2hw[141]),
    .b(net255),
    .c(net244),
    .d(u_gpio_u_reg_masked_oe_lower_data_qs[13]),
    .o1(n3744));
 b15nona23as1n32x5 U5093 (.a(net223),
    .b(n3746),
    .c(n3745),
    .d(n3744),
    .out0(u_gpio_u_reg_u_reg_if_N27));
 b15aoi022as1n06x5 U5094 (.a(u_gpio_reg2hw[110]),
    .b(net278),
    .c(net245),
    .d(u_gpio_u_reg_masked_oe_lower_data_qs[14]),
    .o1(n3750));
 b15aoi022al1n04x5 U5095 (.a(net421),
    .b(u_gpio_reg2hw[174]),
    .c(net267),
    .d(u_gpio_u_reg_data_in_qs[14]),
    .o1(n3749));
 b15aoi022an1n04x5 U5096 (.a(u_gpio_reg2hw[142]),
    .b(net257),
    .c(net392),
    .d(net235),
    .o1(n3748));
 b15aoi022aq1n48x5 U5097 (.a(net414),
    .b(net364),
    .c(net84),
    .d(net231),
    .o1(n3747));
 b15nand04aq1n08x5 U5098 (.a(n3750),
    .b(n3749),
    .c(n3748),
    .d(n3747),
    .o1(n3754));
 b15aoi022an1n24x5 U5099 (.a(u_gpio_reg2hw[78]),
    .b(net433),
    .c(u_gpio_reg2hw[46]),
    .d(net260),
    .o1(n3753));
 b15aoi022ar1n24x5 U5100 (.a(net352),
    .b(net424),
    .c(net457),
    .d(u_gpio_reg2hw[206]),
    .o1(n3752));
 b15nona23ah1n32x5 U5101 (.a(net224),
    .b(n3754),
    .c(n3753),
    .d(n3752),
    .out0(u_gpio_u_reg_u_reg_if_N28));
 b15aoi022ar1n08x5 U5102 (.a(net313),
    .b(net278),
    .c(net421),
    .d(u_gpio_reg2hw[175]),
    .o1(n3759));
 b15aoi022an1n06x5 U5103 (.a(net2181),
    .b(net423),
    .c(net457),
    .d(u_gpio_reg2hw[207]),
    .o1(n3758));
 b15aoi022al1n16x5 U5104 (.a(u_gpio_reg2hw[47]),
    .b(net260),
    .c(net391),
    .d(net235),
    .o1(n3757));
 b15aoi022as1n32x5 U5105 (.a(net85),
    .b(net231),
    .c(net265),
    .d(net438),
    .o1(n3756));
 b15nand04aq1n16x5 U5106 (.a(n3759),
    .b(n3758),
    .c(n3757),
    .d(n3756),
    .o1(n3764));
 b15aoi022al1n48x5 U5107 (.a(net309),
    .b(net433),
    .c(net245),
    .d(u_gpio_u_reg_masked_oe_lower_data_qs[15]),
    .o1(n3763));
 b15aoi022aq1n48x5 U5108 (.a(net287),
    .b(net254),
    .c(net418),
    .d(net103),
    .o1(n3762));
 b15nona23al1n32x5 U5109 (.a(net224),
    .b(n3764),
    .c(n3763),
    .d(n3762),
    .out0(u_gpio_u_reg_u_reg_if_N29));
 b15aoi022ah1n04x5 U5110 (.a(net344),
    .b(net425),
    .c(u_gpio_u_reg_masked_oe_upper_data_qs[3]),
    .d(net247),
    .o1(n3772));
 b15aoi022as1n06x5 U5111 (.a(u_gpio_reg2hw[147]),
    .b(net252),
    .c(net420),
    .d(u_gpio_reg2hw[179]),
    .o1(n3771));
 b15aoi022as1n04x5 U5112 (.a(u_gpio_reg2hw[83]),
    .b(net431),
    .c(net264),
    .d(net2206),
    .o1(n3770));
 b15aoi022ar1n04x5 U5113 (.a(u_gpio_reg2hw[115]),
    .b(net277),
    .c(net272),
    .d(net380),
    .o1(n3767));
 b15aob012ar1n06x5 U5114 (.a(n3767),
    .b(net458),
    .c(u_gpio_reg2hw[211]),
    .out0(n3768));
 b15aoi112aq1n08x5 U5115 (.a(net225),
    .b(n3768),
    .c(u_gpio_reg2hw[51]),
    .d(net259),
    .o1(n3769));
 b15nand04ah1n12x5 U5116 (.a(n3772),
    .b(n3771),
    .c(n3770),
    .d(n3769),
    .o1(u_gpio_u_reg_u_reg_if_N33));
 b15aoi022aq1n12x5 U5117 (.a(u_gpio_reg2hw[154]),
    .b(net255),
    .c(u_gpio_reg2hw[58]),
    .d(net259),
    .o1(n3780));
 b15aoi022as1n06x5 U5118 (.a(u_gpio_reg2hw[90]),
    .b(net430),
    .c(net420),
    .d(u_gpio_reg2hw[186]),
    .o1(n3779));
 b15aoi022ah1n08x5 U5119 (.a(net398),
    .b(net246),
    .c(net263),
    .d(net2161),
    .o1(n3778));
 b15aoi022ar1n02x5 U5120 (.a(net312),
    .b(net279),
    .c(net270),
    .d(net369),
    .o1(n3773));
 b15aob012an1n03x5 U5121 (.a(n3773),
    .b(net455),
    .c(u_gpio_reg2hw[218]),
    .out0(n3774));
 b15aoi112aq1n06x5 U5122 (.a(net225),
    .b(n3774),
    .c(u_gpio_reg2hw[26]),
    .d(net427),
    .o1(n3777));
 b15nand04as1n16x5 U5123 (.a(n3780),
    .b(n3779),
    .c(n3778),
    .d(n3777),
    .o1(u_gpio_u_reg_u_reg_if_N40));
 b15aoi022as1n08x5 U5124 (.a(u_gpio_reg2hw[156]),
    .b(net253),
    .c(net459),
    .d(u_gpio_reg2hw[220]),
    .o1(n3790));
 b15aoi022aq1n16x5 U5125 (.a(u_gpio_reg2hw[28]),
    .b(net427),
    .c(net263),
    .d(u_gpio_u_reg_data_in_qs[28]),
    .o1(n3789));
 b15aoi022ah1n08x5 U5126 (.a(u_gpio_reg2hw[92]),
    .b(net432),
    .c(net394),
    .d(net246),
    .o1(n3788));
 b15aoi022al1n32x5 U5127 (.a(u_gpio_reg2hw[124]),
    .b(net276),
    .c(net420),
    .d(net286),
    .o1(n3784));
 b15aob012an1n16x5 U5128 (.a(n3784),
    .b(net270),
    .c(net99),
    .out0(n3785));
 b15aoi112al1n08x5 U5129 (.a(net225),
    .b(n3785),
    .c(u_gpio_reg2hw[60]),
    .d(net261),
    .o1(n3787));
 b15nand04as1n16x5 U5130 (.a(n3790),
    .b(n3789),
    .c(n3788),
    .d(n3787),
    .o1(u_gpio_u_reg_u_reg_if_N42));
 b15aoi022ar1n12x5 U5131 (.a(u_gpio_reg2hw[157]),
    .b(net253),
    .c(net263),
    .d(net2209),
    .o1(n3807));
 b15aoi022as1n06x5 U5132 (.a(net331),
    .b(net427),
    .c(u_gpio_reg2hw[125]),
    .d(net276),
    .o1(n3806));
 b15aoi022an1n12x5 U5133 (.a(u_gpio_reg2hw[61]),
    .b(net259),
    .c(net420),
    .d(u_gpio_reg2hw[189]),
    .o1(n3805));
 b15aoi022an1n16x5 U5134 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[13]),
    .b(net246),
    .c(net272),
    .d(net367),
    .o1(n3799));
 b15aob012ar1n08x5 U5135 (.a(n3799),
    .b(net455),
    .c(u_gpio_reg2hw[221]),
    .out0(n3801));
 b15aoi112al1n08x5 U5136 (.a(net225),
    .b(n3801),
    .c(u_gpio_reg2hw[93]),
    .d(net432),
    .o1(n3804));
 b15nand04as1n16x5 U5137 (.a(n3807),
    .b(n3806),
    .c(n3805),
    .d(n3804),
    .o1(u_gpio_u_reg_u_reg_if_N43));
 b15nor004al1n04x5 U5138 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .b(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .c(u_gpio_gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .d(n3808),
    .o1(n3810));
 b15nor003an1n03x5 U5139 (.a(n3811),
    .b(n3810),
    .c(n3809),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_ping_set_d));
 b15oab012al1n03x5 U5142 (.a(n3812),
    .b(u_gpio_gen_filter_7__u_filter_diff_ctr_q[3]),
    .c(n3813),
    .out0(u_gpio_gen_filter_7__u_filter_diff_ctr_d[2]));
 b15nano23al1n06x5 U5143 (.a(u_gpio_gen_filter_15__u_filter_diff_ctr_q[2]),
    .b(u_gpio_gen_filter_15__u_filter_diff_ctr_d[0]),
    .c(n3815),
    .d(n3814),
    .out0(eq_x_156_n25));
 b15oab012ah1n03x5 U5144 (.a(n3816),
    .b(u_gpio_gen_filter_27__u_filter_diff_ctr_q[3]),
    .c(n3817),
    .out0(u_gpio_gen_filter_27__u_filter_diff_ctr_d[2]));
 b15nonb02ah1n12x5 U5145 (.a(net230),
    .b(n3818),
    .out0(u_gpio_N38));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_0__u_gpio_cio_gpio_en_q_reg_1_ (.rb(net513),
    .clk(clknet_1_0__leaf_u_gpio_net3604),
    .d1(u_gpio_N114),
    .d2(u_gpio_N115),
    .o1(u_gpio_u_reg_masked_oe_lower_data_qs[0]),
    .o2(u_gpio_u_reg_masked_oe_lower_data_qs[1]),
    .si1(net543),
    .si2(net544),
    .ssb(net1349));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_10__u_gpio_cio_gpio_en_q_reg_11_ (.rb(net513),
    .clk(clknet_1_0__leaf_u_gpio_net3604),
    .d1(u_gpio_N124),
    .d2(u_gpio_N125),
    .o1(u_gpio_u_reg_masked_oe_lower_data_qs[10]),
    .o2(u_gpio_u_reg_masked_oe_lower_data_qs[11]),
    .si1(net545),
    .si2(net546),
    .ssb(net1350));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_12__u_gpio_cio_gpio_en_q_reg_13_ (.rb(net513),
    .clk(clknet_1_1__leaf_u_gpio_net3604),
    .d1(u_gpio_N126),
    .d2(u_gpio_N127),
    .o1(u_gpio_u_reg_masked_oe_lower_data_qs[12]),
    .o2(u_gpio_u_reg_masked_oe_lower_data_qs[13]),
    .si1(net547),
    .si2(net548),
    .ssb(net1351));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_14__u_gpio_cio_gpio_en_q_reg_15_ (.rb(net513),
    .clk(clknet_1_0__leaf_u_gpio_net3604),
    .d1(u_gpio_N128),
    .d2(u_gpio_N129),
    .o1(u_gpio_u_reg_masked_oe_lower_data_qs[14]),
    .o2(u_gpio_u_reg_masked_oe_lower_data_qs[15]),
    .si1(net549),
    .si2(net550),
    .ssb(net1352));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_16__u_gpio_cio_gpio_en_q_reg_17_ (.rb(net524),
    .clk(clknet_1_0__leaf_u_gpio_net3599),
    .d1(u_gpio_N131),
    .d2(u_gpio_N132),
    .o1(u_gpio_u_reg_masked_oe_upper_data_qs[0]),
    .o2(u_gpio_u_reg_masked_oe_upper_data_qs[1]),
    .si1(net551),
    .si2(net552),
    .ssb(net1353));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_18__u_gpio_cio_gpio_en_q_reg_19_ (.rb(net524),
    .clk(clknet_1_1__leaf_u_gpio_net3599),
    .d1(u_gpio_N133),
    .d2(u_gpio_N134),
    .o1(u_gpio_u_reg_masked_oe_upper_data_qs[2]),
    .o2(u_gpio_u_reg_masked_oe_upper_data_qs[3]),
    .si1(net553),
    .si2(net554),
    .ssb(net1354));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_20__u_gpio_cio_gpio_en_q_reg_21_ (.rb(net524),
    .clk(clknet_1_0__leaf_u_gpio_net3599),
    .d1(u_gpio_N135),
    .d2(u_gpio_N136),
    .o1(u_gpio_u_reg_masked_oe_upper_data_qs[4]),
    .o2(u_gpio_u_reg_masked_oe_upper_data_qs[5]),
    .si1(net555),
    .si2(net556),
    .ssb(net1355));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_22__u_gpio_cio_gpio_en_q_reg_23_ (.rb(net525),
    .clk(clknet_1_0__leaf_u_gpio_net3599),
    .d1(u_gpio_N137),
    .d2(u_gpio_N138),
    .o1(u_gpio_u_reg_masked_oe_upper_data_qs[6]),
    .o2(u_gpio_u_reg_masked_oe_upper_data_qs[7]),
    .si1(net557),
    .si2(net558),
    .ssb(net1356));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_24__u_gpio_cio_gpio_en_q_reg_25_ (.rb(net525),
    .clk(clknet_1_1__leaf_u_gpio_net3599),
    .d1(u_gpio_N139),
    .d2(u_gpio_N140),
    .o1(u_gpio_u_reg_masked_oe_upper_data_qs[8]),
    .o2(u_gpio_u_reg_masked_oe_upper_data_qs[9]),
    .si1(net559),
    .si2(net560),
    .ssb(net1357));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_26__u_gpio_cio_gpio_en_q_reg_27_ (.rb(net525),
    .clk(clknet_1_1__leaf_u_gpio_net3599),
    .d1(u_gpio_N141),
    .d2(u_gpio_N142),
    .o1(u_gpio_u_reg_masked_oe_upper_data_qs[10]),
    .o2(u_gpio_u_reg_masked_oe_upper_data_qs[11]),
    .si1(net561),
    .si2(net562),
    .ssb(net1358));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_28__u_gpio_cio_gpio_en_q_reg_29_ (.rb(net525),
    .clk(clknet_1_1__leaf_u_gpio_net3599),
    .d1(u_gpio_N143),
    .d2(u_gpio_N144),
    .o1(u_gpio_u_reg_masked_oe_upper_data_qs[12]),
    .o2(u_gpio_u_reg_masked_oe_upper_data_qs[13]),
    .si1(net563),
    .si2(net564),
    .ssb(net1359));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_2__u_gpio_cio_gpio_en_q_reg_3_ (.rb(net513),
    .clk(clknet_1_1__leaf_u_gpio_net3604),
    .d1(u_gpio_N116),
    .d2(u_gpio_N117),
    .o1(u_gpio_u_reg_masked_oe_lower_data_qs[2]),
    .o2(u_gpio_u_reg_masked_oe_lower_data_qs[3]),
    .si1(net565),
    .si2(net566),
    .ssb(net1360));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_30__u_gpio_cio_gpio_en_q_reg_31_ (.rb(net525),
    .clk(clknet_1_0__leaf_u_gpio_net3599),
    .d1(u_gpio_N145),
    .d2(u_gpio_N146),
    .o1(u_gpio_u_reg_masked_oe_upper_data_qs[14]),
    .o2(u_gpio_u_reg_masked_oe_upper_data_qs[15]),
    .si1(net567),
    .si2(net568),
    .ssb(net1361));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_4__u_gpio_cio_gpio_en_q_reg_5_ (.rb(net513),
    .clk(clknet_1_1__leaf_u_gpio_net3604),
    .d1(u_gpio_N118),
    .d2(u_gpio_N119),
    .o1(u_gpio_u_reg_masked_oe_lower_data_qs[4]),
    .o2(u_gpio_u_reg_masked_oe_lower_data_qs[5]),
    .si1(net569),
    .si2(net570),
    .ssb(net1362));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_6__u_gpio_cio_gpio_en_q_reg_7_ (.rb(net513),
    .clk(clknet_1_0__leaf_u_gpio_net3604),
    .d1(u_gpio_N120),
    .d2(u_gpio_N121),
    .o1(u_gpio_u_reg_masked_oe_lower_data_qs[6]),
    .o2(u_gpio_u_reg_masked_oe_lower_data_qs[7]),
    .si1(net571),
    .si2(net572),
    .ssb(net1363));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_en_q_reg_8__u_gpio_cio_gpio_en_q_reg_9_ (.rb(net513),
    .clk(clknet_1_1__leaf_u_gpio_net3604),
    .d1(u_gpio_N122),
    .d2(u_gpio_N123),
    .o1(u_gpio_u_reg_masked_oe_lower_data_qs[8]),
    .o2(u_gpio_u_reg_masked_oe_lower_data_qs[9]),
    .si1(net573),
    .si2(net574),
    .ssb(net1364));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_0__u_gpio_cio_gpio_q_reg_1_ (.rb(net515),
    .clk(clknet_1_0__leaf_u_gpio_net3594),
    .d1(u_gpio_N39),
    .d2(u_gpio_N40),
    .o1(net79),
    .o2(net90),
    .si1(net575),
    .si2(net576),
    .ssb(net1365));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_10__u_gpio_cio_gpio_q_reg_11_ (.rb(net530),
    .clk(clknet_1_1__leaf_u_gpio_net3594),
    .d1(u_gpio_N49),
    .d2(u_gpio_N50),
    .o1(net80),
    .o2(net81),
    .si1(net577),
    .si2(net578),
    .ssb(net1366));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_12__u_gpio_cio_gpio_q_reg_13_ (.rb(net525),
    .clk(clknet_1_0__leaf_u_gpio_net3594),
    .d1(u_gpio_N51),
    .d2(u_gpio_N52),
    .o1(net82),
    .o2(net83),
    .si1(net579),
    .si2(net580),
    .ssb(net1367));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_14__u_gpio_cio_gpio_q_reg_15_ (.rb(net515),
    .clk(clknet_1_0__leaf_u_gpio_net3594),
    .d1(u_gpio_N53),
    .d2(u_gpio_N54),
    .o1(net84),
    .o2(net85),
    .si1(net581),
    .si2(net582),
    .ssb(net1368));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_16__u_gpio_cio_gpio_q_reg_17_ (.rb(net515),
    .clk(clknet_1_0__leaf_u_gpio_net3588),
    .d1(u_gpio_N56),
    .d2(u_gpio_N57),
    .o1(net86),
    .o2(net87),
    .si1(net583),
    .si2(net584),
    .ssb(net1369));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_18__u_gpio_cio_gpio_q_reg_19_ (.rb(net524),
    .clk(clknet_1_1__leaf_u_gpio_net3588),
    .d1(u_gpio_N58),
    .d2(u_gpio_N59),
    .o1(net88),
    .o2(net89),
    .si1(net585),
    .si2(net586),
    .ssb(net1370));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_20__u_gpio_cio_gpio_q_reg_21_ (.rb(net512),
    .clk(clknet_1_0__leaf_u_gpio_net3588),
    .d1(u_gpio_N60),
    .d2(u_gpio_N61),
    .o1(net91),
    .o2(net92),
    .si1(net587),
    .si2(net588),
    .ssb(net1371));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_22__u_gpio_cio_gpio_q_reg_23_ (.rb(net510),
    .clk(clknet_1_0__leaf_u_gpio_net3588),
    .d1(u_gpio_N62),
    .d2(u_gpio_N63),
    .o1(net93),
    .o2(net94),
    .si1(net589),
    .si2(net590),
    .ssb(net1372));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_24__u_gpio_cio_gpio_q_reg_25_ (.rb(net533),
    .clk(clknet_1_1__leaf_u_gpio_net3588),
    .d1(u_gpio_N64),
    .d2(u_gpio_N65),
    .o1(net95),
    .o2(net96),
    .si1(net591),
    .si2(net592),
    .ssb(net1373));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_26__u_gpio_cio_gpio_q_reg_27_ (.rb(net533),
    .clk(clknet_1_1__leaf_u_gpio_net3588),
    .d1(u_gpio_N66),
    .d2(u_gpio_N67),
    .o1(net97),
    .o2(net98),
    .si1(net593),
    .si2(net594),
    .ssb(net1374));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_28__u_gpio_cio_gpio_q_reg_29_ (.rb(net528),
    .clk(clknet_1_1__leaf_u_gpio_net3588),
    .d1(u_gpio_N68),
    .d2(u_gpio_N69),
    .o1(net99),
    .o2(net100),
    .si1(net595),
    .si2(net596),
    .ssb(net1375));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_2__u_gpio_cio_gpio_q_reg_3_ (.rb(net524),
    .clk(clknet_1_1__leaf_u_gpio_net3594),
    .d1(u_gpio_N41),
    .d2(u_gpio_N42),
    .o1(net101),
    .o2(net104),
    .si1(net597),
    .si2(net598),
    .ssb(net1376));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_30__u_gpio_cio_gpio_q_reg_31_ (.rb(net515),
    .clk(clknet_1_0__leaf_u_gpio_net3588),
    .d1(u_gpio_N70),
    .d2(u_gpio_N71),
    .o1(net102),
    .o2(net103),
    .si1(net599),
    .si2(net600),
    .ssb(net1377));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_4__u_gpio_cio_gpio_q_reg_5_ (.rb(net512),
    .clk(clknet_1_1__leaf_u_gpio_net3594),
    .d1(u_gpio_N43),
    .d2(u_gpio_N44),
    .o1(net105),
    .o2(net106),
    .si1(net601),
    .si2(net602),
    .ssb(net1378));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_6__u_gpio_cio_gpio_q_reg_7_ (.rb(net510),
    .clk(clknet_1_0__leaf_u_gpio_net3594),
    .d1(u_gpio_N45),
    .d2(u_gpio_N46),
    .o1(net107),
    .o2(net108),
    .si1(net603),
    .si2(net604),
    .ssb(net1379));
 b15fqy203ar1n02x5 u_gpio_cio_gpio_q_reg_8__u_gpio_cio_gpio_q_reg_9_ (.rb(net524),
    .clk(clknet_1_1__leaf_u_gpio_net3594),
    .d1(u_gpio_N47),
    .d2(u_gpio_N48),
    .o1(net109),
    .o2(net110),
    .si1(net605),
    .si2(net606),
    .ssb(net1380));
 b15cilb05ah1n02x3 u_gpio_clk_gate_cio_gpio_en_q_reg_0_latch (.clk(clknet_leaf_9_clk_i),
    .clkout(u_gpio_net3604),
    .en(u_gpio_N113),
    .te(net607));
 b15cilb05ah1n02x3 u_gpio_clk_gate_cio_gpio_en_q_reg_latch (.clk(clknet_leaf_8_clk_i),
    .clkout(u_gpio_net3599),
    .en(u_gpio_N130),
    .te(net608));
 b15cilb05ah1n02x3 u_gpio_clk_gate_cio_gpio_q_reg_0_latch (.clk(clknet_leaf_2_clk_i),
    .clkout(u_gpio_net3594),
    .en(u_gpio_N38),
    .te(net609));
 b15cilb05ah1n02x3 u_gpio_clk_gate_cio_gpio_q_reg_latch (.clk(clknet_leaf_11_clk_i),
    .clkout(u_gpio_net3588),
    .en(u_gpio_N55),
    .te(net610));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_0__u_gpio_data_in_q_reg_1_ (.clk(clknet_leaf_10_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[0]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[1]),
    .o1(u_gpio_data_in_q[0]),
    .o2(u_gpio_data_in_q[1]),
    .si1(net611),
    .si2(net612),
    .ssb(net1381));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_10__u_gpio_data_in_q_reg_11_ (.clk(clknet_leaf_2_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[10]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[11]),
    .o1(u_gpio_data_in_q[10]),
    .o2(u_gpio_data_in_q[11]),
    .si1(net613),
    .si2(net614),
    .ssb(net1382));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_12__u_gpio_data_in_q_reg_13_ (.clk(clknet_leaf_11_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[12]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[13]),
    .o1(u_gpio_data_in_q[12]),
    .o2(u_gpio_data_in_q[13]),
    .si1(net615),
    .si2(net616),
    .ssb(net1383));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_14__u_gpio_data_in_q_reg_15_ (.clk(clknet_leaf_11_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[14]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[15]),
    .o1(u_gpio_data_in_q[14]),
    .o2(u_gpio_data_in_q[15]),
    .si1(net617),
    .si2(net618),
    .ssb(net1384));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_16__u_gpio_data_in_q_reg_17_ (.clk(clknet_leaf_8_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[16]),
    .d2(net238),
    .o1(u_gpio_data_in_q[16]),
    .o2(u_gpio_data_in_q[17]),
    .si1(net619),
    .si2(net620),
    .ssb(net1385));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_18__u_gpio_data_in_q_reg_19_ (.clk(clknet_leaf_8_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[18]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[19]),
    .o1(u_gpio_data_in_q[18]),
    .o2(u_gpio_data_in_q[19]),
    .si1(net621),
    .si2(net622),
    .ssb(net1386));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_20__u_gpio_data_in_q_reg_21_ (.clk(clknet_leaf_8_clk_i),
    .d1(net240),
    .d2(u_gpio_u_reg_u_data_in_wr_data[21]),
    .o1(u_gpio_data_in_q[20]),
    .o2(u_gpio_data_in_q[21]),
    .si1(net623),
    .si2(net624),
    .ssb(net1387));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_22__u_gpio_data_in_q_reg_23_ (.clk(clknet_leaf_8_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[22]),
    .d2(net237),
    .o1(u_gpio_data_in_q[22]),
    .o2(u_gpio_data_in_q[23]),
    .si1(net625),
    .si2(net626),
    .ssb(net1388));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_24__u_gpio_data_in_q_reg_25_ (.clk(clknet_leaf_7_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[24]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[25]),
    .o1(u_gpio_data_in_q[24]),
    .o2(u_gpio_data_in_q[25]),
    .si1(net627),
    .si2(net628),
    .ssb(net1389));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_26__u_gpio_data_in_q_reg_27_ (.clk(clknet_leaf_6_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[26]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[27]),
    .o1(u_gpio_data_in_q[26]),
    .o2(u_gpio_data_in_q[27]),
    .si1(net629),
    .si2(net630),
    .ssb(net1390));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_28__u_gpio_data_in_q_reg_29_ (.clk(clknet_leaf_7_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[28]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[29]),
    .o1(u_gpio_data_in_q[28]),
    .o2(u_gpio_data_in_q[29]),
    .si1(net631),
    .si2(net632),
    .ssb(net1391));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_2__u_gpio_data_in_q_reg_3_ (.clk(clknet_leaf_9_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[2]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[3]),
    .o1(u_gpio_data_in_q[2]),
    .o2(u_gpio_data_in_q[3]),
    .si1(net633),
    .si2(net634),
    .ssb(net1392));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_30__u_gpio_data_in_q_reg_31_ (.clk(clknet_leaf_6_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[30]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[31]),
    .o1(u_gpio_data_in_q[30]),
    .o2(u_gpio_data_in_q[31]),
    .si1(net635),
    .si2(net636),
    .ssb(net1393));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_4__u_gpio_data_in_q_reg_5_ (.clk(clknet_leaf_10_clk_i),
    .d1(net2043),
    .d2(u_gpio_u_reg_u_data_in_wr_data[5]),
    .o1(u_gpio_data_in_q[4]),
    .o2(u_gpio_data_in_q[5]),
    .si1(net637),
    .si2(net638),
    .ssb(net1394));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_6__u_gpio_data_in_q_reg_7_ (.clk(clknet_leaf_11_clk_i),
    .d1(net241),
    .d2(u_gpio_u_reg_u_data_in_wr_data[7]),
    .o1(u_gpio_data_in_q[6]),
    .o2(u_gpio_data_in_q[7]),
    .si1(net639),
    .si2(net640),
    .ssb(net1395));
 b15fpy200ar1n02x5 u_gpio_data_in_q_reg_8__u_gpio_data_in_q_reg_9_ (.clk(clknet_leaf_9_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[8]),
    .d2(net239),
    .o1(u_gpio_data_in_q[8]),
    .o2(u_gpio_data_in_q[9]),
    .si1(net641),
    .si2(net642),
    .ssb(net1396));
 b15fqy203ar1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_set_q_reg_u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_0_ (.rb(net510),
    .clk(clknet_leaf_10_clk_i),
    .d1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_req_trigger),
    .d2(u_gpio_gen_filter_4__u_filter_diff_ctr_d[0]),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_n1),
    .o2(u_gpio_gen_filter_4__u_filter_diff_ctr_q[0]),
    .si1(net643),
    .si2(net644),
    .ssb(net1397));
 b15fqy203ar1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q_reg_u_gpio_gen_alert_tx_0__u_prim_alert_sender_ping_set_q_reg (.rb(net534),
    .clk(clknet_leaf_5_clk_i),
    .d1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_test_set_d),
    .d2(u_gpio_gen_alert_tx_0__u_prim_alert_sender_ping_set_d),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q),
    .o2(u_gpio_gen_alert_tx_0__u_prim_alert_sender_ping_set_q),
    .si1(net645),
    .si2(net646),
    .ssb(net1398));
 b15fqy203ar1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_0__u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_1_ (.rb(net534),
    .clk(clknet_leaf_5_clk_i),
    .d1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_d[0]),
    .d2(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_d[1]),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .o2(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .si1(net647),
    .si2(net648),
    .ssb(net1399));
 b15fqy203ar1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_2__u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq_reg (.rb(net534),
    .clk(clknet_leaf_5_clk_i),
    .d1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_d[2]),
    .d2(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .o2(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq),
    .si1(net649),
    .si2(net650),
    .ssb(net1400));
 b15fqy00car1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq_reg (.clk(clknet_leaf_5_clk_i),
    .d(net1959),
    .o(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq),
    .psb(net534),
    .si(net651),
    .ssb(net1401));
 b15fqy00car1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.clk(clknet_leaf_7_clk_i),
    .d(net1402),
    .o(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_intq_0_),
    .psb(net528),
    .si(net652),
    .ssb(net1403));
 b15fqy00car1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.clk(clknet_leaf_7_clk_i),
    .d(net1930),
    .o(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nd),
    .psb(net528),
    .si(net653),
    .ssb(net1404));
 b15fqy203ar1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net536),
    .clk(clknet_leaf_5_clk_i),
    .d1(net654),
    .d2(net655),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_intq_0_),
    .o2(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_intq_0_),
    .si1(net656),
    .si2(net657),
    .ssb(net1405));
 b15fqy203ar1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q_reg (.rb(net534),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2108),
    .d2(u_gpio_gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .o2(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q),
    .si1(net658),
    .si2(net659),
    .ssb(net1406));
 b15fqy043ar1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_0_ (.clk(clknet_leaf_6_clk_i),
    .d(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[0]),
    .den(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39),
    .o(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[0]),
    .rb(net528),
    .si(net660),
    .ssb(net1407));
 b15fqy043ar1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_1_ (.clk(clknet_leaf_6_clk_i),
    .d(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[1]),
    .den(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39),
    .o(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[1]),
    .rb(net534),
    .si(net661),
    .ssb(net1408));
 b15fqy00car1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq_reg (.clk(clknet_leaf_5_clk_i),
    .d(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd),
    .o(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq),
    .psb(net536),
    .si(net662),
    .ssb(net1409));
 b15fqy203ar1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq_reg_u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net536),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2069),
    .d2(net1942),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq),
    .o2(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd),
    .si1(net663),
    .si2(net664),
    .ssb(net1410));
 b15fqy00car1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.clk(clknet_leaf_4_clk_i),
    .d(net1411),
    .o(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_intq_0_),
    .psb(net536),
    .si(net665),
    .ssb(net1412));
 b15fqy00car1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.clk(clknet_leaf_4_clk_i),
    .d(net1935),
    .o(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd),
    .psb(net536),
    .si(net666),
    .ssb(net1413));
 b15fqy043ar1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_0_ (.clk(clknet_leaf_5_clk_i),
    .d(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[0]),
    .den(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39),
    .o(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[0]),
    .rb(net536),
    .si(net667),
    .ssb(net1414));
 b15fqy043ar1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_1_ (.clk(clknet_leaf_5_clk_i),
    .d(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[1]),
    .den(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39),
    .o(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .rb(net534),
    .si(net668),
    .ssb(net1415));
 b15fqy203ar1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q_reg_u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_0_ (.rb(net536),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2123),
    .d2(u_gpio_gen_filter_6__u_filter_diff_ctr_d[0]),
    .o1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q),
    .o2(u_gpio_gen_filter_6__u_filter_diff_ctr_q[0]),
    .si1(net669),
    .si2(net670),
    .ssb(net1416));
 b15fqy203ar1n02x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_16__u_filter_filter_q_reg (.rb(net536),
    .clk(clknet_leaf_4_clk_i),
    .d1(u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_pd),
    .d2(u_gpio_gen_filter_16__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_16__u_filter_filter_q),
    .si1(net671),
    .si2(net672),
    .ssb(net1417));
 b15fqy00car1n06x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_1_ (.clk(clknet_leaf_5_clk_i),
    .d(u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_nd),
    .psb(net534),
    .si(net673),
    .ssb(net1418));
 b15fqy203ar1n02x5 u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_1_ (.rb(net517),
    .clk(clknet_leaf_0_clk_i),
    .d1(u_gpio_gen_filter_0__u_filter_diff_ctr_d[0]),
    .d2(u_gpio_gen_filter_0__u_filter_diff_ctr_d[1]),
    .o1(u_gpio_gen_filter_0__u_filter_diff_ctr_q[0]),
    .o2(u_gpio_gen_filter_0__u_filter_diff_ctr_q[1]),
    .si1(net674),
    .si2(net675),
    .ssb(net1419));
 b15fqy203ar1n02x5 u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_3_ (.rb(net521),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2005),
    .d2(net1992),
    .o1(u_gpio_gen_filter_0__u_filter_diff_ctr_q[2]),
    .o2(u_gpio_gen_filter_0__u_filter_diff_ctr_q[3]),
    .si1(net676),
    .si2(net677),
    .ssb(net1420));
 b15fqy203ar1n02x5 u_gpio_gen_filter_0__u_filter_filter_q_reg_u_gpio_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net519),
    .clk(clknet_leaf_2_clk_i),
    .d1(u_gpio_gen_filter_0__u_filter_filter_synced),
    .d2(net2201),
    .o1(u_gpio_gen_filter_0__u_filter_filter_q),
    .o2(u_gpio_gen_filter_0__u_filter_filter_synced),
    .si1(net678),
    .si2(net679),
    .ssb(net1421));
 b15fqy203ar1n02x5 u_gpio_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net519),
    .clk(clknet_leaf_2_clk_i),
    .d1(net680),
    .d2(net681),
    .o1(u_gpio_gen_filter_0__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_1__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net682),
    .si2(net683),
    .ssb(net1422));
 b15fqy043ar1n02x5 u_gpio_gen_filter_0__u_filter_stored_value_q_reg (.clk(clknet_leaf_0_clk_i),
    .d(u_gpio_gen_filter_0__u_filter_filter_synced),
    .den(eq_x_231_n25),
    .o(u_gpio_gen_filter_0__u_filter_stored_value_q),
    .rb(net519),
    .si(net684),
    .ssb(net1423));
 b15fqy203ar1n02x5 u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_1_ (.rb(net531),
    .clk(clknet_leaf_3_clk_i),
    .d1(net2080),
    .d2(net2191),
    .o1(u_gpio_gen_filter_10__u_filter_diff_ctr_q[0]),
    .o2(u_gpio_gen_filter_10__u_filter_diff_ctr_q[1]),
    .si1(net685),
    .si2(net686),
    .ssb(net1424));
 b15fqy203ar1n02x5 u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_10__u_filter_filter_q_reg (.rb(net531),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2165),
    .d2(u_gpio_gen_filter_10__u_filter_filter_synced),
    .o1(u_gpio_gen_filter_10__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_10__u_filter_filter_q),
    .si1(net687),
    .si2(net688),
    .ssb(net1425));
 b15fqy203ar1n02x5 u_gpio_gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net522),
    .clk(clknet_leaf_2_clk_i),
    .d1(net689),
    .d2(net690),
    .o1(u_gpio_gen_filter_10__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_11__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net691),
    .si2(net692),
    .ssb(net1426));
 b15fqy203ar1n02x5 u_gpio_gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_0_ (.rb(net522),
    .clk(clknet_leaf_2_clk_i),
    .d1(net1947),
    .d2(u_gpio_gen_filter_11__u_filter_diff_ctr_d[0]),
    .o1(u_gpio_gen_filter_10__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_11__u_filter_diff_ctr_q[0]),
    .si1(net693),
    .si2(net694),
    .ssb(net1427));
 b15fqy043ar1n02x5 u_gpio_gen_filter_10__u_filter_stored_value_q_reg (.clk(clknet_leaf_2_clk_i),
    .d(u_gpio_gen_filter_10__u_filter_filter_synced),
    .den(eq_x_181_n25),
    .o(u_gpio_gen_filter_10__u_filter_stored_value_q),
    .rb(net529),
    .si(net695),
    .ssb(net1428));
 b15fqy203ar1n02x5 u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_2_ (.rb(net522),
    .clk(clknet_leaf_1_clk_i),
    .d1(u_gpio_gen_filter_11__u_filter_diff_ctr_d[1]),
    .d2(net2015),
    .o1(u_gpio_gen_filter_11__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_11__u_filter_diff_ctr_q[2]),
    .si1(net696),
    .si2(net697),
    .ssb(net1429));
 b15fqy203ar1n02x5 u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_11__u_filter_filter_q_reg (.rb(net521),
    .clk(clknet_leaf_1_clk_i),
    .d1(u_gpio_gen_filter_11__u_filter_diff_ctr_d[3]),
    .d2(u_gpio_gen_filter_11__u_filter_filter_synced),
    .o1(u_gpio_gen_filter_11__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_11__u_filter_filter_q),
    .si1(net698),
    .si2(net699),
    .ssb(net1430));
 b15fqy043ar1n02x5 u_gpio_gen_filter_11__u_filter_stored_value_q_reg (.clk(clknet_leaf_2_clk_i),
    .d(u_gpio_gen_filter_11__u_filter_filter_synced),
    .den(eq_x_176_n25),
    .o(u_gpio_gen_filter_11__u_filter_stored_value_q),
    .rb(net522),
    .si(net700),
    .ssb(net1431));
 b15fqy203ar1n02x5 u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_2_ (.rb(net515),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2066),
    .d2(net2062),
    .o1(u_gpio_gen_filter_12__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_12__u_filter_diff_ctr_q[2]),
    .si1(net701),
    .si2(net702),
    .ssb(net1432));
 b15fqy203ar1n02x5 u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_12__u_filter_filter_q_reg (.rb(net515),
    .clk(clknet_leaf_0_clk_i),
    .d1(u_gpio_gen_filter_12__u_filter_diff_ctr_d[3]),
    .d2(net452),
    .o1(u_gpio_gen_filter_12__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_12__u_filter_filter_q),
    .si1(net703),
    .si2(net704),
    .ssb(net1433));
 b15fqy203ar1n02x5 u_gpio_gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net517),
    .clk(clknet_leaf_0_clk_i),
    .d1(net705),
    .d2(net706),
    .o1(u_gpio_gen_filter_12__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_13__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net707),
    .si2(net708),
    .ssb(net1434));
 b15fqy203ar1n02x5 u_gpio_gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_0_ (.rb(net517),
    .clk(clknet_leaf_1_clk_i),
    .d1(net1989),
    .d2(u_gpio_gen_filter_22__u_filter_diff_ctr_d[0]),
    .o1(u_gpio_gen_filter_12__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_22__u_filter_diff_ctr_q[0]),
    .si1(net709),
    .si2(net710),
    .ssb(net1435));
 b15fqy043ar1n02x5 u_gpio_gen_filter_12__u_filter_stored_value_q_reg (.clk(clknet_leaf_0_clk_i),
    .d(net452),
    .den(eq_x_171_n25),
    .o(u_gpio_gen_filter_12__u_filter_stored_value_q),
    .rb(net515),
    .si(net711),
    .ssb(net1436));
 b15fqy203ar1n02x5 u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_1_ (.rb(net516),
    .clk(clknet_leaf_0_clk_i),
    .d1(u_gpio_gen_filter_13__u_filter_diff_ctr_d[0]),
    .d2(u_gpio_gen_filter_13__u_filter_diff_ctr_d[1]),
    .o1(u_gpio_gen_filter_13__u_filter_diff_ctr_q[0]),
    .o2(u_gpio_gen_filter_13__u_filter_diff_ctr_q[1]),
    .si1(net712),
    .si2(net713),
    .ssb(net1437));
 b15fqy203ar1n02x5 u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_3_ (.rb(net516),
    .clk(clknet_leaf_0_clk_i),
    .d1(u_gpio_gen_filter_13__u_filter_diff_ctr_d[2]),
    .d2(net1997),
    .o1(u_gpio_gen_filter_13__u_filter_diff_ctr_q[2]),
    .o2(u_gpio_gen_filter_13__u_filter_diff_ctr_q[3]),
    .si1(net714),
    .si2(net715),
    .ssb(net1438));
 b15fqy203ar1n02x5 u_gpio_gen_filter_13__u_filter_filter_q_reg_u_gpio_gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net517),
    .clk(clknet_leaf_0_clk_i),
    .d1(u_gpio_gen_filter_13__u_filter_filter_synced),
    .d2(net1937),
    .o1(u_gpio_gen_filter_13__u_filter_filter_q),
    .o2(u_gpio_gen_filter_13__u_filter_filter_synced),
    .si1(net716),
    .si2(net717),
    .ssb(net1439));
 b15fqy043ar1n02x5 u_gpio_gen_filter_13__u_filter_stored_value_q_reg (.clk(clknet_leaf_0_clk_i),
    .d(u_gpio_gen_filter_13__u_filter_filter_synced),
    .den(eq_x_166_n25),
    .o(u_gpio_gen_filter_13__u_filter_stored_value_q),
    .rb(net516),
    .si(net718),
    .ssb(net1440));
 b15fqy203ar1n02x5 u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_2_ (.rb(net515),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2037),
    .d2(u_gpio_gen_filter_14__u_filter_diff_ctr_d[2]),
    .o1(u_gpio_gen_filter_14__u_filter_diff_ctr_q[0]),
    .o2(u_gpio_gen_filter_14__u_filter_diff_ctr_q[2]),
    .si1(net719),
    .si2(net720),
    .ssb(net1441));
 b15fqy203ar1n02x5 u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_0_ (.rb(net515),
    .clk(clknet_leaf_0_clk_i),
    .d1(u_gpio_gen_filter_14__u_filter_diff_ctr_d[1]),
    .d2(net2007),
    .o1(u_gpio_gen_filter_14__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_15__u_filter_diff_ctr_q[0]),
    .si1(net721),
    .si2(net722),
    .ssb(net1442));
 b15fqy203ar1n02x5 u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_14__u_filter_filter_q_reg (.rb(net515),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2168),
    .d2(net2156),
    .o1(u_gpio_gen_filter_14__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_14__u_filter_filter_q),
    .si1(net723),
    .si2(net724),
    .ssb(net1443));
 b15fqy203ar1n02x5 u_gpio_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net516),
    .clk(clknet_leaf_0_clk_i),
    .d1(net725),
    .d2(net726),
    .o1(u_gpio_gen_filter_14__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_15__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net727),
    .si2(net728),
    .ssb(net1444));
 b15fqy203ar1n02x5 u_gpio_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_0_ (.rb(net516),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2105),
    .d2(net2068),
    .o1(u_gpio_gen_filter_14__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_19__u_filter_diff_ctr_q[0]),
    .si1(net729),
    .si2(net730),
    .ssb(net1445));
 b15fqy043ar1n02x5 u_gpio_gen_filter_14__u_filter_stored_value_q_reg (.clk(clknet_leaf_11_clk_i),
    .d(net451),
    .den(eq_x_161_n25),
    .o(u_gpio_gen_filter_14__u_filter_stored_value_q),
    .rb(net515),
    .si(net731),
    .ssb(net1446));
 b15fqy203ar1n02x5 u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_2_ (.rb(net516),
    .clk(clknet_leaf_0_clk_i),
    .d1(u_gpio_gen_filter_15__u_filter_diff_ctr_d[1]),
    .d2(u_gpio_gen_filter_15__u_filter_diff_ctr_d[2]),
    .o1(u_gpio_gen_filter_15__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_15__u_filter_diff_ctr_q[2]),
    .si1(net732),
    .si2(net733),
    .ssb(net1447));
 b15fqy203ar1n02x5 u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_15__u_filter_filter_q_reg (.rb(net515),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2072),
    .d2(net449),
    .o1(u_gpio_gen_filter_15__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_15__u_filter_filter_q),
    .si1(net734),
    .si2(net735),
    .ssb(net1448));
 b15fqy203ar1n02x5 u_gpio_gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_0_ (.rb(net517),
    .clk(clknet_leaf_1_clk_i),
    .d1(net2130),
    .d2(net1972),
    .o1(u_gpio_gen_filter_15__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_23__u_filter_diff_ctr_q[0]),
    .si1(net736),
    .si2(net737),
    .ssb(net1449));
 b15fqy043ar1n02x5 u_gpio_gen_filter_15__u_filter_stored_value_q_reg (.clk(clknet_leaf_0_clk_i),
    .d(net450),
    .den(eq_x_156_n25),
    .o(u_gpio_gen_filter_15__u_filter_stored_value_q),
    .rb(net515),
    .si(net738),
    .ssb(net1450));
 b15fqy203ar1n02x5 u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_1_ (.rb(net536),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2039),
    .d2(net2018),
    .o1(u_gpio_gen_filter_16__u_filter_diff_ctr_q[0]),
    .o2(u_gpio_gen_filter_16__u_filter_diff_ctr_q[1]),
    .si1(net739),
    .si2(net740),
    .ssb(net1451));
 b15fqy203ar1n02x5 u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_3_ (.rb(net536),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2064),
    .d2(u_gpio_gen_filter_16__u_filter_diff_ctr_d[3]),
    .o1(u_gpio_gen_filter_16__u_filter_diff_ctr_q[2]),
    .o2(u_gpio_gen_filter_16__u_filter_diff_ctr_q[3]),
    .si1(net741),
    .si2(net742),
    .ssb(net1452));
 b15fqy203ar1n02x5 u_gpio_gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net535),
    .clk(clknet_leaf_4_clk_i),
    .d1(net743),
    .d2(net744),
    .o1(u_gpio_gen_filter_16__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_17__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net745),
    .si2(net746),
    .ssb(net1453));
 b15fqy203ar1n02x5 u_gpio_gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_0_ (.rb(net535),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2027),
    .d2(u_gpio_gen_filter_20__u_filter_diff_ctr_d[0]),
    .o1(u_gpio_gen_filter_16__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_20__u_filter_diff_ctr_q[0]),
    .si1(net747),
    .si2(net748),
    .ssb(net1454));
 b15fqy043ar1n02x5 u_gpio_gen_filter_16__u_filter_stored_value_q_reg (.clk(clknet_leaf_5_clk_i),
    .d(u_gpio_gen_filter_16__u_filter_filter_synced),
    .den(eq_x_151_n25),
    .o(u_gpio_gen_filter_16__u_filter_stored_value_q),
    .rb(net536),
    .si(net749),
    .ssb(net1455));
 b15fqy203ar1n02x5 u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_2_ (.rb(net532),
    .clk(clknet_leaf_4_clk_i),
    .d1(net1978),
    .d2(net2059),
    .o1(u_gpio_gen_filter_17__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_17__u_filter_diff_ctr_q[2]),
    .si1(net750),
    .si2(net751),
    .ssb(net1456));
 b15fqy203ar1n02x5 u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_17__u_filter_filter_q_reg (.rb(net532),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2091),
    .d2(u_gpio_gen_filter_17__u_filter_filter_synced),
    .o1(u_gpio_gen_filter_17__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_17__u_filter_filter_q),
    .si1(net752),
    .si2(net753),
    .ssb(net1457));
 b15fqy203ar1n02x5 u_gpio_gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_3_ (.rb(net535),
    .clk(clknet_leaf_4_clk_i),
    .d1(net1940),
    .d2(u_gpio_gen_filter_20__u_filter_diff_ctr_d[3]),
    .o1(u_gpio_gen_filter_17__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_20__u_filter_diff_ctr_q[3]),
    .si1(net754),
    .si2(net755),
    .ssb(net1458));
 b15fqy043ar1n02x5 u_gpio_gen_filter_17__u_filter_stored_value_q_reg (.clk(clknet_leaf_4_clk_i),
    .d(u_gpio_gen_filter_17__u_filter_filter_synced),
    .den(eq_x_146_n25),
    .o(u_gpio_gen_filter_17__u_filter_stored_value_q),
    .rb(net532),
    .si(net756),
    .ssb(net1459));
 b15fqy203ar1n02x5 u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_1_ (.rb(net510),
    .clk(clknet_leaf_11_clk_i),
    .d1(net1974),
    .d2(net2001),
    .o1(u_gpio_gen_filter_18__u_filter_diff_ctr_q[0]),
    .o2(u_gpio_gen_filter_18__u_filter_diff_ctr_q[1]),
    .si1(net757),
    .si2(net758),
    .ssb(net1460));
 b15fqy203ar1n02x5 u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_3_ (.rb(net510),
    .clk(clknet_leaf_11_clk_i),
    .d1(u_gpio_gen_filter_18__u_filter_diff_ctr_d[2]),
    .d2(net2026),
    .o1(u_gpio_gen_filter_18__u_filter_diff_ctr_q[2]),
    .o2(u_gpio_gen_filter_18__u_filter_diff_ctr_q[3]),
    .si1(net759),
    .si2(net760),
    .ssb(net1461));
 b15fqy203ar1n02x5 u_gpio_gen_filter_18__u_filter_filter_q_reg_u_gpio_gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net510),
    .clk(clknet_leaf_11_clk_i),
    .d1(u_gpio_gen_filter_18__u_filter_filter_synced),
    .d2(u_gpio_gen_filter_18__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o1(u_gpio_gen_filter_18__u_filter_filter_q),
    .o2(u_gpio_gen_filter_18__u_filter_filter_synced),
    .si1(net761),
    .si2(net762),
    .ssb(net1462));
 b15fqy203ar1n02x5 u_gpio_gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net516),
    .clk(clknet_leaf_0_clk_i),
    .d1(net763),
    .d2(net764),
    .o1(u_gpio_gen_filter_18__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_19__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net765),
    .si2(net766),
    .ssb(net1463));
 b15fqy043ar1n02x5 u_gpio_gen_filter_18__u_filter_stored_value_q_reg (.clk(clknet_leaf_11_clk_i),
    .d(u_gpio_gen_filter_18__u_filter_filter_synced),
    .den(eq_x_141_n25),
    .o(u_gpio_gen_filter_18__u_filter_stored_value_q),
    .rb(net510),
    .si(net767),
    .ssb(net1464));
 b15fqy203ar1n02x5 u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_2_ (.rb(net515),
    .clk(clknet_leaf_0_clk_i),
    .d1(u_gpio_gen_filter_19__u_filter_diff_ctr_d[1]),
    .d2(net2046),
    .o1(u_gpio_gen_filter_19__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_19__u_filter_diff_ctr_q[2]),
    .si1(net768),
    .si2(net769),
    .ssb(net1465));
 b15fqy203ar1n02x5 u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_19__u_filter_filter_q_reg (.rb(net516),
    .clk(clknet_leaf_0_clk_i),
    .d1(u_gpio_gen_filter_19__u_filter_diff_ctr_d[3]),
    .d2(net446),
    .o1(u_gpio_gen_filter_19__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_19__u_filter_filter_q),
    .si1(net770),
    .si2(net771),
    .ssb(net1466));
 b15fqy203ar1n02x5 u_gpio_gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_2_ (.rb(net521),
    .clk(clknet_leaf_1_clk_i),
    .d1(net2152),
    .d2(net1995),
    .o1(u_gpio_gen_filter_19__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_22__u_filter_diff_ctr_q[2]),
    .si1(net772),
    .si2(net773),
    .ssb(net1467));
 b15fqy043ar1n02x5 u_gpio_gen_filter_19__u_filter_stored_value_q_reg (.clk(clknet_leaf_2_clk_i),
    .d(net447),
    .den(eq_x_136_n25),
    .o(u_gpio_gen_filter_19__u_filter_stored_value_q),
    .rb(net521),
    .si(net774),
    .ssb(net1468));
 b15fqy203ar1n02x5 u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_1_ (.rb(net528),
    .clk(clknet_leaf_7_clk_i),
    .d1(u_gpio_gen_filter_1__u_filter_diff_ctr_d[0]),
    .d2(u_gpio_gen_filter_1__u_filter_diff_ctr_d[1]),
    .o1(u_gpio_gen_filter_1__u_filter_diff_ctr_q[0]),
    .o2(u_gpio_gen_filter_1__u_filter_diff_ctr_q[1]),
    .si1(net775),
    .si2(net776),
    .ssb(net1469));
 b15fqy203ar1n02x5 u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_3_ (.rb(net528),
    .clk(clknet_leaf_7_clk_i),
    .d1(u_gpio_gen_filter_1__u_filter_diff_ctr_d[2]),
    .d2(u_gpio_gen_filter_1__u_filter_diff_ctr_d[3]),
    .o1(u_gpio_gen_filter_1__u_filter_diff_ctr_q[2]),
    .o2(u_gpio_gen_filter_1__u_filter_diff_ctr_q[3]),
    .si1(net777),
    .si2(net778),
    .ssb(net1470));
 b15fqy203ar1n02x5 u_gpio_gen_filter_1__u_filter_filter_q_reg_u_gpio_gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net529),
    .clk(clknet_leaf_3_clk_i),
    .d1(u_gpio_gen_filter_1__u_filter_filter_synced),
    .d2(net1962),
    .o1(u_gpio_gen_filter_1__u_filter_filter_q),
    .o2(u_gpio_gen_filter_1__u_filter_filter_synced),
    .si1(net779),
    .si2(net780),
    .ssb(net1471));
 b15fqy043ar1n02x5 u_gpio_gen_filter_1__u_filter_stored_value_q_reg (.clk(clknet_leaf_3_clk_i),
    .d(u_gpio_gen_filter_1__u_filter_filter_synced),
    .den(eq_x_226_n25),
    .o(u_gpio_gen_filter_1__u_filter_stored_value_q),
    .rb(net529),
    .si(net781),
    .ssb(net1472));
 b15fqy203ar1n02x5 u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_2_ (.rb(net535),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2101),
    .d2(u_gpio_gen_filter_20__u_filter_diff_ctr_d[2]),
    .o1(u_gpio_gen_filter_20__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_20__u_filter_diff_ctr_q[2]),
    .si1(net782),
    .si2(net783),
    .ssb(net1473));
 b15fqy203ar1n02x5 u_gpio_gen_filter_20__u_filter_filter_q_reg_u_gpio_gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net535),
    .clk(clknet_leaf_4_clk_i),
    .d1(u_gpio_gen_filter_20__u_filter_filter_synced),
    .d2(net1931),
    .o1(u_gpio_gen_filter_20__u_filter_filter_q),
    .o2(u_gpio_gen_filter_21__u_filter_filter_synced),
    .si1(net784),
    .si2(net785),
    .ssb(net1474));
 b15fqy203ar1n02x5 u_gpio_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net535),
    .clk(clknet_leaf_4_clk_i),
    .d1(net786),
    .d2(net787),
    .o1(u_gpio_gen_filter_20__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_21__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net788),
    .si2(net789),
    .ssb(net1475));
 b15fqy203ar1n02x5 u_gpio_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_0_ (.rb(net535),
    .clk(clknet_leaf_4_clk_i),
    .d1(net1955),
    .d2(net2031),
    .o1(u_gpio_gen_filter_20__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_25__u_filter_diff_ctr_q[0]),
    .si1(net790),
    .si2(net791),
    .ssb(net1476));
 b15fqy043ar1n02x5 u_gpio_gen_filter_20__u_filter_stored_value_q_reg (.clk(clknet_leaf_4_clk_i),
    .d(u_gpio_gen_filter_20__u_filter_filter_synced),
    .den(eq_x_131_n25),
    .o(u_gpio_gen_filter_20__u_filter_stored_value_q),
    .rb(net532),
    .si(net792),
    .ssb(net1477));
 b15fqy203ar1n02x5 u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_1_ (.rb(net532),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2093),
    .d2(u_gpio_gen_filter_21__u_filter_diff_ctr_d[1]),
    .o1(u_gpio_gen_filter_21__u_filter_diff_ctr_q[0]),
    .o2(u_gpio_gen_filter_21__u_filter_diff_ctr_q[1]),
    .si1(net793),
    .si2(net794),
    .ssb(net1478));
 b15fqy203ar1n02x5 u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_3_ (.rb(net535),
    .clk(clknet_leaf_4_clk_i),
    .d1(u_gpio_gen_filter_21__u_filter_diff_ctr_d[2]),
    .d2(u_gpio_gen_filter_21__u_filter_diff_ctr_d[3]),
    .o1(u_gpio_gen_filter_21__u_filter_diff_ctr_q[2]),
    .o2(u_gpio_gen_filter_21__u_filter_diff_ctr_q[3]),
    .si1(net795),
    .si2(net796),
    .ssb(net1479));
 b15fqy203ar1n02x5 u_gpio_gen_filter_21__u_filter_filter_q_reg_u_gpio_gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net533),
    .clk(clknet_leaf_6_clk_i),
    .d1(u_gpio_gen_filter_21__u_filter_filter_synced),
    .d2(net1943),
    .o1(u_gpio_gen_filter_21__u_filter_filter_q),
    .o2(u_gpio_gen_filter_26__u_filter_filter_synced),
    .si1(net797),
    .si2(net798),
    .ssb(net1480));
 b15fqy043ar1n02x5 u_gpio_gen_filter_21__u_filter_stored_value_q_reg (.clk(clknet_leaf_4_clk_i),
    .d(u_gpio_gen_filter_21__u_filter_filter_synced),
    .den(eq_x_126_n25),
    .o(u_gpio_gen_filter_21__u_filter_stored_value_q),
    .rb(net532),
    .si(net799),
    .ssb(net1481));
 b15fqy203ar1n02x5 u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_3_ (.rb(net521),
    .clk(clknet_leaf_1_clk_i),
    .d1(u_gpio_gen_filter_22__u_filter_diff_ctr_d[1]),
    .d2(u_gpio_gen_filter_22__u_filter_diff_ctr_d[3]),
    .o1(u_gpio_gen_filter_22__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_22__u_filter_diff_ctr_q[3]),
    .si1(net800),
    .si2(net801),
    .ssb(net1482));
 b15fqy203ar1n02x5 u_gpio_gen_filter_22__u_filter_filter_q_reg_u_gpio_gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net535),
    .clk(clknet_leaf_3_clk_i),
    .d1(net2119),
    .d2(net2195),
    .o1(u_gpio_gen_filter_22__u_filter_filter_q),
    .o2(u_gpio_gen_filter_22__u_filter_filter_synced),
    .si1(net802),
    .si2(net803),
    .ssb(net1483));
 b15fqy203ar1n02x5 u_gpio_gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net535),
    .clk(clknet_leaf_5_clk_i),
    .d1(net804),
    .d2(net805),
    .o1(u_gpio_gen_filter_22__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_23__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net806),
    .si2(net807),
    .ssb(net1484));
 b15fqy043ar1n02x5 u_gpio_gen_filter_22__u_filter_stored_value_q_reg (.clk(clknet_leaf_3_clk_i),
    .d(u_gpio_gen_filter_22__u_filter_filter_synced),
    .den(eq_x_121_n25),
    .o(u_gpio_gen_filter_22__u_filter_stored_value_q),
    .rb(net532),
    .si(net808),
    .ssb(net1485));
 b15fqy203ar1n02x5 u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_2_ (.rb(net521),
    .clk(clknet_leaf_1_clk_i),
    .d1(u_gpio_gen_filter_23__u_filter_diff_ctr_d[1]),
    .d2(u_gpio_gen_filter_23__u_filter_diff_ctr_d[2]),
    .o1(u_gpio_gen_filter_23__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_23__u_filter_diff_ctr_q[2]),
    .si1(net809),
    .si2(net810),
    .ssb(net1486));
 b15fqy203ar1n02x5 u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_23__u_filter_filter_q_reg (.rb(net521),
    .clk(clknet_leaf_1_clk_i),
    .d1(net1988),
    .d2(net444),
    .o1(u_gpio_gen_filter_23__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_23__u_filter_filter_q),
    .si1(net811),
    .si2(net812),
    .ssb(net1487));
 b15fqy203ar1n02x5 u_gpio_gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_0_ (.rb(net536),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2011),
    .d2(net2144),
    .o1(u_gpio_gen_filter_23__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_24__u_filter_diff_ctr_q[0]),
    .si1(net813),
    .si2(net814),
    .ssb(net1488));
 b15fqy043ar1n02x5 u_gpio_gen_filter_23__u_filter_stored_value_q_reg (.clk(clknet_leaf_2_clk_i),
    .d(net444),
    .den(eq_x_116_n25),
    .o(u_gpio_gen_filter_23__u_filter_stored_value_q),
    .rb(net531),
    .si(net815),
    .ssb(net1489));
 b15fqy203ar1n02x5 u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_2_ (.rb(net534),
    .clk(clknet_leaf_5_clk_i),
    .d1(u_gpio_gen_filter_24__u_filter_diff_ctr_d[1]),
    .d2(u_gpio_gen_filter_24__u_filter_diff_ctr_d[2]),
    .o1(u_gpio_gen_filter_24__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_24__u_filter_diff_ctr_q[2]),
    .si1(net816),
    .si2(net817),
    .ssb(net1490));
 b15fqy203ar1n02x5 u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_24__u_filter_filter_q_reg (.rb(net536),
    .clk(clknet_leaf_5_clk_i),
    .d1(u_gpio_gen_filter_24__u_filter_diff_ctr_d[3]),
    .d2(net443),
    .o1(u_gpio_gen_filter_24__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_24__u_filter_filter_q),
    .si1(net818),
    .si2(net819),
    .ssb(net1491));
 b15fqy203ar1n02x5 u_gpio_gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net535),
    .clk(clknet_leaf_4_clk_i),
    .d1(net820),
    .d2(net821),
    .o1(u_gpio_gen_filter_24__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_25__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net822),
    .si2(net823),
    .ssb(net1492));
 b15fqy203ar1n02x5 u_gpio_gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_0_ (.rb(net535),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2070),
    .d2(u_gpio_gen_filter_27__u_filter_diff_ctr_d[0]),
    .o1(u_gpio_gen_filter_24__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_27__u_filter_diff_ctr_q[0]),
    .si1(net824),
    .si2(net825),
    .ssb(net1493));
 b15fqy043ar1n02x5 u_gpio_gen_filter_24__u_filter_stored_value_q_reg (.clk(clknet_leaf_5_clk_i),
    .d(net442),
    .den(eq_x_111_n25),
    .o(u_gpio_gen_filter_24__u_filter_stored_value_q),
    .rb(net534),
    .si(net826),
    .ssb(net1494));
 b15fqy203ar1n02x5 u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_2_ (.rb(net535),
    .clk(clknet_leaf_4_clk_i),
    .d1(u_gpio_gen_filter_25__u_filter_diff_ctr_d[1]),
    .d2(net2034),
    .o1(u_gpio_gen_filter_25__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_25__u_filter_diff_ctr_q[2]),
    .si1(net827),
    .si2(net828),
    .ssb(net1495));
 b15fqy203ar1n02x5 u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net535),
    .clk(clknet_leaf_5_clk_i),
    .d1(u_gpio_gen_filter_25__u_filter_diff_ctr_d[3]),
    .d2(net2010),
    .o1(u_gpio_gen_filter_25__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_25__u_filter_filter_synced),
    .si1(net829),
    .si2(net830),
    .ssb(net1496));
 b15fqy203ar1n02x5 u_gpio_gen_filter_25__u_filter_filter_q_reg_u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_0_ (.rb(net530),
    .clk(clknet_leaf_3_clk_i),
    .d1(u_gpio_gen_filter_25__u_filter_filter_synced),
    .d2(net2208),
    .o1(u_gpio_gen_filter_25__u_filter_filter_q),
    .o2(u_gpio_gen_filter_26__u_filter_diff_ctr_q[0]),
    .si1(net831),
    .si2(net832),
    .ssb(net1497));
 b15fqy043ar1n02x5 u_gpio_gen_filter_25__u_filter_stored_value_q_reg (.clk(clknet_leaf_5_clk_i),
    .d(u_gpio_gen_filter_25__u_filter_filter_synced),
    .den(eq_x_106_n25),
    .o(u_gpio_gen_filter_25__u_filter_stored_value_q),
    .rb(net535),
    .si(net833),
    .ssb(net1498));
 b15fqy203ar1n02x5 u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_2_ (.rb(net530),
    .clk(clknet_leaf_3_clk_i),
    .d1(u_gpio_gen_filter_26__u_filter_diff_ctr_d[1]),
    .d2(u_gpio_gen_filter_26__u_filter_diff_ctr_d[2]),
    .o1(u_gpio_gen_filter_26__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_26__u_filter_diff_ctr_q[2]),
    .si1(net834),
    .si2(net835),
    .ssb(net1499));
 b15fqy203ar1n02x5 u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_29__u_filter_filter_q_reg (.rb(net532),
    .clk(clknet_leaf_3_clk_i),
    .d1(net2175),
    .d2(u_gpio_gen_filter_29__u_filter_filter_synced),
    .o1(u_gpio_gen_filter_26__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_29__u_filter_filter_q),
    .si1(net836),
    .si2(net837),
    .ssb(net1500));
 b15fqy203ar1n02x5 u_gpio_gen_filter_26__u_filter_filter_q_reg_u_gpio_intr_hw_intr_o_reg_12_ (.rb(net529),
    .clk(clknet_leaf_3_clk_i),
    .d1(u_gpio_gen_filter_26__u_filter_filter_synced),
    .d2(u_gpio_intr_hw_N20),
    .o1(u_gpio_gen_filter_26__u_filter_filter_q),
    .si1(net838),
    .si2(net839),
    .ssb(net1501));
 b15fqy203ar1n02x5 u_gpio_gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net533),
    .clk(clknet_leaf_6_clk_i),
    .d1(net840),
    .d2(net841),
    .o1(u_gpio_gen_filter_26__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_27__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net842),
    .si2(net843),
    .ssb(net1502));
 b15fqy043ar1n02x5 u_gpio_gen_filter_26__u_filter_stored_value_q_reg (.clk(clknet_leaf_3_clk_i),
    .d(u_gpio_gen_filter_26__u_filter_filter_synced),
    .den(eq_x_101_n25),
    .o(u_gpio_gen_filter_26__u_filter_stored_value_q),
    .rb(net530),
    .si(net844),
    .ssb(net1503));
 b15fqy203ar1n02x5 u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_2_ (.rb(net536),
    .clk(clknet_leaf_5_clk_i),
    .d1(u_gpio_gen_filter_27__u_filter_diff_ctr_d[1]),
    .d2(net2023),
    .o1(u_gpio_gen_filter_27__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_27__u_filter_diff_ctr_q[2]),
    .si1(net845),
    .si2(net846),
    .ssb(net1504));
 b15fqy203ar1n02x5 u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_27__u_filter_filter_q_reg (.rb(net534),
    .clk(clknet_leaf_5_clk_i),
    .d1(u_gpio_gen_filter_27__u_filter_diff_ctr_d[3]),
    .d2(u_gpio_gen_filter_27__u_filter_filter_synced),
    .o1(u_gpio_gen_filter_27__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_27__u_filter_filter_q),
    .si1(net847),
    .si2(net848),
    .ssb(net1505));
 b15fqy203ar1n02x5 u_gpio_gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_intr_hw_intr_o_reg_24_ (.rb(net533),
    .clk(clknet_leaf_6_clk_i),
    .d1(net1936),
    .d2(u_gpio_intr_hw_N8),
    .o1(u_gpio_gen_filter_27__u_filter_filter_synced),
    .si1(net849),
    .si2(net850),
    .ssb(net1506));
 b15fqy043ar1n02x5 u_gpio_gen_filter_27__u_filter_stored_value_q_reg (.clk(clknet_leaf_5_clk_i),
    .d(u_gpio_gen_filter_27__u_filter_filter_synced),
    .den(eq_x_96_n25),
    .o(u_gpio_gen_filter_27__u_filter_stored_value_q),
    .rb(net533),
    .si(net851),
    .ssb(net1507));
 b15fqy203ar1n02x5 u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_1_ (.rb(net531),
    .clk(clknet_leaf_2_clk_i),
    .d1(net1957),
    .d2(u_gpio_gen_filter_28__u_filter_diff_ctr_d[1]),
    .o1(u_gpio_gen_filter_28__u_filter_diff_ctr_q[0]),
    .o2(u_gpio_gen_filter_28__u_filter_diff_ctr_q[1]),
    .si1(net852),
    .si2(net853),
    .ssb(net1508));
 b15fqy203ar1n02x5 u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_3_ (.rb(net529),
    .clk(clknet_leaf_3_clk_i),
    .d1(u_gpio_gen_filter_28__u_filter_diff_ctr_d[2]),
    .d2(u_gpio_gen_filter_28__u_filter_diff_ctr_d[3]),
    .o1(u_gpio_gen_filter_28__u_filter_diff_ctr_q[2]),
    .o2(u_gpio_gen_filter_28__u_filter_diff_ctr_q[3]),
    .si1(net854),
    .si2(net855),
    .ssb(net1509));
 b15fqy203ar1n02x5 u_gpio_gen_filter_28__u_filter_filter_q_reg_u_gpio_gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net531),
    .clk(clknet_leaf_3_clk_i),
    .d1(u_gpio_gen_filter_28__u_filter_filter_synced),
    .d2(net1932),
    .o1(u_gpio_gen_filter_28__u_filter_filter_q),
    .o2(u_gpio_gen_filter_28__u_filter_filter_synced),
    .si1(net856),
    .si2(net857),
    .ssb(net1510));
 b15fqy203ar1n02x5 u_gpio_gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net529),
    .clk(clknet_leaf_3_clk_i),
    .d1(net858),
    .d2(net859),
    .o1(u_gpio_gen_filter_28__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_29__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net860),
    .si2(net861),
    .ssb(net1511));
 b15fqy043ar1n02x5 u_gpio_gen_filter_28__u_filter_stored_value_q_reg (.clk(clknet_leaf_3_clk_i),
    .d(u_gpio_gen_filter_28__u_filter_filter_synced),
    .den(eq_x_91_n25),
    .o(u_gpio_gen_filter_28__u_filter_stored_value_q),
    .rb(net529),
    .si(net862),
    .ssb(net1512));
 b15fqy203ar1n02x5 u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_1_ (.rb(net532),
    .clk(clknet_leaf_3_clk_i),
    .d1(u_gpio_gen_filter_29__u_filter_diff_ctr_d[0]),
    .d2(u_gpio_gen_filter_29__u_filter_diff_ctr_d[1]),
    .o1(u_gpio_gen_filter_29__u_filter_diff_ctr_q[0]),
    .o2(u_gpio_gen_filter_29__u_filter_diff_ctr_q[1]),
    .si1(net863),
    .si2(net864),
    .ssb(net1513));
 b15fqy203ar1n02x5 u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_3_ (.rb(net532),
    .clk(clknet_leaf_4_clk_i),
    .d1(net1950),
    .d2(net1954),
    .o1(u_gpio_gen_filter_29__u_filter_diff_ctr_q[2]),
    .o2(u_gpio_gen_filter_29__u_filter_diff_ctr_q[3]),
    .si1(net865),
    .si2(net866),
    .ssb(net1514));
 b15fqy203ar1n02x5 u_gpio_gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_0_ (.rb(net533),
    .clk(clknet_leaf_5_clk_i),
    .d1(u_gpio_gen_filter_29__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .d2(u_gpio_gen_filter_30__u_filter_diff_ctr_d[0]),
    .o1(u_gpio_gen_filter_29__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_30__u_filter_diff_ctr_q[0]),
    .si1(net867),
    .si2(net868),
    .ssb(net1515));
 b15fqy043ar1n02x5 u_gpio_gen_filter_29__u_filter_stored_value_q_reg (.clk(clknet_leaf_5_clk_i),
    .d(u_gpio_gen_filter_29__u_filter_filter_synced),
    .den(eq_x_86_n25),
    .o(u_gpio_gen_filter_29__u_filter_stored_value_q),
    .rb(net535),
    .si(net869),
    .ssb(net1516));
 b15fqy203ar1n02x5 u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_1_ (.rb(net515),
    .clk(clknet_leaf_0_clk_i),
    .d1(net1976),
    .d2(net2185),
    .o1(u_gpio_gen_filter_2__u_filter_diff_ctr_q[0]),
    .o2(u_gpio_gen_filter_2__u_filter_diff_ctr_q[1]),
    .si1(net870),
    .si2(net871),
    .ssb(net1517));
 b15fqy203ar1n02x5 u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_3_ (.rb(net518),
    .clk(clknet_leaf_0_clk_i),
    .d1(u_gpio_gen_filter_2__u_filter_diff_ctr_d[2]),
    .d2(u_gpio_gen_filter_2__u_filter_diff_ctr_d[3]),
    .o1(u_gpio_gen_filter_2__u_filter_diff_ctr_q[2]),
    .o2(u_gpio_gen_filter_2__u_filter_diff_ctr_q[3]),
    .si1(net872),
    .si2(net873),
    .ssb(net1518));
 b15fqy203ar1n02x5 u_gpio_gen_filter_2__u_filter_filter_q_reg_u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_1_ (.rb(net519),
    .clk(clknet_leaf_2_clk_i),
    .d1(u_gpio_gen_filter_2__u_filter_filter_synced),
    .d2(u_gpio_gen_filter_7__u_filter_diff_ctr_d[1]),
    .o1(u_gpio_gen_filter_2__u_filter_filter_q),
    .o2(u_gpio_gen_filter_7__u_filter_diff_ctr_q[1]),
    .si1(net874),
    .si2(net875),
    .ssb(net1519));
 b15fqy203ar1n02x5 u_gpio_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net521),
    .clk(clknet_leaf_2_clk_i),
    .d1(net876),
    .d2(net877),
    .o1(u_gpio_gen_filter_2__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_3__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net878),
    .si2(net879),
    .ssb(net1520));
 b15fqy203ar1n02x5 u_gpio_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_0_ (.rb(net519),
    .clk(clknet_leaf_2_clk_i),
    .d1(net1945),
    .d2(u_gpio_gen_filter_3__u_filter_diff_ctr_d[0]),
    .o1(u_gpio_gen_filter_2__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_3__u_filter_diff_ctr_q[0]),
    .si1(net880),
    .si2(net881),
    .ssb(net1521));
 b15fqy043ar1n02x5 u_gpio_gen_filter_2__u_filter_stored_value_q_reg (.clk(clknet_leaf_0_clk_i),
    .d(u_gpio_gen_filter_2__u_filter_filter_synced),
    .den(eq_x_221_n25),
    .o(u_gpio_gen_filter_2__u_filter_stored_value_q),
    .rb(net518),
    .si(net882),
    .ssb(net1522));
 b15fqy203ar1n02x5 u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_30__u_filter_filter_q_reg (.rb(net534),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2140),
    .d2(u_gpio_gen_filter_30__u_filter_filter_synced),
    .o1(u_gpio_gen_filter_30__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_30__u_filter_filter_q),
    .si1(net883),
    .si2(net884),
    .ssb(net1523));
 b15fqy203ar1n02x5 u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_3_ (.rb(net534),
    .clk(clknet_leaf_5_clk_i),
    .d1(u_gpio_gen_filter_30__u_filter_diff_ctr_d[2]),
    .d2(u_gpio_gen_filter_30__u_filter_diff_ctr_d[3]),
    .o1(u_gpio_gen_filter_30__u_filter_diff_ctr_q[2]),
    .o2(u_gpio_gen_filter_30__u_filter_diff_ctr_q[3]),
    .si1(net885),
    .si2(net886),
    .ssb(net1524));
 b15fqy203ar1n02x5 u_gpio_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net529),
    .clk(clknet_leaf_3_clk_i),
    .d1(net887),
    .d2(net888),
    .o1(u_gpio_gen_filter_30__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_31__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net889),
    .si2(net890),
    .ssb(net1525));
 b15fqy003ar1n02x5 u_gpio_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net529),
    .clk(clknet_leaf_3_clk_i),
    .d(net1939),
    .o(u_gpio_gen_filter_30__u_filter_filter_synced),
    .si(net891),
    .ssb(net1526));
 b15fqy043ar1n02x5 u_gpio_gen_filter_30__u_filter_stored_value_q_reg (.clk(clknet_leaf_5_clk_i),
    .d(u_gpio_gen_filter_30__u_filter_filter_synced),
    .den(eq_x_81_n25),
    .o(u_gpio_gen_filter_30__u_filter_stored_value_q),
    .rb(net533),
    .si(net892),
    .ssb(net1527));
 b15fqy203ar1n02x5 u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_1_ (.rb(net516),
    .clk(clknet_leaf_0_clk_i),
    .d1(u_gpio_gen_filter_31__u_filter_diff_ctr_d[0]),
    .d2(u_gpio_gen_filter_31__u_filter_diff_ctr_d[1]),
    .o1(u_gpio_gen_filter_31__u_filter_diff_ctr_q[0]),
    .o2(u_gpio_gen_filter_31__u_filter_diff_ctr_q[1]),
    .si1(net893),
    .si2(net894),
    .ssb(net1528));
 b15fqy203ar1n02x5 u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_3_ (.rb(net517),
    .clk(clknet_leaf_0_clk_i),
    .d1(u_gpio_gen_filter_31__u_filter_diff_ctr_d[2]),
    .d2(u_gpio_gen_filter_31__u_filter_diff_ctr_d[3]),
    .o1(u_gpio_gen_filter_31__u_filter_diff_ctr_q[2]),
    .o2(u_gpio_gen_filter_31__u_filter_diff_ctr_q[3]),
    .si1(net895),
    .si2(net896),
    .ssb(net1529));
 b15fqy203ar1n02x5 u_gpio_gen_filter_31__u_filter_filter_q_reg_u_gpio_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net530),
    .clk(clknet_leaf_6_clk_i),
    .d1(u_gpio_gen_filter_31__u_filter_filter_synced),
    .d2(net1933),
    .o1(u_gpio_gen_filter_31__u_filter_filter_q),
    .o2(u_gpio_gen_filter_31__u_filter_filter_synced),
    .si1(net897),
    .si2(net898),
    .ssb(net1530));
 b15fqy043ar1n02x5 u_gpio_gen_filter_31__u_filter_stored_value_q_reg (.clk(clknet_leaf_6_clk_i),
    .d(u_gpio_gen_filter_31__u_filter_filter_synced),
    .den(eq_x_76_n25),
    .o(u_gpio_gen_filter_31__u_filter_stored_value_q),
    .rb(net533),
    .si(net899),
    .ssb(net1531));
 b15fqy203ar1n02x5 u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_2_ (.rb(net521),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2173),
    .d2(u_gpio_gen_filter_3__u_filter_diff_ctr_d[2]),
    .o1(u_gpio_gen_filter_3__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_3__u_filter_diff_ctr_q[2]),
    .si1(net900),
    .si2(net901),
    .ssb(net1532));
 b15fqy203ar1n02x5 u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_3__u_filter_filter_q_reg (.rb(net519),
    .clk(clknet_leaf_0_clk_i),
    .d1(net1984),
    .d2(u_gpio_gen_filter_3__u_filter_filter_synced),
    .o1(u_gpio_gen_filter_3__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_3__u_filter_filter_q),
    .si1(net902),
    .si2(net903),
    .ssb(net1533));
 b15fqy203ar1n02x5 u_gpio_gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_7__u_filter_filter_q_reg (.rb(net522),
    .clk(clknet_leaf_2_clk_i),
    .d1(net1960),
    .d2(net2086),
    .o1(u_gpio_gen_filter_3__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_7__u_filter_filter_q),
    .si1(net904),
    .si2(net905),
    .ssb(net1534));
 b15fqy043ar1n02x5 u_gpio_gen_filter_3__u_filter_stored_value_q_reg (.clk(clknet_leaf_2_clk_i),
    .d(u_gpio_gen_filter_3__u_filter_filter_synced),
    .den(eq_x_216_n25),
    .o(u_gpio_gen_filter_3__u_filter_stored_value_q),
    .rb(net520),
    .si(net906),
    .ssb(net1535));
 b15fqy203ar1n02x5 u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_2_ (.rb(net511),
    .clk(clknet_leaf_10_clk_i),
    .d1(u_gpio_gen_filter_4__u_filter_diff_ctr_d[1]),
    .d2(net2055),
    .o1(u_gpio_gen_filter_4__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_4__u_filter_diff_ctr_q[2]),
    .si1(net907),
    .si2(net908),
    .ssb(net1536));
 b15fqy203ar1n02x5 u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_4__u_filter_filter_q_reg (.rb(net511),
    .clk(clknet_leaf_10_clk_i),
    .d1(u_gpio_gen_filter_4__u_filter_diff_ctr_d[3]),
    .d2(net441),
    .o1(u_gpio_gen_filter_4__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_4__u_filter_filter_q),
    .si1(net909),
    .si2(net910),
    .ssb(net1537));
 b15fqy203ar1n02x5 u_gpio_gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net510),
    .clk(clknet_leaf_11_clk_i),
    .d1(net911),
    .d2(net912),
    .o1(u_gpio_gen_filter_4__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_5__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net913),
    .si2(net914),
    .ssb(net1538));
 b15fqy203ar1n02x5 u_gpio_gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_0_ (.rb(net510),
    .clk(clknet_leaf_11_clk_i),
    .d1(net1944),
    .d2(u_gpio_gen_filter_5__u_filter_diff_ctr_d[0]),
    .o1(u_gpio_gen_filter_4__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_5__u_filter_diff_ctr_q[0]),
    .si1(net915),
    .si2(net916),
    .ssb(net1539));
 b15fqy043ar1n02x5 u_gpio_gen_filter_4__u_filter_stored_value_q_reg (.clk(clknet_leaf_10_clk_i),
    .d(net441),
    .den(eq_x_211_n25),
    .o(u_gpio_gen_filter_4__u_filter_stored_value_q),
    .rb(net511),
    .si(net917),
    .ssb(net1540));
 b15fqy203ar1n02x5 u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_2_ (.rb(net515),
    .clk(clknet_leaf_11_clk_i),
    .d1(net2075),
    .d2(net2099),
    .o1(u_gpio_gen_filter_5__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_5__u_filter_diff_ctr_q[2]),
    .si1(net918),
    .si2(net919),
    .ssb(net1541));
 b15fqy203ar1n02x5 u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_5__u_filter_filter_q_reg (.rb(net510),
    .clk(clknet_leaf_11_clk_i),
    .d1(u_gpio_gen_filter_5__u_filter_diff_ctr_d[3]),
    .d2(net2170),
    .o1(u_gpio_gen_filter_5__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_5__u_filter_filter_q),
    .si1(net920),
    .si2(net921),
    .ssb(net1542));
 b15fqy203ar1n02x5 u_gpio_gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_0_ (.rb(net518),
    .clk(clknet_leaf_11_clk_i),
    .d1(net1958),
    .d2(u_gpio_gen_filter_12__u_filter_diff_ctr_d[0]),
    .o1(u_gpio_gen_filter_5__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_12__u_filter_diff_ctr_q[0]),
    .si1(net922),
    .si2(net923),
    .ssb(net1543));
 b15fqy043ar1n02x5 u_gpio_gen_filter_5__u_filter_stored_value_q_reg (.clk(clknet_leaf_11_clk_i),
    .d(u_gpio_gen_filter_5__u_filter_filter_synced),
    .den(eq_x_206_n25),
    .o(u_gpio_gen_filter_5__u_filter_stored_value_q),
    .rb(net510),
    .si(net924),
    .ssb(net1544));
 b15fqy203ar1n02x5 u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_2_ (.rb(net536),
    .clk(clknet_leaf_4_clk_i),
    .d1(u_gpio_gen_filter_6__u_filter_diff_ctr_d[1]),
    .d2(u_gpio_gen_filter_6__u_filter_diff_ctr_d[2]),
    .o1(u_gpio_gen_filter_6__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_6__u_filter_diff_ctr_q[2]),
    .si1(net925),
    .si2(net926),
    .ssb(net1545));
 b15fqy203ar1n02x5 u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_6__u_filter_filter_q_reg (.rb(net537),
    .clk(clknet_leaf_4_clk_i),
    .d1(u_gpio_gen_filter_6__u_filter_diff_ctr_d[3]),
    .d2(net440),
    .o1(u_gpio_gen_filter_6__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_6__u_filter_filter_q),
    .si1(net927),
    .si2(net928),
    .ssb(net1546));
 b15fqy203ar1n02x5 u_gpio_gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net531),
    .clk(clknet_leaf_3_clk_i),
    .d1(net929),
    .d2(net930),
    .o1(u_gpio_gen_filter_6__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_7__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net931),
    .si2(net932),
    .ssb(net1547));
 b15fqy203ar1n02x5 u_gpio_gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_0_ (.rb(net532),
    .clk(clknet_leaf_3_clk_i),
    .d1(net1938),
    .d2(u_gpio_gen_filter_17__u_filter_diff_ctr_d[0]),
    .o1(u_gpio_gen_filter_6__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_17__u_filter_diff_ctr_q[0]),
    .si1(net933),
    .si2(net934),
    .ssb(net1548));
 b15fqy043ar1n02x5 u_gpio_gen_filter_6__u_filter_stored_value_q_reg (.clk(clknet_leaf_3_clk_i),
    .d(net2094),
    .den(eq_x_201_n25),
    .o(u_gpio_gen_filter_6__u_filter_stored_value_q),
    .rb(net531),
    .si(net935),
    .ssb(net1549));
 b15fqy203ar1n02x5 u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_2_ (.rb(net522),
    .clk(clknet_leaf_2_clk_i),
    .d1(u_gpio_gen_filter_7__u_filter_diff_ctr_d[0]),
    .d2(u_gpio_gen_filter_7__u_filter_diff_ctr_d[2]),
    .o1(u_gpio_gen_filter_7__u_filter_diff_ctr_q[0]),
    .o2(u_gpio_gen_filter_7__u_filter_diff_ctr_q[2]),
    .si1(net936),
    .si2(net937),
    .ssb(net1550));
 b15fqy203ar1n02x5 u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_0_ (.rb(net531),
    .clk(clknet_leaf_2_clk_i),
    .d1(u_gpio_gen_filter_7__u_filter_diff_ctr_d[3]),
    .d2(u_gpio_gen_filter_8__u_filter_diff_ctr_d[0]),
    .o1(u_gpio_gen_filter_7__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_8__u_filter_diff_ctr_q[0]),
    .si1(net938),
    .si2(net939),
    .ssb(net1551));
 b15fqy203ar1n02x5 u_gpio_gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net522),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2166),
    .d2(net1941),
    .o1(u_gpio_gen_filter_7__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_11__u_filter_filter_synced),
    .si1(net940),
    .si2(net941),
    .ssb(net1552));
 b15fqy043ar1n02x5 u_gpio_gen_filter_7__u_filter_stored_value_q_reg (.clk(clknet_leaf_2_clk_i),
    .d(u_gpio_gen_filter_7__u_filter_filter_synced),
    .den(eq_x_196_n25),
    .o(u_gpio_gen_filter_7__u_filter_stored_value_q),
    .rb(net522),
    .si(net942),
    .ssb(net1553));
 b15fqy203ar1n02x5 u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_2_ (.rb(net532),
    .clk(clknet_leaf_4_clk_i),
    .d1(u_gpio_gen_filter_8__u_filter_diff_ctr_d[1]),
    .d2(u_gpio_gen_filter_8__u_filter_diff_ctr_d[2]),
    .o1(u_gpio_gen_filter_8__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_8__u_filter_diff_ctr_q[2]),
    .si1(net943),
    .si2(net944),
    .ssb(net1554));
 b15fqy203ar1n02x5 u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_0_ (.rb(net537),
    .clk(clknet_leaf_4_clk_i),
    .d1(u_gpio_gen_filter_8__u_filter_diff_ctr_d[3]),
    .d2(u_gpio_gen_filter_9__u_filter_diff_ctr_d[0]),
    .o1(u_gpio_gen_filter_8__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_9__u_filter_diff_ctr_q[0]),
    .si1(net945),
    .si2(net946),
    .ssb(net1555));
 b15fqy203ar1n02x5 u_gpio_gen_filter_8__u_filter_filter_q_reg_u_gpio_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net522),
    .clk(clknet_leaf_2_clk_i),
    .d1(u_gpio_gen_filter_8__u_filter_filter_synced),
    .d2(net1934),
    .o1(u_gpio_gen_filter_8__u_filter_filter_q),
    .o2(u_gpio_gen_filter_8__u_filter_filter_synced),
    .si1(net947),
    .si2(net948),
    .ssb(net1556));
 b15fqy203ar1n02x5 u_gpio_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net522),
    .clk(clknet_leaf_2_clk_i),
    .d1(net949),
    .d2(net950),
    .o1(u_gpio_gen_filter_8__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(u_gpio_gen_filter_9__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net951),
    .si2(net952),
    .ssb(net1557));
 b15fqy043ar1n02x5 u_gpio_gen_filter_8__u_filter_stored_value_q_reg (.clk(clknet_leaf_2_clk_i),
    .d(u_gpio_gen_filter_8__u_filter_filter_synced),
    .den(eq_x_191_n25),
    .o(u_gpio_gen_filter_8__u_filter_stored_value_q),
    .rb(net522),
    .si(net953),
    .ssb(net1558));
 b15fqy203ar1n02x5 u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_2_ (.rb(net537),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2041),
    .d2(u_gpio_gen_filter_9__u_filter_diff_ctr_d[2]),
    .o1(u_gpio_gen_filter_9__u_filter_diff_ctr_q[1]),
    .o2(u_gpio_gen_filter_9__u_filter_diff_ctr_q[2]),
    .si1(net954),
    .si2(net955),
    .ssb(net1559));
 b15fqy203ar1n02x5 u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_9__u_filter_filter_q_reg (.rb(net536),
    .clk(clknet_leaf_5_clk_i),
    .d1(u_gpio_gen_filter_9__u_filter_diff_ctr_d[3]),
    .d2(net439),
    .o1(u_gpio_gen_filter_9__u_filter_diff_ctr_q[3]),
    .o2(u_gpio_gen_filter_9__u_filter_filter_q),
    .si1(net956),
    .si2(net957),
    .ssb(net1560));
 b15fqy203ar1n02x5 u_gpio_gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_2_ (.rb(net531),
    .clk(clknet_leaf_3_clk_i),
    .d1(net2021),
    .d2(u_gpio_gen_filter_10__u_filter_diff_ctr_d[2]),
    .o1(u_gpio_gen_filter_9__u_filter_filter_synced),
    .o2(u_gpio_gen_filter_10__u_filter_diff_ctr_q[2]),
    .si1(net958),
    .si2(net959),
    .ssb(net1561));
 b15fqy043ar1n02x5 u_gpio_gen_filter_9__u_filter_stored_value_q_reg (.clk(clknet_leaf_4_clk_i),
    .d(u_gpio_gen_filter_9__u_filter_filter_synced),
    .den(eq_x_186_n25),
    .o(u_gpio_gen_filter_9__u_filter_stored_value_q),
    .rb(net537),
    .si(net960),
    .ssb(net1562));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_0__u_gpio_intr_hw_intr_o_reg_1_ (.rb(net510),
    .clk(clknet_leaf_11_clk_i),
    .d1(u_gpio_intr_hw_N32),
    .d2(u_gpio_intr_hw_N31),
    .si1(net961),
    .si2(net962),
    .ssb(net1563));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_10__u_gpio_intr_hw_intr_o_reg_11_ (.rb(net520),
    .clk(clknet_leaf_2_clk_i),
    .d1(u_gpio_intr_hw_N22),
    .d2(u_gpio_intr_hw_N21),
    .si1(net963),
    .si2(net964),
    .ssb(net1564));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_13__u_gpio_intr_hw_intr_o_reg_14_ (.rb(net520),
    .clk(clknet_leaf_12_clk_i),
    .d1(u_gpio_intr_hw_N19),
    .d2(u_gpio_intr_hw_N18),
    .si1(net965),
    .si2(net966),
    .ssb(net1565));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_15__u_gpio_intr_hw_intr_o_reg_16_ (.rb(net529),
    .clk(clknet_leaf_3_clk_i),
    .d1(u_gpio_intr_hw_N17),
    .d2(u_gpio_intr_hw_N16),
    .si1(net967),
    .si2(net968),
    .ssb(net1566));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_17__u_gpio_intr_hw_intr_o_reg_18_ (.rb(net525),
    .clk(clknet_leaf_8_clk_i),
    .d1(u_gpio_intr_hw_N15),
    .d2(u_gpio_intr_hw_N14),
    .si1(net969),
    .si2(net970),
    .ssb(net1567));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_19__u_gpio_intr_hw_intr_o_reg_20_ (.rb(net524),
    .clk(clknet_leaf_8_clk_i),
    .d1(u_gpio_intr_hw_N13),
    .d2(u_gpio_intr_hw_N12),
    .si1(net971),
    .si2(net972),
    .ssb(net1568));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_21__u_gpio_intr_hw_intr_o_reg_29_ (.rb(net527),
    .clk(clknet_leaf_7_clk_i),
    .d1(u_gpio_intr_hw_N11),
    .d2(u_gpio_intr_hw_N3),
    .si1(net973),
    .si2(net974),
    .ssb(net1569));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_22__u_gpio_intr_hw_intr_o_reg_23_ (.rb(net525),
    .clk(clknet_leaf_6_clk_i),
    .d1(u_gpio_intr_hw_N10),
    .d2(u_gpio_intr_hw_N9),
    .si1(net975),
    .si2(net976),
    .ssb(net1570));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_25__u_gpio_intr_hw_intr_o_reg_26_ (.rb(net533),
    .clk(clknet_leaf_6_clk_i),
    .d1(u_gpio_intr_hw_N7),
    .d2(u_gpio_intr_hw_N6),
    .si1(net977),
    .si2(net978),
    .ssb(net1571));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_27__u_gpio_u_reg_err_q_reg (.rb(net525),
    .clk(clknet_leaf_9_clk_i),
    .d1(u_gpio_intr_hw_N5),
    .d2(net1990),
    .o2(u_gpio_u_reg_err_q),
    .si1(net979),
    .si2(net980),
    .ssb(net1572));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_28__u_gpio_u_reg_u_data_in_q_reg_2_ (.rb(net524),
    .clk(clknet_leaf_8_clk_i),
    .d1(u_gpio_intr_hw_N4),
    .d2(u_gpio_u_reg_u_data_in_wr_data[2]),
    .o2(u_gpio_u_reg_data_in_qs[2]),
    .si1(net981),
    .si2(net982),
    .ssb(net1573));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_2__u_gpio_intr_hw_intr_o_reg_3_ (.rb(net524),
    .clk(clknet_leaf_9_clk_i),
    .d1(u_gpio_intr_hw_N30),
    .d2(u_gpio_intr_hw_N29),
    .si1(net983),
    .si2(net984),
    .ssb(net1574));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_30__u_gpio_intr_hw_intr_o_reg_31_ (.rb(net529),
    .clk(clknet_leaf_3_clk_i),
    .d1(u_gpio_intr_hw_N2),
    .d2(u_gpio_intr_hw_N1),
    .si1(net985),
    .si2(net986),
    .ssb(net1575));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_4__u_gpio_intr_hw_intr_o_reg_5_ (.rb(net511),
    .clk(clknet_leaf_10_clk_i),
    .d1(u_gpio_intr_hw_N28),
    .d2(u_gpio_intr_hw_N27),
    .si1(net987),
    .si2(net988),
    .ssb(net1576));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_6__u_gpio_intr_hw_intr_o_reg_7_ (.rb(net510),
    .clk(clknet_leaf_11_clk_i),
    .d1(u_gpio_intr_hw_N26),
    .d2(u_gpio_intr_hw_N25),
    .si1(net989),
    .si2(net990),
    .ssb(net1577));
 b15fqy203ar1n02x5 u_gpio_intr_hw_intr_o_reg_8__u_gpio_intr_hw_intr_o_reg_9_ (.rb(net529),
    .clk(clknet_leaf_3_clk_i),
    .d1(u_gpio_intr_hw_N24),
    .d2(u_gpio_intr_hw_N23),
    .si1(net991),
    .si2(net992),
    .ssb(net1578));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_ctrl_en_input_filter_clk_gate_q_reg_0_latch (.clk(clknet_leaf_6_clk_i),
    .clkout(u_gpio_u_reg_u_ctrl_en_input_filter_net3627),
    .en(n3942),
    .te(net993));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_ctrl_en_input_filter_clk_gate_q_reg_latch (.clk(clknet_leaf_12_clk_i),
    .clkout(u_gpio_u_reg_u_ctrl_en_input_filter_net3621),
    .en(n3942),
    .te(net994));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_0__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_1_ (.rb(net519),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3621),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[0]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[1]),
    .o1(u_gpio_reg2hw[0]),
    .o2(u_gpio_reg2hw[1]),
    .si1(net995),
    .si2(net996),
    .ssb(net1579));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_10__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_11_ (.rb(net520),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3621),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[10]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[11]),
    .o1(u_gpio_reg2hw[10]),
    .o2(u_gpio_reg2hw[11]),
    .si1(net997),
    .si2(net998),
    .ssb(net1580));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_12__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_13_ (.rb(net519),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3621),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[12]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[13]),
    .o1(u_gpio_reg2hw[12]),
    .o2(u_gpio_reg2hw[13]),
    .si1(net999),
    .si2(net1000),
    .ssb(net1581));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_14__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_15_ (.rb(net519),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3621),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[14]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[15]),
    .o1(u_gpio_reg2hw[14]),
    .o2(u_gpio_reg2hw[15]),
    .si1(net1001),
    .si2(net1002),
    .ssb(net1582));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_16__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_17_ (.rb(net530),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3627),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[16]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[17]),
    .o1(u_gpio_reg2hw[16]),
    .o2(u_gpio_reg2hw[17]),
    .si1(net1003),
    .si2(net1004),
    .ssb(net1583));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_18__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_19_ (.rb(net530),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3627),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[18]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[19]),
    .o1(u_gpio_reg2hw[18]),
    .o2(u_gpio_reg2hw[19]),
    .si1(net1005),
    .si2(net1006),
    .ssb(net1584));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_20__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_21_ (.rb(net530),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3627),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[20]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[21]),
    .o1(u_gpio_reg2hw[20]),
    .o2(u_gpio_reg2hw[21]),
    .si1(net1007),
    .si2(net1008),
    .ssb(net1585));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_22__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_23_ (.rb(net530),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3627),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[22]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[23]),
    .o1(u_gpio_reg2hw[22]),
    .o2(u_gpio_reg2hw[23]),
    .si1(net1009),
    .si2(net1010),
    .ssb(net1586));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_24__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_25_ (.rb(net533),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3627),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[24]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[25]),
    .o1(u_gpio_reg2hw[24]),
    .o2(u_gpio_reg2hw[25]),
    .si1(net1011),
    .si2(net1012),
    .ssb(net1587));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_26__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_27_ (.rb(net533),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3627),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[26]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[27]),
    .o1(u_gpio_reg2hw[26]),
    .o2(u_gpio_reg2hw[27]),
    .si1(net1013),
    .si2(net1014),
    .ssb(net1588));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_28__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_29_ (.rb(net533),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3627),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[28]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[29]),
    .o1(u_gpio_reg2hw[28]),
    .o2(u_gpio_reg2hw[29]),
    .si1(net1015),
    .si2(net1016),
    .ssb(net1589));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_2__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_3_ (.rb(net520),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3621),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[2]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[3]),
    .o1(u_gpio_reg2hw[2]),
    .o2(u_gpio_reg2hw[3]),
    .si1(net1017),
    .si2(net1018),
    .ssb(net1590));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_30__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_31_ (.rb(net533),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3627),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[30]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[31]),
    .o1(u_gpio_reg2hw[30]),
    .o2(u_gpio_reg2hw[31]),
    .si1(net1019),
    .si2(net1020),
    .ssb(net1591));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_4__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_5_ (.rb(net519),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3621),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[4]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[5]),
    .o1(u_gpio_reg2hw[4]),
    .o2(u_gpio_reg2hw[5]),
    .si1(net1021),
    .si2(net1022),
    .ssb(net1592));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_6__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_7_ (.rb(net519),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3621),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[6]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[7]),
    .o1(u_gpio_reg2hw[6]),
    .o2(u_gpio_reg2hw[7]),
    .si1(net1023),
    .si2(net1024),
    .ssb(net1593));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_8__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_9_ (.rb(net520),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3621),
    .d1(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[8]),
    .d2(u_gpio_u_reg_u_ctrl_en_input_filter_wr_data[9]),
    .o1(u_gpio_reg2hw[8]),
    .o2(u_gpio_reg2hw[9]),
    .si1(net1025),
    .si2(net1026),
    .ssb(net1594));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_0__u_gpio_u_reg_u_data_in_q_reg_1_ (.rb(net519),
    .clk(clknet_leaf_0_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[0]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[1]),
    .o1(u_gpio_u_reg_data_in_qs[0]),
    .o2(u_gpio_u_reg_data_in_qs[1]),
    .si1(net1027),
    .si2(net1028),
    .ssb(net1595));
 b15fqy003ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_13_ (.rb(net513),
    .clk(clknet_leaf_11_clk_i),
    .d(u_gpio_u_reg_u_data_in_wr_data[13]),
    .o(u_gpio_u_reg_data_in_qs[13]),
    .si(net1029),
    .ssb(net1596));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_14__u_gpio_u_reg_u_data_in_q_reg_23_ (.rb(net529),
    .clk(clknet_leaf_6_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[14]),
    .d2(net237),
    .o1(u_gpio_u_reg_data_in_qs[14]),
    .o2(u_gpio_u_reg_data_in_qs[23]),
    .si1(net1030),
    .si2(net1031),
    .ssb(net1597));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_15__u_gpio_u_reg_u_data_in_q_reg_16_ (.rb(net520),
    .clk(clknet_leaf_2_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[15]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[16]),
    .o1(u_gpio_u_reg_data_in_qs[15]),
    .o2(u_gpio_u_reg_data_in_qs[16]),
    .si1(net1032),
    .si2(net1033),
    .ssb(net1598));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_17__u_gpio_u_reg_u_data_in_q_reg_18_ (.rb(net524),
    .clk(clknet_leaf_8_clk_i),
    .d1(net238),
    .d2(u_gpio_u_reg_u_data_in_wr_data[18]),
    .o1(u_gpio_u_reg_data_in_qs[17]),
    .o2(u_gpio_u_reg_data_in_qs[18]),
    .si1(net1034),
    .si2(net1035),
    .ssb(net1599));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_19__u_gpio_u_reg_u_data_in_q_reg_20_ (.rb(net524),
    .clk(clknet_leaf_8_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[19]),
    .d2(net240),
    .o1(u_gpio_u_reg_data_in_qs[19]),
    .o2(u_gpio_u_reg_data_in_qs[20]),
    .si1(net1036),
    .si2(net1037),
    .ssb(net1600));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_21__u_gpio_u_reg_u_data_in_q_reg_22_ (.rb(net524),
    .clk(clknet_leaf_8_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[21]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[22]),
    .o1(u_gpio_u_reg_data_in_qs[21]),
    .o2(u_gpio_u_reg_data_in_qs[22]),
    .si1(net1038),
    .si2(net1039),
    .ssb(net1601));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_24__u_gpio_u_reg_u_data_in_q_reg_25_ (.rb(net528),
    .clk(clknet_leaf_6_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[24]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[25]),
    .o1(u_gpio_u_reg_data_in_qs[24]),
    .o2(u_gpio_u_reg_data_in_qs[25]),
    .si1(net1040),
    .si2(net1041),
    .ssb(net1602));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_26__u_gpio_u_reg_u_data_in_q_reg_28_ (.rb(net533),
    .clk(clknet_leaf_6_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[26]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[28]),
    .o1(u_gpio_u_reg_data_in_qs[26]),
    .o2(u_gpio_u_reg_data_in_qs[28]),
    .si1(net1042),
    .si2(net1043),
    .ssb(net1603));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_27__u_gpio_u_reg_u_data_in_q_reg_30_ (.rb(net534),
    .clk(clknet_leaf_6_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[27]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[30]),
    .o1(u_gpio_u_reg_data_in_qs[27]),
    .o2(u_gpio_u_reg_data_in_qs[30]),
    .si1(net1044),
    .si2(net1045),
    .ssb(net1604));
 b15fqy003ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_29_ (.rb(net528),
    .clk(clknet_leaf_7_clk_i),
    .d(u_gpio_u_reg_u_data_in_wr_data[29]),
    .o(u_gpio_u_reg_data_in_qs[29]),
    .si(net1046),
    .ssb(net1605));
 b15fqy003ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_31_ (.rb(net533),
    .clk(clknet_leaf_5_clk_i),
    .d(u_gpio_u_reg_u_data_in_wr_data[31]),
    .o(u_gpio_u_reg_data_in_qs[31]),
    .si(net1047),
    .ssb(net1606));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_3__u_gpio_u_reg_u_data_in_q_reg_4_ (.rb(net512),
    .clk(clknet_leaf_9_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[3]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[4]),
    .o1(u_gpio_u_reg_data_in_qs[3]),
    .o2(u_gpio_u_reg_data_in_qs[4]),
    .si1(net1048),
    .si2(net1049),
    .ssb(net1607));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_5__u_gpio_u_reg_u_data_in_q_reg_12_ (.rb(net513),
    .clk(clknet_leaf_9_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[5]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[12]),
    .o1(u_gpio_u_reg_data_in_qs[5]),
    .o2(u_gpio_u_reg_data_in_qs[12]),
    .si1(net1050),
    .si2(net1051),
    .ssb(net1608));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_6__u_gpio_u_reg_u_data_in_q_reg_7_ (.rb(net510),
    .clk(clknet_leaf_11_clk_i),
    .d1(net241),
    .d2(u_gpio_u_reg_u_data_in_wr_data[7]),
    .o1(u_gpio_u_reg_data_in_qs[6]),
    .o2(u_gpio_u_reg_data_in_qs[7]),
    .si1(net1052),
    .si2(net1053),
    .ssb(net1609));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_8__u_gpio_u_reg_u_data_in_q_reg_11_ (.rb(net520),
    .clk(clknet_leaf_2_clk_i),
    .d1(u_gpio_u_reg_u_data_in_wr_data[8]),
    .d2(u_gpio_u_reg_u_data_in_wr_data[11]),
    .o1(u_gpio_u_reg_data_in_qs[8]),
    .o2(u_gpio_u_reg_data_in_qs[11]),
    .si1(net1054),
    .si2(net1055),
    .ssb(net1610));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_data_in_q_reg_9__u_gpio_u_reg_u_data_in_q_reg_10_ (.rb(net529),
    .clk(clknet_leaf_2_clk_i),
    .d1(net239),
    .d2(u_gpio_u_reg_u_data_in_wr_data[10]),
    .o1(u_gpio_u_reg_data_in_qs[9]),
    .o2(u_gpio_u_reg_data_in_qs[10]),
    .si1(net1056),
    .si2(net1057),
    .ssb(net1611));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_intr_ctrl_en_falling_clk_gate_q_reg_0_latch (.clk(clknet_leaf_8_clk_i),
    .clkout(u_gpio_u_reg_u_intr_ctrl_en_falling_net3627),
    .en(n3940),
    .te(net1058));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_intr_ctrl_en_falling_clk_gate_q_reg_latch (.clk(clknet_leaf_10_clk_i),
    .clkout(u_gpio_u_reg_u_intr_ctrl_en_falling_net3621),
    .en(n3940),
    .te(net1059));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_1_ (.rb(net511),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[0]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[1]),
    .o1(u_gpio_reg2hw[96]),
    .o2(u_gpio_reg2hw[97]),
    .si1(net1060),
    .si2(net1061),
    .ssb(net1612));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_11_ (.rb(net511),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[10]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[11]),
    .o1(u_gpio_reg2hw[106]),
    .o2(u_gpio_reg2hw[107]),
    .si1(net1062),
    .si2(net1063),
    .ssb(net1613));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_13_ (.rb(net512),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[12]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[13]),
    .o1(u_gpio_reg2hw[108]),
    .o2(u_gpio_reg2hw[109]),
    .si1(net1064),
    .si2(net1065),
    .ssb(net1614));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_15_ (.rb(net512),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[14]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[15]),
    .o1(u_gpio_reg2hw[110]),
    .o2(u_gpio_reg2hw[111]),
    .si1(net1066),
    .si2(net1067),
    .ssb(net1615));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_17_ (.rb(net524),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[16]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[17]),
    .o1(u_gpio_reg2hw[112]),
    .o2(u_gpio_reg2hw[113]),
    .si1(net1068),
    .si2(net1069),
    .ssb(net1616));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_19_ (.rb(net524),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[18]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[19]),
    .o1(u_gpio_reg2hw[114]),
    .o2(u_gpio_reg2hw[115]),
    .si1(net1070),
    .si2(net1071),
    .ssb(net1617));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_21_ (.rb(net524),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[20]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[21]),
    .o1(u_gpio_reg2hw[116]),
    .o2(u_gpio_reg2hw[117]),
    .si1(net1072),
    .si2(net1073),
    .ssb(net1618));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_23_ (.rb(net524),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[22]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[23]),
    .o1(u_gpio_reg2hw[118]),
    .o2(u_gpio_reg2hw[119]),
    .si1(net1074),
    .si2(net1075),
    .ssb(net1619));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_25_ (.rb(net527),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[24]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[25]),
    .o1(u_gpio_reg2hw[120]),
    .o2(u_gpio_reg2hw[121]),
    .si1(net1076),
    .si2(net1077),
    .ssb(net1620));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_27_ (.rb(net527),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[26]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[27]),
    .o1(u_gpio_reg2hw[122]),
    .o2(u_gpio_reg2hw[123]),
    .si1(net1078),
    .si2(net1079),
    .ssb(net1621));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_29_ (.rb(net527),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[28]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[29]),
    .o1(u_gpio_reg2hw[124]),
    .o2(u_gpio_reg2hw[125]),
    .si1(net1080),
    .si2(net1081),
    .ssb(net1622));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_3_ (.rb(net512),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[2]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[3]),
    .o1(u_gpio_reg2hw[98]),
    .o2(u_gpio_reg2hw[99]),
    .si1(net1082),
    .si2(net1083),
    .ssb(net1623));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_31_ (.rb(net527),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[30]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[31]),
    .o1(u_gpio_reg2hw[126]),
    .o2(u_gpio_reg2hw[127]),
    .si1(net1084),
    .si2(net1085),
    .ssb(net1624));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_5_ (.rb(net511),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[4]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[5]),
    .o1(u_gpio_reg2hw[100]),
    .o2(u_gpio_reg2hw[101]),
    .si1(net1086),
    .si2(net1087),
    .ssb(net1625));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_7_ (.rb(net511),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[6]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[7]),
    .o1(u_gpio_reg2hw[102]),
    .o2(u_gpio_reg2hw[103]),
    .si1(net1088),
    .si2(net1089),
    .ssb(net1626));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_9_ (.rb(net512),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[8]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_falling_wr_data[9]),
    .o1(u_gpio_reg2hw[104]),
    .o2(u_gpio_reg2hw[105]),
    .si1(net1090),
    .si2(net1091),
    .ssb(net1627));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_clk_gate_q_reg_0_latch (.clk(clknet_leaf_7_clk_i),
    .clkout(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627),
    .en(n3943),
    .te(net1092));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_clk_gate_q_reg_latch (.clk(clknet_leaf_10_clk_i),
    .clkout(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621),
    .en(net197),
    .te(net1093));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_1_ (.rb(net510),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[0]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[1]),
    .o1(u_gpio_reg2hw[64]),
    .o2(u_gpio_reg2hw[65]),
    .si1(net1094),
    .si2(net1095),
    .ssb(net1628));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_11_ (.rb(net510),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[10]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[11]),
    .o1(u_gpio_reg2hw[74]),
    .o2(u_gpio_reg2hw[75]),
    .si1(net1096),
    .si2(net1097),
    .ssb(net1629));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_13_ (.rb(net542),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[12]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[13]),
    .o1(u_gpio_reg2hw[76]),
    .o2(u_gpio_reg2hw[77]),
    .si1(net1098),
    .si2(net1099),
    .ssb(net1630));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_15_ (.rb(net542),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[14]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[15]),
    .o1(u_gpio_reg2hw[78]),
    .o2(u_gpio_reg2hw[79]),
    .si1(net1100),
    .si2(net1101),
    .ssb(net1631));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_17_ (.rb(net528),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[16]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[17]),
    .o1(u_gpio_reg2hw[80]),
    .o2(u_gpio_reg2hw[81]),
    .si1(net1102),
    .si2(net1103),
    .ssb(net1632));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_19_ (.rb(net528),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[18]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[19]),
    .o1(u_gpio_reg2hw[82]),
    .o2(u_gpio_reg2hw[83]),
    .si1(net1104),
    .si2(net1105),
    .ssb(net1633));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_21_ (.rb(net528),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[20]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[21]),
    .o1(u_gpio_reg2hw[84]),
    .o2(u_gpio_reg2hw[85]),
    .si1(net1106),
    .si2(net1107),
    .ssb(net1634));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_23_ (.rb(net528),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[22]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[23]),
    .o1(u_gpio_reg2hw[86]),
    .o2(u_gpio_reg2hw[87]),
    .si1(net1108),
    .si2(net1109),
    .ssb(net1635));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_25_ (.rb(net528),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[24]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[25]),
    .o1(u_gpio_reg2hw[88]),
    .o2(u_gpio_reg2hw[89]),
    .si1(net1110),
    .si2(net1111),
    .ssb(net1636));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_27_ (.rb(net528),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[26]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[27]),
    .o1(u_gpio_reg2hw[90]),
    .o2(u_gpio_reg2hw[91]),
    .si1(net1112),
    .si2(net1113),
    .ssb(net1637));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_29_ (.rb(net539),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[28]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[29]),
    .o1(u_gpio_reg2hw[92]),
    .o2(u_gpio_reg2hw[93]),
    .si1(net1114),
    .si2(net1115),
    .ssb(net1638));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_3_ (.rb(net542),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[2]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[3]),
    .o1(u_gpio_reg2hw[66]),
    .o2(u_gpio_reg2hw[67]),
    .si1(net1116),
    .si2(net1117),
    .ssb(net1639));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_31_ (.rb(net539),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[30]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[31]),
    .o1(u_gpio_reg2hw[94]),
    .o2(u_gpio_reg2hw[95]),
    .si1(net1118),
    .si2(net1119),
    .ssb(net1640));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_5_ (.rb(net511),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[4]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[5]),
    .o1(u_gpio_reg2hw[68]),
    .o2(u_gpio_reg2hw[69]),
    .si1(net1120),
    .si2(net1121),
    .ssb(net1641));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_7_ (.rb(net511),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[6]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[7]),
    .o1(u_gpio_reg2hw[70]),
    .o2(u_gpio_reg2hw[71]),
    .si1(net1122),
    .si2(net1123),
    .ssb(net1642));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_9_ (.rb(net511),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[8]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_wr_data[9]),
    .o1(u_gpio_reg2hw[72]),
    .o2(u_gpio_reg2hw[73]),
    .si1(net1124),
    .si2(net1125),
    .ssb(net1643));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_intr_ctrl_en_lvllow_clk_gate_q_reg_0_latch (.clk(clknet_leaf_7_clk_i),
    .clkout(u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627),
    .en(net179),
    .te(net1126));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_intr_ctrl_en_lvllow_clk_gate_q_reg_latch (.clk(clknet_leaf_10_clk_i),
    .clkout(u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621),
    .en(net179),
    .te(net1127));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_1_ (.rb(net512),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[0]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[1]),
    .o1(u_gpio_reg2hw[32]),
    .o2(u_gpio_reg2hw[33]),
    .si1(net1128),
    .si2(net1129),
    .ssb(net1644));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_11_ (.rb(net512),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[10]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[11]),
    .o1(u_gpio_reg2hw[42]),
    .o2(u_gpio_reg2hw[43]),
    .si1(net1130),
    .si2(net1131),
    .ssb(net1645));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_13_ (.rb(net514),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[12]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[13]),
    .o1(u_gpio_reg2hw[44]),
    .o2(u_gpio_reg2hw[45]),
    .si1(net1132),
    .si2(net1133),
    .ssb(net1646));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_15_ (.rb(net512),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[14]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[15]),
    .o1(u_gpio_reg2hw[46]),
    .o2(u_gpio_reg2hw[47]),
    .si1(net1134),
    .si2(net1135),
    .ssb(net1647));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_17_ (.rb(net527),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[16]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[17]),
    .o1(u_gpio_reg2hw[48]),
    .o2(u_gpio_reg2hw[49]),
    .si1(net1136),
    .si2(net1137),
    .ssb(net1648));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_19_ (.rb(net527),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[18]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[19]),
    .o1(u_gpio_reg2hw[50]),
    .o2(u_gpio_reg2hw[51]),
    .si1(net1138),
    .si2(net1139),
    .ssb(net1649));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_21_ (.rb(net527),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[20]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[21]),
    .o1(u_gpio_reg2hw[52]),
    .o2(u_gpio_reg2hw[53]),
    .si1(net1140),
    .si2(net1141),
    .ssb(net1650));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_23_ (.rb(net527),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[22]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[23]),
    .o1(u_gpio_reg2hw[54]),
    .o2(u_gpio_reg2hw[55]),
    .si1(net1142),
    .si2(net1143),
    .ssb(net1651));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_25_ (.rb(net527),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[24]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[25]),
    .o1(u_gpio_reg2hw[56]),
    .o2(u_gpio_reg2hw[57]),
    .si1(net1144),
    .si2(net1145),
    .ssb(net1652));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_27_ (.rb(net527),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[26]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[27]),
    .o1(u_gpio_reg2hw[58]),
    .o2(u_gpio_reg2hw[59]),
    .si1(net1146),
    .si2(net1147),
    .ssb(net1653));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_29_ (.rb(net528),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[28]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[29]),
    .o1(u_gpio_reg2hw[60]),
    .o2(u_gpio_reg2hw[61]),
    .si1(net1148),
    .si2(net1149),
    .ssb(net1654));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_3_ (.rb(net514),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[2]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[3]),
    .o1(u_gpio_reg2hw[34]),
    .o2(u_gpio_reg2hw[35]),
    .si1(net1150),
    .si2(net1151),
    .ssb(net1655));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_31_ (.rb(net527),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[30]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[31]),
    .o1(u_gpio_reg2hw[62]),
    .o2(u_gpio_reg2hw[63]),
    .si1(net1152),
    .si2(net1153),
    .ssb(net1656));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_5_ (.rb(net512),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[4]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[5]),
    .o1(u_gpio_reg2hw[36]),
    .o2(u_gpio_reg2hw[37]),
    .si1(net1154),
    .si2(net1155),
    .ssb(net1657));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_7_ (.rb(net512),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[6]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[7]),
    .o1(u_gpio_reg2hw[38]),
    .o2(u_gpio_reg2hw[39]),
    .si1(net1156),
    .si2(net1157),
    .ssb(net1658));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_9_ (.rb(net514),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[8]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_lvllow_wr_data[9]),
    .o1(u_gpio_reg2hw[40]),
    .o2(u_gpio_reg2hw[41]),
    .si1(net1158),
    .si2(net1159),
    .ssb(net1659));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_intr_ctrl_en_rising_clk_gate_q_reg_0_latch (.clk(clknet_leaf_8_clk_i),
    .clkout(u_gpio_u_reg_u_intr_ctrl_en_rising_net3627),
    .en(n3941),
    .te(net1160));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_intr_ctrl_en_rising_clk_gate_q_reg_latch (.clk(clknet_leaf_10_clk_i),
    .clkout(u_gpio_u_reg_u_intr_ctrl_en_rising_net3621),
    .en(n3941),
    .te(net1161));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_1_ (.rb(net511),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[0]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[1]),
    .o1(u_gpio_reg2hw[128]),
    .o2(u_gpio_reg2hw[129]),
    .si1(net1162),
    .si2(net1163),
    .ssb(net1660));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_11_ (.rb(net512),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[10]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[11]),
    .o1(u_gpio_reg2hw[138]),
    .o2(u_gpio_reg2hw[139]),
    .si1(net1164),
    .si2(net1165),
    .ssb(net1661));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_13_ (.rb(net512),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[12]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[13]),
    .o1(u_gpio_reg2hw[140]),
    .o2(u_gpio_reg2hw[141]),
    .si1(net1166),
    .si2(net1167),
    .ssb(net1662));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_15_ (.rb(net511),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[14]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[15]),
    .o1(u_gpio_reg2hw[142]),
    .o2(u_gpio_reg2hw[143]),
    .si1(net1168),
    .si2(net1169),
    .ssb(net1663));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_17_ (.rb(net526),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[16]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[17]),
    .o1(u_gpio_reg2hw[144]),
    .o2(u_gpio_reg2hw[145]),
    .si1(net1170),
    .si2(net1171),
    .ssb(net1664));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_19_ (.rb(net526),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[18]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[19]),
    .o1(u_gpio_reg2hw[146]),
    .o2(u_gpio_reg2hw[147]),
    .si1(net1172),
    .si2(net1173),
    .ssb(net1665));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_21_ (.rb(net526),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[20]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[21]),
    .o1(u_gpio_reg2hw[148]),
    .o2(u_gpio_reg2hw[149]),
    .si1(net1174),
    .si2(net1175),
    .ssb(net1666));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_23_ (.rb(net526),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[22]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[23]),
    .o1(u_gpio_reg2hw[150]),
    .o2(u_gpio_reg2hw[151]),
    .si1(net1176),
    .si2(net1177),
    .ssb(net1667));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_25_ (.rb(net527),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[24]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[25]),
    .o1(u_gpio_reg2hw[152]),
    .o2(u_gpio_reg2hw[153]),
    .si1(net1178),
    .si2(net1179),
    .ssb(net1668));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_27_ (.rb(net527),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[26]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[27]),
    .o1(u_gpio_reg2hw[154]),
    .o2(u_gpio_reg2hw[155]),
    .si1(net1180),
    .si2(net1181),
    .ssb(net1669));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_29_ (.rb(net527),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[28]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[29]),
    .o1(u_gpio_reg2hw[156]),
    .o2(u_gpio_reg2hw[157]),
    .si1(net1182),
    .si2(net1183),
    .ssb(net1670));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_3_ (.rb(net511),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[2]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[3]),
    .o1(u_gpio_reg2hw[130]),
    .o2(u_gpio_reg2hw[131]),
    .si1(net1184),
    .si2(net1185),
    .ssb(net1671));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_31_ (.rb(net527),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[30]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[31]),
    .o1(u_gpio_reg2hw[158]),
    .o2(u_gpio_reg2hw[159]),
    .si1(net1186),
    .si2(net1187),
    .ssb(net1672));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_5_ (.rb(net512),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[4]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[5]),
    .o1(u_gpio_reg2hw[132]),
    .o2(u_gpio_reg2hw[133]),
    .si1(net1188),
    .si2(net1189),
    .ssb(net1673));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_7_ (.rb(net511),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[6]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[7]),
    .o1(u_gpio_reg2hw[134]),
    .o2(u_gpio_reg2hw[135]),
    .si1(net1190),
    .si2(net1191),
    .ssb(net1674));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_9_ (.rb(net512),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621),
    .d1(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[8]),
    .d2(u_gpio_u_reg_u_intr_ctrl_en_rising_wr_data[9]),
    .o1(u_gpio_reg2hw[136]),
    .o2(u_gpio_reg2hw[137]),
    .si1(net1192),
    .si2(net1193),
    .ssb(net1675));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_intr_enable_clk_gate_q_reg_0_latch (.clk(clknet_leaf_6_clk_i),
    .clkout(u_gpio_u_reg_u_intr_enable_net3627),
    .en(n3939),
    .te(net1194));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_intr_enable_clk_gate_q_reg_latch (.clk(clknet_leaf_11_clk_i),
    .clkout(u_gpio_u_reg_u_intr_enable_net3621),
    .en(n3939),
    .te(net1195));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_0__u_gpio_u_reg_u_intr_enable_q_reg_1_ (.rb(net519),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_enable_net3621),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[0]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[1]),
    .o1(u_gpio_reg2hw[160]),
    .o2(u_gpio_reg2hw[161]),
    .si1(net1196),
    .si2(net1197),
    .ssb(net1676));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_10__u_gpio_u_reg_u_intr_enable_q_reg_11_ (.rb(net519),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_enable_net3621),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[10]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[11]),
    .o1(u_gpio_reg2hw[170]),
    .o2(u_gpio_reg2hw[171]),
    .si1(net1198),
    .si2(net1199),
    .ssb(net1677));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_12__u_gpio_u_reg_u_intr_enable_q_reg_13_ (.rb(net513),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_enable_net3621),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[12]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[13]),
    .o1(u_gpio_reg2hw[172]),
    .o2(u_gpio_reg2hw[173]),
    .si1(net1200),
    .si2(net1201),
    .ssb(net1678));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_14__u_gpio_u_reg_u_intr_enable_q_reg_15_ (.rb(net519),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_enable_net3621),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[14]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[15]),
    .o1(u_gpio_reg2hw[174]),
    .o2(u_gpio_reg2hw[175]),
    .si1(net1202),
    .si2(net1203),
    .ssb(net1679));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_16__u_gpio_u_reg_u_intr_enable_q_reg_17_ (.rb(net529),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_enable_net3627),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[16]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[17]),
    .o1(u_gpio_reg2hw[176]),
    .o2(u_gpio_reg2hw[177]),
    .si1(net1204),
    .si2(net1205),
    .ssb(net1680));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_18__u_gpio_u_reg_u_intr_enable_q_reg_19_ (.rb(net525),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_enable_net3627),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[18]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[19]),
    .o1(u_gpio_reg2hw[178]),
    .o2(u_gpio_reg2hw[179]),
    .si1(net1206),
    .si2(net1207),
    .ssb(net1681));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_20__u_gpio_u_reg_u_intr_enable_q_reg_21_ (.rb(net525),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_enable_net3627),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[20]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[21]),
    .o1(u_gpio_reg2hw[180]),
    .o2(u_gpio_reg2hw[181]),
    .si1(net1208),
    .si2(net1209),
    .ssb(net1682));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_22__u_gpio_u_reg_u_intr_enable_q_reg_23_ (.rb(net525),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_enable_net3627),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[22]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[23]),
    .o1(u_gpio_reg2hw[182]),
    .o2(u_gpio_reg2hw[183]),
    .si1(net1210),
    .si2(net1211),
    .ssb(net1683));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_24__u_gpio_u_reg_u_intr_enable_q_reg_25_ (.rb(net530),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_enable_net3627),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[24]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[25]),
    .o1(u_gpio_reg2hw[184]),
    .o2(u_gpio_reg2hw[185]),
    .si1(net1212),
    .si2(net1213),
    .ssb(net1684));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_26__u_gpio_u_reg_u_intr_enable_q_reg_27_ (.rb(net530),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_enable_net3627),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[26]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[27]),
    .o1(u_gpio_reg2hw[186]),
    .o2(u_gpio_reg2hw[187]),
    .si1(net1214),
    .si2(net1215),
    .ssb(net1685));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_28__u_gpio_u_reg_u_intr_enable_q_reg_29_ (.rb(net525),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_enable_net3627),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[28]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[29]),
    .o1(u_gpio_reg2hw[188]),
    .o2(u_gpio_reg2hw[189]),
    .si1(net1216),
    .si2(net1217),
    .ssb(net1686));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_2__u_gpio_u_reg_u_intr_enable_q_reg_3_ (.rb(net513),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_enable_net3621),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[2]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[3]),
    .o1(u_gpio_reg2hw[162]),
    .o2(u_gpio_reg2hw[163]),
    .si1(net1218),
    .si2(net1219),
    .ssb(net1687));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_30__u_gpio_u_reg_u_intr_enable_q_reg_31_ (.rb(net529),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_enable_net3627),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[30]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[31]),
    .o1(u_gpio_reg2hw[190]),
    .o2(u_gpio_reg2hw[191]),
    .si1(net1220),
    .si2(net1221),
    .ssb(net1688));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_4__u_gpio_u_reg_u_intr_enable_q_reg_5_ (.rb(net513),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_enable_net3621),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[4]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[5]),
    .o1(u_gpio_reg2hw[164]),
    .o2(u_gpio_reg2hw[165]),
    .si1(net1222),
    .si2(net1223),
    .ssb(net1689));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_6__u_gpio_u_reg_u_intr_enable_q_reg_7_ (.rb(net513),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_enable_net3621),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[6]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[7]),
    .o1(u_gpio_reg2hw[166]),
    .o2(u_gpio_reg2hw[167]),
    .si1(net1224),
    .si2(net1225),
    .ssb(net1690));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_enable_q_reg_8__u_gpio_u_reg_u_intr_enable_q_reg_9_ (.rb(net519),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_enable_net3621),
    .d1(u_gpio_u_reg_u_intr_enable_wr_data[8]),
    .d2(u_gpio_u_reg_u_intr_enable_wr_data[9]),
    .o1(u_gpio_reg2hw[168]),
    .o2(u_gpio_reg2hw[169]),
    .si1(net1226),
    .si2(net1227),
    .ssb(net1691));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_intr_state_clk_gate_q_reg_0_latch (.clk(clknet_leaf_6_clk_i),
    .clkout(u_gpio_u_reg_u_intr_state_net3650),
    .en(u_gpio_u_reg_u_intr_state_n1),
    .te(net1228));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_intr_state_clk_gate_q_reg_latch (.clk(clknet_leaf_9_clk_i),
    .clkout(u_gpio_u_reg_u_intr_state_net3644),
    .en(u_gpio_u_reg_u_intr_state_n1),
    .te(net1229));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_0__u_gpio_u_reg_u_intr_state_q_reg_1_ (.rb(net513),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_state_net3644),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[0]),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[1]),
    .o1(u_gpio_reg2hw[192]),
    .o2(u_gpio_reg2hw[193]),
    .si1(net1230),
    .si2(net1231),
    .ssb(net1692));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_10__u_gpio_u_reg_u_intr_state_q_reg_11_ (.rb(net513),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_state_net3644),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[10]),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[11]),
    .o1(u_gpio_reg2hw[202]),
    .o2(u_gpio_reg2hw[203]),
    .si1(net1232),
    .si2(net1233),
    .ssb(net1693));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_12__u_gpio_u_reg_u_intr_state_q_reg_13_ (.rb(net514),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_state_net3644),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[12]),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[13]),
    .o1(u_gpio_reg2hw[204]),
    .o2(u_gpio_reg2hw[205]),
    .si1(net1234),
    .si2(net1235),
    .ssb(net1694));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_14__u_gpio_u_reg_u_intr_state_q_reg_15_ (.rb(net514),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_state_net3644),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[14]),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[15]),
    .o1(u_gpio_reg2hw[206]),
    .o2(u_gpio_reg2hw[207]),
    .si1(net1236),
    .si2(net1237),
    .ssb(net1695));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_16__u_gpio_u_reg_u_intr_state_q_reg_17_ (.rb(net525),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_state_net3650),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[16]),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[17]),
    .o1(u_gpio_reg2hw[208]),
    .o2(u_gpio_reg2hw[209]),
    .si1(net1238),
    .si2(net1239),
    .ssb(net1696));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_18__u_gpio_u_reg_u_intr_state_q_reg_19_ (.rb(net526),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_state_net3650),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[18]),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[19]),
    .o1(u_gpio_reg2hw[210]),
    .o2(u_gpio_reg2hw[211]),
    .si1(net1240),
    .si2(net1241),
    .ssb(net1697));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_20__u_gpio_u_reg_u_intr_state_q_reg_21_ (.rb(net526),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_state_net3650),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[20]),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[21]),
    .o1(u_gpio_reg2hw[212]),
    .o2(u_gpio_reg2hw[213]),
    .si1(net1242),
    .si2(net1243),
    .ssb(net1698));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_22__u_gpio_u_reg_u_intr_state_q_reg_23_ (.rb(net526),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_state_net3650),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[22]),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[23]),
    .o1(u_gpio_reg2hw[214]),
    .o2(u_gpio_reg2hw[215]),
    .si1(net1244),
    .si2(net1245),
    .ssb(net1699));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_24__u_gpio_u_reg_u_intr_state_q_reg_25_ (.rb(net526),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_state_net3650),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[24]),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[25]),
    .o1(u_gpio_reg2hw[216]),
    .o2(u_gpio_reg2hw[217]),
    .si1(net1246),
    .si2(net1247),
    .ssb(net1700));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_26__u_gpio_u_reg_u_intr_state_q_reg_27_ (.rb(net526),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_state_net3650),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[26]),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[27]),
    .o1(u_gpio_reg2hw[218]),
    .o2(u_gpio_reg2hw[219]),
    .si1(net1248),
    .si2(net1249),
    .ssb(net1701));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_28__u_gpio_u_reg_u_intr_state_q_reg_29_ (.rb(net526),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_state_net3650),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[28]),
    .d2(net1967),
    .o1(u_gpio_reg2hw[220]),
    .o2(u_gpio_reg2hw[221]),
    .si1(net1250),
    .si2(net1251),
    .ssb(net1702));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_2__u_gpio_u_reg_u_intr_state_q_reg_3_ (.rb(net525),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_state_net3644),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[2]),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[3]),
    .o1(u_gpio_reg2hw[194]),
    .o2(u_gpio_reg2hw[195]),
    .si1(net1252),
    .si2(net1253),
    .ssb(net1703));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_30__u_gpio_u_reg_u_intr_state_q_reg_31_ (.rb(net526),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_state_net3650),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[30]),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[31]),
    .o1(u_gpio_reg2hw[222]),
    .o2(u_gpio_reg2hw[223]),
    .si1(net1254),
    .si2(net1255),
    .ssb(net1704));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_4__u_gpio_u_reg_u_intr_state_q_reg_5_ (.rb(net514),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_state_net3644),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[4]),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[5]),
    .o1(u_gpio_reg2hw[196]),
    .o2(u_gpio_reg2hw[197]),
    .si1(net1256),
    .si2(net1257),
    .ssb(net1705));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_6__u_gpio_u_reg_u_intr_state_q_reg_7_ (.rb(net514),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_intr_state_net3644),
    .d1(net2154),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[7]),
    .o1(u_gpio_reg2hw[198]),
    .o2(u_gpio_reg2hw[199]),
    .si1(net1258),
    .si2(net1259),
    .ssb(net1706));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_intr_state_q_reg_8__u_gpio_u_reg_u_intr_state_q_reg_9_ (.rb(net525),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_intr_state_net3644),
    .d1(u_gpio_u_reg_u_intr_state_wr_data[8]),
    .d2(u_gpio_u_reg_u_intr_state_wr_data[9]),
    .o1(u_gpio_reg2hw[200]),
    .o2(u_gpio_reg2hw[201]),
    .si1(net1260),
    .si2(net1261),
    .ssb(net1707));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_reg_if_clk_gate_rdata_reg_0_latch (.clk(clknet_leaf_2_clk_i),
    .clkout(u_gpio_u_reg_u_reg_if_net3678),
    .en(n3831),
    .te(net1262));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_reg_if_clk_gate_rdata_reg_latch (.clk(clknet_leaf_1_clk_i),
    .clkout(u_gpio_u_reg_u_reg_if_net3673),
    .en(n3831),
    .te(net1263));
 b15cilb05ah1n02x3 u_gpio_u_reg_u_reg_if_clk_gate_reqid_reg_latch (.clk(clknet_leaf_1_clk_i),
    .clkout(u_gpio_u_reg_u_reg_if_net3667),
    .en(n3831),
    .te(net1264));
 b15fqy043ar1n02x5 u_gpio_u_reg_u_reg_if_error_reg (.clk(clknet_leaf_1_clk_i),
    .d(u_gpio_u_reg_u_reg_if_N46),
    .den(n3831),
    .o(u_xbar_periph_u_s1n_6_tl_u_i[10]),
    .rb(net517),
    .si(net1265),
    .ssb(net1708));
 b15fqy043ar1n02x5 u_gpio_u_reg_u_reg_if_outstanding_reg (.clk(clknet_leaf_1_clk_i),
    .d(n3831),
    .den(u_gpio_u_reg_u_reg_if_N7),
    .o(u_xbar_periph_u_s1n_6_tl_u_i[24]),
    .rb(net517),
    .si(net1266),
    .ssb(net1709));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_0__u_gpio_u_reg_u_reg_if_rdata_reg_1_ (.rb(net522),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3673),
    .d1(u_gpio_u_reg_u_reg_if_N14),
    .d2(u_gpio_u_reg_u_reg_if_N15),
    .o1(gpio_2_xbar[0]),
    .o2(gpio_2_xbar[1]),
    .si1(net1267),
    .si2(net1268),
    .ssb(net1710));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_10__u_gpio_u_reg_u_reg_if_rdata_reg_11_ (.rb(net522),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3673),
    .d1(u_gpio_u_reg_u_reg_if_N24),
    .d2(u_gpio_u_reg_u_reg_if_N25),
    .o1(gpio_2_xbar[10]),
    .o2(gpio_2_xbar[11]),
    .si1(net1269),
    .si2(net1270),
    .ssb(net1711));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_12__u_gpio_u_reg_u_reg_if_rdata_reg_13_ (.rb(net522),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3673),
    .d1(u_gpio_u_reg_u_reg_if_N26),
    .d2(u_gpio_u_reg_u_reg_if_N27),
    .o1(gpio_2_xbar[12]),
    .o2(gpio_2_xbar[13]),
    .si1(net1271),
    .si2(net1272),
    .ssb(net1712));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_14__u_gpio_u_reg_u_reg_if_rdata_reg_15_ (.rb(net522),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3673),
    .d1(u_gpio_u_reg_u_reg_if_N28),
    .d2(u_gpio_u_reg_u_reg_if_N29),
    .o1(gpio_2_xbar[14]),
    .o2(gpio_2_xbar[15]),
    .si1(net1273),
    .si2(net1274),
    .ssb(net1713));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_16__u_gpio_u_reg_u_reg_if_rdata_reg_17_ (.rb(net531),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3678),
    .d1(u_gpio_u_reg_u_reg_if_N30),
    .d2(u_gpio_u_reg_u_reg_if_N31),
    .o1(gpio_2_xbar[16]),
    .o2(gpio_2_xbar[17]),
    .si1(net1275),
    .si2(net1276),
    .ssb(net1714));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_18__u_gpio_u_reg_u_reg_if_rdata_reg_19_ (.rb(net531),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3678),
    .d1(u_gpio_u_reg_u_reg_if_N32),
    .d2(net177),
    .o1(gpio_2_xbar[18]),
    .o2(gpio_2_xbar[19]),
    .si1(net1277),
    .si2(net1278),
    .ssb(net1715));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_20__u_gpio_u_reg_u_reg_if_rdata_reg_21_ (.rb(net531),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3678),
    .d1(net185),
    .d2(net187),
    .o1(gpio_2_xbar[20]),
    .o2(gpio_2_xbar[21]),
    .si1(net1279),
    .si2(net1280),
    .ssb(net1716));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_22__u_gpio_u_reg_u_reg_if_rdata_reg_23_ (.rb(net531),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3678),
    .d1(u_gpio_u_reg_u_reg_if_N36),
    .d2(u_gpio_u_reg_u_reg_if_N37),
    .o1(gpio_2_xbar[22]),
    .o2(gpio_2_xbar[23]),
    .si1(net1281),
    .si2(net1282),
    .ssb(net1717));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_24__u_gpio_u_reg_u_reg_if_rdata_reg_25_ (.rb(net531),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3678),
    .d1(net186),
    .d2(net188),
    .o1(gpio_2_xbar[24]),
    .o2(gpio_2_xbar[25]),
    .si1(net1283),
    .si2(net1284),
    .ssb(net1718));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_26__u_gpio_u_reg_u_reg_if_rdata_reg_27_ (.rb(net531),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3678),
    .d1(u_gpio_u_reg_u_reg_if_N40),
    .d2(u_gpio_u_reg_u_reg_if_N41),
    .o1(gpio_2_xbar[26]),
    .o2(gpio_2_xbar[27]),
    .si1(net1285),
    .si2(net1286),
    .ssb(net1719));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_28__u_gpio_u_reg_u_reg_if_rdata_reg_29_ (.rb(net531),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3678),
    .d1(net176),
    .d2(net175),
    .o1(gpio_2_xbar[28]),
    .o2(gpio_2_xbar[29]),
    .si1(net1287),
    .si2(net1288),
    .ssb(net1720));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_2__u_gpio_u_reg_u_reg_if_rdata_reg_3_ (.rb(net522),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3673),
    .d1(net193),
    .d2(net192),
    .o1(gpio_2_xbar[2]),
    .o2(gpio_2_xbar[3]),
    .si1(net1289),
    .si2(net1290),
    .ssb(net1721));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_30__u_gpio_u_reg_u_reg_if_rdata_reg_31_ (.rb(net540),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3678),
    .d1(net178),
    .d2(u_gpio_u_reg_u_reg_if_N45),
    .o1(gpio_2_xbar[30]),
    .o2(gpio_2_xbar[31]),
    .si1(net1291),
    .si2(net1292),
    .ssb(net1722));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_4__u_gpio_u_reg_u_reg_if_rdata_reg_5_ (.rb(net523),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3673),
    .d1(net191),
    .d2(net190),
    .o1(gpio_2_xbar[4]),
    .o2(gpio_2_xbar[5]),
    .si1(net1293),
    .si2(net1294),
    .ssb(net1723));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_6__u_gpio_u_reg_u_reg_if_rdata_reg_7_ (.rb(net523),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3673),
    .d1(net189),
    .d2(u_gpio_u_reg_u_reg_if_N21),
    .o1(gpio_2_xbar[6]),
    .o2(gpio_2_xbar[7]),
    .si1(net1295),
    .si2(net1296),
    .ssb(net1724));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rdata_reg_8__u_gpio_u_reg_u_reg_if_rdata_reg_9_ (.rb(net523),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3673),
    .d1(u_gpio_u_reg_u_reg_if_N22),
    .d2(u_gpio_u_reg_u_reg_if_N23),
    .o1(gpio_2_xbar[8]),
    .o2(gpio_2_xbar[9]),
    .si1(net1297),
    .si2(net1298),
    .ssb(net1725));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_reqid_reg_0__u_gpio_u_reg_u_reg_if_reqid_reg_1_ (.rb(net521),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3667),
    .d1(net71),
    .d2(net72),
    .o1(u_xbar_periph_u_s1n_6_tl_u_i[11]),
    .o2(u_xbar_periph_u_s1n_6_tl_u_i[12]),
    .si1(net1299),
    .si2(net1300),
    .ssb(net1726));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_reqid_reg_2__u_gpio_u_reg_u_reg_if_reqid_reg_3_ (.rb(net521),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3667),
    .d1(net73),
    .d2(net74),
    .o1(u_xbar_periph_u_s1n_6_tl_u_i[13]),
    .o2(u_xbar_periph_u_s1n_6_tl_u_i[14]),
    .si1(net1301),
    .si2(net1302),
    .ssb(net1727));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_reqid_reg_4__u_gpio_u_reg_u_reg_if_reqid_reg_5_ (.rb(net521),
    .clk(clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3667),
    .d1(net75),
    .d2(net76),
    .o1(u_xbar_periph_u_s1n_6_tl_u_i[15]),
    .o2(u_xbar_periph_u_s1n_6_tl_u_i[16]),
    .si1(net1303),
    .si2(net1304),
    .ssb(net1728));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_reqid_reg_6__u_gpio_u_reg_u_reg_if_reqid_reg_7_ (.rb(net521),
    .clk(clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3667),
    .d1(net77),
    .d2(net78),
    .o1(u_xbar_periph_u_s1n_6_tl_u_i[17]),
    .o2(u_xbar_periph_u_s1n_6_tl_u_i[18]),
    .si1(net1305),
    .si2(net1306),
    .ssb(net1729));
 b15fqy043ar1n02x5 u_gpio_u_reg_u_reg_if_reqsz_reg_0_ (.clk(clknet_leaf_1_clk_i),
    .d(net3),
    .den(n3831),
    .o(u_xbar_periph_u_s1n_6_tl_u_i[19]),
    .rb(net517),
    .si(net1307),
    .ssb(net1730));
 b15fqy043ar1n02x5 u_gpio_u_reg_u_reg_if_reqsz_reg_1_ (.clk(clknet_leaf_1_clk_i),
    .d(net4),
    .den(n3831),
    .o(u_xbar_periph_u_s1n_6_tl_u_i[20]),
    .rb(net517),
    .si(net1308),
    .ssb(net1731));
 b15fqy043ar1n02x5 u_gpio_u_reg_u_reg_if_rspop_reg_0_ (.clk(clknet_leaf_1_clk_i),
    .d(u_gpio_u_reg_u_reg_if_rd_req),
    .den(n3831),
    .o(u_xbar_periph_u_s1n_6_tl_u_i[21]),
    .rb(net517),
    .si(net1309),
    .ssb(net1732));
 b15fqy203ar1n02x5 u_gpio_u_reg_u_reg_if_rspop_reg_1__u_gpio_u_reg_u_reg_if_rspop_reg_2_ (.rb(net517),
    .clk(clknet_leaf_1_clk_i),
    .d1(n1527),
    .d2(n1530),
    .o1(u_xbar_periph_u_s1n_6_tl_u_i[22]),
    .o2(u_xbar_periph_u_s1n_6_tl_u_i[23]),
    .si1(net1310),
    .si2(net1311),
    .ssb(net1733));
 b15cilb05ah1n02x3 u_xbar_periph_u_s1n_6_clk_gate_num_req_outstanding_reg_latch (.clk(clknet_leaf_4_clk_i),
    .clkout(u_xbar_periph_u_s1n_6_net3695),
    .en(u_xbar_periph_u_s1n_6_N59),
    .te(net1312));
 b15fqy043ar1n02x5 u_xbar_periph_u_s1n_6_dev_select_outstanding_reg_0_ (.clk(clknet_leaf_1_clk_i),
    .d(u_xbar_periph_u_s1n_6_dev_select_t[0]),
    .den(net111),
    .o(u_xbar_periph_u_s1n_6_dev_select_outstanding[0]),
    .rb(net517),
    .si(net1313),
    .ssb(net1734));
 b15fqy043ar1n02x5 u_xbar_periph_u_s1n_6_dev_select_outstanding_reg_1_ (.clk(clknet_leaf_1_clk_i),
    .d(u_xbar_periph_u_s1n_6_dev_select_t[1]),
    .den(net111),
    .o(u_xbar_periph_u_s1n_6_dev_select_outstanding[1]),
    .rb(net517),
    .si(net1314),
    .ssb(net1735));
 b15fqy043ar1n02x5 u_xbar_periph_u_s1n_6_dev_select_outstanding_reg_2_ (.clk(clknet_leaf_1_clk_i),
    .d(u_xbar_periph_u_s1n_6_dev_select_t[2]),
    .den(net111),
    .o(u_xbar_periph_u_s1n_6_dev_select_outstanding[2]),
    .rb(net517),
    .si(net1315),
    .ssb(net1736));
 b15cilb05ah1n02x3 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_clk_gate_err_source_reg_latch (.clk(clknet_leaf_1_clk_i),
    .clkout(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713),
    .en(n3829),
    .te(net1316));
 b15fqy043ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type_reg_0_ (.clk(clknet_leaf_1_clk_i),
    .d(n1443),
    .den(n3829),
    .o(n1446),
    .rb(net516),
    .si(net1317),
    .ssb(net1737));
 b15fqy043ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type_reg_1_ (.clk(clknet_leaf_0_clk_i),
    .d(net10),
    .den(n3829),
    .o(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type[1]),
    .rb(net516),
    .si(net1318),
    .ssb(net1738));
 b15fqy043ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type_reg_2_ (.clk(clknet_leaf_1_clk_i),
    .d(net11),
    .den(n3829),
    .o(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type[2]),
    .rb(net516),
    .si(net1319),
    .ssb(net1739));
 b15fqy043ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type_reg_3_ (.clk(clknet_leaf_1_clk_i),
    .d(n1435),
    .den(n3829),
    .o(n1438),
    .rb(net516),
    .si(net1320),
    .ssb(net1740));
 b15fqy043ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_opcode_reg_0_ (.clk(clknet_leaf_1_clk_i),
    .d(net5),
    .den(n3829),
    .o(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_opcode[0]),
    .rb(net516),
    .si(net1321),
    .ssb(net1741));
 b15fqy043ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_opcode_reg_1_ (.clk(clknet_leaf_1_clk_i),
    .d(net6),
    .den(n3829),
    .o(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_opcode[1]),
    .rb(net516),
    .si(net1322),
    .ssb(net1742));
 b15fqy043ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_opcode_reg_2_ (.clk(clknet_leaf_1_clk_i),
    .d(n1451),
    .den(n3829),
    .o(n1454),
    .rb(net516),
    .si(net1323),
    .ssb(net1743));
 b15fqy043ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_req_pending_reg (.clk(clknet_leaf_1_clk_i),
    .d(n3829),
    .den(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_N8),
    .o(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_req_pending),
    .rb(net517),
    .si(net1324),
    .ssb(net1744));
 b15fqy003ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_rsp_pending_reg (.rb(net518),
    .clk(clknet_leaf_1_clk_i),
    .d(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_N12),
    .o(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_rsp_pending),
    .si(net1325),
    .ssb(net1745));
 b15fqy043ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_size_reg_0_ (.clk(clknet_leaf_1_clk_i),
    .d(net3),
    .den(n3829),
    .o(u_xbar_periph_u_s1n_6_tl_u_i[8]),
    .rb(net518),
    .si(net1326),
    .ssb(net1746));
 b15fqy043ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_size_reg_1_ (.clk(clknet_leaf_1_clk_i),
    .d(net4),
    .den(n3829),
    .o(u_xbar_periph_u_s1n_6_tl_u_i[9]),
    .rb(net518),
    .si(net1327),
    .ssb(net1747));
 b15fqy203ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_0__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_1_ (.rb(net521),
    .clk(clknet_1_0__leaf_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713),
    .d1(net71),
    .d2(net72),
    .o1(u_xbar_periph_u_s1n_6_tl_u_i[0]),
    .o2(u_xbar_periph_u_s1n_6_tl_u_i[1]),
    .si1(net1328),
    .si2(net1329),
    .ssb(net1748));
 b15fqy203ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_2__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_3_ (.rb(net521),
    .clk(clknet_1_1__leaf_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713),
    .d1(net73),
    .d2(net74),
    .o1(u_xbar_periph_u_s1n_6_tl_u_i[2]),
    .o2(u_xbar_periph_u_s1n_6_tl_u_i[3]),
    .si1(net1330),
    .si2(net1331),
    .ssb(net1749));
 b15fqy203ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_4__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_5_ (.rb(net521),
    .clk(clknet_1_0__leaf_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713),
    .d1(net75),
    .d2(net76),
    .o1(u_xbar_periph_u_s1n_6_tl_u_i[4]),
    .o2(u_xbar_periph_u_s1n_6_tl_u_i[5]),
    .si1(net1332),
    .si2(net1333),
    .ssb(net1750));
 b15fqy203ar1n02x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_6__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_7_ (.rb(net523),
    .clk(clknet_1_1__leaf_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713),
    .d1(net77),
    .d2(net78),
    .o1(u_xbar_periph_u_s1n_6_tl_u_i[6]),
    .o2(u_xbar_periph_u_s1n_6_tl_u_i[7]),
    .si1(net1334),
    .si2(net1335),
    .ssb(net1751));
 b15fqy203ar1n02x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_0__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_1_ (.rb(net532),
    .clk(clknet_1_1__leaf_u_xbar_periph_u_s1n_6_net3695),
    .d1(u_xbar_periph_u_s1n_6_N60),
    .d2(u_xbar_periph_u_s1n_6_N61),
    .o1(u_xbar_periph_u_s1n_6_num_req_outstanding[0]),
    .o2(u_xbar_periph_u_s1n_6_num_req_outstanding[1]),
    .si1(net1336),
    .si2(net1337),
    .ssb(net1752));
 b15fqy203ar1n02x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_2__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_3_ (.rb(net532),
    .clk(clknet_1_0__leaf_u_xbar_periph_u_s1n_6_net3695),
    .d1(u_xbar_periph_u_s1n_6_N62),
    .d2(u_xbar_periph_u_s1n_6_N63),
    .o1(u_xbar_periph_u_s1n_6_num_req_outstanding[2]),
    .o2(u_xbar_periph_u_s1n_6_num_req_outstanding[3]),
    .si1(net1338),
    .si2(net1339),
    .ssb(net1753));
 b15fqy203ar1n02x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_4__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_5_ (.rb(net532),
    .clk(clknet_1_0__leaf_u_xbar_periph_u_s1n_6_net3695),
    .d1(u_xbar_periph_u_s1n_6_N64),
    .d2(u_xbar_periph_u_s1n_6_N65),
    .o1(u_xbar_periph_u_s1n_6_num_req_outstanding[4]),
    .o2(u_xbar_periph_u_s1n_6_num_req_outstanding[5]),
    .si1(net1340),
    .si2(net1341),
    .ssb(net1754));
 b15fqy203ar1n02x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_6__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_7_ (.rb(net532),
    .clk(clknet_1_1__leaf_u_xbar_periph_u_s1n_6_net3695),
    .d1(u_xbar_periph_u_s1n_6_N66),
    .d2(u_xbar_periph_u_s1n_6_N67),
    .o1(u_xbar_periph_u_s1n_6_num_req_outstanding[6]),
    .o2(u_xbar_periph_u_s1n_6_num_req_outstanding[7]),
    .si1(net1342),
    .si2(net1343),
    .ssb(net1755));
 b15fqy003ar1n02x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_8_ (.rb(net538),
    .clk(clknet_1_1__leaf_u_xbar_periph_u_s1n_6_net3695),
    .d(u_xbar_periph_u_s1n_6_N68),
    .o(u_xbar_periph_u_s1n_6_num_req_outstanding[8]),
    .si(net1344),
    .ssb(net1756));
 b15tihi00an1n03x5 U3303_1345 (.o(net1345));
 b15cbf000an1n16x5 clkbuf_leaf_0_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_0_clk_i));
 b15ztpn00an1n08x5 PHY_95 ();
 b15ztpn00an1n08x5 PHY_96 ();
 b15ztpn00an1n08x5 PHY_97 ();
 b15ztpn00an1n08x5 PHY_98 ();
 b15ztpn00an1n08x5 PHY_99 ();
 b15ztpn00an1n08x5 PHY_100 ();
 b15ztpn00an1n08x5 PHY_101 ();
 b15ztpn00an1n08x5 PHY_102 ();
 b15ztpn00an1n08x5 PHY_103 ();
 b15ztpn00an1n08x5 PHY_104 ();
 b15ztpn00an1n08x5 PHY_105 ();
 b15ztpn00an1n08x5 PHY_106 ();
 b15ztpn00an1n08x5 PHY_107 ();
 b15ztpn00an1n08x5 PHY_108 ();
 b15ztpn00an1n08x5 PHY_109 ();
 b15ztpn00an1n08x5 PHY_110 ();
 b15ztpn00an1n08x5 PHY_111 ();
 b15ztpn00an1n08x5 PHY_112 ();
 b15ztpn00an1n08x5 PHY_113 ();
 b15ztpn00an1n08x5 PHY_114 ();
 b15ztpn00an1n08x5 PHY_115 ();
 b15ztpn00an1n08x5 PHY_116 ();
 b15ztpn00an1n08x5 PHY_117 ();
 b15ztpn00an1n08x5 PHY_118 ();
 b15ztpn00an1n08x5 PHY_119 ();
 b15ztpn00an1n08x5 PHY_120 ();
 b15ztpn00an1n08x5 PHY_121 ();
 b15ztpn00an1n08x5 PHY_122 ();
 b15ztpn00an1n08x5 PHY_123 ();
 b15ztpn00an1n08x5 PHY_124 ();
 b15ztpn00an1n08x5 PHY_125 ();
 b15ztpn00an1n08x5 PHY_126 ();
 b15ztpn00an1n08x5 PHY_127 ();
 b15ztpn00an1n08x5 PHY_128 ();
 b15ztpn00an1n08x5 PHY_129 ();
 b15ztpn00an1n08x5 PHY_130 ();
 b15ztpn00an1n08x5 PHY_131 ();
 b15ztpn00an1n08x5 PHY_132 ();
 b15ztpn00an1n08x5 PHY_133 ();
 b15ztpn00an1n08x5 PHY_134 ();
 b15ztpn00an1n08x5 PHY_135 ();
 b15ztpn00an1n08x5 PHY_136 ();
 b15ztpn00an1n08x5 PHY_137 ();
 b15ztpn00an1n08x5 PHY_138 ();
 b15ztpn00an1n08x5 PHY_139 ();
 b15ztpn00an1n08x5 PHY_140 ();
 b15ztpn00an1n08x5 PHY_141 ();
 b15ztpn00an1n08x5 PHY_142 ();
 b15ztpn00an1n08x5 PHY_143 ();
 b15ztpn00an1n08x5 PHY_144 ();
 b15ztpn00an1n08x5 PHY_145 ();
 b15ztpn00an1n08x5 PHY_146 ();
 b15ztpn00an1n08x5 PHY_147 ();
 b15ztpn00an1n08x5 PHY_148 ();
 b15ztpn00an1n08x5 PHY_149 ();
 b15ztpn00an1n08x5 PHY_150 ();
 b15ztpn00an1n08x5 PHY_151 ();
 b15ztpn00an1n08x5 PHY_152 ();
 b15ztpn00an1n08x5 PHY_153 ();
 b15ztpn00an1n08x5 PHY_154 ();
 b15ztpn00an1n08x5 PHY_155 ();
 b15ztpn00an1n08x5 PHY_156 ();
 b15ztpn00an1n08x5 PHY_157 ();
 b15ztpn00an1n08x5 PHY_158 ();
 b15ztpn00an1n08x5 PHY_159 ();
 b15ztpn00an1n08x5 PHY_160 ();
 b15ztpn00an1n08x5 PHY_161 ();
 b15ztpn00an1n08x5 PHY_162 ();
 b15ztpn00an1n08x5 PHY_163 ();
 b15ztpn00an1n08x5 PHY_164 ();
 b15ztpn00an1n08x5 PHY_165 ();
 b15ztpn00an1n08x5 PHY_166 ();
 b15ztpn00an1n08x5 PHY_167 ();
 b15ztpn00an1n08x5 PHY_168 ();
 b15ztpn00an1n08x5 PHY_169 ();
 b15ztpn00an1n08x5 PHY_170 ();
 b15ztpn00an1n08x5 PHY_171 ();
 b15ztpn00an1n08x5 PHY_172 ();
 b15ztpn00an1n08x5 PHY_173 ();
 b15ztpn00an1n08x5 PHY_174 ();
 b15ztpn00an1n08x5 PHY_175 ();
 b15ztpn00an1n08x5 PHY_176 ();
 b15ztpn00an1n08x5 PHY_177 ();
 b15ztpn00an1n08x5 PHY_178 ();
 b15ztpn00an1n08x5 PHY_179 ();
 b15ztpn00an1n08x5 PHY_180 ();
 b15ztpn00an1n08x5 PHY_181 ();
 b15ztpn00an1n08x5 PHY_182 ();
 b15ztpn00an1n08x5 PHY_183 ();
 b15ztpn00an1n08x5 PHY_184 ();
 b15ztpn00an1n08x5 PHY_185 ();
 b15ztpn00an1n08x5 PHY_186 ();
 b15ztpn00an1n08x5 PHY_187 ();
 b15ztpn00an1n08x5 PHY_188 ();
 b15ztpn00an1n08x5 PHY_189 ();
 b15ztpn00an1n08x5 PHY_190 ();
 b15ztpn00an1n08x5 PHY_191 ();
 b15ztpn00an1n08x5 PHY_192 ();
 b15ztpn00an1n08x5 PHY_193 ();
 b15ztpn00an1n08x5 PHY_194 ();
 b15ztpn00an1n08x5 PHY_195 ();
 b15ztpn00an1n08x5 PHY_196 ();
 b15ztpn00an1n08x5 PHY_197 ();
 b15ztpn00an1n08x5 PHY_198 ();
 b15ztpn00an1n08x5 PHY_199 ();
 b15ztpn00an1n08x5 PHY_200 ();
 b15ztpn00an1n08x5 PHY_201 ();
 b15ztpn00an1n08x5 PHY_202 ();
 b15ztpn00an1n08x5 PHY_203 ();
 b15ztpn00an1n08x5 PHY_204 ();
 b15ztpn00an1n08x5 PHY_205 ();
 b15ztpn00an1n08x5 PHY_206 ();
 b15ztpn00an1n08x5 PHY_207 ();
 b15ztpn00an1n08x5 PHY_208 ();
 b15ztpn00an1n08x5 PHY_209 ();
 b15ztpn00an1n08x5 PHY_210 ();
 b15ztpn00an1n08x5 PHY_211 ();
 b15ztpn00an1n08x5 PHY_212 ();
 b15ztpn00an1n08x5 PHY_213 ();
 b15ztpn00an1n08x5 PHY_214 ();
 b15ztpn00an1n08x5 PHY_215 ();
 b15ztpn00an1n08x5 PHY_216 ();
 b15ztpn00an1n08x5 PHY_217 ();
 b15ztpn00an1n08x5 PHY_218 ();
 b15ztpn00an1n08x5 PHY_219 ();
 b15ztpn00an1n08x5 PHY_220 ();
 b15ztpn00an1n08x5 PHY_221 ();
 b15ztpn00an1n08x5 PHY_222 ();
 b15ztpn00an1n08x5 PHY_223 ();
 b15ztpn00an1n08x5 PHY_224 ();
 b15ztpn00an1n08x5 PHY_225 ();
 b15ztpn00an1n08x5 PHY_226 ();
 b15ztpn00an1n08x5 PHY_227 ();
 b15ztpn00an1n08x5 PHY_228 ();
 b15ztpn00an1n08x5 PHY_229 ();
 b15ztpn00an1n08x5 PHY_230 ();
 b15ztpn00an1n08x5 PHY_231 ();
 b15ztpn00an1n08x5 PHY_232 ();
 b15ztpn00an1n08x5 PHY_233 ();
 b15ztpn00an1n08x5 PHY_234 ();
 b15ztpn00an1n08x5 PHY_235 ();
 b15ztpn00an1n08x5 PHY_236 ();
 b15ztpn00an1n08x5 PHY_237 ();
 b15ztpn00an1n08x5 PHY_238 ();
 b15ztpn00an1n08x5 PHY_239 ();
 b15ztpn00an1n08x5 PHY_240 ();
 b15ztpn00an1n08x5 PHY_241 ();
 b15ztpn00an1n08x5 PHY_242 ();
 b15ztpn00an1n08x5 PHY_243 ();
 b15ztpn00an1n08x5 PHY_244 ();
 b15ztpn00an1n08x5 PHY_245 ();
 b15ztpn00an1n08x5 PHY_246 ();
 b15ztpn00an1n08x5 PHY_247 ();
 b15ztpn00an1n08x5 PHY_248 ();
 b15ztpn00an1n08x5 PHY_249 ();
 b15ztpn00an1n08x5 PHY_250 ();
 b15ztpn00an1n08x5 PHY_251 ();
 b15ztpn00an1n08x5 PHY_252 ();
 b15ztpn00an1n08x5 PHY_253 ();
 b15ztpn00an1n08x5 PHY_254 ();
 b15ztpn00an1n08x5 PHY_255 ();
 b15ztpn00an1n08x5 PHY_256 ();
 b15ztpn00an1n08x5 PHY_257 ();
 b15ztpn00an1n08x5 PHY_258 ();
 b15ztpn00an1n08x5 PHY_259 ();
 b15ztpn00an1n08x5 PHY_260 ();
 b15ztpn00an1n08x5 PHY_261 ();
 b15ztpn00an1n08x5 PHY_262 ();
 b15ztpn00an1n08x5 PHY_263 ();
 b15ztpn00an1n08x5 PHY_264 ();
 b15ztpn00an1n08x5 PHY_265 ();
 b15ztpn00an1n08x5 PHY_266 ();
 b15ztpn00an1n08x5 PHY_267 ();
 b15ztpn00an1n08x5 PHY_268 ();
 b15ztpn00an1n08x5 PHY_269 ();
 b15ztpn00an1n08x5 PHY_270 ();
 b15ztpn00an1n08x5 PHY_271 ();
 b15ztpn00an1n08x5 PHY_272 ();
 b15ztpn00an1n08x5 PHY_273 ();
 b15ztpn00an1n08x5 PHY_274 ();
 b15ztpn00an1n08x5 PHY_275 ();
 b15ztpn00an1n08x5 PHY_276 ();
 b15ztpn00an1n08x5 PHY_277 ();
 b15ztpn00an1n08x5 PHY_278 ();
 b15ztpn00an1n08x5 PHY_279 ();
 b15ztpn00an1n08x5 PHY_280 ();
 b15ztpn00an1n08x5 PHY_281 ();
 b15ztpn00an1n08x5 PHY_282 ();
 b15ztpn00an1n08x5 PHY_283 ();
 b15ztpn00an1n08x5 PHY_284 ();
 b15ztpn00an1n08x5 PHY_285 ();
 b15ztpn00an1n08x5 PHY_286 ();
 b15ztpn00an1n08x5 PHY_287 ();
 b15ztpn00an1n08x5 PHY_288 ();
 b15ztpn00an1n08x5 PHY_289 ();
 b15ztpn00an1n08x5 PHY_290 ();
 b15ztpn00an1n08x5 PHY_291 ();
 b15ztpn00an1n08x5 PHY_292 ();
 b15ztpn00an1n08x5 PHY_293 ();
 b15ztpn00an1n08x5 PHY_294 ();
 b15ztpn00an1n08x5 PHY_295 ();
 b15ztpn00an1n08x5 PHY_296 ();
 b15ztpn00an1n08x5 PHY_297 ();
 b15ztpn00an1n08x5 PHY_298 ();
 b15ztpn00an1n08x5 PHY_299 ();
 b15ztpn00an1n08x5 PHY_300 ();
 b15ztpn00an1n08x5 PHY_301 ();
 b15ztpn00an1n08x5 PHY_302 ();
 b15ztpn00an1n08x5 PHY_303 ();
 b15ztpn00an1n08x5 PHY_304 ();
 b15ztpn00an1n08x5 PHY_305 ();
 b15ztpn00an1n08x5 PHY_306 ();
 b15ztpn00an1n08x5 PHY_307 ();
 b15ztpn00an1n08x5 PHY_308 ();
 b15ztpn00an1n08x5 PHY_309 ();
 b15ztpn00an1n08x5 PHY_310 ();
 b15ztpn00an1n08x5 PHY_311 ();
 b15ztpn00an1n08x5 PHY_312 ();
 b15ztpn00an1n08x5 PHY_313 ();
 b15ztpn00an1n08x5 PHY_314 ();
 b15ztpn00an1n08x5 PHY_315 ();
 b15ztpn00an1n08x5 PHY_316 ();
 b15ztpn00an1n08x5 PHY_317 ();
 b15ztpn00an1n08x5 PHY_318 ();
 b15ztpn00an1n08x5 PHY_319 ();
 b15ztpn00an1n08x5 PHY_320 ();
 b15ztpn00an1n08x5 PHY_321 ();
 b15ztpn00an1n08x5 PHY_322 ();
 b15ztpn00an1n08x5 PHY_323 ();
 b15ztpn00an1n08x5 PHY_324 ();
 b15ztpn00an1n08x5 PHY_325 ();
 b15ztpn00an1n08x5 PHY_326 ();
 b15ztpn00an1n08x5 PHY_327 ();
 b15ztpn00an1n08x5 PHY_328 ();
 b15ztpn00an1n08x5 PHY_329 ();
 b15ztpn00an1n08x5 PHY_330 ();
 b15ztpn00an1n08x5 PHY_331 ();
 b15ztpn00an1n08x5 PHY_332 ();
 b15ztpn00an1n08x5 PHY_333 ();
 b15ztpn00an1n08x5 PHY_334 ();
 b15ztpn00an1n08x5 PHY_335 ();
 b15ztpn00an1n08x5 PHY_336 ();
 b15ztpn00an1n08x5 PHY_337 ();
 b15ztpn00an1n08x5 PHY_338 ();
 b15ztpn00an1n08x5 PHY_339 ();
 b15ztpn00an1n08x5 PHY_340 ();
 b15ztpn00an1n08x5 PHY_341 ();
 b15ztpn00an1n08x5 PHY_342 ();
 b15ztpn00an1n08x5 PHY_343 ();
 b15ztpn00an1n08x5 PHY_344 ();
 b15ztpn00an1n08x5 PHY_345 ();
 b15ztpn00an1n08x5 PHY_346 ();
 b15ztpn00an1n08x5 PHY_347 ();
 b15ztpn00an1n08x5 PHY_348 ();
 b15ztpn00an1n08x5 PHY_349 ();
 b15ztpn00an1n08x5 PHY_350 ();
 b15ztpn00an1n08x5 PHY_351 ();
 b15ztpn00an1n08x5 PHY_352 ();
 b15ztpn00an1n08x5 PHY_353 ();
 b15ztpn00an1n08x5 PHY_354 ();
 b15ztpn00an1n08x5 PHY_355 ();
 b15ztpn00an1n08x5 PHY_356 ();
 b15ztpn00an1n08x5 PHY_357 ();
 b15ztpn00an1n08x5 PHY_358 ();
 b15ztpn00an1n08x5 PHY_359 ();
 b15ztpn00an1n08x5 PHY_360 ();
 b15ztpn00an1n08x5 PHY_361 ();
 b15ztpn00an1n08x5 PHY_362 ();
 b15ztpn00an1n08x5 PHY_363 ();
 b15ztpn00an1n08x5 PHY_364 ();
 b15ztpn00an1n08x5 PHY_365 ();
 b15ztpn00an1n08x5 PHY_366 ();
 b15ztpn00an1n08x5 PHY_367 ();
 b15ztpn00an1n08x5 PHY_368 ();
 b15ztpn00an1n08x5 PHY_369 ();
 b15ztpn00an1n08x5 PHY_370 ();
 b15ztpn00an1n08x5 PHY_371 ();
 b15ztpn00an1n08x5 PHY_372 ();
 b15ztpn00an1n08x5 PHY_373 ();
 b15ztpn00an1n08x5 PHY_374 ();
 b15ztpn00an1n08x5 PHY_375 ();
 b15ztpn00an1n08x5 PHY_376 ();
 b15ztpn00an1n08x5 PHY_377 ();
 b15ztpn00an1n08x5 PHY_378 ();
 b15ztpn00an1n08x5 PHY_379 ();
 b15ztpn00an1n08x5 PHY_380 ();
 b15ztpn00an1n08x5 PHY_381 ();
 b15ztpn00an1n08x5 PHY_382 ();
 b15ztpn00an1n08x5 PHY_383 ();
 b15ztpn00an1n08x5 PHY_384 ();
 b15ztpn00an1n08x5 PHY_385 ();
 b15ztpn00an1n08x5 PHY_386 ();
 b15ztpn00an1n08x5 PHY_387 ();
 b15ztpn00an1n08x5 PHY_388 ();
 b15ztpn00an1n08x5 PHY_389 ();
 b15ztpn00an1n08x5 TAP_390 ();
 b15ztpn00an1n08x5 TAP_391 ();
 b15ztpn00an1n08x5 TAP_392 ();
 b15ztpn00an1n08x5 TAP_393 ();
 b15ztpn00an1n08x5 TAP_394 ();
 b15ztpn00an1n08x5 TAP_395 ();
 b15ztpn00an1n08x5 TAP_396 ();
 b15ztpn00an1n08x5 TAP_397 ();
 b15ztpn00an1n08x5 TAP_398 ();
 b15ztpn00an1n08x5 TAP_399 ();
 b15ztpn00an1n08x5 TAP_400 ();
 b15ztpn00an1n08x5 TAP_401 ();
 b15ztpn00an1n08x5 TAP_402 ();
 b15ztpn00an1n08x5 TAP_403 ();
 b15ztpn00an1n08x5 TAP_404 ();
 b15ztpn00an1n08x5 TAP_405 ();
 b15ztpn00an1n08x5 TAP_406 ();
 b15ztpn00an1n08x5 TAP_407 ();
 b15ztpn00an1n08x5 TAP_408 ();
 b15ztpn00an1n08x5 TAP_409 ();
 b15ztpn00an1n08x5 TAP_410 ();
 b15ztpn00an1n08x5 TAP_411 ();
 b15ztpn00an1n08x5 TAP_412 ();
 b15ztpn00an1n08x5 TAP_413 ();
 b15ztpn00an1n08x5 TAP_414 ();
 b15ztpn00an1n08x5 TAP_415 ();
 b15ztpn00an1n08x5 TAP_416 ();
 b15ztpn00an1n08x5 TAP_417 ();
 b15ztpn00an1n08x5 TAP_418 ();
 b15ztpn00an1n08x5 TAP_419 ();
 b15ztpn00an1n08x5 TAP_420 ();
 b15ztpn00an1n08x5 TAP_421 ();
 b15ztpn00an1n08x5 TAP_422 ();
 b15ztpn00an1n08x5 TAP_423 ();
 b15ztpn00an1n08x5 TAP_424 ();
 b15ztpn00an1n08x5 TAP_425 ();
 b15ztpn00an1n08x5 TAP_426 ();
 b15ztpn00an1n08x5 TAP_427 ();
 b15ztpn00an1n08x5 TAP_428 ();
 b15ztpn00an1n08x5 TAP_429 ();
 b15ztpn00an1n08x5 TAP_430 ();
 b15ztpn00an1n08x5 TAP_431 ();
 b15ztpn00an1n08x5 TAP_432 ();
 b15ztpn00an1n08x5 TAP_433 ();
 b15ztpn00an1n08x5 TAP_434 ();
 b15ztpn00an1n08x5 TAP_435 ();
 b15ztpn00an1n08x5 TAP_436 ();
 b15ztpn00an1n08x5 TAP_437 ();
 b15ztpn00an1n08x5 TAP_438 ();
 b15ztpn00an1n08x5 TAP_439 ();
 b15ztpn00an1n08x5 TAP_440 ();
 b15ztpn00an1n08x5 TAP_441 ();
 b15ztpn00an1n08x5 TAP_442 ();
 b15ztpn00an1n08x5 TAP_443 ();
 b15ztpn00an1n08x5 TAP_444 ();
 b15ztpn00an1n08x5 TAP_445 ();
 b15ztpn00an1n08x5 TAP_446 ();
 b15ztpn00an1n08x5 TAP_447 ();
 b15ztpn00an1n08x5 TAP_448 ();
 b15ztpn00an1n08x5 TAP_449 ();
 b15ztpn00an1n08x5 TAP_450 ();
 b15ztpn00an1n08x5 TAP_451 ();
 b15ztpn00an1n08x5 TAP_452 ();
 b15ztpn00an1n08x5 TAP_453 ();
 b15ztpn00an1n08x5 TAP_454 ();
 b15ztpn00an1n08x5 TAP_455 ();
 b15ztpn00an1n08x5 TAP_456 ();
 b15ztpn00an1n08x5 TAP_457 ();
 b15ztpn00an1n08x5 TAP_458 ();
 b15ztpn00an1n08x5 TAP_459 ();
 b15ztpn00an1n08x5 TAP_460 ();
 b15ztpn00an1n08x5 TAP_461 ();
 b15ztpn00an1n08x5 TAP_462 ();
 b15ztpn00an1n08x5 TAP_463 ();
 b15ztpn00an1n08x5 TAP_464 ();
 b15ztpn00an1n08x5 TAP_465 ();
 b15ztpn00an1n08x5 TAP_466 ();
 b15ztpn00an1n08x5 TAP_467 ();
 b15ztpn00an1n08x5 TAP_468 ();
 b15ztpn00an1n08x5 TAP_469 ();
 b15ztpn00an1n08x5 TAP_470 ();
 b15ztpn00an1n08x5 TAP_471 ();
 b15ztpn00an1n08x5 TAP_472 ();
 b15ztpn00an1n08x5 TAP_473 ();
 b15ztpn00an1n08x5 TAP_474 ();
 b15ztpn00an1n08x5 TAP_475 ();
 b15ztpn00an1n08x5 TAP_476 ();
 b15ztpn00an1n08x5 TAP_477 ();
 b15ztpn00an1n08x5 TAP_478 ();
 b15ztpn00an1n08x5 TAP_479 ();
 b15ztpn00an1n08x5 TAP_480 ();
 b15ztpn00an1n08x5 TAP_481 ();
 b15ztpn00an1n08x5 TAP_482 ();
 b15ztpn00an1n08x5 TAP_483 ();
 b15ztpn00an1n08x5 TAP_484 ();
 b15ztpn00an1n08x5 TAP_485 ();
 b15ztpn00an1n08x5 TAP_486 ();
 b15ztpn00an1n08x5 TAP_487 ();
 b15ztpn00an1n08x5 TAP_488 ();
 b15ztpn00an1n08x5 TAP_489 ();
 b15ztpn00an1n08x5 TAP_490 ();
 b15ztpn00an1n08x5 TAP_491 ();
 b15ztpn00an1n08x5 TAP_492 ();
 b15ztpn00an1n08x5 TAP_493 ();
 b15ztpn00an1n08x5 TAP_494 ();
 b15ztpn00an1n08x5 TAP_495 ();
 b15ztpn00an1n08x5 TAP_496 ();
 b15ztpn00an1n08x5 TAP_497 ();
 b15ztpn00an1n08x5 TAP_498 ();
 b15ztpn00an1n08x5 TAP_499 ();
 b15ztpn00an1n08x5 TAP_500 ();
 b15ztpn00an1n08x5 TAP_501 ();
 b15ztpn00an1n08x5 TAP_502 ();
 b15ztpn00an1n08x5 TAP_503 ();
 b15ztpn00an1n08x5 TAP_504 ();
 b15ztpn00an1n08x5 TAP_505 ();
 b15ztpn00an1n08x5 TAP_506 ();
 b15ztpn00an1n08x5 TAP_507 ();
 b15ztpn00an1n08x5 TAP_508 ();
 b15ztpn00an1n08x5 TAP_509 ();
 b15ztpn00an1n08x5 TAP_510 ();
 b15ztpn00an1n08x5 TAP_511 ();
 b15ztpn00an1n08x5 TAP_512 ();
 b15ztpn00an1n08x5 TAP_513 ();
 b15ztpn00an1n08x5 TAP_514 ();
 b15ztpn00an1n08x5 TAP_515 ();
 b15ztpn00an1n08x5 TAP_516 ();
 b15ztpn00an1n08x5 TAP_517 ();
 b15ztpn00an1n08x5 TAP_518 ();
 b15ztpn00an1n08x5 TAP_519 ();
 b15ztpn00an1n08x5 TAP_520 ();
 b15ztpn00an1n08x5 TAP_521 ();
 b15ztpn00an1n08x5 TAP_522 ();
 b15ztpn00an1n08x5 TAP_523 ();
 b15ztpn00an1n08x5 TAP_524 ();
 b15ztpn00an1n08x5 TAP_525 ();
 b15ztpn00an1n08x5 TAP_526 ();
 b15ztpn00an1n08x5 TAP_527 ();
 b15ztpn00an1n08x5 TAP_528 ();
 b15ztpn00an1n08x5 TAP_529 ();
 b15ztpn00an1n08x5 TAP_530 ();
 b15ztpn00an1n08x5 TAP_531 ();
 b15ztpn00an1n08x5 TAP_532 ();
 b15ztpn00an1n08x5 TAP_533 ();
 b15ztpn00an1n08x5 TAP_534 ();
 b15ztpn00an1n08x5 TAP_535 ();
 b15ztpn00an1n08x5 TAP_536 ();
 b15ztpn00an1n08x5 TAP_537 ();
 b15ztpn00an1n08x5 TAP_538 ();
 b15ztpn00an1n08x5 TAP_539 ();
 b15ztpn00an1n08x5 TAP_540 ();
 b15ztpn00an1n08x5 TAP_541 ();
 b15ztpn00an1n08x5 TAP_542 ();
 b15ztpn00an1n08x5 TAP_543 ();
 b15ztpn00an1n08x5 TAP_544 ();
 b15ztpn00an1n08x5 TAP_545 ();
 b15ztpn00an1n08x5 TAP_546 ();
 b15ztpn00an1n08x5 TAP_547 ();
 b15ztpn00an1n08x5 TAP_548 ();
 b15ztpn00an1n08x5 TAP_549 ();
 b15ztpn00an1n08x5 TAP_550 ();
 b15ztpn00an1n08x5 TAP_551 ();
 b15ztpn00an1n08x5 TAP_552 ();
 b15ztpn00an1n08x5 TAP_553 ();
 b15ztpn00an1n08x5 TAP_554 ();
 b15ztpn00an1n08x5 TAP_555 ();
 b15ztpn00an1n08x5 TAP_556 ();
 b15ztpn00an1n08x5 TAP_557 ();
 b15ztpn00an1n08x5 TAP_558 ();
 b15ztpn00an1n08x5 TAP_559 ();
 b15ztpn00an1n08x5 TAP_560 ();
 b15ztpn00an1n08x5 TAP_561 ();
 b15ztpn00an1n08x5 TAP_562 ();
 b15ztpn00an1n08x5 TAP_563 ();
 b15ztpn00an1n08x5 TAP_564 ();
 b15ztpn00an1n08x5 TAP_565 ();
 b15ztpn00an1n08x5 TAP_566 ();
 b15ztpn00an1n08x5 TAP_567 ();
 b15ztpn00an1n08x5 TAP_568 ();
 b15ztpn00an1n08x5 TAP_569 ();
 b15ztpn00an1n08x5 TAP_570 ();
 b15ztpn00an1n08x5 TAP_571 ();
 b15ztpn00an1n08x5 TAP_572 ();
 b15ztpn00an1n08x5 TAP_573 ();
 b15ztpn00an1n08x5 TAP_574 ();
 b15ztpn00an1n08x5 TAP_575 ();
 b15ztpn00an1n08x5 TAP_576 ();
 b15ztpn00an1n08x5 TAP_577 ();
 b15ztpn00an1n08x5 TAP_578 ();
 b15ztpn00an1n08x5 TAP_579 ();
 b15ztpn00an1n08x5 TAP_580 ();
 b15ztpn00an1n08x5 TAP_581 ();
 b15ztpn00an1n08x5 TAP_582 ();
 b15ztpn00an1n08x5 TAP_583 ();
 b15ztpn00an1n08x5 TAP_584 ();
 b15ztpn00an1n08x5 TAP_585 ();
 b15ztpn00an1n08x5 TAP_586 ();
 b15ztpn00an1n08x5 TAP_587 ();
 b15ztpn00an1n08x5 TAP_588 ();
 b15ztpn00an1n08x5 TAP_589 ();
 b15ztpn00an1n08x5 TAP_590 ();
 b15ztpn00an1n08x5 TAP_591 ();
 b15ztpn00an1n08x5 TAP_592 ();
 b15ztpn00an1n08x5 TAP_593 ();
 b15ztpn00an1n08x5 TAP_594 ();
 b15ztpn00an1n08x5 TAP_595 ();
 b15ztpn00an1n08x5 TAP_596 ();
 b15ztpn00an1n08x5 TAP_597 ();
 b15ztpn00an1n08x5 TAP_598 ();
 b15ztpn00an1n08x5 TAP_599 ();
 b15ztpn00an1n08x5 TAP_600 ();
 b15ztpn00an1n08x5 TAP_601 ();
 b15ztpn00an1n08x5 TAP_602 ();
 b15ztpn00an1n08x5 TAP_603 ();
 b15ztpn00an1n08x5 TAP_604 ();
 b15ztpn00an1n08x5 TAP_605 ();
 b15ztpn00an1n08x5 TAP_606 ();
 b15ztpn00an1n08x5 TAP_607 ();
 b15ztpn00an1n08x5 TAP_608 ();
 b15ztpn00an1n08x5 TAP_609 ();
 b15ztpn00an1n08x5 TAP_610 ();
 b15ztpn00an1n08x5 TAP_611 ();
 b15ztpn00an1n08x5 TAP_612 ();
 b15ztpn00an1n08x5 TAP_613 ();
 b15ztpn00an1n08x5 TAP_614 ();
 b15ztpn00an1n08x5 TAP_615 ();
 b15ztpn00an1n08x5 TAP_616 ();
 b15ztpn00an1n08x5 TAP_617 ();
 b15ztpn00an1n08x5 TAP_618 ();
 b15ztpn00an1n08x5 TAP_619 ();
 b15ztpn00an1n08x5 TAP_620 ();
 b15ztpn00an1n08x5 TAP_621 ();
 b15ztpn00an1n08x5 TAP_622 ();
 b15ztpn00an1n08x5 TAP_623 ();
 b15ztpn00an1n08x5 TAP_624 ();
 b15ztpn00an1n08x5 TAP_625 ();
 b15ztpn00an1n08x5 TAP_626 ();
 b15ztpn00an1n08x5 TAP_627 ();
 b15ztpn00an1n08x5 TAP_628 ();
 b15ztpn00an1n08x5 TAP_629 ();
 b15ztpn00an1n08x5 TAP_630 ();
 b15ztpn00an1n08x5 TAP_631 ();
 b15ztpn00an1n08x5 TAP_632 ();
 b15ztpn00an1n08x5 TAP_633 ();
 b15ztpn00an1n08x5 TAP_634 ();
 b15ztpn00an1n08x5 TAP_635 ();
 b15ztpn00an1n08x5 TAP_636 ();
 b15ztpn00an1n08x5 TAP_637 ();
 b15ztpn00an1n08x5 TAP_638 ();
 b15ztpn00an1n08x5 TAP_639 ();
 b15ztpn00an1n08x5 TAP_640 ();
 b15ztpn00an1n08x5 TAP_641 ();
 b15ztpn00an1n08x5 TAP_642 ();
 b15ztpn00an1n08x5 TAP_643 ();
 b15ztpn00an1n08x5 TAP_644 ();
 b15ztpn00an1n08x5 TAP_645 ();
 b15ztpn00an1n08x5 TAP_646 ();
 b15ztpn00an1n08x5 TAP_647 ();
 b15ztpn00an1n08x5 TAP_648 ();
 b15ztpn00an1n08x5 TAP_649 ();
 b15ztpn00an1n08x5 TAP_650 ();
 b15ztpn00an1n08x5 TAP_651 ();
 b15ztpn00an1n08x5 TAP_652 ();
 b15ztpn00an1n08x5 TAP_653 ();
 b15ztpn00an1n08x5 TAP_654 ();
 b15ztpn00an1n08x5 TAP_655 ();
 b15ztpn00an1n08x5 TAP_656 ();
 b15ztpn00an1n08x5 TAP_657 ();
 b15ztpn00an1n08x5 TAP_658 ();
 b15ztpn00an1n08x5 TAP_659 ();
 b15ztpn00an1n08x5 TAP_660 ();
 b15ztpn00an1n08x5 TAP_661 ();
 b15ztpn00an1n08x5 TAP_662 ();
 b15ztpn00an1n08x5 TAP_663 ();
 b15ztpn00an1n08x5 TAP_664 ();
 b15ztpn00an1n08x5 TAP_665 ();
 b15ztpn00an1n08x5 TAP_666 ();
 b15ztpn00an1n08x5 TAP_667 ();
 b15ztpn00an1n08x5 TAP_668 ();
 b15ztpn00an1n08x5 TAP_669 ();
 b15ztpn00an1n08x5 TAP_670 ();
 b15ztpn00an1n08x5 TAP_671 ();
 b15ztpn00an1n08x5 TAP_672 ();
 b15ztpn00an1n08x5 TAP_673 ();
 b15ztpn00an1n08x5 TAP_674 ();
 b15ztpn00an1n08x5 TAP_675 ();
 b15ztpn00an1n08x5 TAP_676 ();
 b15ztpn00an1n08x5 TAP_677 ();
 b15ztpn00an1n08x5 TAP_678 ();
 b15ztpn00an1n08x5 TAP_679 ();
 b15ztpn00an1n08x5 TAP_680 ();
 b15ztpn00an1n08x5 TAP_681 ();
 b15ztpn00an1n08x5 TAP_682 ();
 b15ztpn00an1n08x5 TAP_683 ();
 b15ztpn00an1n08x5 TAP_684 ();
 b15ztpn00an1n08x5 TAP_685 ();
 b15ztpn00an1n08x5 TAP_686 ();
 b15ztpn00an1n08x5 TAP_687 ();
 b15ztpn00an1n08x5 TAP_688 ();
 b15ztpn00an1n08x5 TAP_689 ();
 b15ztpn00an1n08x5 TAP_690 ();
 b15ztpn00an1n08x5 TAP_691 ();
 b15ztpn00an1n08x5 TAP_692 ();
 b15ztpn00an1n08x5 TAP_693 ();
 b15ztpn00an1n08x5 TAP_694 ();
 b15ztpn00an1n08x5 TAP_695 ();
 b15ztpn00an1n08x5 TAP_696 ();
 b15ztpn00an1n08x5 TAP_697 ();
 b15ztpn00an1n08x5 TAP_698 ();
 b15ztpn00an1n08x5 TAP_699 ();
 b15ztpn00an1n08x5 TAP_700 ();
 b15ztpn00an1n08x5 TAP_701 ();
 b15ztpn00an1n08x5 TAP_702 ();
 b15ztpn00an1n08x5 TAP_703 ();
 b15ztpn00an1n08x5 TAP_704 ();
 b15ztpn00an1n08x5 TAP_705 ();
 b15ztpn00an1n08x5 TAP_706 ();
 b15ztpn00an1n08x5 TAP_707 ();
 b15ztpn00an1n08x5 TAP_708 ();
 b15ztpn00an1n08x5 TAP_709 ();
 b15ztpn00an1n08x5 TAP_710 ();
 b15ztpn00an1n08x5 TAP_711 ();
 b15ztpn00an1n08x5 TAP_712 ();
 b15ztpn00an1n08x5 TAP_713 ();
 b15ztpn00an1n08x5 TAP_714 ();
 b15ztpn00an1n08x5 TAP_715 ();
 b15ztpn00an1n08x5 TAP_716 ();
 b15ztpn00an1n08x5 TAP_717 ();
 b15ztpn00an1n08x5 TAP_718 ();
 b15ztpn00an1n08x5 TAP_719 ();
 b15ztpn00an1n08x5 TAP_720 ();
 b15ztpn00an1n08x5 TAP_721 ();
 b15ztpn00an1n08x5 TAP_722 ();
 b15ztpn00an1n08x5 TAP_723 ();
 b15ztpn00an1n08x5 TAP_724 ();
 b15ztpn00an1n08x5 TAP_725 ();
 b15ztpn00an1n08x5 TAP_726 ();
 b15ztpn00an1n08x5 TAP_727 ();
 b15ztpn00an1n08x5 TAP_728 ();
 b15ztpn00an1n08x5 TAP_729 ();
 b15ztpn00an1n08x5 TAP_730 ();
 b15ztpn00an1n08x5 TAP_731 ();
 b15ztpn00an1n08x5 TAP_732 ();
 b15ztpn00an1n08x5 TAP_733 ();
 b15ztpn00an1n08x5 TAP_734 ();
 b15ztpn00an1n08x5 TAP_735 ();
 b15ztpn00an1n08x5 TAP_736 ();
 b15ztpn00an1n08x5 TAP_737 ();
 b15ztpn00an1n08x5 TAP_738 ();
 b15ztpn00an1n08x5 TAP_739 ();
 b15ztpn00an1n08x5 TAP_740 ();
 b15ztpn00an1n08x5 TAP_741 ();
 b15ztpn00an1n08x5 TAP_742 ();
 b15ztpn00an1n08x5 TAP_743 ();
 b15ztpn00an1n08x5 TAP_744 ();
 b15ztpn00an1n08x5 TAP_745 ();
 b15ztpn00an1n08x5 TAP_746 ();
 b15ztpn00an1n08x5 TAP_747 ();
 b15ztpn00an1n08x5 TAP_748 ();
 b15ztpn00an1n08x5 TAP_749 ();
 b15ztpn00an1n08x5 TAP_750 ();
 b15ztpn00an1n08x5 TAP_751 ();
 b15ztpn00an1n08x5 TAP_752 ();
 b15ztpn00an1n08x5 TAP_753 ();
 b15ztpn00an1n08x5 TAP_754 ();
 b15ztpn00an1n08x5 TAP_755 ();
 b15ztpn00an1n08x5 TAP_756 ();
 b15ztpn00an1n08x5 TAP_757 ();
 b15ztpn00an1n08x5 TAP_758 ();
 b15ztpn00an1n08x5 TAP_759 ();
 b15ztpn00an1n08x5 TAP_760 ();
 b15ztpn00an1n08x5 TAP_761 ();
 b15ztpn00an1n08x5 TAP_762 ();
 b15ztpn00an1n08x5 TAP_763 ();
 b15ztpn00an1n08x5 TAP_764 ();
 b15ztpn00an1n08x5 TAP_765 ();
 b15ztpn00an1n08x5 TAP_766 ();
 b15ztpn00an1n08x5 TAP_767 ();
 b15ztpn00an1n08x5 TAP_768 ();
 b15ztpn00an1n08x5 TAP_769 ();
 b15ztpn00an1n08x5 TAP_770 ();
 b15ztpn00an1n08x5 TAP_771 ();
 b15ztpn00an1n08x5 TAP_772 ();
 b15ztpn00an1n08x5 TAP_773 ();
 b15ztpn00an1n08x5 TAP_774 ();
 b15ztpn00an1n08x5 TAP_775 ();
 b15ztpn00an1n08x5 TAP_776 ();
 b15ztpn00an1n08x5 TAP_777 ();
 b15ztpn00an1n08x5 TAP_778 ();
 b15ztpn00an1n08x5 TAP_779 ();
 b15ztpn00an1n08x5 TAP_780 ();
 b15bfn001as1n08x5 input1 (.a(net2200),
    .o(net1));
 b15bfn001ah1n12x5 input2 (.a(tl_peri_device_i[0]),
    .o(net2));
 b15bfn001as1n16x5 input3 (.a(tl_peri_device_i[100]),
    .o(net3));
 b15bfn001ah1n12x5 input4 (.a(tl_peri_device_i[101]),
    .o(net4));
 b15bfn001ah1n08x5 input5 (.a(tl_peri_device_i[105]),
    .o(net5));
 b15bfn000as1n06x5 input6 (.a(tl_peri_device_i[106]),
    .o(net6));
 b15bfn000as1n04x5 input7 (.a(tl_peri_device_i[107]),
    .o(net7));
 b15bfn001as1n08x5 input8 (.a(tl_peri_device_i[108]),
    .o(net8));
 b15bfn000ah1n03x5 input9 (.a(tl_peri_device_i[15]),
    .o(net9));
 b15bfn001ah1n08x5 input10 (.a(tl_peri_device_i[16]),
    .o(net10));
 b15bfn001as1n06x5 input11 (.a(tl_peri_device_i[17]),
    .o(net11));
 b15bfn001aq1n06x5 input12 (.a(tl_peri_device_i[18]),
    .o(net12));
 b15bfn001as1n32x5 input13 (.a(tl_peri_device_i[24]),
    .o(net13));
 b15bfn001as1n16x5 input14 (.a(tl_peri_device_i[25]),
    .o(net14));
 b15bfn001as1n12x5 input15 (.a(tl_peri_device_i[26]),
    .o(net15));
 b15bfn001ah1n16x5 input16 (.a(tl_peri_device_i[27]),
    .o(net16));
 b15bfn001as1n12x5 input17 (.a(tl_peri_device_i[28]),
    .o(net17));
 b15bfn001as1n12x5 input18 (.a(tl_peri_device_i[29]),
    .o(net18));
 b15bfn001ah1n24x5 input19 (.a(tl_peri_device_i[30]),
    .o(net19));
 b15bfn001ah1n32x5 input20 (.a(tl_peri_device_i[31]),
    .o(net20));
 b15bfn001as1n16x5 input21 (.a(tl_peri_device_i[32]),
    .o(net21));
 b15bfn001as1n16x5 input22 (.a(tl_peri_device_i[33]),
    .o(net22));
 b15bfn001as1n24x5 input23 (.a(tl_peri_device_i[34]),
    .o(net23));
 b15bfn001ah1n24x5 input24 (.a(tl_peri_device_i[35]),
    .o(net24));
 b15bfn001as1n24x5 input25 (.a(tl_peri_device_i[36]),
    .o(net25));
 b15bfn001ah1n24x5 input26 (.a(tl_peri_device_i[37]),
    .o(net26));
 b15bfn001as1n24x5 input27 (.a(tl_peri_device_i[38]),
    .o(net27));
 b15bfn001as1n24x5 input28 (.a(tl_peri_device_i[39]),
    .o(net28));
 b15bfn001as1n16x5 input29 (.a(tl_peri_device_i[40]),
    .o(net29));
 b15bfn001as1n16x5 input30 (.a(tl_peri_device_i[41]),
    .o(net30));
 b15bfn001as1n16x5 input31 (.a(tl_peri_device_i[42]),
    .o(net31));
 b15bfn001ah1n16x5 input32 (.a(tl_peri_device_i[43]),
    .o(net32));
 b15bfn001as1n16x5 input33 (.a(tl_peri_device_i[44]),
    .o(net33));
 b15bfn001as1n24x5 input34 (.a(tl_peri_device_i[45]),
    .o(net34));
 b15bfn001ah1n24x5 input35 (.a(tl_peri_device_i[46]),
    .o(net35));
 b15bfn000as1n24x5 input36 (.a(tl_peri_device_i[47]),
    .o(net36));
 b15bfn001as1n06x5 input37 (.a(tl_peri_device_i[48]),
    .o(net37));
 b15bfn001as1n16x5 input38 (.a(tl_peri_device_i[49]),
    .o(net38));
 b15bfn001ah1n32x5 input39 (.a(tl_peri_device_i[50]),
    .o(net39));
 b15bfn001ah1n32x5 input40 (.a(tl_peri_device_i[51]),
    .o(net40));
 b15bfn001ah1n24x5 input41 (.a(tl_peri_device_i[52]),
    .o(net41));
 b15bfn001ah1n24x5 input42 (.a(tl_peri_device_i[53]),
    .o(net42));
 b15bfn001as1n32x5 input43 (.a(tl_peri_device_i[54]),
    .o(net43));
 b15bfn001as1n32x5 input44 (.a(tl_peri_device_i[55]),
    .o(net44));
 b15bfn001ah1n06x5 input45 (.a(tl_peri_device_i[56]),
    .o(net45));
 b15bfn001aq1n06x5 input46 (.a(tl_peri_device_i[57]),
    .o(net46));
 b15bfn001al1n08x5 input47 (.a(tl_peri_device_i[58]),
    .o(net47));
 b15bfn001aq1n06x5 input48 (.a(tl_peri_device_i[59]),
    .o(net48));
 b15bfn000as1n06x5 input49 (.a(tl_peri_device_i[60]),
    .o(net49));
 b15qgbbf1an1n05x5 input50 (.a(tl_peri_device_i[61]),
    .o(net50));
 b15bfn001ah1n48x5 input51 (.a(tl_peri_device_i[62]),
    .o(net51));
 b15bfn001ah1n48x5 input52 (.a(tl_peri_device_i[63]),
    .o(net52));
 b15bfn001as1n32x5 input53 (.a(tl_peri_device_i[64]),
    .o(net53));
 b15bfn001as1n24x5 input54 (.a(tl_peri_device_i[65]),
    .o(net54));
 b15bfn000ah1n04x5 input55 (.a(tl_peri_device_i[76]),
    .o(net55));
 b15bfn001aq1n06x5 input56 (.a(tl_peri_device_i[77]),
    .o(net56));
 b15bfn000ah1n02x5 input57 (.a(tl_peri_device_i[78]),
    .o(net57));
 b15bfn000ar1n02x5 input58 (.a(tl_peri_device_i[79]),
    .o(net58));
 b15bfn000al1n02x5 input59 (.a(tl_peri_device_i[80]),
    .o(net59));
 b15bfn000ar1n02x5 input60 (.a(tl_peri_device_i[81]),
    .o(net60));
 b15bfn000ar1n02x5 input61 (.a(tl_peri_device_i[82]),
    .o(net61));
 b15bfn000an1n02x5 input62 (.a(tl_peri_device_i[83]),
    .o(net62));
 b15bfn000ar1n02x5 input63 (.a(tl_peri_device_i[84]),
    .o(net63));
 b15bfn000ar1n02x5 input64 (.a(tl_peri_device_i[85]),
    .o(net64));
 b15bfn000ar1n02x5 input65 (.a(tl_peri_device_i[86]),
    .o(net65));
 b15bfn000ar1n02x5 input66 (.a(tl_peri_device_i[87]),
    .o(net66));
 b15bfn000al1n02x5 input67 (.a(tl_peri_device_i[88]),
    .o(net67));
 b15bfn000ar1n02x5 input68 (.a(tl_peri_device_i[89]),
    .o(net68));
 b15bfn000al1n02x5 input69 (.a(tl_peri_device_i[90]),
    .o(net69));
 b15bfn000al1n02x5 input70 (.a(tl_peri_device_i[91]),
    .o(net70));
 b15bfn001ah1n08x5 input71 (.a(tl_peri_device_i[92]),
    .o(net71));
 b15bfn001ah1n08x5 input72 (.a(tl_peri_device_i[93]),
    .o(net72));
 b15bfn001ah1n08x5 input73 (.a(tl_peri_device_i[94]),
    .o(net73));
 b15bfn001ah1n08x5 input74 (.a(tl_peri_device_i[95]),
    .o(net74));
 b15bfn001ah1n08x5 input75 (.a(tl_peri_device_i[96]),
    .o(net75));
 b15bfn001ah1n08x5 input76 (.a(tl_peri_device_i[97]),
    .o(net76));
 b15bfn001as1n06x5 input77 (.a(tl_peri_device_i[98]),
    .o(net77));
 b15bfn001as1n06x5 input78 (.a(tl_peri_device_i[99]),
    .o(net78));
 b15bfn000ah1n03x5 output79 (.a(net79),
    .o(gpio_o[0]));
 b15bfn000ah1n03x5 output80 (.a(net389),
    .o(gpio_o[10]));
 b15bfn000ah1n03x5 output81 (.a(net388),
    .o(gpio_o[11]));
 b15bfn000ah1n03x5 output82 (.a(net386),
    .o(gpio_o[12]));
 b15bfn000ah1n03x5 output83 (.a(net385),
    .o(gpio_o[13]));
 b15bfn000ah1n03x5 output84 (.a(net84),
    .o(gpio_o[14]));
 b15bfn000ah1n03x5 output85 (.a(net85),
    .o(gpio_o[15]));
 b15bfn000ah1n03x5 output86 (.a(net86),
    .o(gpio_o[16]));
 b15bfn000ah1n03x5 output87 (.a(net87),
    .o(gpio_o[17]));
 b15bfn000ah1n03x5 output88 (.a(net88),
    .o(gpio_o[18]));
 b15bfn000ah1n03x5 output89 (.a(net2126),
    .o(gpio_o[19]));
 b15bfn000ah1n03x5 output90 (.a(net90),
    .o(gpio_o[1]));
 b15bfn000ah1n03x5 output91 (.a(net2192),
    .o(gpio_o[20]));
 b15bfn000ah1n03x5 output92 (.a(net1985),
    .o(gpio_o[21]));
 b15bfn000ah1n03x5 output93 (.a(net2087),
    .o(gpio_o[22]));
 b15bfn000ah1n03x5 output94 (.a(net2095),
    .o(gpio_o[23]));
 b15bfn000ah1n03x5 output95 (.a(net2106),
    .o(gpio_o[24]));
 b15bfn000ah1n03x5 output96 (.a(net96),
    .o(gpio_o[25]));
 b15bfn000ah1n03x5 output97 (.a(net2178),
    .o(gpio_o[26]));
 b15bfn000ah1n03x5 output98 (.a(net98),
    .o(gpio_o[27]));
 b15bfn000ah1n03x5 output99 (.a(net99),
    .o(gpio_o[28]));
 b15bfn000ah1n03x5 output100 (.a(net2020),
    .o(gpio_o[29]));
 b15bfn000ah1n03x5 output101 (.a(net2103),
    .o(gpio_o[2]));
 b15bfn000ah1n03x5 output102 (.a(net2052),
    .o(gpio_o[30]));
 b15bfn000ah1n03x5 output103 (.a(net363),
    .o(gpio_o[31]));
 b15bfn000ah1n03x5 output104 (.a(net2158),
    .o(gpio_o[3]));
 b15bfn000ah1n03x5 output105 (.a(net1964),
    .o(gpio_o[4]));
 b15bfn000ah1n03x5 output106 (.a(net2097),
    .o(gpio_o[5]));
 b15bfn000ah1n03x5 output107 (.a(net2053),
    .o(gpio_o[6]));
 b15bfn000ah1n03x5 output108 (.a(net108),
    .o(gpio_o[7]));
 b15bfn000ah1n03x5 output109 (.a(net361),
    .o(gpio_o[8]));
 b15bfn000ah1n03x5 output110 (.a(net358),
    .o(gpio_o[9]));
 b15bfn000ah1n03x5 output111 (.a(net1868),
    .o(tl_peri_device_o[0]));
 b15bfn000ah1n03x5 output112 (.a(net1808),
    .o(net1809));
 b15bfn000ah1n03x5 output113 (.a(net1850),
    .o(net1851));
 b15bfn000ah1n03x5 output114 (.a(net1892),
    .o(tl_peri_device_o[12]));
 b15bfn000ah1n03x5 output115 (.a(net1782),
    .o(net1783));
 b15bfn000ah1n03x5 output116 (.a(net116),
    .o(tl_peri_device_o[14]));
 b15bfn000ah1n03x5 output117 (.a(net1862),
    .o(tl_peri_device_o[15]));
 b15bfn000ah1n03x5 output118 (.a(net118),
    .o(tl_peri_device_o[16]));
 b15bfn000ah1n03x5 output119 (.a(net119),
    .o(tl_peri_device_o[17]));
 b15bfn000ah1n03x5 output120 (.a(net120),
    .o(tl_peri_device_o[18]));
 b15bfn000ah1n03x5 output121 (.a(net121),
    .o(tl_peri_device_o[19]));
 b15bfn000ah1n03x5 output122 (.a(net1917),
    .o(tl_peri_device_o[1]));
 b15bfn000ah1n03x5 output123 (.a(net123),
    .o(tl_peri_device_o[20]));
 b15bfn000ah1n03x5 output124 (.a(net124),
    .o(tl_peri_device_o[21]));
 b15bfn000ah1n03x5 output125 (.a(net125),
    .o(tl_peri_device_o[22]));
 b15bfn000ah1n03x5 output126 (.a(net126),
    .o(tl_peri_device_o[23]));
 b15bfn000ah1n03x5 output127 (.a(net127),
    .o(tl_peri_device_o[24]));
 b15bfn000ah1n03x5 output128 (.a(net128),
    .o(tl_peri_device_o[25]));
 b15bfn000ah1n03x5 output129 (.a(net129),
    .o(tl_peri_device_o[26]));
 b15bfn000ah1n03x5 output130 (.a(net1804),
    .o(tl_peri_device_o[27]));
 b15bfn000ah1n03x5 output131 (.a(net131),
    .o(tl_peri_device_o[28]));
 b15bfn000ah1n03x5 output132 (.a(net132),
    .o(tl_peri_device_o[29]));
 b15bfn000ah1n03x5 output133 (.a(net1879),
    .o(tl_peri_device_o[2]));
 b15bfn000ah1n03x5 output134 (.a(net134),
    .o(tl_peri_device_o[30]));
 b15bfn000ah1n03x5 output135 (.a(net1794),
    .o(tl_peri_device_o[31]));
 b15bfn000ah1n03x5 output136 (.a(net136),
    .o(tl_peri_device_o[32]));
 b15bfn000ah1n03x5 output137 (.a(net1821),
    .o(tl_peri_device_o[33]));
 b15bfn000ah1n03x5 output138 (.a(net138),
    .o(tl_peri_device_o[34]));
 b15bfn000ah1n03x5 output139 (.a(net139),
    .o(tl_peri_device_o[35]));
 b15bfn000ah1n03x5 output140 (.a(net140),
    .o(tl_peri_device_o[36]));
 b15bfn000ah1n03x5 output141 (.a(net1825),
    .o(tl_peri_device_o[37]));
 b15bfn000ah1n03x5 output142 (.a(net1856),
    .o(tl_peri_device_o[38]));
 b15bfn000ah1n03x5 output143 (.a(net143),
    .o(tl_peri_device_o[39]));
 b15bfn000ah1n03x5 output144 (.a(net1872),
    .o(tl_peri_device_o[3]));
 b15bfn000ah1n03x5 output145 (.a(net145),
    .o(tl_peri_device_o[40]));
 b15bfn000ah1n03x5 output146 (.a(net1779),
    .o(tl_peri_device_o[41]));
 b15bfn000ah1n03x5 output147 (.a(net147),
    .o(tl_peri_device_o[42]));
 b15bfn000ah1n03x5 output148 (.a(net148),
    .o(tl_peri_device_o[43]));
 b15bfn000ah1n03x5 output149 (.a(net149),
    .o(tl_peri_device_o[44]));
 b15bfn000ah1n03x5 output150 (.a(net150),
    .o(tl_peri_device_o[45]));
 b15bfn000ah1n03x5 output151 (.a(net151),
    .o(tl_peri_device_o[46]));
 b15bfn000ah1n03x5 output152 (.a(net152),
    .o(tl_peri_device_o[47]));
 b15bfn000ah1n03x5 output153 (.a(net1845),
    .o(net1846));
 b15bfn000ah1n03x5 output154 (.a(net1927),
    .o(tl_peri_device_o[4]));
 b15bfn000ah1n03x5 output155 (.a(net1833),
    .o(net1834));
 b15bfn000ah1n03x5 output156 (.a(net1817),
    .o(net1818));
 b15bfn000ah1n03x5 output157 (.a(net1836),
    .o(net1837));
 b15bfn000ah1n03x5 output158 (.a(net1800),
    .o(net1801));
 b15bfn000ah1n03x5 output159 (.a(net1814),
    .o(net1815));
 b15bfn000ah1n03x5 output160 (.a(net1763),
    .o(net1764));
 b15bfn000ah1n03x5 output161 (.a(net1811),
    .o(net1812));
 b15bfn000ah1n03x5 output162 (.a(net1797),
    .o(net1798));
 b15bfn000ah1n03x5 output163 (.a(net1787),
    .o(tl_peri_device_o[58]));
 b15bfn000ah1n03x5 output164 (.a(net1876),
    .o(tl_peri_device_o[5]));
 b15bfn000ah1n03x5 output165 (.a(net1768),
    .o(net1769));
 b15bfn000ah1n03x5 output166 (.a(net1790),
    .o(net1791));
 b15bfn000ah1n03x5 output167 (.a(net1896),
    .o(tl_peri_device_o[64]));
 b15bfn000ah1n03x5 output168 (.a(net1760),
    .o(net1761));
 b15bfn000ah1n03x5 output169 (.a(net1924),
    .o(tl_peri_device_o[6]));
 b15bfn000ah1n03x5 output170 (.a(net170),
    .o(tl_peri_device_o[7]));
 b15bfn000ah1n03x5 output171 (.a(net1920),
    .o(tl_peri_device_o[8]));
 b15bfn000ah1n03x5 output172 (.a(net1774),
    .o(net1775));
 b15bfn001as1n16x5 fanout173 (.a(n3944),
    .o(net173));
 b15bfn001ah1n16x5 fanout174 (.a(n3944),
    .o(net174));
 b15bfn001as1n24x5 wire175 (.a(u_gpio_u_reg_u_reg_if_N43),
    .o(net175));
 b15bfn000as1n24x5 wire176 (.a(u_gpio_u_reg_u_reg_if_N42),
    .o(net176));
 b15bfn001as1n16x5 wire177 (.a(u_gpio_u_reg_u_reg_if_N33),
    .o(net177));
 b15bfn001ah1n24x5 wire178 (.a(u_gpio_u_reg_u_reg_if_N44),
    .o(net178));
 b15bfn001as1n32x5 wire179 (.a(u_gpio_u_reg_reg_we_check_14_),
    .o(net179));
 b15bfn001ah1n64x5 fanout180 (.a(net181),
    .o(net180));
 b15bfn001as1n80x5 fanout181 (.a(n3343),
    .o(net181));
 b15bfn001as1n32x5 fanout182 (.a(net183),
    .o(net182));
 b15bfn001ah1n48x5 fanout183 (.a(n3296),
    .o(net183));
 b15bfn001ah1n48x5 fanout184 (.a(n3330),
    .o(net184));
 b15bfn001ah1n24x5 wire185 (.a(u_gpio_u_reg_u_reg_if_N34),
    .o(net185));
 b15bfn001as1n16x5 wire186 (.a(u_gpio_u_reg_u_reg_if_N38),
    .o(net186));
 b15bfn001as1n16x5 wire187 (.a(u_gpio_u_reg_u_reg_if_N35),
    .o(net187));
 b15bfn001as1n16x5 wire188 (.a(u_gpio_u_reg_u_reg_if_N39),
    .o(net188));
 b15bfn001as1n16x5 wire189 (.a(u_gpio_u_reg_u_reg_if_N20),
    .o(net189));
 b15bfn001as1n16x5 wire190 (.a(u_gpio_u_reg_u_reg_if_N19),
    .o(net190));
 b15bfn001as1n16x5 wire191 (.a(u_gpio_u_reg_u_reg_if_N18),
    .o(net191));
 b15bfn001as1n16x5 wire192 (.a(u_gpio_u_reg_u_reg_if_N17),
    .o(net192));
 b15bfn001as1n16x5 wire193 (.a(u_gpio_u_reg_u_reg_if_N16),
    .o(net193));
 b15bfn001ah1n48x5 wire194 (.a(n3292),
    .o(net194));
 b15bfn001ah1n32x5 wire195 (.a(net196),
    .o(net195));
 b15bfn001ah1n32x5 max_length196 (.a(n3292),
    .o(net196));
 b15bfn001as1n16x5 wire197 (.a(n3943),
    .o(net197));
 b15bfn001as1n32x5 wire198 (.a(n3938),
    .o(net198));
 b15bfn001ah1n24x5 wire199 (.a(net200),
    .o(net199));
 b15bfn001as1n24x5 max_length200 (.a(n3938),
    .o(net200));
 b15bfn001as1n24x5 fanout201 (.a(net202),
    .o(net201));
 b15bfn001as1n24x5 fanout202 (.a(n3429),
    .o(net202));
 b15bfn001as1n48x5 fanout203 (.a(net206),
    .o(net203));
 b15bfn001ah1n24x5 wire204 (.a(net205),
    .o(net204));
 b15bfn001as1n32x5 max_length205 (.a(net203),
    .o(net205));
 b15bfn001as1n48x5 fanout206 (.a(n3237),
    .o(net206));
 b15bfn001as1n48x5 wire207 (.a(net208),
    .o(net207));
 b15bfn001as1n32x5 wire208 (.a(net206),
    .o(net208));
 b15bfn001ah1n32x5 wire209 (.a(n3237),
    .o(net209));
 b15bfn001as1n24x5 fanout210 (.a(n3129),
    .o(net210));
 b15bfn000as1n24x5 fanout211 (.a(n3129),
    .o(net211));
 b15bfn000as1n24x5 fanout212 (.a(n3034),
    .o(net212));
 b15bfn001as1n16x5 fanout213 (.a(n3034),
    .o(net213));
 b15bfn001ah1n32x5 fanout214 (.a(n3032),
    .o(net214));
 b15bfn001ah1n24x5 fanout215 (.a(n3032),
    .o(net215));
 b15bfn000as1n24x5 fanout216 (.a(net217),
    .o(net216));
 b15bfn001as1n16x5 fanout217 (.a(n3030),
    .o(net217));
 b15bfn000as1n32x5 wire218 (.a(net217),
    .o(net218));
 b15bfn001as1n16x5 fanout219 (.a(net221),
    .o(net219));
 b15bfn001ah1n24x5 fanout220 (.a(n3028),
    .o(net220));
 b15bfn001ah1n24x5 wire221 (.a(n3028),
    .o(net221));
 b15bfn001as1n48x5 fanout222 (.a(net226),
    .o(net222));
 b15bfn001as1n32x5 wire223 (.a(net222),
    .o(net223));
 b15bfn001as1n32x5 max_length224 (.a(net222),
    .o(net224));
 b15bfn001ah1n64x5 fanout225 (.a(net226),
    .o(net225));
 b15bfn001ah1n32x5 wire226 (.a(n3936),
    .o(net226));
 b15bfn001ah1n48x5 load_slew227 (.a(n3256),
    .o(net227));
 b15bfn001ah1n16x5 fanout228 (.a(net229),
    .o(net228));
 b15bfn001as1n16x5 fanout229 (.a(net1824),
    .o(net229));
 b15bfn001as1n64x5 fanout230 (.a(n3819),
    .o(net230));
 b15bfn001as1n48x5 load_slew231 (.a(net230),
    .o(net231));
 b15bfn001ah1n48x5 max_length232 (.a(net230),
    .o(net232));
 b15bfn001as1n32x5 wire233 (.a(n3819),
    .o(net233));
 b15bfn001ah1n48x5 load_slew234 (.a(net235),
    .o(net234));
 b15bfn001as1n32x5 max_length235 (.a(net236),
    .o(net235));
 b15bfn001ah1n32x5 wire236 (.a(n3755),
    .o(net236));
 b15bfn001as1n24x5 wire237 (.a(u_gpio_u_reg_u_data_in_wr_data[23]),
    .o(net237));
 b15bfn001ah1n24x5 wire238 (.a(u_gpio_u_reg_u_data_in_wr_data[17]),
    .o(net238));
 b15bfn001as1n24x5 wire239 (.a(u_gpio_u_reg_u_data_in_wr_data[9]),
    .o(net239));
 b15bfn001ah1n24x5 wire240 (.a(u_gpio_u_reg_u_data_in_wr_data[20]),
    .o(net240));
 b15bfn001ah1n24x5 wire241 (.a(u_gpio_u_reg_u_data_in_wr_data[6]),
    .o(net241));
 b15bfn001as1n48x5 fanout242 (.a(n3760),
    .o(net242));
 b15bfn001ah1n32x5 max_length243 (.a(net245),
    .o(net243));
 b15bfn001ah1n48x5 max_length244 (.a(net245),
    .o(net244));
 b15bfn001ah1n48x5 load_slew245 (.a(net242),
    .o(net245));
 b15bfn001as1n32x5 wire246 (.a(net247),
    .o(net246));
 b15bfn001ah1n48x5 wire247 (.a(n3798),
    .o(net247));
 b15bfn000ah1n24x5 wire248 (.a(n3142),
    .o(net248));
 b15bfn001as1n12x5 fanout249 (.a(net250),
    .o(net249));
 b15bfn001as1n16x5 fanout250 (.a(net1778),
    .o(net250));
 b15bfn001as1n32x5 fanout251 (.a(net257),
    .o(net251));
 b15bfn001as1n32x5 wire252 (.a(net253),
    .o(net252));
 b15bfn001as1n32x5 wire253 (.a(net251),
    .o(net253));
 b15bfn001as1n48x5 fanout254 (.a(n3031),
    .o(net254));
 b15bfn001as1n48x5 max_length255 (.a(net256),
    .o(net255));
 b15bfn001as1n48x5 max_length256 (.a(net257),
    .o(net256));
 b15bfn001ah1n32x5 wire257 (.a(net254),
    .o(net257));
 b15bfn001as1n24x5 wire258 (.a(n3031),
    .o(net258));
 b15bfn001ah1n80x5 fanout259 (.a(net260),
    .o(net259));
 b15bfn001as1n80x5 fanout260 (.a(n3133),
    .o(net260));
 b15bfn001ah1n24x5 wire261 (.a(n3133),
    .o(net261));
 b15bfn001as1n48x5 fanout262 (.a(net267),
    .o(net262));
 b15bfn000ah1n48x5 wire263 (.a(net262),
    .o(net263));
 b15bfn001ah1n32x5 max_length264 (.a(net262),
    .o(net264));
 b15bfn001as1n64x5 fanout265 (.a(n3132),
    .o(net265));
 b15bfn001as1n24x5 wire266 (.a(net265),
    .o(net266));
 b15bfn001as1n48x5 max_length267 (.a(net265),
    .o(net267));
 b15bfn000ah1n24x5 wire268 (.a(n3132),
    .o(net268));
 b15bfn001as1n64x5 fanout269 (.a(n3797),
    .o(net269));
 b15bfn001ah1n24x5 wire270 (.a(net272),
    .o(net270));
 b15bfn001as1n32x5 max_length271 (.a(net273),
    .o(net271));
 b15bfn001as1n32x5 max_length272 (.a(net273),
    .o(net272));
 b15bfn001as1n32x5 max_length273 (.a(net269),
    .o(net273));
 b15bfn001as1n24x5 wire274 (.a(n3797),
    .o(net274));
 b15bfn001as1n24x5 fanout275 (.a(net278),
    .o(net275));
 b15bfn001ah1n48x5 load_slew276 (.a(net277),
    .o(net276));
 b15bfn001as1n32x5 wire277 (.a(net275),
    .o(net277));
 b15bfn001as1n80x5 fanout278 (.a(n3033),
    .o(net278));
 b15bfn000as1n24x5 wire279 (.a(n3033),
    .o(net279));
 b15bfn001ah1n16x5 wire280 (.a(net1819),
    .o(net280));
 b15bfn001ah1n16x5 wire281 (.a(u_gpio_reg2hw[198]),
    .o(net281));
 b15bfn001as1n12x5 wire282 (.a(u_gpio_reg2hw[222]),
    .o(net282));
 b15bfn001as1n08x5 wire283 (.a(net284),
    .o(net283));
 b15bfn001as1n16x5 wire284 (.a(u_gpio_reg2hw[163]),
    .o(net284));
 b15bfn001as1n16x5 wire285 (.a(u_gpio_reg2hw[162]),
    .o(net285));
 b15bfn001ah1n16x5 wire286 (.a(u_gpio_reg2hw[188]),
    .o(net286));
 b15bfn001ah1n24x5 wire287 (.a(net288),
    .o(net287));
 b15bfn001ah1n12x5 wire288 (.a(u_gpio_reg2hw[143]),
    .o(net288));
 b15bfn001ah1n12x5 wire289 (.a(u_gpio_reg2hw[143]),
    .o(net289));
 b15bfn001ah1n16x5 wire290 (.a(u_gpio_reg2hw[139]),
    .o(net290));
 b15bfn001as1n16x5 wire291 (.a(u_gpio_reg2hw[138]),
    .o(net291));
 b15bfn001ah1n16x5 wire292 (.a(u_gpio_reg2hw[59]),
    .o(net292));
 b15bfn001ah1n12x5 load_slew293 (.a(u_gpio_reg2hw[54]),
    .o(net293));
 b15bfn001ah1n12x5 wire294 (.a(u_gpio_reg2hw[45]),
    .o(net294));
 b15bfn001as1n12x5 wire295 (.a(u_gpio_reg2hw[45]),
    .o(net295));
 b15bfn001ah1n16x5 wire296 (.a(u_gpio_reg2hw[44]),
    .o(net296));
 b15bfn001ah1n16x5 wire297 (.a(u_gpio_reg2hw[43]),
    .o(net297));
 b15bfn001ah1n16x5 wire298 (.a(u_gpio_reg2hw[42]),
    .o(net298));
 b15bfn001ah1n16x5 wire299 (.a(u_gpio_reg2hw[73]),
    .o(net299));
 b15bfn001ah1n16x5 wire300 (.a(u_gpio_reg2hw[72]),
    .o(net300));
 b15bfn001as1n24x5 wire301 (.a(net302),
    .o(net301));
 b15bfn001ah1n16x5 wire302 (.a(net303),
    .o(net302));
 b15bfn001ah1n12x5 wire303 (.a(u_gpio_reg2hw[95]),
    .o(net303));
 b15bfn000ah1n24x5 wire304 (.a(u_gpio_reg2hw[66]),
    .o(net304));
 b15bfn001ah1n16x5 wire305 (.a(u_gpio_reg2hw[87]),
    .o(net305));
 b15bfn001as1n16x5 wire306 (.a(u_gpio_reg2hw[82]),
    .o(net306));
 b15bfn001ah1n12x5 wire307 (.a(net308),
    .o(net307));
 b15bfn001as1n08x5 wire308 (.a(u_gpio_reg2hw[80]),
    .o(net308));
 b15bfn001ah1n16x5 wire309 (.a(u_gpio_reg2hw[79]),
    .o(net309));
 b15bfn001ah1n16x5 wire310 (.a(u_gpio_reg2hw[75]),
    .o(net310));
 b15bfn001as1n16x5 wire311 (.a(u_gpio_reg2hw[74]),
    .o(net311));
 b15bfn001ah1n16x5 wire312 (.a(u_gpio_reg2hw[122]),
    .o(net312));
 b15bfn001as1n16x5 wire313 (.a(u_gpio_reg2hw[111]),
    .o(net313));
 b15bfn001as1n16x5 wire314 (.a(u_gpio_reg2hw[107]),
    .o(net314));
 b15bfn001ah1n24x5 wire315 (.a(u_gpio_reg2hw[106]),
    .o(net315));
 b15bfn001ah1n24x5 wire316 (.a(net317),
    .o(net316));
 b15bfn001ah1n12x5 wire317 (.a(u_gpio_reg2hw[96]),
    .o(net317));
 b15bfn001ah1n12x5 wire318 (.a(u_gpio_reg2hw[9]),
    .o(net318));
 b15bfn001ah1n12x5 wire319 (.a(u_gpio_reg2hw[8]),
    .o(net319));
 b15bfn001ah1n12x5 load_slew320 (.a(u_gpio_reg2hw[7]),
    .o(net320));
 b15bfn001as1n12x5 load_slew321 (.a(u_gpio_reg2hw[7]),
    .o(net321));
 b15bfn001ah1n16x5 max_cap322 (.a(u_gpio_reg2hw[6]),
    .o(net322));
 b15bfn001ah1n16x5 wire323 (.a(u_gpio_reg2hw[5]),
    .o(net323));
 b15bfn001as1n16x5 wire324 (.a(u_gpio_reg2hw[5]),
    .o(net324));
 b15bfn001ah1n12x5 wire325 (.a(net326),
    .o(net325));
 b15bfn001as1n12x5 wire326 (.a(u_gpio_reg2hw[4]),
    .o(net326));
 b15bfn000as1n12x5 wire327 (.a(u_gpio_reg2hw[3]),
    .o(net327));
 b15bfn001ah1n12x5 load_slew328 (.a(u_gpio_reg2hw[3]),
    .o(net328));
 b15bfn001as1n12x5 wire329 (.a(u_gpio_reg2hw[2]),
    .o(net329));
 b15bfn001ah1n12x5 wire330 (.a(u_gpio_reg2hw[2]),
    .o(net330));
 b15bfn001ah1n16x5 max_cap331 (.a(u_gpio_reg2hw[29]),
    .o(net331));
 b15bfn001ah1n12x5 load_slew332 (.a(net333),
    .o(net332));
 b15bfn001ah1n12x5 wire333 (.a(u_gpio_reg2hw[28]),
    .o(net333));
 b15bfn001as1n12x5 max_cap334 (.a(u_gpio_reg2hw[27]),
    .o(net334));
 b15bfn001as1n12x5 max_cap335 (.a(u_gpio_reg2hw[25]),
    .o(net335));
 b15bfn001as1n08x5 load_slew336 (.a(net337),
    .o(net336));
 b15bfn001as1n08x5 wire337 (.a(u_gpio_reg2hw[24]),
    .o(net337));
 b15bfn000ah1n12x5 wire338 (.a(u_gpio_reg2hw[23]),
    .o(net338));
 b15bfn001ah1n12x5 load_slew339 (.a(u_gpio_reg2hw[22]),
    .o(net339));
 b15bfn001as1n08x5 load_slew340 (.a(u_gpio_reg2hw[22]),
    .o(net340));
 b15bfn001ah1n12x5 wire341 (.a(u_gpio_reg2hw[21]),
    .o(net341));
 b15bfn001as1n12x5 wire342 (.a(u_gpio_reg2hw[21]),
    .o(net342));
 b15bfn001as1n12x5 wire343 (.a(u_gpio_reg2hw[20]),
    .o(net343));
 b15bfn001as1n12x5 wire344 (.a(net345),
    .o(net344));
 b15bfn001ah1n16x5 wire345 (.a(u_gpio_reg2hw[19]),
    .o(net345));
 b15bfn001ah1n12x5 load_slew346 (.a(net347),
    .o(net346));
 b15bfn001ah1n12x5 wire347 (.a(u_gpio_reg2hw[18]),
    .o(net347));
 b15bfn001as1n12x5 wire348 (.a(u_gpio_reg2hw[16]),
    .o(net348));
 b15bfn001ah1n12x5 load_slew349 (.a(net350),
    .o(net349));
 b15bfn001as1n08x5 load_slew350 (.a(net2212),
    .o(net350));
 b15bfn001as1n16x5 wire351 (.a(net352),
    .o(net351));
 b15bfn001as1n12x5 wire352 (.a(net1948),
    .o(net352));
 b15bfn001ah1n12x5 wire353 (.a(net2127),
    .o(net353));
 b15bfn001ah1n16x5 wire354 (.a(u_gpio_reg2hw[13]),
    .o(net354));
 b15bfn001as1n08x5 wire355 (.a(net2216),
    .o(net355));
 b15bfn001ah1n12x5 wire356 (.a(net1986),
    .o(net356));
 b15bfn001as1n12x5 wire357 (.a(net2211),
    .o(net357));
 b15bfn001ah1n12x5 wire358 (.a(net359),
    .o(net358));
 b15bfn001ah1n16x5 wire359 (.a(net110),
    .o(net359));
 b15bfn001ah1n12x5 wire360 (.a(net109),
    .o(net360));
 b15bfn001as1n08x5 wire361 (.a(net362),
    .o(net361));
 b15bfn001ah1n16x5 wire362 (.a(net109),
    .o(net362));
 b15bfn001as1n12x5 load_slew363 (.a(net103),
    .o(net363));
 b15bfn001as1n08x5 load_slew364 (.a(net102),
    .o(net364));
 b15bfn001as1n12x5 wire365 (.a(net366),
    .o(net365));
 b15bfn001ah1n12x5 load_slew366 (.a(net102),
    .o(net366));
 b15bfn001ah1n16x5 wire367 (.a(net100),
    .o(net367));
 b15bfn001as1n16x5 wire368 (.a(net98),
    .o(net368));
 b15bfn001ah1n16x5 wire369 (.a(net97),
    .o(net369));
 b15bfn001ah1n16x5 wire370 (.a(net96),
    .o(net370));
 b15bfn001as1n12x5 wire371 (.a(net372),
    .o(net371));
 b15bfn001ah1n12x5 load_slew372 (.a(net95),
    .o(net372));
 b15bfn001as1n16x5 wire373 (.a(net374),
    .o(net373));
 b15bfn001as1n06x5 load_slew374 (.a(net94),
    .o(net374));
 b15bfn001as1n12x5 wire375 (.a(net376),
    .o(net375));
 b15bfn001ah1n12x5 load_slew376 (.a(net93),
    .o(net376));
 b15bfn001as1n12x5 wire377 (.a(net92),
    .o(net377));
 b15bfn001ah1n16x5 max_cap378 (.a(net91),
    .o(net378));
 b15bfn001ah1n12x5 load_slew379 (.a(net89),
    .o(net379));
 b15bfn001ah1n12x5 load_slew380 (.a(net89),
    .o(net380));
 b15bfn001as1n08x5 load_slew381 (.a(net382),
    .o(net381));
 b15bfn001as1n12x5 wire382 (.a(net87),
    .o(net382));
 b15bfn001ah1n16x5 wire383 (.a(net384),
    .o(net383));
 b15bfn001ah1n12x5 load_slew384 (.a(net86),
    .o(net384));
 b15bfn001ah1n16x5 wire385 (.a(net2204),
    .o(net385));
 b15bfn001ah1n16x5 wire386 (.a(net2121),
    .o(net386));
 b15bfn001as1n06x5 load_slew387 (.a(net82),
    .o(net387));
 b15bfn001ah1n16x5 wire388 (.a(net81),
    .o(net388));
 b15bfn001ah1n16x5 wire389 (.a(net80),
    .o(net389));
 b15bfn001ah1n12x5 wire390 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[15]),
    .o(net390));
 b15bfn001as1n12x5 wire391 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[15]),
    .o(net391));
 b15bfn001as1n12x5 wire392 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[14]),
    .o(net392));
 b15bfn001ah1n12x5 wire393 (.a(u_gpio_u_reg_masked_oe_lower_data_qs[2]),
    .o(net393));
 b15bfn001ah1n16x5 max_cap394 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[12]),
    .o(net394));
 b15bfn001ah1n16x5 max_cap395 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[12]),
    .o(net395));
 b15bfn001ah1n16x5 wire396 (.a(net397),
    .o(net396));
 b15bfn001ah1n16x5 wire397 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[11]),
    .o(net397));
 b15bfn001as1n12x5 load_slew398 (.a(net399),
    .o(net398));
 b15bfn001ah1n12x5 wire399 (.a(net2146),
    .o(net399));
 b15bfn001ah1n12x5 wire400 (.a(net401),
    .o(net400));
 b15bfn001ah1n12x5 wire401 (.a(net2125),
    .o(net401));
 b15bfn001ah1n12x5 load_slew402 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[8]),
    .o(net402));
 b15bfn001as1n08x5 load_slew403 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[8]),
    .o(net403));
 b15bfn001as1n12x5 wire404 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[7]),
    .o(net404));
 b15bfn001ah1n12x5 load_slew405 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[7]),
    .o(net405));
 b15bfn001as1n12x5 wire406 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[6]),
    .o(net406));
 b15bfn001ah1n24x5 wire407 (.a(net408),
    .o(net407));
 b15bfn001ah1n12x5 load_slew408 (.a(net409),
    .o(net408));
 b15bfn001ah1n12x5 load_slew409 (.a(net410),
    .o(net409));
 b15bfn001ah1n12x5 wire410 (.a(net2197),
    .o(net410));
 b15bfn001ah1n16x5 wire411 (.a(u_gpio_u_reg_masked_oe_upper_data_qs[0]),
    .o(net411));
 b15bfn001as1n16x5 wire412 (.a(net413),
    .o(net412));
 b15bfn001ah1n16x5 wire413 (.a(u_gpio_u_reg_masked_oe_lower_data_qs[11]),
    .o(net413));
 b15bfn001as1n48x5 fanout414 (.a(n3761),
    .o(net414));
 b15bfn001as1n32x5 wire415 (.a(net417),
    .o(net415));
 b15bfn001as1n32x5 wire416 (.a(net418),
    .o(net416));
 b15bfn001ah1n32x5 max_length417 (.a(net418),
    .o(net417));
 b15bfn001ah1n48x5 load_slew418 (.a(net414),
    .o(net418));
 b15bfn001as1n32x5 wire419 (.a(n3761),
    .o(net419));
 b15bfn001ah1n64x5 fanout420 (.a(n3665),
    .o(net420));
 b15bfn001as1n48x5 fanout421 (.a(n3665),
    .o(net421));
 b15bfn001ah1n24x5 max_length422 (.a(net421),
    .o(net422));
 b15bfn001as1n48x5 fanout423 (.a(net426),
    .o(net423));
 b15bfn001as1n32x5 wire424 (.a(net425),
    .o(net424));
 b15bfn001ah1n48x5 load_slew425 (.a(net423),
    .o(net425));
 b15bfn001as1n64x5 fanout426 (.a(n3029),
    .o(net426));
 b15bfn001ah1n48x5 max_length427 (.a(net428),
    .o(net427));
 b15bfn001aq1n48x5 wire428 (.a(net426),
    .o(net428));
 b15bfn001as1n24x5 wire429 (.a(n3029),
    .o(net429));
 b15bfn001as1n48x5 fanout430 (.a(net433),
    .o(net430));
 b15bfn001ah1n32x5 max_length431 (.a(net430),
    .o(net431));
 b15bfn001ah1n32x5 max_length432 (.a(net430),
    .o(net432));
 b15bfn001as1n80x5 fanout433 (.a(n3027),
    .o(net433));
 b15bfn001ah1n16x5 wire434 (.a(net1765),
    .o(net434));
 b15bfn001ah1n16x5 wire435 (.a(u_gpio_u_reg_data_in_qs[7]),
    .o(net435));
 b15bfn001as1n24x5 wire436 (.a(net437),
    .o(net436));
 b15bfn001ah1n16x5 wire437 (.a(u_gpio_u_reg_data_in_qs[12]),
    .o(net437));
 b15bfn001ah1n24x5 wire438 (.a(u_gpio_u_reg_data_in_qs[15]),
    .o(net438));
 b15bfn001as1n08x5 wire439 (.a(u_gpio_gen_filter_9__u_filter_filter_synced),
    .o(net439));
 b15bfn001as1n12x5 wire440 (.a(net2094),
    .o(net440));
 b15bfn001ah1n16x5 wire441 (.a(net2047),
    .o(net441));
 b15bfn001as1n08x5 load_slew442 (.a(net443),
    .o(net442));
 b15bfn001as1n08x5 wire443 (.a(net1961),
    .o(net443));
 b15bfn001as1n12x5 wire444 (.a(net445),
    .o(net444));
 b15bfn001as1n12x5 wire445 (.a(net2162),
    .o(net445));
 b15bfn001ah1n12x5 wire446 (.a(net1998),
    .o(net446));
 b15bfn001ah1n12x5 wire447 (.a(u_gpio_gen_filter_19__u_filter_filter_synced),
    .o(net447));
 b15bfn001as1n12x5 wire448 (.a(u_gpio_gen_filter_18__u_filter_filter_synced),
    .o(net448));
 b15bfn001as1n08x5 load_slew449 (.a(net450),
    .o(net449));
 b15bfn001as1n08x5 wire450 (.a(net1979),
    .o(net450));
 b15bfn001as1n08x5 load_slew451 (.a(u_gpio_gen_filter_14__u_filter_filter_synced),
    .o(net451));
 b15bfn001as1n08x5 load_slew452 (.a(u_gpio_gen_filter_12__u_filter_filter_synced),
    .o(net452));
 b15bfn001ah1n16x5 wire453 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q),
    .o(net453));
 b15bfn001as1n16x5 wire454 (.a(u_gpio_gen_alert_tx_0__u_prim_alert_sender_n1),
    .o(net454));
 b15bfn001ah1n64x5 fanout455 (.a(net457),
    .o(net455));
 b15bfn001as1n48x5 fanout456 (.a(n3135),
    .o(net456));
 b15bfn001as1n48x5 max_length457 (.a(net458),
    .o(net457));
 b15bfn001ah1n32x5 wire458 (.a(net456),
    .o(net458));
 b15bfn001ah1n32x5 wire459 (.a(n3135),
    .o(net459));
 b15bfn000as1n24x5 wire460 (.a(net461),
    .o(net460));
 b15bfn001as1n32x5 wire461 (.a(n3548),
    .o(net461));
 b15bfn001ah1n32x5 max_length462 (.a(net463),
    .o(net462));
 b15bfn001as1n24x5 wire463 (.a(n3551),
    .o(net463));
 b15bfn001ah1n24x5 wire464 (.a(n3553),
    .o(net464));
 b15bfn001as1n24x5 wire465 (.a(n3553),
    .o(net465));
 b15bfn001as1n24x5 wire466 (.a(net467),
    .o(net466));
 b15bfn000as1n24x5 wire467 (.a(n3547),
    .o(net467));
 b15bfn001as1n24x5 wire468 (.a(net469),
    .o(net468));
 b15bfn001as1n32x5 wire469 (.a(n3552),
    .o(net469));
 b15bfn001ah1n24x5 wire470 (.a(net471),
    .o(net470));
 b15bfn001as1n32x5 max_length471 (.a(n3549),
    .o(net471));
 b15bfn001as1n24x5 wire472 (.a(net473),
    .o(net472));
 b15bfn001as1n24x5 max_length473 (.a(n3545),
    .o(net473));
 b15bfn000as1n24x5 wire474 (.a(net475),
    .o(net474));
 b15bfn001ah1n32x5 wire475 (.a(n3542),
    .o(net475));
 b15bfn001ah1n24x5 wire476 (.a(n3550),
    .o(net476));
 b15bfn001ah1n24x5 wire477 (.a(n3550),
    .o(net477));
 b15bfn001as1n16x5 max_length478 (.a(net479),
    .o(net478));
 b15bfn001as1n24x5 wire479 (.a(net480),
    .o(net479));
 b15bfn001as1n32x5 max_length480 (.a(n3906),
    .o(net480));
 b15bfn001as1n24x5 wire481 (.a(n3905),
    .o(net481));
 b15bfn001ah1n24x5 max_length482 (.a(n3905),
    .o(net482));
 b15bfn001as1n24x5 max_length483 (.a(n3905),
    .o(net483));
 b15bfn001as1n24x5 wire484 (.a(net485),
    .o(net484));
 b15bfn001ah1n32x5 max_length485 (.a(n3903),
    .o(net485));
 b15bfn001ah1n24x5 max_length486 (.a(net487),
    .o(net486));
 b15bfn001as1n32x5 wire487 (.a(n3898),
    .o(net487));
 b15bfn001ah1n24x5 max_length488 (.a(net489),
    .o(net488));
 b15bfn001ah1n32x5 wire489 (.a(n3897),
    .o(net489));
 b15bfn001ah1n32x5 max_length490 (.a(net491),
    .o(net490));
 b15bfn001ah1n32x5 max_length491 (.a(n3896),
    .o(net491));
 b15bfn001ah1n24x5 max_length492 (.a(n3895),
    .o(net492));
 b15bfn001ah1n24x5 max_length493 (.a(n3895),
    .o(net493));
 b15bfn001as1n16x5 max_length494 (.a(n3894),
    .o(net494));
 b15bfn000as1n24x5 wire495 (.a(n3894),
    .o(net495));
 b15bfn001ah1n24x5 wire496 (.a(n3892),
    .o(net496));
 b15bfn001as1n24x5 wire497 (.a(net498),
    .o(net497));
 b15bfn001ah1n32x5 max_length498 (.a(n3892),
    .o(net498));
 b15bfn001ah1n32x5 max_length499 (.a(net500),
    .o(net499));
 b15bfn001ah1n24x5 max_length500 (.a(net501),
    .o(net500));
 b15bfn001ah1n24x5 wire501 (.a(n3891),
    .o(net501));
 b15bfn001as1n32x5 wire502 (.a(net38),
    .o(net502));
 b15bfn000as1n32x5 wire503 (.a(net37),
    .o(net503));
 b15bfn001as1n32x5 wire504 (.a(net30),
    .o(net504));
 b15bfn001as1n32x5 wire505 (.a(net29),
    .o(net505));
 b15bfn001as1n32x5 wire506 (.a(net22),
    .o(net506));
 b15bfn001as1n32x5 wire507 (.a(net21),
    .o(net507));
 b15bfn001as1n32x5 wire508 (.a(net14),
    .o(net508));
 b15bfn001ah1n16x5 max_length509 (.a(net13),
    .o(net509));
 b15bfn001as1n48x5 fanout510 (.a(net511),
    .o(net510));
 b15bfn001ah1n64x5 fanout511 (.a(net542),
    .o(net511));
 b15bfn001ah1n64x5 fanout512 (.a(net514),
    .o(net512));
 b15bfn001ah1n64x5 fanout513 (.a(net514),
    .o(net513));
 b15bfn001as1n48x5 fanout514 (.a(net542),
    .o(net514));
 b15bfn001ah1n64x5 fanout515 (.a(net518),
    .o(net515));
 b15bfn001as1n32x5 fanout516 (.a(net518),
    .o(net516));
 b15bfn001as1n32x5 fanout517 (.a(net518),
    .o(net517));
 b15bfn001as1n48x5 fanout518 (.a(net541),
    .o(net518));
 b15bfn001as1n48x5 fanout519 (.a(net523),
    .o(net519));
 b15bfn001as1n24x5 fanout520 (.a(net523),
    .o(net520));
 b15bfn001as1n48x5 fanout521 (.a(net523),
    .o(net521));
 b15bfn001ah1n48x5 fanout522 (.a(net523),
    .o(net522));
 b15bfn001ah1n48x5 fanout523 (.a(net541),
    .o(net523));
 b15bfn001as1n48x5 fanout524 (.a(net526),
    .o(net524));
 b15bfn001ah1n64x5 fanout525 (.a(net526),
    .o(net525));
 b15bfn001as1n48x5 fanout526 (.a(net539),
    .o(net526));
 b15bfn001ah1n48x5 fanout527 (.a(net528),
    .o(net527));
 b15bfn001ah1n64x5 fanout528 (.a(net539),
    .o(net528));
 b15bfn001ah1n48x5 fanout529 (.a(net540),
    .o(net529));
 b15bfn001as1n32x5 fanout530 (.a(net540),
    .o(net530));
 b15bfn001ah1n48x5 fanout531 (.a(net540),
    .o(net531));
 b15bfn001ah1n48x5 fanout532 (.a(net538),
    .o(net532));
 b15bfn001as1n48x5 fanout533 (.a(net537),
    .o(net533));
 b15bfn001ah1n48x5 fanout534 (.a(net537),
    .o(net534));
 b15bfn001as1n48x5 fanout535 (.a(net537),
    .o(net535));
 b15bfn001ah1n48x5 fanout536 (.a(net537),
    .o(net536));
 b15bfn001ah1n48x5 fanout537 (.a(net538),
    .o(net537));
 b15bfn001as1n64x5 fanout538 (.a(net541),
    .o(net538));
 b15bfn001as1n32x5 wire539 (.a(net540),
    .o(net539));
 b15bfn001as1n32x5 load_slew540 (.a(net538),
    .o(net540));
 b15bfn001as1n48x5 fanout541 (.a(net1),
    .o(net541));
 b15bfn001ah1n48x5 wire542 (.a(net541),
    .o(net542));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_0__u_gpio_cio_gpio_en_q_reg_1__543 (.o(net543));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_0__u_gpio_cio_gpio_en_q_reg_1__544 (.o(net544));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_10__u_gpio_cio_gpio_en_q_reg_11__545 (.o(net545));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_10__u_gpio_cio_gpio_en_q_reg_11__546 (.o(net546));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_12__u_gpio_cio_gpio_en_q_reg_13__547 (.o(net547));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_12__u_gpio_cio_gpio_en_q_reg_13__548 (.o(net548));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_14__u_gpio_cio_gpio_en_q_reg_15__549 (.o(net549));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_14__u_gpio_cio_gpio_en_q_reg_15__550 (.o(net550));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_16__u_gpio_cio_gpio_en_q_reg_17__551 (.o(net551));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_16__u_gpio_cio_gpio_en_q_reg_17__552 (.o(net552));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_18__u_gpio_cio_gpio_en_q_reg_19__553 (.o(net553));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_18__u_gpio_cio_gpio_en_q_reg_19__554 (.o(net554));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_20__u_gpio_cio_gpio_en_q_reg_21__555 (.o(net555));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_20__u_gpio_cio_gpio_en_q_reg_21__556 (.o(net556));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_22__u_gpio_cio_gpio_en_q_reg_23__557 (.o(net557));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_22__u_gpio_cio_gpio_en_q_reg_23__558 (.o(net558));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_24__u_gpio_cio_gpio_en_q_reg_25__559 (.o(net559));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_24__u_gpio_cio_gpio_en_q_reg_25__560 (.o(net560));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_26__u_gpio_cio_gpio_en_q_reg_27__561 (.o(net561));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_26__u_gpio_cio_gpio_en_q_reg_27__562 (.o(net562));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_28__u_gpio_cio_gpio_en_q_reg_29__563 (.o(net563));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_28__u_gpio_cio_gpio_en_q_reg_29__564 (.o(net564));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_2__u_gpio_cio_gpio_en_q_reg_3__565 (.o(net565));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_2__u_gpio_cio_gpio_en_q_reg_3__566 (.o(net566));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_30__u_gpio_cio_gpio_en_q_reg_31__567 (.o(net567));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_30__u_gpio_cio_gpio_en_q_reg_31__568 (.o(net568));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_4__u_gpio_cio_gpio_en_q_reg_5__569 (.o(net569));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_4__u_gpio_cio_gpio_en_q_reg_5__570 (.o(net570));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_6__u_gpio_cio_gpio_en_q_reg_7__571 (.o(net571));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_6__u_gpio_cio_gpio_en_q_reg_7__572 (.o(net572));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_8__u_gpio_cio_gpio_en_q_reg_9__573 (.o(net573));
 b15tilo00an1n03x5 u_gpio_cio_gpio_en_q_reg_8__u_gpio_cio_gpio_en_q_reg_9__574 (.o(net574));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_0__u_gpio_cio_gpio_q_reg_1__575 (.o(net575));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_0__u_gpio_cio_gpio_q_reg_1__576 (.o(net576));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_10__u_gpio_cio_gpio_q_reg_11__577 (.o(net577));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_10__u_gpio_cio_gpio_q_reg_11__578 (.o(net578));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_12__u_gpio_cio_gpio_q_reg_13__579 (.o(net579));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_12__u_gpio_cio_gpio_q_reg_13__580 (.o(net580));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_14__u_gpio_cio_gpio_q_reg_15__581 (.o(net581));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_14__u_gpio_cio_gpio_q_reg_15__582 (.o(net582));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_16__u_gpio_cio_gpio_q_reg_17__583 (.o(net583));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_16__u_gpio_cio_gpio_q_reg_17__584 (.o(net584));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_18__u_gpio_cio_gpio_q_reg_19__585 (.o(net585));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_18__u_gpio_cio_gpio_q_reg_19__586 (.o(net586));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_20__u_gpio_cio_gpio_q_reg_21__587 (.o(net587));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_20__u_gpio_cio_gpio_q_reg_21__588 (.o(net588));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_22__u_gpio_cio_gpio_q_reg_23__589 (.o(net589));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_22__u_gpio_cio_gpio_q_reg_23__590 (.o(net590));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_24__u_gpio_cio_gpio_q_reg_25__591 (.o(net591));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_24__u_gpio_cio_gpio_q_reg_25__592 (.o(net592));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_26__u_gpio_cio_gpio_q_reg_27__593 (.o(net593));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_26__u_gpio_cio_gpio_q_reg_27__594 (.o(net594));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_28__u_gpio_cio_gpio_q_reg_29__595 (.o(net595));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_28__u_gpio_cio_gpio_q_reg_29__596 (.o(net596));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_2__u_gpio_cio_gpio_q_reg_3__597 (.o(net597));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_2__u_gpio_cio_gpio_q_reg_3__598 (.o(net598));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_30__u_gpio_cio_gpio_q_reg_31__599 (.o(net599));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_30__u_gpio_cio_gpio_q_reg_31__600 (.o(net600));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_4__u_gpio_cio_gpio_q_reg_5__601 (.o(net601));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_4__u_gpio_cio_gpio_q_reg_5__602 (.o(net602));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_6__u_gpio_cio_gpio_q_reg_7__603 (.o(net603));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_6__u_gpio_cio_gpio_q_reg_7__604 (.o(net604));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_8__u_gpio_cio_gpio_q_reg_9__605 (.o(net605));
 b15tilo00an1n03x5 u_gpio_cio_gpio_q_reg_8__u_gpio_cio_gpio_q_reg_9__606 (.o(net606));
 b15tilo00an1n03x5 u_gpio_clk_gate_cio_gpio_en_q_reg_0_latch_607 (.o(net607));
 b15tilo00an1n03x5 u_gpio_clk_gate_cio_gpio_en_q_reg_latch_608 (.o(net608));
 b15tilo00an1n03x5 u_gpio_clk_gate_cio_gpio_q_reg_0_latch_609 (.o(net609));
 b15tilo00an1n03x5 u_gpio_clk_gate_cio_gpio_q_reg_latch_610 (.o(net610));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_0__u_gpio_data_in_q_reg_1__611 (.o(net611));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_0__u_gpio_data_in_q_reg_1__612 (.o(net612));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_10__u_gpio_data_in_q_reg_11__613 (.o(net613));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_10__u_gpio_data_in_q_reg_11__614 (.o(net614));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_12__u_gpio_data_in_q_reg_13__615 (.o(net615));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_12__u_gpio_data_in_q_reg_13__616 (.o(net616));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_14__u_gpio_data_in_q_reg_15__617 (.o(net617));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_14__u_gpio_data_in_q_reg_15__618 (.o(net618));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_16__u_gpio_data_in_q_reg_17__619 (.o(net619));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_16__u_gpio_data_in_q_reg_17__620 (.o(net620));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_18__u_gpio_data_in_q_reg_19__621 (.o(net621));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_18__u_gpio_data_in_q_reg_19__622 (.o(net622));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_20__u_gpio_data_in_q_reg_21__623 (.o(net623));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_20__u_gpio_data_in_q_reg_21__624 (.o(net624));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_22__u_gpio_data_in_q_reg_23__625 (.o(net625));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_22__u_gpio_data_in_q_reg_23__626 (.o(net626));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_24__u_gpio_data_in_q_reg_25__627 (.o(net627));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_24__u_gpio_data_in_q_reg_25__628 (.o(net628));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_26__u_gpio_data_in_q_reg_27__629 (.o(net629));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_26__u_gpio_data_in_q_reg_27__630 (.o(net630));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_28__u_gpio_data_in_q_reg_29__631 (.o(net631));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_28__u_gpio_data_in_q_reg_29__632 (.o(net632));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_2__u_gpio_data_in_q_reg_3__633 (.o(net633));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_2__u_gpio_data_in_q_reg_3__634 (.o(net634));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_30__u_gpio_data_in_q_reg_31__635 (.o(net635));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_30__u_gpio_data_in_q_reg_31__636 (.o(net636));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_4__u_gpio_data_in_q_reg_5__637 (.o(net637));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_4__u_gpio_data_in_q_reg_5__638 (.o(net638));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_6__u_gpio_data_in_q_reg_7__639 (.o(net639));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_6__u_gpio_data_in_q_reg_7__640 (.o(net640));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_8__u_gpio_data_in_q_reg_9__641 (.o(net641));
 b15tilo00an1n03x5 u_gpio_data_in_q_reg_8__u_gpio_data_in_q_reg_9__642 (.o(net642));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_set_q_reg_u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_0__643 (.o(net643));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_set_q_reg_u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_0__644 (.o(net644));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q_reg_u_gpio_gen_alert_tx_0__u_prim_alert_sender_ping_set_q_reg_645 (.o(net645));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q_reg_u_gpio_gen_alert_tx_0__u_prim_alert_sender_ping_set_q_reg_646 (.o(net646));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_0__u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_1__647 (.o(net647));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_0__u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_1__648 (.o(net648));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_2__u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq_reg_649 (.o(net649));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_2__u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq_reg_650 (.o(net650));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq_reg_651 (.o(net651));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__652 (.o(net652));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__653 (.o(net653));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__654 (.o(net654));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__655 (.o(net655));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__656 (.o(net656));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__657 (.o(net657));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q_reg_658 (.o(net658));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q_reg_659 (.o(net659));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_0__660 (.o(net660));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_1__661 (.o(net661));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq_reg_662 (.o(net662));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq_reg_u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__663 (.o(net663));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq_reg_u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__664 (.o(net664));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__665 (.o(net665));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__666 (.o(net666));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_0__667 (.o(net667));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_1__668 (.o(net668));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q_reg_u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_0__669 (.o(net669));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q_reg_u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_0__670 (.o(net670));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_16__u_filter_filter_q_reg_671 (.o(net671));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_16__u_filter_filter_q_reg_672 (.o(net672));
 b15tilo00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_1__673 (.o(net673));
 b15tilo00an1n03x5 u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_1__674 (.o(net674));
 b15tilo00an1n03x5 u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_1__675 (.o(net675));
 b15tilo00an1n03x5 u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_3__676 (.o(net676));
 b15tilo00an1n03x5 u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_3__677 (.o(net677));
 b15tilo00an1n03x5 u_gpio_gen_filter_0__u_filter_filter_q_reg_u_gpio_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__678 (.o(net678));
 b15tilo00an1n03x5 u_gpio_gen_filter_0__u_filter_filter_q_reg_u_gpio_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__679 (.o(net679));
 b15tilo00an1n03x5 u_gpio_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__680 (.o(net680));
 b15tilo00an1n03x5 u_gpio_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__681 (.o(net681));
 b15tilo00an1n03x5 u_gpio_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__682 (.o(net682));
 b15tilo00an1n03x5 u_gpio_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__683 (.o(net683));
 b15tilo00an1n03x5 u_gpio_gen_filter_0__u_filter_stored_value_q_reg_684 (.o(net684));
 b15tilo00an1n03x5 u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_1__685 (.o(net685));
 b15tilo00an1n03x5 u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_1__686 (.o(net686));
 b15tilo00an1n03x5 u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_10__u_filter_filter_q_reg_687 (.o(net687));
 b15tilo00an1n03x5 u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_10__u_filter_filter_q_reg_688 (.o(net688));
 b15tilo00an1n03x5 u_gpio_gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__689 (.o(net689));
 b15tilo00an1n03x5 u_gpio_gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__690 (.o(net690));
 b15tilo00an1n03x5 u_gpio_gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__691 (.o(net691));
 b15tilo00an1n03x5 u_gpio_gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__692 (.o(net692));
 b15tilo00an1n03x5 u_gpio_gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_0__693 (.o(net693));
 b15tilo00an1n03x5 u_gpio_gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_0__694 (.o(net694));
 b15tilo00an1n03x5 u_gpio_gen_filter_10__u_filter_stored_value_q_reg_695 (.o(net695));
 b15tilo00an1n03x5 u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_2__696 (.o(net696));
 b15tilo00an1n03x5 u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_2__697 (.o(net697));
 b15tilo00an1n03x5 u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_11__u_filter_filter_q_reg_698 (.o(net698));
 b15tilo00an1n03x5 u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_11__u_filter_filter_q_reg_699 (.o(net699));
 b15tilo00an1n03x5 u_gpio_gen_filter_11__u_filter_stored_value_q_reg_700 (.o(net700));
 b15tilo00an1n03x5 u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_2__701 (.o(net701));
 b15tilo00an1n03x5 u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_2__702 (.o(net702));
 b15tilo00an1n03x5 u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_12__u_filter_filter_q_reg_703 (.o(net703));
 b15tilo00an1n03x5 u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_12__u_filter_filter_q_reg_704 (.o(net704));
 b15tilo00an1n03x5 u_gpio_gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__705 (.o(net705));
 b15tilo00an1n03x5 u_gpio_gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__706 (.o(net706));
 b15tilo00an1n03x5 u_gpio_gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__707 (.o(net707));
 b15tilo00an1n03x5 u_gpio_gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__708 (.o(net708));
 b15tilo00an1n03x5 u_gpio_gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_0__709 (.o(net709));
 b15tilo00an1n03x5 u_gpio_gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_0__710 (.o(net710));
 b15tilo00an1n03x5 u_gpio_gen_filter_12__u_filter_stored_value_q_reg_711 (.o(net711));
 b15tilo00an1n03x5 u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_1__712 (.o(net712));
 b15tilo00an1n03x5 u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_1__713 (.o(net713));
 b15tilo00an1n03x5 u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_3__714 (.o(net714));
 b15tilo00an1n03x5 u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_3__715 (.o(net715));
 b15tilo00an1n03x5 u_gpio_gen_filter_13__u_filter_filter_q_reg_u_gpio_gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__716 (.o(net716));
 b15tilo00an1n03x5 u_gpio_gen_filter_13__u_filter_filter_q_reg_u_gpio_gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__717 (.o(net717));
 b15tilo00an1n03x5 u_gpio_gen_filter_13__u_filter_stored_value_q_reg_718 (.o(net718));
 b15tilo00an1n03x5 u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_2__719 (.o(net719));
 b15tilo00an1n03x5 u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_2__720 (.o(net720));
 b15tilo00an1n03x5 u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_0__721 (.o(net721));
 b15tilo00an1n03x5 u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_0__722 (.o(net722));
 b15tilo00an1n03x5 u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_14__u_filter_filter_q_reg_723 (.o(net723));
 b15tilo00an1n03x5 u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_14__u_filter_filter_q_reg_724 (.o(net724));
 b15tilo00an1n03x5 u_gpio_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__725 (.o(net725));
 b15tilo00an1n03x5 u_gpio_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__726 (.o(net726));
 b15tilo00an1n03x5 u_gpio_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__727 (.o(net727));
 b15tilo00an1n03x5 u_gpio_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__728 (.o(net728));
 b15tilo00an1n03x5 u_gpio_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_0__729 (.o(net729));
 b15tilo00an1n03x5 u_gpio_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_0__730 (.o(net730));
 b15tilo00an1n03x5 u_gpio_gen_filter_14__u_filter_stored_value_q_reg_731 (.o(net731));
 b15tilo00an1n03x5 u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_2__732 (.o(net732));
 b15tilo00an1n03x5 u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_2__733 (.o(net733));
 b15tilo00an1n03x5 u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_15__u_filter_filter_q_reg_734 (.o(net734));
 b15tilo00an1n03x5 u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_15__u_filter_filter_q_reg_735 (.o(net735));
 b15tilo00an1n03x5 u_gpio_gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_0__736 (.o(net736));
 b15tilo00an1n03x5 u_gpio_gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_0__737 (.o(net737));
 b15tilo00an1n03x5 u_gpio_gen_filter_15__u_filter_stored_value_q_reg_738 (.o(net738));
 b15tilo00an1n03x5 u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_1__739 (.o(net739));
 b15tilo00an1n03x5 u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_1__740 (.o(net740));
 b15tilo00an1n03x5 u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_3__741 (.o(net741));
 b15tilo00an1n03x5 u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_3__742 (.o(net742));
 b15tilo00an1n03x5 u_gpio_gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__743 (.o(net743));
 b15tilo00an1n03x5 u_gpio_gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__744 (.o(net744));
 b15tilo00an1n03x5 u_gpio_gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__745 (.o(net745));
 b15tilo00an1n03x5 u_gpio_gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__746 (.o(net746));
 b15tilo00an1n03x5 u_gpio_gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_0__747 (.o(net747));
 b15tilo00an1n03x5 u_gpio_gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_0__748 (.o(net748));
 b15tilo00an1n03x5 u_gpio_gen_filter_16__u_filter_stored_value_q_reg_749 (.o(net749));
 b15tilo00an1n03x5 u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_2__750 (.o(net750));
 b15tilo00an1n03x5 u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_2__751 (.o(net751));
 b15tilo00an1n03x5 u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_17__u_filter_filter_q_reg_752 (.o(net752));
 b15tilo00an1n03x5 u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_17__u_filter_filter_q_reg_753 (.o(net753));
 b15tilo00an1n03x5 u_gpio_gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_3__754 (.o(net754));
 b15tilo00an1n03x5 u_gpio_gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_3__755 (.o(net755));
 b15tilo00an1n03x5 u_gpio_gen_filter_17__u_filter_stored_value_q_reg_756 (.o(net756));
 b15tilo00an1n03x5 u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_1__757 (.o(net757));
 b15tilo00an1n03x5 u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_1__758 (.o(net758));
 b15tilo00an1n03x5 u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_3__759 (.o(net759));
 b15tilo00an1n03x5 u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_3__760 (.o(net760));
 b15tilo00an1n03x5 u_gpio_gen_filter_18__u_filter_filter_q_reg_u_gpio_gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__761 (.o(net761));
 b15tilo00an1n03x5 u_gpio_gen_filter_18__u_filter_filter_q_reg_u_gpio_gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__762 (.o(net762));
 b15tilo00an1n03x5 u_gpio_gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__763 (.o(net763));
 b15tilo00an1n03x5 u_gpio_gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__764 (.o(net764));
 b15tilo00an1n03x5 u_gpio_gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__765 (.o(net765));
 b15tilo00an1n03x5 u_gpio_gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__766 (.o(net766));
 b15tilo00an1n03x5 u_gpio_gen_filter_18__u_filter_stored_value_q_reg_767 (.o(net767));
 b15tilo00an1n03x5 u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_2__768 (.o(net768));
 b15tilo00an1n03x5 u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_2__769 (.o(net769));
 b15tilo00an1n03x5 u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_19__u_filter_filter_q_reg_770 (.o(net770));
 b15tilo00an1n03x5 u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_19__u_filter_filter_q_reg_771 (.o(net771));
 b15tilo00an1n03x5 u_gpio_gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_2__772 (.o(net772));
 b15tilo00an1n03x5 u_gpio_gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_2__773 (.o(net773));
 b15tilo00an1n03x5 u_gpio_gen_filter_19__u_filter_stored_value_q_reg_774 (.o(net774));
 b15tilo00an1n03x5 u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_1__775 (.o(net775));
 b15tilo00an1n03x5 u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_1__776 (.o(net776));
 b15tilo00an1n03x5 u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_3__777 (.o(net777));
 b15tilo00an1n03x5 u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_3__778 (.o(net778));
 b15tilo00an1n03x5 u_gpio_gen_filter_1__u_filter_filter_q_reg_u_gpio_gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__779 (.o(net779));
 b15tilo00an1n03x5 u_gpio_gen_filter_1__u_filter_filter_q_reg_u_gpio_gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__780 (.o(net780));
 b15tilo00an1n03x5 u_gpio_gen_filter_1__u_filter_stored_value_q_reg_781 (.o(net781));
 b15tilo00an1n03x5 u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_2__782 (.o(net782));
 b15tilo00an1n03x5 u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_2__783 (.o(net783));
 b15tilo00an1n03x5 u_gpio_gen_filter_20__u_filter_filter_q_reg_u_gpio_gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__784 (.o(net784));
 b15tilo00an1n03x5 u_gpio_gen_filter_20__u_filter_filter_q_reg_u_gpio_gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__785 (.o(net785));
 b15tilo00an1n03x5 u_gpio_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__786 (.o(net786));
 b15tilo00an1n03x5 u_gpio_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__787 (.o(net787));
 b15tilo00an1n03x5 u_gpio_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__788 (.o(net788));
 b15tilo00an1n03x5 u_gpio_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__789 (.o(net789));
 b15tilo00an1n03x5 u_gpio_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_0__790 (.o(net790));
 b15tilo00an1n03x5 u_gpio_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_0__791 (.o(net791));
 b15tilo00an1n03x5 u_gpio_gen_filter_20__u_filter_stored_value_q_reg_792 (.o(net792));
 b15tilo00an1n03x5 u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_1__793 (.o(net793));
 b15tilo00an1n03x5 u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_1__794 (.o(net794));
 b15tilo00an1n03x5 u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_3__795 (.o(net795));
 b15tilo00an1n03x5 u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_3__796 (.o(net796));
 b15tilo00an1n03x5 u_gpio_gen_filter_21__u_filter_filter_q_reg_u_gpio_gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__797 (.o(net797));
 b15tilo00an1n03x5 u_gpio_gen_filter_21__u_filter_filter_q_reg_u_gpio_gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__798 (.o(net798));
 b15tilo00an1n03x5 u_gpio_gen_filter_21__u_filter_stored_value_q_reg_799 (.o(net799));
 b15tilo00an1n03x5 u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_3__800 (.o(net800));
 b15tilo00an1n03x5 u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_3__801 (.o(net801));
 b15tilo00an1n03x5 u_gpio_gen_filter_22__u_filter_filter_q_reg_u_gpio_gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__802 (.o(net802));
 b15tilo00an1n03x5 u_gpio_gen_filter_22__u_filter_filter_q_reg_u_gpio_gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__803 (.o(net803));
 b15tilo00an1n03x5 u_gpio_gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__804 (.o(net804));
 b15tilo00an1n03x5 u_gpio_gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__805 (.o(net805));
 b15tilo00an1n03x5 u_gpio_gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__806 (.o(net806));
 b15tilo00an1n03x5 u_gpio_gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__807 (.o(net807));
 b15tilo00an1n03x5 u_gpio_gen_filter_22__u_filter_stored_value_q_reg_808 (.o(net808));
 b15tilo00an1n03x5 u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_2__809 (.o(net809));
 b15tilo00an1n03x5 u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_2__810 (.o(net810));
 b15tilo00an1n03x5 u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_23__u_filter_filter_q_reg_811 (.o(net811));
 b15tilo00an1n03x5 u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_23__u_filter_filter_q_reg_812 (.o(net812));
 b15tilo00an1n03x5 u_gpio_gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_0__813 (.o(net813));
 b15tilo00an1n03x5 u_gpio_gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_0__814 (.o(net814));
 b15tilo00an1n03x5 u_gpio_gen_filter_23__u_filter_stored_value_q_reg_815 (.o(net815));
 b15tilo00an1n03x5 u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_2__816 (.o(net816));
 b15tilo00an1n03x5 u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_2__817 (.o(net817));
 b15tilo00an1n03x5 u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_24__u_filter_filter_q_reg_818 (.o(net818));
 b15tilo00an1n03x5 u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_24__u_filter_filter_q_reg_819 (.o(net819));
 b15tilo00an1n03x5 u_gpio_gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__820 (.o(net820));
 b15tilo00an1n03x5 u_gpio_gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__821 (.o(net821));
 b15tilo00an1n03x5 u_gpio_gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__822 (.o(net822));
 b15tilo00an1n03x5 u_gpio_gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__823 (.o(net823));
 b15tilo00an1n03x5 u_gpio_gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_0__824 (.o(net824));
 b15tilo00an1n03x5 u_gpio_gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_0__825 (.o(net825));
 b15tilo00an1n03x5 u_gpio_gen_filter_24__u_filter_stored_value_q_reg_826 (.o(net826));
 b15tilo00an1n03x5 u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_2__827 (.o(net827));
 b15tilo00an1n03x5 u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_2__828 (.o(net828));
 b15tilo00an1n03x5 u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__829 (.o(net829));
 b15tilo00an1n03x5 u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__830 (.o(net830));
 b15tilo00an1n03x5 u_gpio_gen_filter_25__u_filter_filter_q_reg_u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_0__831 (.o(net831));
 b15tilo00an1n03x5 u_gpio_gen_filter_25__u_filter_filter_q_reg_u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_0__832 (.o(net832));
 b15tilo00an1n03x5 u_gpio_gen_filter_25__u_filter_stored_value_q_reg_833 (.o(net833));
 b15tilo00an1n03x5 u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_2__834 (.o(net834));
 b15tilo00an1n03x5 u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_2__835 (.o(net835));
 b15tilo00an1n03x5 u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_29__u_filter_filter_q_reg_836 (.o(net836));
 b15tilo00an1n03x5 u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_29__u_filter_filter_q_reg_837 (.o(net837));
 b15tilo00an1n03x5 u_gpio_gen_filter_26__u_filter_filter_q_reg_u_gpio_intr_hw_intr_o_reg_12__838 (.o(net838));
 b15tilo00an1n03x5 u_gpio_gen_filter_26__u_filter_filter_q_reg_u_gpio_intr_hw_intr_o_reg_12__839 (.o(net839));
 b15tilo00an1n03x5 u_gpio_gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__840 (.o(net840));
 b15tilo00an1n03x5 u_gpio_gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__841 (.o(net841));
 b15tilo00an1n03x5 u_gpio_gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__842 (.o(net842));
 b15tilo00an1n03x5 u_gpio_gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__843 (.o(net843));
 b15tilo00an1n03x5 u_gpio_gen_filter_26__u_filter_stored_value_q_reg_844 (.o(net844));
 b15tilo00an1n03x5 u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_2__845 (.o(net845));
 b15tilo00an1n03x5 u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_2__846 (.o(net846));
 b15tilo00an1n03x5 u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_27__u_filter_filter_q_reg_847 (.o(net847));
 b15tilo00an1n03x5 u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_27__u_filter_filter_q_reg_848 (.o(net848));
 b15tilo00an1n03x5 u_gpio_gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_intr_hw_intr_o_reg_24__849 (.o(net849));
 b15tilo00an1n03x5 u_gpio_gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_intr_hw_intr_o_reg_24__850 (.o(net850));
 b15tilo00an1n03x5 u_gpio_gen_filter_27__u_filter_stored_value_q_reg_851 (.o(net851));
 b15tilo00an1n03x5 u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_1__852 (.o(net852));
 b15tilo00an1n03x5 u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_1__853 (.o(net853));
 b15tilo00an1n03x5 u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_3__854 (.o(net854));
 b15tilo00an1n03x5 u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_3__855 (.o(net855));
 b15tilo00an1n03x5 u_gpio_gen_filter_28__u_filter_filter_q_reg_u_gpio_gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__856 (.o(net856));
 b15tilo00an1n03x5 u_gpio_gen_filter_28__u_filter_filter_q_reg_u_gpio_gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__857 (.o(net857));
 b15tilo00an1n03x5 u_gpio_gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__858 (.o(net858));
 b15tilo00an1n03x5 u_gpio_gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__859 (.o(net859));
 b15tilo00an1n03x5 u_gpio_gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__860 (.o(net860));
 b15tilo00an1n03x5 u_gpio_gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__861 (.o(net861));
 b15tilo00an1n03x5 u_gpio_gen_filter_28__u_filter_stored_value_q_reg_862 (.o(net862));
 b15tilo00an1n03x5 u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_1__863 (.o(net863));
 b15tilo00an1n03x5 u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_1__864 (.o(net864));
 b15tilo00an1n03x5 u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_3__865 (.o(net865));
 b15tilo00an1n03x5 u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_3__866 (.o(net866));
 b15tilo00an1n03x5 u_gpio_gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_0__867 (.o(net867));
 b15tilo00an1n03x5 u_gpio_gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_0__868 (.o(net868));
 b15tilo00an1n03x5 u_gpio_gen_filter_29__u_filter_stored_value_q_reg_869 (.o(net869));
 b15tilo00an1n03x5 u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_1__870 (.o(net870));
 b15tilo00an1n03x5 u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_1__871 (.o(net871));
 b15tilo00an1n03x5 u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_3__872 (.o(net872));
 b15tilo00an1n03x5 u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_3__873 (.o(net873));
 b15tilo00an1n03x5 u_gpio_gen_filter_2__u_filter_filter_q_reg_u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_1__874 (.o(net874));
 b15tilo00an1n03x5 u_gpio_gen_filter_2__u_filter_filter_q_reg_u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_1__875 (.o(net875));
 b15tilo00an1n03x5 u_gpio_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__876 (.o(net876));
 b15tilo00an1n03x5 u_gpio_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__877 (.o(net877));
 b15tilo00an1n03x5 u_gpio_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__878 (.o(net878));
 b15tilo00an1n03x5 u_gpio_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__879 (.o(net879));
 b15tilo00an1n03x5 u_gpio_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_0__880 (.o(net880));
 b15tilo00an1n03x5 u_gpio_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_0__881 (.o(net881));
 b15tilo00an1n03x5 u_gpio_gen_filter_2__u_filter_stored_value_q_reg_882 (.o(net882));
 b15tilo00an1n03x5 u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_30__u_filter_filter_q_reg_883 (.o(net883));
 b15tilo00an1n03x5 u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_30__u_filter_filter_q_reg_884 (.o(net884));
 b15tilo00an1n03x5 u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_3__885 (.o(net885));
 b15tilo00an1n03x5 u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_3__886 (.o(net886));
 b15tilo00an1n03x5 u_gpio_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__887 (.o(net887));
 b15tilo00an1n03x5 u_gpio_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__888 (.o(net888));
 b15tilo00an1n03x5 u_gpio_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__889 (.o(net889));
 b15tilo00an1n03x5 u_gpio_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__890 (.o(net890));
 b15tilo00an1n03x5 u_gpio_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__891 (.o(net891));
 b15tilo00an1n03x5 u_gpio_gen_filter_30__u_filter_stored_value_q_reg_892 (.o(net892));
 b15tilo00an1n03x5 u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_1__893 (.o(net893));
 b15tilo00an1n03x5 u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_1__894 (.o(net894));
 b15tilo00an1n03x5 u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_3__895 (.o(net895));
 b15tilo00an1n03x5 u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_3__896 (.o(net896));
 b15tilo00an1n03x5 u_gpio_gen_filter_31__u_filter_filter_q_reg_u_gpio_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__897 (.o(net897));
 b15tilo00an1n03x5 u_gpio_gen_filter_31__u_filter_filter_q_reg_u_gpio_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__898 (.o(net898));
 b15tilo00an1n03x5 u_gpio_gen_filter_31__u_filter_stored_value_q_reg_899 (.o(net899));
 b15tilo00an1n03x5 u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_2__900 (.o(net900));
 b15tilo00an1n03x5 u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_2__901 (.o(net901));
 b15tilo00an1n03x5 u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_3__u_filter_filter_q_reg_902 (.o(net902));
 b15tilo00an1n03x5 u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_3__u_filter_filter_q_reg_903 (.o(net903));
 b15tilo00an1n03x5 u_gpio_gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_7__u_filter_filter_q_reg_904 (.o(net904));
 b15tilo00an1n03x5 u_gpio_gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_7__u_filter_filter_q_reg_905 (.o(net905));
 b15tilo00an1n03x5 u_gpio_gen_filter_3__u_filter_stored_value_q_reg_906 (.o(net906));
 b15tilo00an1n03x5 u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_2__907 (.o(net907));
 b15tilo00an1n03x5 u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_2__908 (.o(net908));
 b15tilo00an1n03x5 u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_4__u_filter_filter_q_reg_909 (.o(net909));
 b15tilo00an1n03x5 u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_4__u_filter_filter_q_reg_910 (.o(net910));
 b15tilo00an1n03x5 u_gpio_gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__911 (.o(net911));
 b15tilo00an1n03x5 u_gpio_gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__912 (.o(net912));
 b15tilo00an1n03x5 u_gpio_gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__913 (.o(net913));
 b15tilo00an1n03x5 u_gpio_gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__914 (.o(net914));
 b15tilo00an1n03x5 u_gpio_gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_0__915 (.o(net915));
 b15tilo00an1n03x5 u_gpio_gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_0__916 (.o(net916));
 b15tilo00an1n03x5 u_gpio_gen_filter_4__u_filter_stored_value_q_reg_917 (.o(net917));
 b15tilo00an1n03x5 u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_2__918 (.o(net918));
 b15tilo00an1n03x5 u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_2__919 (.o(net919));
 b15tilo00an1n03x5 u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_5__u_filter_filter_q_reg_920 (.o(net920));
 b15tilo00an1n03x5 u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_5__u_filter_filter_q_reg_921 (.o(net921));
 b15tilo00an1n03x5 u_gpio_gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_0__922 (.o(net922));
 b15tilo00an1n03x5 u_gpio_gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_0__923 (.o(net923));
 b15tilo00an1n03x5 u_gpio_gen_filter_5__u_filter_stored_value_q_reg_924 (.o(net924));
 b15tilo00an1n03x5 u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_2__925 (.o(net925));
 b15tilo00an1n03x5 u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_2__926 (.o(net926));
 b15tilo00an1n03x5 u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_6__u_filter_filter_q_reg_927 (.o(net927));
 b15tilo00an1n03x5 u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_6__u_filter_filter_q_reg_928 (.o(net928));
 b15tilo00an1n03x5 u_gpio_gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__929 (.o(net929));
 b15tilo00an1n03x5 u_gpio_gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__930 (.o(net930));
 b15tilo00an1n03x5 u_gpio_gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__931 (.o(net931));
 b15tilo00an1n03x5 u_gpio_gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__932 (.o(net932));
 b15tilo00an1n03x5 u_gpio_gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_0__933 (.o(net933));
 b15tilo00an1n03x5 u_gpio_gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_0__934 (.o(net934));
 b15tilo00an1n03x5 u_gpio_gen_filter_6__u_filter_stored_value_q_reg_935 (.o(net935));
 b15tilo00an1n03x5 u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_2__936 (.o(net936));
 b15tilo00an1n03x5 u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_2__937 (.o(net937));
 b15tilo00an1n03x5 u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_0__938 (.o(net938));
 b15tilo00an1n03x5 u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_0__939 (.o(net939));
 b15tilo00an1n03x5 u_gpio_gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__940 (.o(net940));
 b15tilo00an1n03x5 u_gpio_gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__941 (.o(net941));
 b15tilo00an1n03x5 u_gpio_gen_filter_7__u_filter_stored_value_q_reg_942 (.o(net942));
 b15tilo00an1n03x5 u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_2__943 (.o(net943));
 b15tilo00an1n03x5 u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_2__944 (.o(net944));
 b15tilo00an1n03x5 u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_0__945 (.o(net945));
 b15tilo00an1n03x5 u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_0__946 (.o(net946));
 b15tilo00an1n03x5 u_gpio_gen_filter_8__u_filter_filter_q_reg_u_gpio_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__947 (.o(net947));
 b15tilo00an1n03x5 u_gpio_gen_filter_8__u_filter_filter_q_reg_u_gpio_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__948 (.o(net948));
 b15tilo00an1n03x5 u_gpio_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__949 (.o(net949));
 b15tilo00an1n03x5 u_gpio_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__950 (.o(net950));
 b15tilo00an1n03x5 u_gpio_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__951 (.o(net951));
 b15tilo00an1n03x5 u_gpio_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__952 (.o(net952));
 b15tilo00an1n03x5 u_gpio_gen_filter_8__u_filter_stored_value_q_reg_953 (.o(net953));
 b15tilo00an1n03x5 u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_2__954 (.o(net954));
 b15tilo00an1n03x5 u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_2__955 (.o(net955));
 b15tilo00an1n03x5 u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_9__u_filter_filter_q_reg_956 (.o(net956));
 b15tilo00an1n03x5 u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_9__u_filter_filter_q_reg_957 (.o(net957));
 b15tilo00an1n03x5 u_gpio_gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_2__958 (.o(net958));
 b15tilo00an1n03x5 u_gpio_gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_2__959 (.o(net959));
 b15tilo00an1n03x5 u_gpio_gen_filter_9__u_filter_stored_value_q_reg_960 (.o(net960));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_0__u_gpio_intr_hw_intr_o_reg_1__961 (.o(net961));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_0__u_gpio_intr_hw_intr_o_reg_1__962 (.o(net962));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_10__u_gpio_intr_hw_intr_o_reg_11__963 (.o(net963));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_10__u_gpio_intr_hw_intr_o_reg_11__964 (.o(net964));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_13__u_gpio_intr_hw_intr_o_reg_14__965 (.o(net965));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_13__u_gpio_intr_hw_intr_o_reg_14__966 (.o(net966));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_15__u_gpio_intr_hw_intr_o_reg_16__967 (.o(net967));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_15__u_gpio_intr_hw_intr_o_reg_16__968 (.o(net968));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_17__u_gpio_intr_hw_intr_o_reg_18__969 (.o(net969));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_17__u_gpio_intr_hw_intr_o_reg_18__970 (.o(net970));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_19__u_gpio_intr_hw_intr_o_reg_20__971 (.o(net971));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_19__u_gpio_intr_hw_intr_o_reg_20__972 (.o(net972));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_21__u_gpio_intr_hw_intr_o_reg_29__973 (.o(net973));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_21__u_gpio_intr_hw_intr_o_reg_29__974 (.o(net974));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_22__u_gpio_intr_hw_intr_o_reg_23__975 (.o(net975));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_22__u_gpio_intr_hw_intr_o_reg_23__976 (.o(net976));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_25__u_gpio_intr_hw_intr_o_reg_26__977 (.o(net977));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_25__u_gpio_intr_hw_intr_o_reg_26__978 (.o(net978));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_27__u_gpio_u_reg_err_q_reg_979 (.o(net979));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_27__u_gpio_u_reg_err_q_reg_980 (.o(net980));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_28__u_gpio_u_reg_u_data_in_q_reg_2__981 (.o(net981));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_28__u_gpio_u_reg_u_data_in_q_reg_2__982 (.o(net982));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_2__u_gpio_intr_hw_intr_o_reg_3__983 (.o(net983));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_2__u_gpio_intr_hw_intr_o_reg_3__984 (.o(net984));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_30__u_gpio_intr_hw_intr_o_reg_31__985 (.o(net985));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_30__u_gpio_intr_hw_intr_o_reg_31__986 (.o(net986));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_4__u_gpio_intr_hw_intr_o_reg_5__987 (.o(net987));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_4__u_gpio_intr_hw_intr_o_reg_5__988 (.o(net988));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_6__u_gpio_intr_hw_intr_o_reg_7__989 (.o(net989));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_6__u_gpio_intr_hw_intr_o_reg_7__990 (.o(net990));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_8__u_gpio_intr_hw_intr_o_reg_9__991 (.o(net991));
 b15tilo00an1n03x5 u_gpio_intr_hw_intr_o_reg_8__u_gpio_intr_hw_intr_o_reg_9__992 (.o(net992));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_clk_gate_q_reg_0_latch_993 (.o(net993));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_clk_gate_q_reg_latch_994 (.o(net994));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_0__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_1__995 (.o(net995));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_0__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_1__996 (.o(net996));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_10__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_11__997 (.o(net997));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_10__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_11__998 (.o(net998));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_12__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_13__999 (.o(net999));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_12__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_13__1000 (.o(net1000));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_14__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_15__1001 (.o(net1001));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_14__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_15__1002 (.o(net1002));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_16__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_17__1003 (.o(net1003));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_16__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_17__1004 (.o(net1004));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_18__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_19__1005 (.o(net1005));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_18__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_19__1006 (.o(net1006));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_20__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_21__1007 (.o(net1007));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_20__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_21__1008 (.o(net1008));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_22__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_23__1009 (.o(net1009));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_22__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_23__1010 (.o(net1010));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_24__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_25__1011 (.o(net1011));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_24__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_25__1012 (.o(net1012));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_26__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_27__1013 (.o(net1013));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_26__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_27__1014 (.o(net1014));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_28__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_29__1015 (.o(net1015));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_28__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_29__1016 (.o(net1016));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_2__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_3__1017 (.o(net1017));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_2__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_3__1018 (.o(net1018));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_30__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_31__1019 (.o(net1019));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_30__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_31__1020 (.o(net1020));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_4__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_5__1021 (.o(net1021));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_4__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_5__1022 (.o(net1022));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_6__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_7__1023 (.o(net1023));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_6__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_7__1024 (.o(net1024));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_8__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_9__1025 (.o(net1025));
 b15tilo00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_8__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_9__1026 (.o(net1026));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_0__u_gpio_u_reg_u_data_in_q_reg_1__1027 (.o(net1027));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_0__u_gpio_u_reg_u_data_in_q_reg_1__1028 (.o(net1028));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_13__1029 (.o(net1029));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_14__u_gpio_u_reg_u_data_in_q_reg_23__1030 (.o(net1030));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_14__u_gpio_u_reg_u_data_in_q_reg_23__1031 (.o(net1031));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_15__u_gpio_u_reg_u_data_in_q_reg_16__1032 (.o(net1032));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_15__u_gpio_u_reg_u_data_in_q_reg_16__1033 (.o(net1033));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_17__u_gpio_u_reg_u_data_in_q_reg_18__1034 (.o(net1034));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_17__u_gpio_u_reg_u_data_in_q_reg_18__1035 (.o(net1035));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_19__u_gpio_u_reg_u_data_in_q_reg_20__1036 (.o(net1036));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_19__u_gpio_u_reg_u_data_in_q_reg_20__1037 (.o(net1037));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_21__u_gpio_u_reg_u_data_in_q_reg_22__1038 (.o(net1038));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_21__u_gpio_u_reg_u_data_in_q_reg_22__1039 (.o(net1039));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_24__u_gpio_u_reg_u_data_in_q_reg_25__1040 (.o(net1040));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_24__u_gpio_u_reg_u_data_in_q_reg_25__1041 (.o(net1041));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_26__u_gpio_u_reg_u_data_in_q_reg_28__1042 (.o(net1042));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_26__u_gpio_u_reg_u_data_in_q_reg_28__1043 (.o(net1043));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_27__u_gpio_u_reg_u_data_in_q_reg_30__1044 (.o(net1044));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_27__u_gpio_u_reg_u_data_in_q_reg_30__1045 (.o(net1045));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_29__1046 (.o(net1046));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_31__1047 (.o(net1047));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_3__u_gpio_u_reg_u_data_in_q_reg_4__1048 (.o(net1048));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_3__u_gpio_u_reg_u_data_in_q_reg_4__1049 (.o(net1049));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_5__u_gpio_u_reg_u_data_in_q_reg_12__1050 (.o(net1050));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_5__u_gpio_u_reg_u_data_in_q_reg_12__1051 (.o(net1051));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_6__u_gpio_u_reg_u_data_in_q_reg_7__1052 (.o(net1052));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_6__u_gpio_u_reg_u_data_in_q_reg_7__1053 (.o(net1053));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_8__u_gpio_u_reg_u_data_in_q_reg_11__1054 (.o(net1054));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_8__u_gpio_u_reg_u_data_in_q_reg_11__1055 (.o(net1055));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_9__u_gpio_u_reg_u_data_in_q_reg_10__1056 (.o(net1056));
 b15tilo00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_9__u_gpio_u_reg_u_data_in_q_reg_10__1057 (.o(net1057));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_clk_gate_q_reg_0_latch_1058 (.o(net1058));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_clk_gate_q_reg_latch_1059 (.o(net1059));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_1__1060 (.o(net1060));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_1__1061 (.o(net1061));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_11__1062 (.o(net1062));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_11__1063 (.o(net1063));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_13__1064 (.o(net1064));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_13__1065 (.o(net1065));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_15__1066 (.o(net1066));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_15__1067 (.o(net1067));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_17__1068 (.o(net1068));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_17__1069 (.o(net1069));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_19__1070 (.o(net1070));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_19__1071 (.o(net1071));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_21__1072 (.o(net1072));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_21__1073 (.o(net1073));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_23__1074 (.o(net1074));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_23__1075 (.o(net1075));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_25__1076 (.o(net1076));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_25__1077 (.o(net1077));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_27__1078 (.o(net1078));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_27__1079 (.o(net1079));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_29__1080 (.o(net1080));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_29__1081 (.o(net1081));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_3__1082 (.o(net1082));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_3__1083 (.o(net1083));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_31__1084 (.o(net1084));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_31__1085 (.o(net1085));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_5__1086 (.o(net1086));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_5__1087 (.o(net1087));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_7__1088 (.o(net1088));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_7__1089 (.o(net1089));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_9__1090 (.o(net1090));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_9__1091 (.o(net1091));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_clk_gate_q_reg_0_latch_1092 (.o(net1092));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_clk_gate_q_reg_latch_1093 (.o(net1093));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_1__1094 (.o(net1094));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_1__1095 (.o(net1095));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_11__1096 (.o(net1096));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_11__1097 (.o(net1097));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_13__1098 (.o(net1098));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_13__1099 (.o(net1099));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_15__1100 (.o(net1100));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_15__1101 (.o(net1101));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_17__1102 (.o(net1102));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_17__1103 (.o(net1103));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_19__1104 (.o(net1104));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_19__1105 (.o(net1105));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_21__1106 (.o(net1106));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_21__1107 (.o(net1107));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_23__1108 (.o(net1108));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_23__1109 (.o(net1109));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_25__1110 (.o(net1110));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_25__1111 (.o(net1111));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_27__1112 (.o(net1112));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_27__1113 (.o(net1113));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_29__1114 (.o(net1114));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_29__1115 (.o(net1115));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_3__1116 (.o(net1116));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_3__1117 (.o(net1117));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_31__1118 (.o(net1118));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_31__1119 (.o(net1119));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_5__1120 (.o(net1120));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_5__1121 (.o(net1121));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_7__1122 (.o(net1122));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_7__1123 (.o(net1123));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_9__1124 (.o(net1124));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_9__1125 (.o(net1125));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_clk_gate_q_reg_0_latch_1126 (.o(net1126));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_clk_gate_q_reg_latch_1127 (.o(net1127));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_1__1128 (.o(net1128));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_1__1129 (.o(net1129));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_11__1130 (.o(net1130));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_11__1131 (.o(net1131));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_13__1132 (.o(net1132));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_13__1133 (.o(net1133));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_15__1134 (.o(net1134));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_15__1135 (.o(net1135));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_17__1136 (.o(net1136));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_17__1137 (.o(net1137));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_19__1138 (.o(net1138));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_19__1139 (.o(net1139));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_21__1140 (.o(net1140));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_21__1141 (.o(net1141));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_23__1142 (.o(net1142));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_23__1143 (.o(net1143));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_25__1144 (.o(net1144));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_25__1145 (.o(net1145));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_27__1146 (.o(net1146));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_27__1147 (.o(net1147));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_29__1148 (.o(net1148));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_29__1149 (.o(net1149));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_3__1150 (.o(net1150));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_3__1151 (.o(net1151));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_31__1152 (.o(net1152));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_31__1153 (.o(net1153));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_5__1154 (.o(net1154));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_5__1155 (.o(net1155));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_7__1156 (.o(net1156));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_7__1157 (.o(net1157));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_9__1158 (.o(net1158));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_9__1159 (.o(net1159));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_clk_gate_q_reg_0_latch_1160 (.o(net1160));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_clk_gate_q_reg_latch_1161 (.o(net1161));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_1__1162 (.o(net1162));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_1__1163 (.o(net1163));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_11__1164 (.o(net1164));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_11__1165 (.o(net1165));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_13__1166 (.o(net1166));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_13__1167 (.o(net1167));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_15__1168 (.o(net1168));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_15__1169 (.o(net1169));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_17__1170 (.o(net1170));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_17__1171 (.o(net1171));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_19__1172 (.o(net1172));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_19__1173 (.o(net1173));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_21__1174 (.o(net1174));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_21__1175 (.o(net1175));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_23__1176 (.o(net1176));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_23__1177 (.o(net1177));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_25__1178 (.o(net1178));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_25__1179 (.o(net1179));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_27__1180 (.o(net1180));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_27__1181 (.o(net1181));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_29__1182 (.o(net1182));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_29__1183 (.o(net1183));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_3__1184 (.o(net1184));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_3__1185 (.o(net1185));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_31__1186 (.o(net1186));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_31__1187 (.o(net1187));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_5__1188 (.o(net1188));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_5__1189 (.o(net1189));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_7__1190 (.o(net1190));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_7__1191 (.o(net1191));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_9__1192 (.o(net1192));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_9__1193 (.o(net1193));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_clk_gate_q_reg_0_latch_1194 (.o(net1194));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_clk_gate_q_reg_latch_1195 (.o(net1195));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_0__u_gpio_u_reg_u_intr_enable_q_reg_1__1196 (.o(net1196));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_0__u_gpio_u_reg_u_intr_enable_q_reg_1__1197 (.o(net1197));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_10__u_gpio_u_reg_u_intr_enable_q_reg_11__1198 (.o(net1198));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_10__u_gpio_u_reg_u_intr_enable_q_reg_11__1199 (.o(net1199));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_12__u_gpio_u_reg_u_intr_enable_q_reg_13__1200 (.o(net1200));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_12__u_gpio_u_reg_u_intr_enable_q_reg_13__1201 (.o(net1201));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_14__u_gpio_u_reg_u_intr_enable_q_reg_15__1202 (.o(net1202));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_14__u_gpio_u_reg_u_intr_enable_q_reg_15__1203 (.o(net1203));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_16__u_gpio_u_reg_u_intr_enable_q_reg_17__1204 (.o(net1204));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_16__u_gpio_u_reg_u_intr_enable_q_reg_17__1205 (.o(net1205));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_18__u_gpio_u_reg_u_intr_enable_q_reg_19__1206 (.o(net1206));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_18__u_gpio_u_reg_u_intr_enable_q_reg_19__1207 (.o(net1207));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_20__u_gpio_u_reg_u_intr_enable_q_reg_21__1208 (.o(net1208));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_20__u_gpio_u_reg_u_intr_enable_q_reg_21__1209 (.o(net1209));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_22__u_gpio_u_reg_u_intr_enable_q_reg_23__1210 (.o(net1210));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_22__u_gpio_u_reg_u_intr_enable_q_reg_23__1211 (.o(net1211));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_24__u_gpio_u_reg_u_intr_enable_q_reg_25__1212 (.o(net1212));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_24__u_gpio_u_reg_u_intr_enable_q_reg_25__1213 (.o(net1213));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_26__u_gpio_u_reg_u_intr_enable_q_reg_27__1214 (.o(net1214));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_26__u_gpio_u_reg_u_intr_enable_q_reg_27__1215 (.o(net1215));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_28__u_gpio_u_reg_u_intr_enable_q_reg_29__1216 (.o(net1216));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_28__u_gpio_u_reg_u_intr_enable_q_reg_29__1217 (.o(net1217));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_2__u_gpio_u_reg_u_intr_enable_q_reg_3__1218 (.o(net1218));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_2__u_gpio_u_reg_u_intr_enable_q_reg_3__1219 (.o(net1219));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_30__u_gpio_u_reg_u_intr_enable_q_reg_31__1220 (.o(net1220));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_30__u_gpio_u_reg_u_intr_enable_q_reg_31__1221 (.o(net1221));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_4__u_gpio_u_reg_u_intr_enable_q_reg_5__1222 (.o(net1222));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_4__u_gpio_u_reg_u_intr_enable_q_reg_5__1223 (.o(net1223));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_6__u_gpio_u_reg_u_intr_enable_q_reg_7__1224 (.o(net1224));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_6__u_gpio_u_reg_u_intr_enable_q_reg_7__1225 (.o(net1225));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_8__u_gpio_u_reg_u_intr_enable_q_reg_9__1226 (.o(net1226));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_8__u_gpio_u_reg_u_intr_enable_q_reg_9__1227 (.o(net1227));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_clk_gate_q_reg_0_latch_1228 (.o(net1228));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_clk_gate_q_reg_latch_1229 (.o(net1229));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_0__u_gpio_u_reg_u_intr_state_q_reg_1__1230 (.o(net1230));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_0__u_gpio_u_reg_u_intr_state_q_reg_1__1231 (.o(net1231));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_10__u_gpio_u_reg_u_intr_state_q_reg_11__1232 (.o(net1232));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_10__u_gpio_u_reg_u_intr_state_q_reg_11__1233 (.o(net1233));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_12__u_gpio_u_reg_u_intr_state_q_reg_13__1234 (.o(net1234));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_12__u_gpio_u_reg_u_intr_state_q_reg_13__1235 (.o(net1235));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_14__u_gpio_u_reg_u_intr_state_q_reg_15__1236 (.o(net1236));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_14__u_gpio_u_reg_u_intr_state_q_reg_15__1237 (.o(net1237));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_16__u_gpio_u_reg_u_intr_state_q_reg_17__1238 (.o(net1238));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_16__u_gpio_u_reg_u_intr_state_q_reg_17__1239 (.o(net1239));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_18__u_gpio_u_reg_u_intr_state_q_reg_19__1240 (.o(net1240));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_18__u_gpio_u_reg_u_intr_state_q_reg_19__1241 (.o(net1241));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_20__u_gpio_u_reg_u_intr_state_q_reg_21__1242 (.o(net1242));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_20__u_gpio_u_reg_u_intr_state_q_reg_21__1243 (.o(net1243));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_22__u_gpio_u_reg_u_intr_state_q_reg_23__1244 (.o(net1244));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_22__u_gpio_u_reg_u_intr_state_q_reg_23__1245 (.o(net1245));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_24__u_gpio_u_reg_u_intr_state_q_reg_25__1246 (.o(net1246));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_24__u_gpio_u_reg_u_intr_state_q_reg_25__1247 (.o(net1247));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_26__u_gpio_u_reg_u_intr_state_q_reg_27__1248 (.o(net1248));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_26__u_gpio_u_reg_u_intr_state_q_reg_27__1249 (.o(net1249));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_28__u_gpio_u_reg_u_intr_state_q_reg_29__1250 (.o(net1250));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_28__u_gpio_u_reg_u_intr_state_q_reg_29__1251 (.o(net1251));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_2__u_gpio_u_reg_u_intr_state_q_reg_3__1252 (.o(net1252));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_2__u_gpio_u_reg_u_intr_state_q_reg_3__1253 (.o(net1253));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_30__u_gpio_u_reg_u_intr_state_q_reg_31__1254 (.o(net1254));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_30__u_gpio_u_reg_u_intr_state_q_reg_31__1255 (.o(net1255));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_4__u_gpio_u_reg_u_intr_state_q_reg_5__1256 (.o(net1256));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_4__u_gpio_u_reg_u_intr_state_q_reg_5__1257 (.o(net1257));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_6__u_gpio_u_reg_u_intr_state_q_reg_7__1258 (.o(net1258));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_6__u_gpio_u_reg_u_intr_state_q_reg_7__1259 (.o(net1259));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_8__u_gpio_u_reg_u_intr_state_q_reg_9__1260 (.o(net1260));
 b15tilo00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_8__u_gpio_u_reg_u_intr_state_q_reg_9__1261 (.o(net1261));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_clk_gate_rdata_reg_0_latch_1262 (.o(net1262));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_clk_gate_rdata_reg_latch_1263 (.o(net1263));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_clk_gate_reqid_reg_latch_1264 (.o(net1264));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_error_reg_1265 (.o(net1265));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_outstanding_reg_1266 (.o(net1266));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_0__u_gpio_u_reg_u_reg_if_rdata_reg_1__1267 (.o(net1267));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_0__u_gpio_u_reg_u_reg_if_rdata_reg_1__1268 (.o(net1268));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_10__u_gpio_u_reg_u_reg_if_rdata_reg_11__1269 (.o(net1269));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_10__u_gpio_u_reg_u_reg_if_rdata_reg_11__1270 (.o(net1270));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_12__u_gpio_u_reg_u_reg_if_rdata_reg_13__1271 (.o(net1271));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_12__u_gpio_u_reg_u_reg_if_rdata_reg_13__1272 (.o(net1272));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_14__u_gpio_u_reg_u_reg_if_rdata_reg_15__1273 (.o(net1273));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_14__u_gpio_u_reg_u_reg_if_rdata_reg_15__1274 (.o(net1274));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_16__u_gpio_u_reg_u_reg_if_rdata_reg_17__1275 (.o(net1275));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_16__u_gpio_u_reg_u_reg_if_rdata_reg_17__1276 (.o(net1276));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_18__u_gpio_u_reg_u_reg_if_rdata_reg_19__1277 (.o(net1277));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_18__u_gpio_u_reg_u_reg_if_rdata_reg_19__1278 (.o(net1278));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_20__u_gpio_u_reg_u_reg_if_rdata_reg_21__1279 (.o(net1279));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_20__u_gpio_u_reg_u_reg_if_rdata_reg_21__1280 (.o(net1280));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_22__u_gpio_u_reg_u_reg_if_rdata_reg_23__1281 (.o(net1281));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_22__u_gpio_u_reg_u_reg_if_rdata_reg_23__1282 (.o(net1282));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_24__u_gpio_u_reg_u_reg_if_rdata_reg_25__1283 (.o(net1283));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_24__u_gpio_u_reg_u_reg_if_rdata_reg_25__1284 (.o(net1284));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_26__u_gpio_u_reg_u_reg_if_rdata_reg_27__1285 (.o(net1285));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_26__u_gpio_u_reg_u_reg_if_rdata_reg_27__1286 (.o(net1286));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_28__u_gpio_u_reg_u_reg_if_rdata_reg_29__1287 (.o(net1287));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_28__u_gpio_u_reg_u_reg_if_rdata_reg_29__1288 (.o(net1288));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_2__u_gpio_u_reg_u_reg_if_rdata_reg_3__1289 (.o(net1289));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_2__u_gpio_u_reg_u_reg_if_rdata_reg_3__1290 (.o(net1290));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_30__u_gpio_u_reg_u_reg_if_rdata_reg_31__1291 (.o(net1291));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_30__u_gpio_u_reg_u_reg_if_rdata_reg_31__1292 (.o(net1292));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_4__u_gpio_u_reg_u_reg_if_rdata_reg_5__1293 (.o(net1293));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_4__u_gpio_u_reg_u_reg_if_rdata_reg_5__1294 (.o(net1294));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_6__u_gpio_u_reg_u_reg_if_rdata_reg_7__1295 (.o(net1295));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_6__u_gpio_u_reg_u_reg_if_rdata_reg_7__1296 (.o(net1296));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_8__u_gpio_u_reg_u_reg_if_rdata_reg_9__1297 (.o(net1297));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_8__u_gpio_u_reg_u_reg_if_rdata_reg_9__1298 (.o(net1298));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_reqid_reg_0__u_gpio_u_reg_u_reg_if_reqid_reg_1__1299 (.o(net1299));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_reqid_reg_0__u_gpio_u_reg_u_reg_if_reqid_reg_1__1300 (.o(net1300));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_reqid_reg_2__u_gpio_u_reg_u_reg_if_reqid_reg_3__1301 (.o(net1301));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_reqid_reg_2__u_gpio_u_reg_u_reg_if_reqid_reg_3__1302 (.o(net1302));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_reqid_reg_4__u_gpio_u_reg_u_reg_if_reqid_reg_5__1303 (.o(net1303));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_reqid_reg_4__u_gpio_u_reg_u_reg_if_reqid_reg_5__1304 (.o(net1304));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_reqid_reg_6__u_gpio_u_reg_u_reg_if_reqid_reg_7__1305 (.o(net1305));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_reqid_reg_6__u_gpio_u_reg_u_reg_if_reqid_reg_7__1306 (.o(net1306));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_reqsz_reg_0__1307 (.o(net1307));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_reqsz_reg_1__1308 (.o(net1308));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rspop_reg_0__1309 (.o(net1309));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rspop_reg_1__u_gpio_u_reg_u_reg_if_rspop_reg_2__1310 (.o(net1310));
 b15tilo00an1n03x5 u_gpio_u_reg_u_reg_if_rspop_reg_1__u_gpio_u_reg_u_reg_if_rspop_reg_2__1311 (.o(net1311));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_clk_gate_num_req_outstanding_reg_latch_1312 (.o(net1312));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_dev_select_outstanding_reg_0__1313 (.o(net1313));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_dev_select_outstanding_reg_1__1314 (.o(net1314));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_dev_select_outstanding_reg_2__1315 (.o(net1315));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_clk_gate_err_source_reg_latch_1316 (.o(net1316));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type_reg_0__1317 (.o(net1317));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type_reg_1__1318 (.o(net1318));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type_reg_2__1319 (.o(net1319));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type_reg_3__1320 (.o(net1320));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_opcode_reg_0__1321 (.o(net1321));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_opcode_reg_1__1322 (.o(net1322));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_opcode_reg_2__1323 (.o(net1323));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_req_pending_reg_1324 (.o(net1324));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_rsp_pending_reg_1325 (.o(net1325));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_size_reg_0__1326 (.o(net1326));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_size_reg_1__1327 (.o(net1327));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_0__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_1__1328 (.o(net1328));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_0__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_1__1329 (.o(net1329));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_2__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_3__1330 (.o(net1330));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_2__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_3__1331 (.o(net1331));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_4__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_5__1332 (.o(net1332));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_4__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_5__1333 (.o(net1333));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_6__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_7__1334 (.o(net1334));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_6__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_7__1335 (.o(net1335));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_0__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_1__1336 (.o(net1336));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_0__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_1__1337 (.o(net1337));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_2__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_3__1338 (.o(net1338));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_2__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_3__1339 (.o(net1339));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_4__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_5__1340 (.o(net1340));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_4__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_5__1341 (.o(net1341));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_6__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_7__1342 (.o(net1342));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_6__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_7__1343 (.o(net1343));
 b15tilo00an1n03x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_8__1344 (.o(net1344));
 b15tihi00an1n03x5 U3305_1346 (.o(net1346));
 b15tihi00an1n03x5 U3307_1347 (.o(net1347));
 b15tihi00an1n03x5 U3309_1348 (.o(net1348));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_0__u_gpio_cio_gpio_en_q_reg_1__1349 (.o(net1349));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_10__u_gpio_cio_gpio_en_q_reg_11__1350 (.o(net1350));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_12__u_gpio_cio_gpio_en_q_reg_13__1351 (.o(net1351));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_14__u_gpio_cio_gpio_en_q_reg_15__1352 (.o(net1352));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_16__u_gpio_cio_gpio_en_q_reg_17__1353 (.o(net1353));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_18__u_gpio_cio_gpio_en_q_reg_19__1354 (.o(net1354));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_20__u_gpio_cio_gpio_en_q_reg_21__1355 (.o(net1355));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_22__u_gpio_cio_gpio_en_q_reg_23__1356 (.o(net1356));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_24__u_gpio_cio_gpio_en_q_reg_25__1357 (.o(net1357));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_26__u_gpio_cio_gpio_en_q_reg_27__1358 (.o(net1358));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_28__u_gpio_cio_gpio_en_q_reg_29__1359 (.o(net1359));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_2__u_gpio_cio_gpio_en_q_reg_3__1360 (.o(net1360));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_30__u_gpio_cio_gpio_en_q_reg_31__1361 (.o(net1361));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_4__u_gpio_cio_gpio_en_q_reg_5__1362 (.o(net1362));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_6__u_gpio_cio_gpio_en_q_reg_7__1363 (.o(net1363));
 b15tihi00an1n03x5 u_gpio_cio_gpio_en_q_reg_8__u_gpio_cio_gpio_en_q_reg_9__1364 (.o(net1364));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_0__u_gpio_cio_gpio_q_reg_1__1365 (.o(net1365));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_10__u_gpio_cio_gpio_q_reg_11__1366 (.o(net1366));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_12__u_gpio_cio_gpio_q_reg_13__1367 (.o(net1367));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_14__u_gpio_cio_gpio_q_reg_15__1368 (.o(net1368));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_16__u_gpio_cio_gpio_q_reg_17__1369 (.o(net1369));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_18__u_gpio_cio_gpio_q_reg_19__1370 (.o(net1370));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_20__u_gpio_cio_gpio_q_reg_21__1371 (.o(net1371));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_22__u_gpio_cio_gpio_q_reg_23__1372 (.o(net1372));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_24__u_gpio_cio_gpio_q_reg_25__1373 (.o(net1373));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_26__u_gpio_cio_gpio_q_reg_27__1374 (.o(net1374));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_28__u_gpio_cio_gpio_q_reg_29__1375 (.o(net1375));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_2__u_gpio_cio_gpio_q_reg_3__1376 (.o(net1376));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_30__u_gpio_cio_gpio_q_reg_31__1377 (.o(net1377));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_4__u_gpio_cio_gpio_q_reg_5__1378 (.o(net1378));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_6__u_gpio_cio_gpio_q_reg_7__1379 (.o(net1379));
 b15tihi00an1n03x5 u_gpio_cio_gpio_q_reg_8__u_gpio_cio_gpio_q_reg_9__1380 (.o(net1380));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_0__u_gpio_data_in_q_reg_1__1381 (.o(net1381));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_10__u_gpio_data_in_q_reg_11__1382 (.o(net1382));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_12__u_gpio_data_in_q_reg_13__1383 (.o(net1383));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_14__u_gpio_data_in_q_reg_15__1384 (.o(net1384));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_16__u_gpio_data_in_q_reg_17__1385 (.o(net1385));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_18__u_gpio_data_in_q_reg_19__1386 (.o(net1386));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_20__u_gpio_data_in_q_reg_21__1387 (.o(net1387));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_22__u_gpio_data_in_q_reg_23__1388 (.o(net1388));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_24__u_gpio_data_in_q_reg_25__1389 (.o(net1389));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_26__u_gpio_data_in_q_reg_27__1390 (.o(net1390));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_28__u_gpio_data_in_q_reg_29__1391 (.o(net1391));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_2__u_gpio_data_in_q_reg_3__1392 (.o(net1392));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_30__u_gpio_data_in_q_reg_31__1393 (.o(net1393));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_4__u_gpio_data_in_q_reg_5__1394 (.o(net1394));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_6__u_gpio_data_in_q_reg_7__1395 (.o(net1395));
 b15tihi00an1n03x5 u_gpio_data_in_q_reg_8__u_gpio_data_in_q_reg_9__1396 (.o(net1396));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_set_q_reg_u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_0__1397 (.o(net1397));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q_reg_u_gpio_gen_alert_tx_0__u_prim_alert_sender_ping_set_q_reg_1398 (.o(net1398));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_0__u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_1__1399 (.o(net1399));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_2__u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq_reg_1400 (.o(net1400));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq_reg_1401 (.o(net1401));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1402 (.o(net1402));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1403 (.o(net1403));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1404 (.o(net1404));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1405 (.o(net1405));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q_reg_1406 (.o(net1406));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_0__1407 (.o(net1407));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_1__1408 (.o(net1408));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq_reg_1409 (.o(net1409));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq_reg_u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1410 (.o(net1410));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1411 (.o(net1411));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1412 (.o(net1412));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1413 (.o(net1413));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_0__1414 (.o(net1414));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_1__1415 (.o(net1415));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q_reg_u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_0__1416 (.o(net1416));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_16__u_filter_filter_q_reg_1417 (.o(net1417));
 b15tihi00an1n03x5 u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_1__1418 (.o(net1418));
 b15tihi00an1n03x5 u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_1__1419 (.o(net1419));
 b15tihi00an1n03x5 u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_0__u_filter_diff_ctr_q_reg_3__1420 (.o(net1420));
 b15tihi00an1n03x5 u_gpio_gen_filter_0__u_filter_filter_q_reg_u_gpio_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1421 (.o(net1421));
 b15tihi00an1n03x5 u_gpio_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1422 (.o(net1422));
 b15tihi00an1n03x5 u_gpio_gen_filter_0__u_filter_stored_value_q_reg_1423 (.o(net1423));
 b15tihi00an1n03x5 u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_1__1424 (.o(net1424));
 b15tihi00an1n03x5 u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_10__u_filter_filter_q_reg_1425 (.o(net1425));
 b15tihi00an1n03x5 u_gpio_gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1426 (.o(net1426));
 b15tihi00an1n03x5 u_gpio_gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_0__1427 (.o(net1427));
 b15tihi00an1n03x5 u_gpio_gen_filter_10__u_filter_stored_value_q_reg_1428 (.o(net1428));
 b15tihi00an1n03x5 u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_2__1429 (.o(net1429));
 b15tihi00an1n03x5 u_gpio_gen_filter_11__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_11__u_filter_filter_q_reg_1430 (.o(net1430));
 b15tihi00an1n03x5 u_gpio_gen_filter_11__u_filter_stored_value_q_reg_1431 (.o(net1431));
 b15tihi00an1n03x5 u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_2__1432 (.o(net1432));
 b15tihi00an1n03x5 u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_12__u_filter_filter_q_reg_1433 (.o(net1433));
 b15tihi00an1n03x5 u_gpio_gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1434 (.o(net1434));
 b15tihi00an1n03x5 u_gpio_gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_0__1435 (.o(net1435));
 b15tihi00an1n03x5 u_gpio_gen_filter_12__u_filter_stored_value_q_reg_1436 (.o(net1436));
 b15tihi00an1n03x5 u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_1__1437 (.o(net1437));
 b15tihi00an1n03x5 u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_13__u_filter_diff_ctr_q_reg_3__1438 (.o(net1438));
 b15tihi00an1n03x5 u_gpio_gen_filter_13__u_filter_filter_q_reg_u_gpio_gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1439 (.o(net1439));
 b15tihi00an1n03x5 u_gpio_gen_filter_13__u_filter_stored_value_q_reg_1440 (.o(net1440));
 b15tihi00an1n03x5 u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_2__1441 (.o(net1441));
 b15tihi00an1n03x5 u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_0__1442 (.o(net1442));
 b15tihi00an1n03x5 u_gpio_gen_filter_14__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_14__u_filter_filter_q_reg_1443 (.o(net1443));
 b15tihi00an1n03x5 u_gpio_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1444 (.o(net1444));
 b15tihi00an1n03x5 u_gpio_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_0__1445 (.o(net1445));
 b15tihi00an1n03x5 u_gpio_gen_filter_14__u_filter_stored_value_q_reg_1446 (.o(net1446));
 b15tihi00an1n03x5 u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_2__1447 (.o(net1447));
 b15tihi00an1n03x5 u_gpio_gen_filter_15__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_15__u_filter_filter_q_reg_1448 (.o(net1448));
 b15tihi00an1n03x5 u_gpio_gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_0__1449 (.o(net1449));
 b15tihi00an1n03x5 u_gpio_gen_filter_15__u_filter_stored_value_q_reg_1450 (.o(net1450));
 b15tihi00an1n03x5 u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_1__1451 (.o(net1451));
 b15tihi00an1n03x5 u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_16__u_filter_diff_ctr_q_reg_3__1452 (.o(net1452));
 b15tihi00an1n03x5 u_gpio_gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1453 (.o(net1453));
 b15tihi00an1n03x5 u_gpio_gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_0__1454 (.o(net1454));
 b15tihi00an1n03x5 u_gpio_gen_filter_16__u_filter_stored_value_q_reg_1455 (.o(net1455));
 b15tihi00an1n03x5 u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_2__1456 (.o(net1456));
 b15tihi00an1n03x5 u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_17__u_filter_filter_q_reg_1457 (.o(net1457));
 b15tihi00an1n03x5 u_gpio_gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_3__1458 (.o(net1458));
 b15tihi00an1n03x5 u_gpio_gen_filter_17__u_filter_stored_value_q_reg_1459 (.o(net1459));
 b15tihi00an1n03x5 u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_1__1460 (.o(net1460));
 b15tihi00an1n03x5 u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_18__u_filter_diff_ctr_q_reg_3__1461 (.o(net1461));
 b15tihi00an1n03x5 u_gpio_gen_filter_18__u_filter_filter_q_reg_u_gpio_gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1462 (.o(net1462));
 b15tihi00an1n03x5 u_gpio_gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1463 (.o(net1463));
 b15tihi00an1n03x5 u_gpio_gen_filter_18__u_filter_stored_value_q_reg_1464 (.o(net1464));
 b15tihi00an1n03x5 u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_2__1465 (.o(net1465));
 b15tihi00an1n03x5 u_gpio_gen_filter_19__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_19__u_filter_filter_q_reg_1466 (.o(net1466));
 b15tihi00an1n03x5 u_gpio_gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_2__1467 (.o(net1467));
 b15tihi00an1n03x5 u_gpio_gen_filter_19__u_filter_stored_value_q_reg_1468 (.o(net1468));
 b15tihi00an1n03x5 u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_1__1469 (.o(net1469));
 b15tihi00an1n03x5 u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_1__u_filter_diff_ctr_q_reg_3__1470 (.o(net1470));
 b15tihi00an1n03x5 u_gpio_gen_filter_1__u_filter_filter_q_reg_u_gpio_gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1471 (.o(net1471));
 b15tihi00an1n03x5 u_gpio_gen_filter_1__u_filter_stored_value_q_reg_1472 (.o(net1472));
 b15tihi00an1n03x5 u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_20__u_filter_diff_ctr_q_reg_2__1473 (.o(net1473));
 b15tihi00an1n03x5 u_gpio_gen_filter_20__u_filter_filter_q_reg_u_gpio_gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1474 (.o(net1474));
 b15tihi00an1n03x5 u_gpio_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1475 (.o(net1475));
 b15tihi00an1n03x5 u_gpio_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_0__1476 (.o(net1476));
 b15tihi00an1n03x5 u_gpio_gen_filter_20__u_filter_stored_value_q_reg_1477 (.o(net1477));
 b15tihi00an1n03x5 u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_1__1478 (.o(net1478));
 b15tihi00an1n03x5 u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_21__u_filter_diff_ctr_q_reg_3__1479 (.o(net1479));
 b15tihi00an1n03x5 u_gpio_gen_filter_21__u_filter_filter_q_reg_u_gpio_gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1480 (.o(net1480));
 b15tihi00an1n03x5 u_gpio_gen_filter_21__u_filter_stored_value_q_reg_1481 (.o(net1481));
 b15tihi00an1n03x5 u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_22__u_filter_diff_ctr_q_reg_3__1482 (.o(net1482));
 b15tihi00an1n03x5 u_gpio_gen_filter_22__u_filter_filter_q_reg_u_gpio_gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1483 (.o(net1483));
 b15tihi00an1n03x5 u_gpio_gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1484 (.o(net1484));
 b15tihi00an1n03x5 u_gpio_gen_filter_22__u_filter_stored_value_q_reg_1485 (.o(net1485));
 b15tihi00an1n03x5 u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_2__1486 (.o(net1486));
 b15tihi00an1n03x5 u_gpio_gen_filter_23__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_23__u_filter_filter_q_reg_1487 (.o(net1487));
 b15tihi00an1n03x5 u_gpio_gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_0__1488 (.o(net1488));
 b15tihi00an1n03x5 u_gpio_gen_filter_23__u_filter_stored_value_q_reg_1489 (.o(net1489));
 b15tihi00an1n03x5 u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_2__1490 (.o(net1490));
 b15tihi00an1n03x5 u_gpio_gen_filter_24__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_24__u_filter_filter_q_reg_1491 (.o(net1491));
 b15tihi00an1n03x5 u_gpio_gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1492 (.o(net1492));
 b15tihi00an1n03x5 u_gpio_gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_0__1493 (.o(net1493));
 b15tihi00an1n03x5 u_gpio_gen_filter_24__u_filter_stored_value_q_reg_1494 (.o(net1494));
 b15tihi00an1n03x5 u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_2__1495 (.o(net1495));
 b15tihi00an1n03x5 u_gpio_gen_filter_25__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1496 (.o(net1496));
 b15tihi00an1n03x5 u_gpio_gen_filter_25__u_filter_filter_q_reg_u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_0__1497 (.o(net1497));
 b15tihi00an1n03x5 u_gpio_gen_filter_25__u_filter_stored_value_q_reg_1498 (.o(net1498));
 b15tihi00an1n03x5 u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_2__1499 (.o(net1499));
 b15tihi00an1n03x5 u_gpio_gen_filter_26__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_29__u_filter_filter_q_reg_1500 (.o(net1500));
 b15tihi00an1n03x5 u_gpio_gen_filter_26__u_filter_filter_q_reg_u_gpio_intr_hw_intr_o_reg_12__1501 (.o(net1501));
 b15tihi00an1n03x5 u_gpio_gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1502 (.o(net1502));
 b15tihi00an1n03x5 u_gpio_gen_filter_26__u_filter_stored_value_q_reg_1503 (.o(net1503));
 b15tihi00an1n03x5 u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_2__1504 (.o(net1504));
 b15tihi00an1n03x5 u_gpio_gen_filter_27__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_27__u_filter_filter_q_reg_1505 (.o(net1505));
 b15tihi00an1n03x5 u_gpio_gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_intr_hw_intr_o_reg_24__1506 (.o(net1506));
 b15tihi00an1n03x5 u_gpio_gen_filter_27__u_filter_stored_value_q_reg_1507 (.o(net1507));
 b15tihi00an1n03x5 u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_1__1508 (.o(net1508));
 b15tihi00an1n03x5 u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_28__u_filter_diff_ctr_q_reg_3__1509 (.o(net1509));
 b15tihi00an1n03x5 u_gpio_gen_filter_28__u_filter_filter_q_reg_u_gpio_gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1510 (.o(net1510));
 b15tihi00an1n03x5 u_gpio_gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1511 (.o(net1511));
 b15tihi00an1n03x5 u_gpio_gen_filter_28__u_filter_stored_value_q_reg_1512 (.o(net1512));
 b15tihi00an1n03x5 u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_1__1513 (.o(net1513));
 b15tihi00an1n03x5 u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_29__u_filter_diff_ctr_q_reg_3__1514 (.o(net1514));
 b15tihi00an1n03x5 u_gpio_gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_0__1515 (.o(net1515));
 b15tihi00an1n03x5 u_gpio_gen_filter_29__u_filter_stored_value_q_reg_1516 (.o(net1516));
 b15tihi00an1n03x5 u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_1__1517 (.o(net1517));
 b15tihi00an1n03x5 u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_2__u_filter_diff_ctr_q_reg_3__1518 (.o(net1518));
 b15tihi00an1n03x5 u_gpio_gen_filter_2__u_filter_filter_q_reg_u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_1__1519 (.o(net1519));
 b15tihi00an1n03x5 u_gpio_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1520 (.o(net1520));
 b15tihi00an1n03x5 u_gpio_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_0__1521 (.o(net1521));
 b15tihi00an1n03x5 u_gpio_gen_filter_2__u_filter_stored_value_q_reg_1522 (.o(net1522));
 b15tihi00an1n03x5 u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_30__u_filter_filter_q_reg_1523 (.o(net1523));
 b15tihi00an1n03x5 u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_30__u_filter_diff_ctr_q_reg_3__1524 (.o(net1524));
 b15tihi00an1n03x5 u_gpio_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1525 (.o(net1525));
 b15tihi00an1n03x5 u_gpio_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1526 (.o(net1526));
 b15tihi00an1n03x5 u_gpio_gen_filter_30__u_filter_stored_value_q_reg_1527 (.o(net1527));
 b15tihi00an1n03x5 u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_1__1528 (.o(net1528));
 b15tihi00an1n03x5 u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_2__u_gpio_gen_filter_31__u_filter_diff_ctr_q_reg_3__1529 (.o(net1529));
 b15tihi00an1n03x5 u_gpio_gen_filter_31__u_filter_filter_q_reg_u_gpio_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1530 (.o(net1530));
 b15tihi00an1n03x5 u_gpio_gen_filter_31__u_filter_stored_value_q_reg_1531 (.o(net1531));
 b15tihi00an1n03x5 u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_2__1532 (.o(net1532));
 b15tihi00an1n03x5 u_gpio_gen_filter_3__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_3__u_filter_filter_q_reg_1533 (.o(net1533));
 b15tihi00an1n03x5 u_gpio_gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_7__u_filter_filter_q_reg_1534 (.o(net1534));
 b15tihi00an1n03x5 u_gpio_gen_filter_3__u_filter_stored_value_q_reg_1535 (.o(net1535));
 b15tihi00an1n03x5 u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_2__1536 (.o(net1536));
 b15tihi00an1n03x5 u_gpio_gen_filter_4__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_4__u_filter_filter_q_reg_1537 (.o(net1537));
 b15tihi00an1n03x5 u_gpio_gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1538 (.o(net1538));
 b15tihi00an1n03x5 u_gpio_gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_0__1539 (.o(net1539));
 b15tihi00an1n03x5 u_gpio_gen_filter_4__u_filter_stored_value_q_reg_1540 (.o(net1540));
 b15tihi00an1n03x5 u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_2__1541 (.o(net1541));
 b15tihi00an1n03x5 u_gpio_gen_filter_5__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_5__u_filter_filter_q_reg_1542 (.o(net1542));
 b15tihi00an1n03x5 u_gpio_gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_12__u_filter_diff_ctr_q_reg_0__1543 (.o(net1543));
 b15tihi00an1n03x5 u_gpio_gen_filter_5__u_filter_stored_value_q_reg_1544 (.o(net1544));
 b15tihi00an1n03x5 u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_2__1545 (.o(net1545));
 b15tihi00an1n03x5 u_gpio_gen_filter_6__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_6__u_filter_filter_q_reg_1546 (.o(net1546));
 b15tihi00an1n03x5 u_gpio_gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1547 (.o(net1547));
 b15tihi00an1n03x5 u_gpio_gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_17__u_filter_diff_ctr_q_reg_0__1548 (.o(net1548));
 b15tihi00an1n03x5 u_gpio_gen_filter_6__u_filter_stored_value_q_reg_1549 (.o(net1549));
 b15tihi00an1n03x5 u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_0__u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_2__1550 (.o(net1550));
 b15tihi00an1n03x5 u_gpio_gen_filter_7__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_0__1551 (.o(net1551));
 b15tihi00an1n03x5 u_gpio_gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1552 (.o(net1552));
 b15tihi00an1n03x5 u_gpio_gen_filter_7__u_filter_stored_value_q_reg_1553 (.o(net1553));
 b15tihi00an1n03x5 u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_2__1554 (.o(net1554));
 b15tihi00an1n03x5 u_gpio_gen_filter_8__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_0__1555 (.o(net1555));
 b15tihi00an1n03x5 u_gpio_gen_filter_8__u_filter_filter_q_reg_u_gpio_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1556 (.o(net1556));
 b15tihi00an1n03x5 u_gpio_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1557 (.o(net1557));
 b15tihi00an1n03x5 u_gpio_gen_filter_8__u_filter_stored_value_q_reg_1558 (.o(net1558));
 b15tihi00an1n03x5 u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_1__u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_2__1559 (.o(net1559));
 b15tihi00an1n03x5 u_gpio_gen_filter_9__u_filter_diff_ctr_q_reg_3__u_gpio_gen_filter_9__u_filter_filter_q_reg_1560 (.o(net1560));
 b15tihi00an1n03x5 u_gpio_gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_gpio_gen_filter_10__u_filter_diff_ctr_q_reg_2__1561 (.o(net1561));
 b15tihi00an1n03x5 u_gpio_gen_filter_9__u_filter_stored_value_q_reg_1562 (.o(net1562));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_0__u_gpio_intr_hw_intr_o_reg_1__1563 (.o(net1563));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_10__u_gpio_intr_hw_intr_o_reg_11__1564 (.o(net1564));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_13__u_gpio_intr_hw_intr_o_reg_14__1565 (.o(net1565));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_15__u_gpio_intr_hw_intr_o_reg_16__1566 (.o(net1566));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_17__u_gpio_intr_hw_intr_o_reg_18__1567 (.o(net1567));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_19__u_gpio_intr_hw_intr_o_reg_20__1568 (.o(net1568));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_21__u_gpio_intr_hw_intr_o_reg_29__1569 (.o(net1569));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_22__u_gpio_intr_hw_intr_o_reg_23__1570 (.o(net1570));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_25__u_gpio_intr_hw_intr_o_reg_26__1571 (.o(net1571));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_27__u_gpio_u_reg_err_q_reg_1572 (.o(net1572));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_28__u_gpio_u_reg_u_data_in_q_reg_2__1573 (.o(net1573));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_2__u_gpio_intr_hw_intr_o_reg_3__1574 (.o(net1574));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_30__u_gpio_intr_hw_intr_o_reg_31__1575 (.o(net1575));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_4__u_gpio_intr_hw_intr_o_reg_5__1576 (.o(net1576));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_6__u_gpio_intr_hw_intr_o_reg_7__1577 (.o(net1577));
 b15tihi00an1n03x5 u_gpio_intr_hw_intr_o_reg_8__u_gpio_intr_hw_intr_o_reg_9__1578 (.o(net1578));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_0__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_1__1579 (.o(net1579));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_10__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_11__1580 (.o(net1580));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_12__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_13__1581 (.o(net1581));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_14__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_15__1582 (.o(net1582));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_16__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_17__1583 (.o(net1583));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_18__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_19__1584 (.o(net1584));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_20__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_21__1585 (.o(net1585));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_22__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_23__1586 (.o(net1586));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_24__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_25__1587 (.o(net1587));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_26__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_27__1588 (.o(net1588));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_28__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_29__1589 (.o(net1589));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_2__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_3__1590 (.o(net1590));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_30__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_31__1591 (.o(net1591));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_4__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_5__1592 (.o(net1592));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_6__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_7__1593 (.o(net1593));
 b15tihi00an1n03x5 u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_8__u_gpio_u_reg_u_ctrl_en_input_filter_q_reg_9__1594 (.o(net1594));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_0__u_gpio_u_reg_u_data_in_q_reg_1__1595 (.o(net1595));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_13__1596 (.o(net1596));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_14__u_gpio_u_reg_u_data_in_q_reg_23__1597 (.o(net1597));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_15__u_gpio_u_reg_u_data_in_q_reg_16__1598 (.o(net1598));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_17__u_gpio_u_reg_u_data_in_q_reg_18__1599 (.o(net1599));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_19__u_gpio_u_reg_u_data_in_q_reg_20__1600 (.o(net1600));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_21__u_gpio_u_reg_u_data_in_q_reg_22__1601 (.o(net1601));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_24__u_gpio_u_reg_u_data_in_q_reg_25__1602 (.o(net1602));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_26__u_gpio_u_reg_u_data_in_q_reg_28__1603 (.o(net1603));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_27__u_gpio_u_reg_u_data_in_q_reg_30__1604 (.o(net1604));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_29__1605 (.o(net1605));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_31__1606 (.o(net1606));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_3__u_gpio_u_reg_u_data_in_q_reg_4__1607 (.o(net1607));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_5__u_gpio_u_reg_u_data_in_q_reg_12__1608 (.o(net1608));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_6__u_gpio_u_reg_u_data_in_q_reg_7__1609 (.o(net1609));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_8__u_gpio_u_reg_u_data_in_q_reg_11__1610 (.o(net1610));
 b15tihi00an1n03x5 u_gpio_u_reg_u_data_in_q_reg_9__u_gpio_u_reg_u_data_in_q_reg_10__1611 (.o(net1611));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_1__1612 (.o(net1612));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_11__1613 (.o(net1613));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_13__1614 (.o(net1614));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_15__1615 (.o(net1615));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_17__1616 (.o(net1616));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_19__1617 (.o(net1617));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_21__1618 (.o(net1618));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_23__1619 (.o(net1619));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_25__1620 (.o(net1620));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_27__1621 (.o(net1621));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_29__1622 (.o(net1622));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_3__1623 (.o(net1623));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_31__1624 (.o(net1624));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_5__1625 (.o(net1625));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_7__1626 (.o(net1626));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_falling_q_reg_9__1627 (.o(net1627));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_1__1628 (.o(net1628));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_11__1629 (.o(net1629));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_13__1630 (.o(net1630));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_15__1631 (.o(net1631));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_17__1632 (.o(net1632));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_19__1633 (.o(net1633));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_21__1634 (.o(net1634));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_23__1635 (.o(net1635));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_25__1636 (.o(net1636));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_27__1637 (.o(net1637));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_29__1638 (.o(net1638));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_3__1639 (.o(net1639));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_31__1640 (.o(net1640));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_5__1641 (.o(net1641));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_7__1642 (.o(net1642));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_q_reg_9__1643 (.o(net1643));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_1__1644 (.o(net1644));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_11__1645 (.o(net1645));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_13__1646 (.o(net1646));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_15__1647 (.o(net1647));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_17__1648 (.o(net1648));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_19__1649 (.o(net1649));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_21__1650 (.o(net1650));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_23__1651 (.o(net1651));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_25__1652 (.o(net1652));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_27__1653 (.o(net1653));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_29__1654 (.o(net1654));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_3__1655 (.o(net1655));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_31__1656 (.o(net1656));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_5__1657 (.o(net1657));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_7__1658 (.o(net1658));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_lvllow_q_reg_9__1659 (.o(net1659));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_0__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_1__1660 (.o(net1660));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_10__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_11__1661 (.o(net1661));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_12__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_13__1662 (.o(net1662));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_14__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_15__1663 (.o(net1663));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_16__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_17__1664 (.o(net1664));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_18__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_19__1665 (.o(net1665));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_20__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_21__1666 (.o(net1666));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_22__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_23__1667 (.o(net1667));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_24__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_25__1668 (.o(net1668));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_26__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_27__1669 (.o(net1669));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_28__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_29__1670 (.o(net1670));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_2__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_3__1671 (.o(net1671));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_30__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_31__1672 (.o(net1672));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_4__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_5__1673 (.o(net1673));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_6__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_7__1674 (.o(net1674));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_8__u_gpio_u_reg_u_intr_ctrl_en_rising_q_reg_9__1675 (.o(net1675));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_0__u_gpio_u_reg_u_intr_enable_q_reg_1__1676 (.o(net1676));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_10__u_gpio_u_reg_u_intr_enable_q_reg_11__1677 (.o(net1677));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_12__u_gpio_u_reg_u_intr_enable_q_reg_13__1678 (.o(net1678));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_14__u_gpio_u_reg_u_intr_enable_q_reg_15__1679 (.o(net1679));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_16__u_gpio_u_reg_u_intr_enable_q_reg_17__1680 (.o(net1680));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_18__u_gpio_u_reg_u_intr_enable_q_reg_19__1681 (.o(net1681));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_20__u_gpio_u_reg_u_intr_enable_q_reg_21__1682 (.o(net1682));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_22__u_gpio_u_reg_u_intr_enable_q_reg_23__1683 (.o(net1683));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_24__u_gpio_u_reg_u_intr_enable_q_reg_25__1684 (.o(net1684));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_26__u_gpio_u_reg_u_intr_enable_q_reg_27__1685 (.o(net1685));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_28__u_gpio_u_reg_u_intr_enable_q_reg_29__1686 (.o(net1686));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_2__u_gpio_u_reg_u_intr_enable_q_reg_3__1687 (.o(net1687));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_30__u_gpio_u_reg_u_intr_enable_q_reg_31__1688 (.o(net1688));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_4__u_gpio_u_reg_u_intr_enable_q_reg_5__1689 (.o(net1689));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_6__u_gpio_u_reg_u_intr_enable_q_reg_7__1690 (.o(net1690));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_enable_q_reg_8__u_gpio_u_reg_u_intr_enable_q_reg_9__1691 (.o(net1691));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_0__u_gpio_u_reg_u_intr_state_q_reg_1__1692 (.o(net1692));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_10__u_gpio_u_reg_u_intr_state_q_reg_11__1693 (.o(net1693));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_12__u_gpio_u_reg_u_intr_state_q_reg_13__1694 (.o(net1694));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_14__u_gpio_u_reg_u_intr_state_q_reg_15__1695 (.o(net1695));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_16__u_gpio_u_reg_u_intr_state_q_reg_17__1696 (.o(net1696));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_18__u_gpio_u_reg_u_intr_state_q_reg_19__1697 (.o(net1697));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_20__u_gpio_u_reg_u_intr_state_q_reg_21__1698 (.o(net1698));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_22__u_gpio_u_reg_u_intr_state_q_reg_23__1699 (.o(net1699));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_24__u_gpio_u_reg_u_intr_state_q_reg_25__1700 (.o(net1700));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_26__u_gpio_u_reg_u_intr_state_q_reg_27__1701 (.o(net1701));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_28__u_gpio_u_reg_u_intr_state_q_reg_29__1702 (.o(net1702));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_2__u_gpio_u_reg_u_intr_state_q_reg_3__1703 (.o(net1703));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_30__u_gpio_u_reg_u_intr_state_q_reg_31__1704 (.o(net1704));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_4__u_gpio_u_reg_u_intr_state_q_reg_5__1705 (.o(net1705));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_6__u_gpio_u_reg_u_intr_state_q_reg_7__1706 (.o(net1706));
 b15tihi00an1n03x5 u_gpio_u_reg_u_intr_state_q_reg_8__u_gpio_u_reg_u_intr_state_q_reg_9__1707 (.o(net1707));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_error_reg_1708 (.o(net1708));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_outstanding_reg_1709 (.o(net1709));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_0__u_gpio_u_reg_u_reg_if_rdata_reg_1__1710 (.o(net1710));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_10__u_gpio_u_reg_u_reg_if_rdata_reg_11__1711 (.o(net1711));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_12__u_gpio_u_reg_u_reg_if_rdata_reg_13__1712 (.o(net1712));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_14__u_gpio_u_reg_u_reg_if_rdata_reg_15__1713 (.o(net1713));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_16__u_gpio_u_reg_u_reg_if_rdata_reg_17__1714 (.o(net1714));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_18__u_gpio_u_reg_u_reg_if_rdata_reg_19__1715 (.o(net1715));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_20__u_gpio_u_reg_u_reg_if_rdata_reg_21__1716 (.o(net1716));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_22__u_gpio_u_reg_u_reg_if_rdata_reg_23__1717 (.o(net1717));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_24__u_gpio_u_reg_u_reg_if_rdata_reg_25__1718 (.o(net1718));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_26__u_gpio_u_reg_u_reg_if_rdata_reg_27__1719 (.o(net1719));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_28__u_gpio_u_reg_u_reg_if_rdata_reg_29__1720 (.o(net1720));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_2__u_gpio_u_reg_u_reg_if_rdata_reg_3__1721 (.o(net1721));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_30__u_gpio_u_reg_u_reg_if_rdata_reg_31__1722 (.o(net1722));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_4__u_gpio_u_reg_u_reg_if_rdata_reg_5__1723 (.o(net1723));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_6__u_gpio_u_reg_u_reg_if_rdata_reg_7__1724 (.o(net1724));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rdata_reg_8__u_gpio_u_reg_u_reg_if_rdata_reg_9__1725 (.o(net1725));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_reqid_reg_0__u_gpio_u_reg_u_reg_if_reqid_reg_1__1726 (.o(net1726));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_reqid_reg_2__u_gpio_u_reg_u_reg_if_reqid_reg_3__1727 (.o(net1727));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_reqid_reg_4__u_gpio_u_reg_u_reg_if_reqid_reg_5__1728 (.o(net1728));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_reqid_reg_6__u_gpio_u_reg_u_reg_if_reqid_reg_7__1729 (.o(net1729));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_reqsz_reg_0__1730 (.o(net1730));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_reqsz_reg_1__1731 (.o(net1731));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rspop_reg_0__1732 (.o(net1732));
 b15tihi00an1n03x5 u_gpio_u_reg_u_reg_if_rspop_reg_1__u_gpio_u_reg_u_reg_if_rspop_reg_2__1733 (.o(net1733));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_dev_select_outstanding_reg_0__1734 (.o(net1734));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_dev_select_outstanding_reg_1__1735 (.o(net1735));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_dev_select_outstanding_reg_2__1736 (.o(net1736));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type_reg_0__1737 (.o(net1737));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type_reg_1__1738 (.o(net1738));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type_reg_2__1739 (.o(net1739));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_instr_type_reg_3__1740 (.o(net1740));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_opcode_reg_0__1741 (.o(net1741));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_opcode_reg_1__1742 (.o(net1742));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_opcode_reg_2__1743 (.o(net1743));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_req_pending_reg_1744 (.o(net1744));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_rsp_pending_reg_1745 (.o(net1745));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_size_reg_0__1746 (.o(net1746));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_size_reg_1__1747 (.o(net1747));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_0__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_1__1748 (.o(net1748));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_2__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_3__1749 (.o(net1749));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_4__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_5__1750 (.o(net1750));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_6__u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_source_reg_7__1751 (.o(net1751));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_0__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_1__1752 (.o(net1752));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_2__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_3__1753 (.o(net1753));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_4__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_5__1754 (.o(net1754));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_6__u_xbar_periph_u_s1n_6_num_req_outstanding_reg_7__1755 (.o(net1755));
 b15tihi00an1n03x5 u_xbar_periph_u_s1n_6_num_req_outstanding_reg_8__1756 (.o(net1756));
 b15cbf000an1n16x5 clkbuf_leaf_1_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_1_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_2_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_2_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_3_clk_i (.clk(clknet_1_1__leaf_clk_i),
    .clkout(clknet_leaf_3_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_4_clk_i (.clk(clknet_1_1__leaf_clk_i),
    .clkout(clknet_leaf_4_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_5_clk_i (.clk(clknet_1_1__leaf_clk_i),
    .clkout(clknet_leaf_5_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_6_clk_i (.clk(clknet_1_1__leaf_clk_i),
    .clkout(clknet_leaf_6_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_7_clk_i (.clk(clknet_1_1__leaf_clk_i),
    .clkout(clknet_leaf_7_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_8_clk_i (.clk(clknet_1_1__leaf_clk_i),
    .clkout(clknet_leaf_8_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_9_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_9_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_10_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_10_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_11_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_11_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_12_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_12_clk_i));
 b15cbf000an1n16x5 clkbuf_0_clk_i (.clk(net1757),
    .clkout(clknet_0_clk_i));
 b15cbf000an1n16x5 clkbuf_1_0__f_clk_i (.clk(clknet_0_clk_i),
    .clkout(clknet_1_0__leaf_clk_i));
 b15cbf000an1n16x5 clkbuf_1_1__f_clk_i (.clk(clknet_0_clk_i),
    .clkout(clknet_1_1__leaf_clk_i));
 b15cbf000an1n16x5 clkbuf_0_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713 (.clk(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713),
    .clkout(clknet_0_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713 (.clk(clknet_0_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713),
    .clkout(clknet_1_0__leaf_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713 (.clk(clknet_0_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713),
    .clkout(clknet_1_1__leaf_u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_net3713));
 b15cbf000an1n16x5 clkbuf_0_u_xbar_periph_u_s1n_6_net3695 (.clk(u_xbar_periph_u_s1n_6_net3695),
    .clkout(clknet_0_u_xbar_periph_u_s1n_6_net3695));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_xbar_periph_u_s1n_6_net3695 (.clk(clknet_0_u_xbar_periph_u_s1n_6_net3695),
    .clkout(clknet_1_0__leaf_u_xbar_periph_u_s1n_6_net3695));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_xbar_periph_u_s1n_6_net3695 (.clk(clknet_0_u_xbar_periph_u_s1n_6_net3695),
    .clkout(clknet_1_1__leaf_u_xbar_periph_u_s1n_6_net3695));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_reg_if_net3667 (.clk(u_gpio_u_reg_u_reg_if_net3667),
    .clkout(clknet_0_u_gpio_u_reg_u_reg_if_net3667));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_reg_if_net3667 (.clk(clknet_0_u_gpio_u_reg_u_reg_if_net3667),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3667));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_reg_if_net3667 (.clk(clknet_0_u_gpio_u_reg_u_reg_if_net3667),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3667));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_reg_if_net3673 (.clk(u_gpio_u_reg_u_reg_if_net3673),
    .clkout(clknet_0_u_gpio_u_reg_u_reg_if_net3673));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_reg_if_net3673 (.clk(clknet_0_u_gpio_u_reg_u_reg_if_net3673),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3673));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_reg_if_net3673 (.clk(clknet_0_u_gpio_u_reg_u_reg_if_net3673),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3673));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_reg_if_net3678 (.clk(u_gpio_u_reg_u_reg_if_net3678),
    .clkout(clknet_0_u_gpio_u_reg_u_reg_if_net3678));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_reg_if_net3678 (.clk(clknet_0_u_gpio_u_reg_u_reg_if_net3678),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_reg_if_net3678));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_reg_if_net3678 (.clk(clknet_0_u_gpio_u_reg_u_reg_if_net3678),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_reg_if_net3678));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_intr_state_net3644 (.clk(u_gpio_u_reg_u_intr_state_net3644),
    .clkout(clknet_0_u_gpio_u_reg_u_intr_state_net3644));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_intr_state_net3644 (.clk(clknet_0_u_gpio_u_reg_u_intr_state_net3644),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_intr_state_net3644));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_intr_state_net3644 (.clk(clknet_0_u_gpio_u_reg_u_intr_state_net3644),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_intr_state_net3644));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_intr_state_net3650 (.clk(u_gpio_u_reg_u_intr_state_net3650),
    .clkout(clknet_0_u_gpio_u_reg_u_intr_state_net3650));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_intr_state_net3650 (.clk(clknet_0_u_gpio_u_reg_u_intr_state_net3650),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_intr_state_net3650));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_intr_state_net3650 (.clk(clknet_0_u_gpio_u_reg_u_intr_state_net3650),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_intr_state_net3650));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_intr_enable_net3621 (.clk(u_gpio_u_reg_u_intr_enable_net3621),
    .clkout(clknet_0_u_gpio_u_reg_u_intr_enable_net3621));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_intr_enable_net3621 (.clk(clknet_0_u_gpio_u_reg_u_intr_enable_net3621),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_intr_enable_net3621));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_intr_enable_net3621 (.clk(clknet_0_u_gpio_u_reg_u_intr_enable_net3621),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_intr_enable_net3621));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_intr_enable_net3627 (.clk(u_gpio_u_reg_u_intr_enable_net3627),
    .clkout(clknet_0_u_gpio_u_reg_u_intr_enable_net3627));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_intr_enable_net3627 (.clk(clknet_0_u_gpio_u_reg_u_intr_enable_net3627),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_intr_enable_net3627));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_intr_enable_net3627 (.clk(clknet_0_u_gpio_u_reg_u_intr_enable_net3627),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_intr_enable_net3627));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621 (.clk(u_gpio_u_reg_u_intr_ctrl_en_rising_net3621),
    .clkout(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3621));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627 (.clk(u_gpio_u_reg_u_intr_ctrl_en_rising_net3627),
    .clkout(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_rising_net3627));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621 (.clk(u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621),
    .clkout(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3621));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627 (.clk(u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627),
    .clkout(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvllow_net3627));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621 (.clk(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621),
    .clkout(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3621));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627 (.clk(u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627),
    .clkout(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_lvlhigh_net3627));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621 (.clk(u_gpio_u_reg_u_intr_ctrl_en_falling_net3621),
    .clkout(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3621));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627 (.clk(u_gpio_u_reg_u_intr_ctrl_en_falling_net3627),
    .clkout(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627 (.clk(clknet_0_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_intr_ctrl_en_falling_net3627));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_ctrl_en_input_filter_net3621 (.clk(u_gpio_u_reg_u_ctrl_en_input_filter_net3621),
    .clkout(clknet_0_u_gpio_u_reg_u_ctrl_en_input_filter_net3621));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_ctrl_en_input_filter_net3621 (.clk(clknet_0_u_gpio_u_reg_u_ctrl_en_input_filter_net3621),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3621));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_ctrl_en_input_filter_net3621 (.clk(clknet_0_u_gpio_u_reg_u_ctrl_en_input_filter_net3621),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3621));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_u_reg_u_ctrl_en_input_filter_net3627 (.clk(u_gpio_u_reg_u_ctrl_en_input_filter_net3627),
    .clkout(clknet_0_u_gpio_u_reg_u_ctrl_en_input_filter_net3627));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_u_reg_u_ctrl_en_input_filter_net3627 (.clk(clknet_0_u_gpio_u_reg_u_ctrl_en_input_filter_net3627),
    .clkout(clknet_1_0__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3627));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_u_reg_u_ctrl_en_input_filter_net3627 (.clk(clknet_0_u_gpio_u_reg_u_ctrl_en_input_filter_net3627),
    .clkout(clknet_1_1__leaf_u_gpio_u_reg_u_ctrl_en_input_filter_net3627));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_net3588 (.clk(u_gpio_net3588),
    .clkout(clknet_0_u_gpio_net3588));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_net3588 (.clk(clknet_0_u_gpio_net3588),
    .clkout(clknet_1_0__leaf_u_gpio_net3588));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_net3588 (.clk(clknet_0_u_gpio_net3588),
    .clkout(clknet_1_1__leaf_u_gpio_net3588));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_net3594 (.clk(u_gpio_net3594),
    .clkout(clknet_0_u_gpio_net3594));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_net3594 (.clk(clknet_0_u_gpio_net3594),
    .clkout(clknet_1_0__leaf_u_gpio_net3594));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_net3594 (.clk(clknet_0_u_gpio_net3594),
    .clkout(clknet_1_1__leaf_u_gpio_net3594));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_net3599 (.clk(u_gpio_net3599),
    .clkout(clknet_0_u_gpio_net3599));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_net3599 (.clk(clknet_0_u_gpio_net3599),
    .clkout(clknet_1_0__leaf_u_gpio_net3599));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_net3599 (.clk(clknet_0_u_gpio_net3599),
    .clkout(clknet_1_1__leaf_u_gpio_net3599));
 b15cbf000an1n16x5 clkbuf_0_u_gpio_net3604 (.clk(u_gpio_net3604),
    .clkout(clknet_0_u_gpio_net3604));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_gpio_net3604 (.clk(clknet_0_u_gpio_net3604),
    .clkout(clknet_1_0__leaf_u_gpio_net3604));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_gpio_net3604 (.clk(clknet_0_u_gpio_net3604),
    .clkout(clknet_1_1__leaf_u_gpio_net3604));
 b15bfn001ah1n32x5 wire1 (.a(clk_i),
    .o(net1757));
 b15cbf034ar1n64x5 hold2 (.clk(u_xbar_periph_u_s1n_6_gen_err_resp_err_resp_err_req_pending),
    .clkout(net1758));
 b15cbf034ar1n64x5 hold3 (.clk(n3618),
    .clkout(net1759));
 b15cbf034ar1n64x5 hold4 (.clk(net168),
    .clkout(net1760));
 b15cbf034ar1n64x5 hold5 (.clk(net1761),
    .clkout(tl_peri_device_o[65]));
 b15cbf034ar1n64x5 hold6 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[6]),
    .clkout(net1762));
 b15cbf034ar1n64x5 hold7 (.clk(net160),
    .clkout(net1763));
 b15cbf034ar1n64x5 hold8 (.clk(net1764),
    .clkout(tl_peri_device_o[55]));
 b15cbf034ar1n64x5 hold9 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[21]),
    .clkout(net1765));
 b15cbf034ar1n64x5 hold10 (.clk(net434),
    .clkout(net1766));
 b15cbf034ar1n64x5 hold11 (.clk(n2944),
    .clkout(net1767));
 b15cbf034ar1n64x5 hold12 (.clk(net165),
    .clkout(net1768));
 b15cbf034ar1n64x5 hold13 (.clk(net1769),
    .clkout(tl_peri_device_o[62]));
 b15cbf034ar1n64x5 hold14 (.clk(net1788),
    .clkout(net1770));
 b15cbf034ar1n64x5 hold15 (.clk(n2916),
    .clkout(net1771));
 b15cbf034ar1n64x5 hold16 (.clk(n2917),
    .clkout(net1772));
 b15cbf034ar1n64x5 hold17 (.clk(n2941),
    .clkout(net1773));
 b15cbf034ar1n64x5 hold18 (.clk(net172),
    .clkout(net1774));
 b15cbf034ar1n64x5 hold19 (.clk(net1775),
    .clkout(tl_peri_device_o[9]));
 b15cbf034ar1n64x5 hold20 (.clk(n1446),
    .clkout(net1776));
 b15cbf034ar1n64x5 hold21 (.clk(n3047),
    .clkout(net1777));
 b15cbf034ar1n64x5 hold22 (.clk(n3050),
    .clkout(net1778));
 b15cbf034ar1n64x5 hold23 (.clk(net146),
    .clkout(net1779));
 b15cbf034ar1n64x5 hold24 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[9]),
    .clkout(net1780));
 b15cbf034ar1n64x5 hold25 (.clk(n2993),
    .clkout(net1781));
 b15cbf034ar1n64x5 hold26 (.clk(net115),
    .clkout(net1782));
 b15cbf034ar1n64x5 hold27 (.clk(net1783),
    .clkout(tl_peri_device_o[13]));
 b15cbf034ar1n64x5 hold28 (.clk(u_xbar_periph_u_s1n_6_dev_select_outstanding[0]),
    .clkout(net1784));
 b15cbf034ar1n64x5 hold29 (.clk(n2895),
    .clkout(net1785));
 b15cbf034ar1n64x5 hold30 (.clk(n3063),
    .clkout(net1786));
 b15cbf034ar1n64x5 hold31 (.clk(net163),
    .clkout(net1787));
 b15cbf034ar1n64x5 hold32 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[22]),
    .clkout(net1788));
 b15cbf034ar1n64x5 hold33 (.clk(net1770),
    .clkout(net1789));
 b15cbf034ar1n64x5 hold34 (.clk(net1861),
    .clkout(net1790));
 b15cbf034ar1n64x5 hold35 (.clk(net1791),
    .clkout(tl_peri_device_o[63]));
 b15cbf034ar1n64x5 hold36 (.clk(gpio_2_xbar[15]),
    .clkout(net1792));
 b15cbf034ar1n64x5 hold37 (.clk(n3105),
    .clkout(net1793));
 b15cbf034ar1n64x5 hold38 (.clk(net135),
    .clkout(net1794));
 b15cbf034ar1n64x5 hold39 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[8]),
    .clkout(net1795));
 b15cbf034ar1n64x5 hold40 (.clk(n2918),
    .clkout(net1796));
 b15cbf034ar1n64x5 hold41 (.clk(net162),
    .clkout(net1797));
 b15cbf034ar1n64x5 hold42 (.clk(net1798),
    .clkout(tl_peri_device_o[57]));
 b15cbf034ar1n64x5 hold43 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[15]),
    .clkout(net1799));
 b15cbf034ar1n64x5 hold44 (.clk(net158),
    .clkout(net1800));
 b15cbf034ar1n64x5 hold45 (.clk(net1801),
    .clkout(tl_peri_device_o[53]));
 b15cbf034ar1n64x5 hold46 (.clk(gpio_2_xbar[11]),
    .clkout(net1802));
 b15cbf034ar1n64x5 hold47 (.clk(n3086),
    .clkout(net1803));
 b15cbf034ar1n64x5 hold48 (.clk(net130),
    .clkout(net1804));
 b15cbf034ar1n64x5 hold49 (.clk(n1454),
    .clkout(net1805));
 b15cbf034ar1n64x5 hold50 (.clk(n3049),
    .clkout(net1806));
 b15cbf034ar1n64x5 hold51 (.clk(n2943),
    .clkout(net1807));
 b15cbf034ar1n64x5 hold52 (.clk(net112),
    .clkout(net1808));
 b15cbf034ar1n64x5 hold53 (.clk(net1809),
    .clkout(tl_peri_device_o[10]));
 b15cbf034ar1n64x5 hold54 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[7]),
    .clkout(net1810));
 b15cbf034ar1n64x5 hold55 (.clk(net161),
    .clkout(net1811));
 b15cbf034ar1n64x5 hold56 (.clk(net1812),
    .clkout(tl_peri_device_o[56]));
 b15cbf034ar1n64x5 hold57 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[16]),
    .clkout(net1813));
 b15cbf034ar1n64x5 hold58 (.clk(net159),
    .clkout(net1814));
 b15cbf034ar1n64x5 hold59 (.clk(net1815),
    .clkout(tl_peri_device_o[54]));
 b15cbf034ar1n64x5 hold60 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[2]),
    .clkout(net1816));
 b15cbf034ar1n64x5 hold61 (.clk(net156),
    .clkout(net1817));
 b15cbf034ar1n64x5 hold62 (.clk(net1818),
    .clkout(tl_peri_device_o[51]));
 b15cbf034ar1n64x5 hold63 (.clk(gpio_2_xbar[17]),
    .clkout(net1819));
 b15cbf034ar1n64x5 hold64 (.clk(net280),
    .clkout(net1820));
 b15cbf034ar1n64x5 hold65 (.clk(net137),
    .clkout(net1821));
 b15cbf034ar1n64x5 hold66 (.clk(net1895),
    .clkout(net1822));
 b15cbf034ar1n64x5 hold67 (.clk(n3045),
    .clkout(net1823));
 b15cbf034ar1n64x5 hold68 (.clk(n3046),
    .clkout(net1824));
 b15cbf034ar1n64x5 hold69 (.clk(net141),
    .clkout(net1825));
 b15cbf034ar1n64x5 hold70 (.clk(gpio_2_xbar[0]),
    .clkout(net1826));
 b15cbf034ar1n64x5 hold71 (.clk(n3096),
    .clkout(net1827));
 b15cbf034ar1n64x5 hold72 (.clk(net1918),
    .clkout(net1828));
 b15cbf034ar1n64x5 hold73 (.clk(n3089),
    .clkout(net1829));
 b15cbf034ar1n64x5 hold74 (.clk(gpio_2_xbar[29]),
    .clkout(net1830));
 b15cbf034ar1n64x5 hold75 (.clk(n3087),
    .clkout(net1831));
 b15cbf034ar1n64x5 hold76 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[1]),
    .clkout(net1832));
 b15cbf034ar1n64x5 hold77 (.clk(net155),
    .clkout(net1833));
 b15cbf034ar1n64x5 hold78 (.clk(net1834),
    .clkout(tl_peri_device_o[50]));
 b15cbf034ar1n64x5 hold79 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[3]),
    .clkout(net1835));
 b15cbf034ar1n64x5 hold80 (.clk(net157),
    .clkout(net1836));
 b15cbf034ar1n64x5 hold81 (.clk(net1837),
    .clkout(tl_peri_device_o[52]));
 b15cbf034ar1n64x5 hold82 (.clk(gpio_2_xbar[5]),
    .clkout(net1838));
 b15cbf034ar1n64x5 hold83 (.clk(n3069),
    .clkout(net1839));
 b15cbf034ar1n64x5 hold84 (.clk(gpio_2_xbar[31]),
    .clkout(net1840));
 b15cbf034ar1n64x5 hold85 (.clk(n3082),
    .clkout(net1841));
 b15cbf034ar1n64x5 hold86 (.clk(gpio_2_xbar[4]),
    .clkout(net1842));
 b15cbf034ar1n64x5 hold87 (.clk(n3067),
    .clkout(net1843));
 b15cbf034ar1n64x5 hold88 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[0]),
    .clkout(net1844));
 b15cbf034ar1n64x5 hold89 (.clk(net153),
    .clkout(net1845));
 b15cbf034ar1n64x5 hold90 (.clk(net1846),
    .clkout(tl_peri_device_o[49]));
 b15cbf034ar1n64x5 hold91 (.clk(gpio_2_xbar[30]),
    .clkout(net1847));
 b15cbf034ar1n64x5 hold92 (.clk(n3085),
    .clkout(net1848));
 b15cbf034ar1n64x5 hold93 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[10]),
    .clkout(net1849));
 b15cbf034ar1n64x5 hold94 (.clk(net113),
    .clkout(net1850));
 b15cbf034ar1n64x5 hold95 (.clk(net1851),
    .clkout(tl_peri_device_o[11]));
 b15cbf034ar1n64x5 hold96 (.clk(gpio_2_xbar[16]),
    .clkout(net1852));
 b15cbf034ar1n64x5 hold97 (.clk(n3080),
    .clkout(net1853));
 b15cbf034ar1n64x5 hold98 (.clk(net1921),
    .clkout(net1854));
 b15cbf034ar1n64x5 hold99 (.clk(n3098),
    .clkout(net1855));
 b15cbf034ar1n64x5 hold100 (.clk(net142),
    .clkout(net1856));
 b15cbf034ar1n64x5 hold101 (.clk(gpio_2_xbar[14]),
    .clkout(net1857));
 b15cbf034ar1n64x5 hold102 (.clk(n3083),
    .clkout(net1858));
 b15cbf034ar1n64x5 hold103 (.clk(net1877),
    .clkout(net1859));
 b15cbf034ar1n64x5 hold104 (.clk(n3620),
    .clkout(net1860));
 b15cbf034ar1n64x5 hold105 (.clk(net166),
    .clkout(net1861));
 b15cbf034ar1n64x5 hold106 (.clk(net117),
    .clkout(net1862));
 b15cbf034ar1n64x5 hold107 (.clk(gpio_2_xbar[24]),
    .clkout(net1863));
 b15cbf034ar1n64x5 hold108 (.clk(n3095),
    .clkout(net1864));
 b15cbf034ar1n64x5 hold109 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[24]),
    .clkout(net1865));
 b15cbf034ar1n64x5 hold110 (.clk(n3612),
    .clkout(net1866));
 b15cbf034ar1n64x5 hold111 (.clk(n3615),
    .clkout(net1867));
 b15cbf034ar1n64x5 hold112 (.clk(net111),
    .clkout(net1868));
 b15cbf034ar1n64x5 hold113 (.clk(net1886),
    .clkout(net1869));
 b15cbf034ar1n64x5 hold114 (.clk(n2930),
    .clkout(net1870));
 b15cbf034ar1n64x5 hold115 (.clk(n2953),
    .clkout(net1871));
 b15cbf034ar1n64x5 hold116 (.clk(net144),
    .clkout(net1872));
 b15cbf034ar1n64x5 hold117 (.clk(net1910),
    .clkout(net1873));
 b15cbf034ar1n64x5 hold118 (.clk(n3059),
    .clkout(net1874));
 b15cbf034ar1n64x5 hold119 (.clk(n2963),
    .clkout(net1875));
 b15cbf034ar1n64x5 hold120 (.clk(net164),
    .clkout(net1876));
 b15cbf034ar1n64x5 hold121 (.clk(u_xbar_periph_u_s1n_6_dev_select_outstanding[1]),
    .clkout(net1877));
 b15cbf034ar1n64x5 hold122 (.clk(n2896),
    .clkout(net1878));
 b15cbf034ar1n64x5 hold123 (.clk(net133),
    .clkout(net1879));
 b15cbf034ar1n64x5 hold124 (.clk(gpio_2_xbar[6]),
    .clkout(net1880));
 b15cbf034ar1n64x5 hold125 (.clk(n3051),
    .clkout(net1881));
 b15cbf034ar1n64x5 hold126 (.clk(gpio_2_xbar[1]),
    .clkout(net1882));
 b15cbf034ar1n64x5 hold127 (.clk(n3070),
    .clkout(net1883));
 b15cbf034ar1n64x5 hold128 (.clk(gpio_2_xbar[23]),
    .clkout(net1884));
 b15cbf034ar1n64x5 hold129 (.clk(n3073),
    .clkout(net1885));
 b15cbf034ar1n64x5 hold130 (.clk(gpio_2_xbar[19]),
    .clkout(net1886));
 b15cbf034ar1n64x5 hold131 (.clk(net1869),
    .clkout(net1887));
 b15cbf034ar1n64x5 hold132 (.clk(gpio_2_xbar[20]),
    .clkout(net1888));
 b15cbf034ar1n64x5 hold133 (.clk(n3076),
    .clkout(net1889));
 b15cbf034ar1n64x5 hold134 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[19]),
    .clkout(net1890));
 b15cbf034ar1n64x5 hold135 (.clk(n2922),
    .clkout(net1891));
 b15cbf034ar1n64x5 hold136 (.clk(net114),
    .clkout(net1892));
 b15cbf034ar1n64x5 hold137 (.clk(gpio_2_xbar[3]),
    .clkout(net1893));
 b15cbf034ar1n64x5 hold138 (.clk(n3068),
    .clkout(net1894));
 b15cbf034ar1n64x5 hold139 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[23]),
    .clkout(net1895));
 b15cbf034ar1n64x5 hold140 (.clk(net167),
    .clkout(net1896));
 b15cbf034ar1n64x5 hold141 (.clk(gpio_2_xbar[8]),
    .clkout(net1897));
 b15cbf034ar1n64x5 hold142 (.clk(n3102),
    .clkout(net1898));
 b15cbf034ar1n64x5 hold143 (.clk(gpio_2_xbar[18]),
    .clkout(net1899));
 b15cbf034ar1n64x5 hold144 (.clk(n3078),
    .clkout(net1900));
 b15cbf034ar1n64x5 hold145 (.clk(gpio_2_xbar[2]),
    .clkout(net1901));
 b15cbf034ar1n64x5 hold146 (.clk(gpio_2_xbar[7]),
    .clkout(net1902));
 b15cbf034ar1n64x5 hold147 (.clk(n3090),
    .clkout(net1903));
 b15cbf034ar1n64x5 hold148 (.clk(gpio_2_xbar[26]),
    .clkout(net1904));
 b15cbf034ar1n64x5 hold149 (.clk(n3092),
    .clkout(net1905));
 b15cbf034ar1n64x5 hold150 (.clk(gpio_2_xbar[12]),
    .clkout(net1906));
 b15cbf034ar1n64x5 hold151 (.clk(n3099),
    .clkout(net1907));
 b15cbf034ar1n64x5 hold152 (.clk(gpio_2_xbar[27]),
    .clkout(net1908));
 b15cbf034ar1n64x5 hold153 (.clk(n3091),
    .clkout(net1909));
 b15cbf034ar1n64x5 hold154 (.clk(gpio_2_xbar[9]),
    .clkout(net1910));
 b15cbf034ar1n64x5 hold155 (.clk(net1928),
    .clkout(net1911));
 b15cbf034ar1n64x5 hold156 (.clk(n3084),
    .clkout(net1912));
 b15cbf034ar1n64x5 hold157 (.clk(gpio_2_xbar[10]),
    .clkout(net1913));
 b15cbf034ar1n64x5 hold158 (.clk(n3100),
    .clkout(net1914));
 b15cbf034ar1n64x5 hold159 (.clk(net2223),
    .clkout(net1915));
 b15cbf034ar1n64x5 hold160 (.clk(n3617),
    .clkout(net1916));
 b15cbf034ar1n64x5 hold161 (.clk(net122),
    .clkout(net1917));
 b15cbf034ar1n64x5 hold162 (.clk(gpio_2_xbar[28]),
    .clkout(net1918));
 b15cbf034ar1n64x5 hold163 (.clk(n3023),
    .clkout(net1919));
 b15cbf034ar1n64x5 hold164 (.clk(net171),
    .clkout(net1920));
 b15cbf034ar1n64x5 hold165 (.clk(gpio_2_xbar[22]),
    .clkout(net1921));
 b15cbf034ar1n64x5 hold166 (.clk(n3060),
    .clkout(net1922));
 b15cbf034ar1n64x5 hold167 (.clk(n3066),
    .clkout(net1923));
 b15cbf034ar1n64x5 hold168 (.clk(net169),
    .clkout(net1924));
 b15cbf034ar1n64x5 hold169 (.clk(gpio_2_xbar[21]),
    .clkout(net1925));
 b15cbf034ar1n64x5 hold170 (.clk(n3003),
    .clkout(net1926));
 b15cbf034ar1n64x5 hold171 (.clk(net154),
    .clkout(net1927));
 b15cbf034ar1n64x5 hold172 (.clk(gpio_2_xbar[13]),
    .clkout(net1928));
 b15cbf034ar1n64x5 hold173 (.clk(n2949),
    .clkout(net1929));
 b15cbf034ar1n64x5 hold174 (.clk(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_intq_0_),
    .clkout(net1930));
 b15cbf034ar1n64x5 hold175 (.clk(u_gpio_gen_filter_21__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1931));
 b15cbf034ar1n64x5 hold176 (.clk(u_gpio_gen_filter_28__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1932));
 b15cbf034ar1n64x5 hold177 (.clk(u_gpio_gen_filter_31__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1933));
 b15cbf034ar1n64x5 hold178 (.clk(u_gpio_gen_filter_8__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1934));
 b15cbf034ar1n64x5 hold179 (.clk(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_intq_0_),
    .clkout(net1935));
 b15cbf034ar1n64x5 hold180 (.clk(u_gpio_gen_filter_27__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1936));
 b15cbf034ar1n64x5 hold181 (.clk(u_gpio_gen_filter_13__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1937));
 b15cbf034ar1n64x5 hold182 (.clk(u_gpio_gen_filter_6__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1938));
 b15cbf034ar1n64x5 hold183 (.clk(u_gpio_gen_filter_30__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1939));
 b15cbf034ar1n64x5 hold184 (.clk(u_gpio_gen_filter_17__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1940));
 b15cbf034ar1n64x5 hold185 (.clk(u_gpio_gen_filter_11__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1941));
 b15cbf034ar1n64x5 hold186 (.clk(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_intq_0_),
    .clkout(net1942));
 b15cbf034ar1n64x5 hold187 (.clk(u_gpio_gen_filter_26__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1943));
 b15cbf034ar1n64x5 hold188 (.clk(u_gpio_gen_filter_4__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1944));
 b15cbf034ar1n64x5 hold189 (.clk(u_gpio_gen_filter_2__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1945));
 b15cbf034ar1n64x5 hold190 (.clk(u_gpio_data_in_q[28]),
    .clkout(net1946));
 b15cbf034ar1n64x5 hold191 (.clk(u_gpio_gen_filter_10__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1947));
 b15cbf034ar1n64x5 hold192 (.clk(u_gpio_reg2hw[14]),
    .clkout(net1948));
 b15cbf034ar1n64x5 hold193 (.clk(u_gpio_gen_filter_29__u_filter_filter_q),
    .clkout(net1949));
 b15cbf034ar1n64x5 hold194 (.clk(u_gpio_gen_filter_29__u_filter_diff_ctr_d[2]),
    .clkout(net1950));
 b15cbf034ar1n64x5 hold195 (.clk(u_gpio_data_in_q[24]),
    .clkout(net1951));
 b15cbf034ar1n64x5 hold196 (.clk(u_gpio_gen_filter_29__u_filter_diff_ctr_q[1]),
    .clkout(net1952));
 b15cbf034ar1n64x5 hold197 (.clk(n2859),
    .clkout(net1953));
 b15cbf034ar1n64x5 hold198 (.clk(u_gpio_gen_filter_29__u_filter_diff_ctr_d[3]),
    .clkout(net1954));
 b15cbf034ar1n64x5 hold199 (.clk(u_gpio_gen_filter_20__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1955));
 b15cbf034ar1n64x5 hold200 (.clk(u_gpio_gen_filter_28__u_filter_filter_q),
    .clkout(net1956));
 b15cbf034ar1n64x5 hold201 (.clk(u_gpio_gen_filter_28__u_filter_diff_ctr_d[0]),
    .clkout(net1957));
 b15cbf034ar1n64x5 hold202 (.clk(u_gpio_gen_filter_5__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1958));
 b15cbf034ar1n64x5 hold203 (.clk(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nd),
    .clkout(net1959));
 b15cbf034ar1n64x5 hold204 (.clk(u_gpio_gen_filter_3__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1960));
 b15cbf034ar1n64x5 hold205 (.clk(u_gpio_gen_filter_24__u_filter_filter_synced),
    .clkout(net1961));
 b15cbf034ar1n64x5 hold206 (.clk(u_gpio_gen_filter_1__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1962));
 b15cbf034ar1n64x5 hold207 (.clk(u_gpio_gen_filter_10__u_filter_stored_value_q),
    .clkout(net1963));
 b15cbf034ar1n64x5 hold208 (.clk(net105),
    .clkout(net1964));
 b15cbf034ar1n64x5 hold209 (.clk(u_gpio_data_in_q[29]),
    .clkout(net1965));
 b15cbf034ar1n64x5 hold210 (.clk(n3593),
    .clkout(net1966));
 b15cbf034ar1n64x5 hold211 (.clk(u_gpio_u_reg_u_intr_state_wr_data[29]),
    .clkout(net1967));
 b15cbf034ar1n64x5 hold212 (.clk(u_gpio_gen_filter_28__u_filter_diff_ctr_q[3]),
    .clkout(net1968));
 b15cbf034ar1n64x5 hold213 (.clk(u_gpio_data_in_q[22]),
    .clkout(net1969));
 b15cbf034ar1n64x5 hold214 (.clk(n3594),
    .clkout(net1970));
 b15cbf034ar1n64x5 hold215 (.clk(u_gpio_gen_filter_23__u_filter_diff_ctr_q[0]),
    .clkout(net1971));
 b15cbf034ar1n64x5 hold216 (.clk(u_gpio_gen_filter_23__u_filter_diff_ctr_d[0]),
    .clkout(net1972));
 b15cbf034ar1n64x5 hold217 (.clk(u_gpio_gen_filter_18__u_filter_diff_ctr_q[0]),
    .clkout(net1973));
 b15cbf034ar1n64x5 hold218 (.clk(u_gpio_gen_filter_18__u_filter_diff_ctr_d[0]),
    .clkout(net1974));
 b15cbf034ar1n64x5 hold219 (.clk(u_gpio_gen_filter_2__u_filter_diff_ctr_q[0]),
    .clkout(net1975));
 b15cbf034ar1n64x5 hold220 (.clk(u_gpio_gen_filter_2__u_filter_diff_ctr_d[0]),
    .clkout(net1976));
 b15cbf034ar1n64x5 hold221 (.clk(u_gpio_gen_filter_17__u_filter_diff_ctr_q[0]),
    .clkout(net1977));
 b15cbf034ar1n64x5 hold222 (.clk(u_gpio_gen_filter_17__u_filter_diff_ctr_d[1]),
    .clkout(net1978));
 b15cbf034ar1n64x5 hold223 (.clk(u_gpio_gen_filter_15__u_filter_filter_synced),
    .clkout(net1979));
 b15cbf034ar1n64x5 hold224 (.clk(u_gpio_data_in_q[25]),
    .clkout(net1980));
 b15cbf034ar1n64x5 hold225 (.clk(n3589),
    .clkout(net1981));
 b15cbf034ar1n64x5 hold226 (.clk(u_gpio_gen_filter_3__u_filter_diff_ctr_q[2]),
    .clkout(net1982));
 b15cbf034ar1n64x5 hold227 (.clk(n2853),
    .clkout(net1983));
 b15cbf034ar1n64x5 hold228 (.clk(u_gpio_gen_filter_3__u_filter_diff_ctr_d[3]),
    .clkout(net1984));
 b15cbf034ar1n64x5 hold229 (.clk(net92),
    .clkout(net1985));
 b15cbf034ar1n64x5 hold230 (.clk(u_gpio_reg2hw[12]),
    .clkout(net1986));
 b15cbf034ar1n64x5 hold231 (.clk(u_gpio_gen_filter_23__u_filter_filter_q),
    .clkout(net1987));
 b15cbf034ar1n64x5 hold232 (.clk(u_gpio_gen_filter_23__u_filter_diff_ctr_d[3]),
    .clkout(net1988));
 b15cbf034ar1n64x5 hold233 (.clk(u_gpio_gen_filter_12__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net1989));
 b15cbf034ar1n64x5 hold234 (.clk(u_gpio_u_reg_err_q),
    .clkout(net1990));
 b15cbf034ar1n64x5 hold235 (.clk(u_gpio_gen_filter_0__u_filter_filter_q),
    .clkout(net1991));
 b15cbf034ar1n64x5 hold236 (.clk(u_gpio_gen_filter_0__u_filter_diff_ctr_d[3]),
    .clkout(net1992));
 b15cbf034ar1n64x5 hold237 (.clk(u_gpio_gen_filter_22__u_filter_diff_ctr_q[3]),
    .clkout(net1993));
 b15cbf034ar1n64x5 hold238 (.clk(n2886),
    .clkout(net1994));
 b15cbf034ar1n64x5 hold239 (.clk(u_gpio_gen_filter_22__u_filter_diff_ctr_d[2]),
    .clkout(net1995));
 b15cbf034ar1n64x5 hold240 (.clk(u_gpio_gen_filter_13__u_filter_diff_ctr_q[3]),
    .clkout(net1996));
 b15cbf034ar1n64x5 hold241 (.clk(u_gpio_gen_filter_13__u_filter_diff_ctr_d[3]),
    .clkout(net1997));
 b15cbf034ar1n64x5 hold242 (.clk(u_gpio_gen_filter_19__u_filter_filter_synced),
    .clkout(net1998));
 b15cbf034ar1n64x5 hold243 (.clk(u_gpio_u_reg_data_in_qs[8]),
    .clkout(net1999));
 b15cbf034ar1n64x5 hold244 (.clk(u_gpio_gen_filter_18__u_filter_filter_q),
    .clkout(net2000));
 b15cbf034ar1n64x5 hold245 (.clk(u_gpio_gen_filter_18__u_filter_diff_ctr_d[1]),
    .clkout(net2001));
 b15cbf034ar1n64x5 hold246 (.clk(u_gpio_gen_filter_1__u_filter_stored_value_q),
    .clkout(net2002));
 b15cbf034ar1n64x5 hold247 (.clk(u_gpio_gen_filter_22__u_filter_filter_q),
    .clkout(net2003));
 b15cbf034ar1n64x5 hold248 (.clk(u_gpio_gen_filter_0__u_filter_diff_ctr_q[2]),
    .clkout(net2004));
 b15cbf034ar1n64x5 hold249 (.clk(u_gpio_gen_filter_0__u_filter_diff_ctr_d[2]),
    .clkout(net2005));
 b15cbf034ar1n64x5 hold250 (.clk(u_gpio_gen_filter_15__u_filter_diff_ctr_q[0]),
    .clkout(net2006));
 b15cbf034ar1n64x5 hold251 (.clk(u_gpio_gen_filter_15__u_filter_diff_ctr_d[0]),
    .clkout(net2007));
 b15cbf034ar1n64x5 hold252 (.clk(u_gpio_gen_filter_6__u_filter_filter_q),
    .clkout(net2008));
 b15cbf034ar1n64x5 hold253 (.clk(n2739),
    .clkout(net2009));
 b15cbf034ar1n64x5 hold254 (.clk(u_gpio_gen_filter_25__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2010));
 b15cbf034ar1n64x5 hold255 (.clk(u_gpio_gen_filter_23__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2011));
 b15cbf034ar1n64x5 hold256 (.clk(u_gpio_data_in_q[17]),
    .clkout(net2012));
 b15cbf034ar1n64x5 hold257 (.clk(n3590),
    .clkout(net2013));
 b15cbf034ar1n64x5 hold258 (.clk(u_gpio_gen_filter_11__u_filter_filter_q),
    .clkout(net2014));
 b15cbf034ar1n64x5 hold259 (.clk(u_gpio_gen_filter_11__u_filter_diff_ctr_d[2]),
    .clkout(net2015));
 b15cbf034ar1n64x5 hold260 (.clk(u_gpio_gen_filter_16__u_filter_diff_ctr_q[2]),
    .clkout(net2016));
 b15cbf034ar1n64x5 hold261 (.clk(n2784),
    .clkout(net2017));
 b15cbf034ar1n64x5 hold262 (.clk(u_gpio_gen_filter_16__u_filter_diff_ctr_d[1]),
    .clkout(net2018));
 b15cbf034ar1n64x5 hold263 (.clk(u_gpio_gen_filter_11__u_filter_diff_ctr_q[3]),
    .clkout(net2019));
 b15cbf034ar1n64x5 hold264 (.clk(net100),
    .clkout(net2020));
 b15cbf034ar1n64x5 hold265 (.clk(u_gpio_gen_filter_9__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2021));
 b15cbf034ar1n64x5 hold266 (.clk(u_gpio_gen_filter_27__u_filter_filter_q),
    .clkout(net2022));
 b15cbf034ar1n64x5 hold267 (.clk(u_gpio_gen_filter_27__u_filter_diff_ctr_d[2]),
    .clkout(net2023));
 b15cbf034ar1n64x5 hold268 (.clk(u_gpio_data_in_q[15]),
    .clkout(net2024));
 b15cbf034ar1n64x5 hold269 (.clk(u_gpio_gen_filter_18__u_filter_diff_ctr_q[3]),
    .clkout(net2025));
 b15cbf034ar1n64x5 hold270 (.clk(u_gpio_gen_filter_18__u_filter_diff_ctr_d[3]),
    .clkout(net2026));
 b15cbf034ar1n64x5 hold271 (.clk(u_gpio_gen_filter_16__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2027));
 b15cbf034ar1n64x5 hold272 (.clk(u_gpio_gen_filter_8__u_filter_filter_q),
    .clkout(net2028));
 b15cbf034ar1n64x5 hold273 (.clk(u_gpio_gen_alert_tx_0__u_prim_alert_sender_ping_set_q),
    .clkout(net2029));
 b15cbf034ar1n64x5 hold274 (.clk(u_gpio_gen_filter_25__u_filter_filter_q),
    .clkout(net2030));
 b15cbf034ar1n64x5 hold275 (.clk(u_gpio_gen_filter_25__u_filter_diff_ctr_d[0]),
    .clkout(net2031));
 b15cbf034ar1n64x5 hold276 (.clk(u_gpio_gen_filter_25__u_filter_diff_ctr_q[2]),
    .clkout(net2032));
 b15cbf034ar1n64x5 hold277 (.clk(n2797),
    .clkout(net2033));
 b15cbf034ar1n64x5 hold278 (.clk(u_gpio_gen_filter_25__u_filter_diff_ctr_d[2]),
    .clkout(net2034));
 b15cbf034ar1n64x5 hold279 (.clk(u_gpio_gen_filter_18__u_filter_diff_ctr_q[0]),
    .clkout(net2035));
 b15cbf034ar1n64x5 hold280 (.clk(u_gpio_gen_filter_14__u_filter_diff_ctr_q[0]),
    .clkout(net2036));
 b15cbf034ar1n64x5 hold281 (.clk(u_gpio_gen_filter_14__u_filter_diff_ctr_d[0]),
    .clkout(net2037));
 b15cbf034ar1n64x5 hold282 (.clk(u_gpio_gen_filter_16__u_filter_diff_ctr_q[0]),
    .clkout(net2038));
 b15cbf034ar1n64x5 hold283 (.clk(u_gpio_gen_filter_16__u_filter_diff_ctr_d[0]),
    .clkout(net2039));
 b15cbf034ar1n64x5 hold284 (.clk(u_gpio_gen_filter_9__u_filter_filter_q),
    .clkout(net2040));
 b15cbf034ar1n64x5 hold285 (.clk(u_gpio_gen_filter_9__u_filter_diff_ctr_d[1]),
    .clkout(net2041));
 b15cbf034ar1n64x5 hold286 (.clk(u_gpio_gen_filter_4__u_filter_stored_value_q),
    .clkout(net2042));
 b15cbf034ar1n64x5 hold287 (.clk(u_gpio_u_reg_u_data_in_wr_data[4]),
    .clkout(net2043));
 b15cbf034ar1n64x5 hold288 (.clk(u_gpio_gen_filter_19__u_filter_diff_ctr_q[2]),
    .clkout(net2044));
 b15cbf034ar1n64x5 hold289 (.clk(n2712),
    .clkout(net2045));
 b15cbf034ar1n64x5 hold290 (.clk(u_gpio_gen_filter_19__u_filter_diff_ctr_d[2]),
    .clkout(net2046));
 b15cbf034ar1n64x5 hold291 (.clk(u_gpio_gen_filter_4__u_filter_filter_synced),
    .clkout(net2047));
 b15cbf034ar1n64x5 hold292 (.clk(u_gpio_gen_filter_7__u_filter_filter_q),
    .clkout(net2048));
 b15cbf034ar1n64x5 hold293 (.clk(u_gpio_gen_filter_23__u_filter_diff_ctr_q[2]),
    .clkout(net2049));
 b15cbf034ar1n64x5 hold294 (.clk(n2631),
    .clkout(net2050));
 b15cbf034ar1n64x5 hold295 (.clk(u_gpio_gen_filter_13__u_filter_diff_ctr_q[2]),
    .clkout(net2051));
 b15cbf034ar1n64x5 hold296 (.clk(net102),
    .clkout(net2052));
 b15cbf034ar1n64x5 hold297 (.clk(net107),
    .clkout(net2053));
 b15cbf034ar1n64x5 hold298 (.clk(u_gpio_gen_filter_4__u_filter_diff_ctr_q[3]),
    .clkout(net2054));
 b15cbf034ar1n64x5 hold299 (.clk(u_gpio_gen_filter_4__u_filter_diff_ctr_d[2]),
    .clkout(net2055));
 b15cbf034ar1n64x5 hold300 (.clk(u_gpio_gen_filter_13__u_filter_filter_q),
    .clkout(net2056));
 b15cbf034ar1n64x5 hold301 (.clk(u_gpio_gen_filter_17__u_filter_diff_ctr_q[2]),
    .clkout(net2057));
 b15cbf034ar1n64x5 hold302 (.clk(n2805),
    .clkout(net2058));
 b15cbf034ar1n64x5 hold303 (.clk(u_gpio_gen_filter_17__u_filter_diff_ctr_d[2]),
    .clkout(net2059));
 b15cbf034ar1n64x5 hold304 (.clk(u_gpio_data_in_q[18]),
    .clkout(net2060));
 b15cbf034ar1n64x5 hold305 (.clk(u_gpio_gen_filter_12__u_filter_diff_ctr_q[3]),
    .clkout(net2061));
 b15cbf034ar1n64x5 hold306 (.clk(u_gpio_gen_filter_12__u_filter_diff_ctr_d[2]),
    .clkout(net2062));
 b15cbf034ar1n64x5 hold307 (.clk(u_gpio_gen_filter_16__u_filter_filter_q),
    .clkout(net2063));
 b15cbf034ar1n64x5 hold308 (.clk(u_gpio_gen_filter_16__u_filter_diff_ctr_d[2]),
    .clkout(net2064));
 b15cbf034ar1n64x5 hold309 (.clk(u_gpio_gen_filter_12__u_filter_diff_ctr_q[2]),
    .clkout(net2065));
 b15cbf034ar1n64x5 hold310 (.clk(u_gpio_gen_filter_12__u_filter_diff_ctr_d[1]),
    .clkout(net2066));
 b15cbf034ar1n64x5 hold311 (.clk(u_gpio_gen_filter_19__u_filter_filter_q),
    .clkout(net2067));
 b15cbf034ar1n64x5 hold312 (.clk(u_gpio_gen_filter_19__u_filter_diff_ctr_d[0]),
    .clkout(net2068));
 b15cbf034ar1n64x5 hold313 (.clk(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd),
    .clkout(net2069));
 b15cbf034ar1n64x5 hold314 (.clk(u_gpio_gen_filter_24__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2070));
 b15cbf034ar1n64x5 hold315 (.clk(u_gpio_gen_filter_15__u_filter_filter_q),
    .clkout(net2071));
 b15cbf034ar1n64x5 hold316 (.clk(u_gpio_gen_filter_15__u_filter_diff_ctr_d[3]),
    .clkout(net2072));
 b15cbf034ar1n64x5 hold317 (.clk(u_gpio_gen_filter_9__u_filter_diff_ctr_q[3]),
    .clkout(net2073));
 b15cbf034ar1n64x5 hold318 (.clk(u_gpio_gen_filter_5__u_filter_filter_q),
    .clkout(net2074));
 b15cbf034ar1n64x5 hold319 (.clk(u_gpio_gen_filter_5__u_filter_diff_ctr_d[1]),
    .clkout(net2075));
 b15cbf034ar1n64x5 hold320 (.clk(u_gpio_data_in_q[14]),
    .clkout(net2076));
 b15cbf034ar1n64x5 hold321 (.clk(u_gpio_gen_filter_30__u_filter_stored_value_q),
    .clkout(net2077));
 b15cbf034ar1n64x5 hold322 (.clk(u_gpio_gen_filter_19__u_filter_diff_ctr_q[3]),
    .clkout(net2078));
 b15cbf034ar1n64x5 hold323 (.clk(u_gpio_gen_filter_10__u_filter_diff_ctr_q[0]),
    .clkout(net2079));
 b15cbf034ar1n64x5 hold324 (.clk(u_gpio_gen_filter_10__u_filter_diff_ctr_d[0]),
    .clkout(net2080));
 b15cbf034ar1n64x5 hold325 (.clk(u_gpio_data_in_q[2]),
    .clkout(net2081));
 b15cbf034ar1n64x5 hold326 (.clk(n3588),
    .clkout(net2082));
 b15cbf034ar1n64x5 hold327 (.clk(u_gpio_gen_filter_25__u_filter_diff_ctr_q[3]),
    .clkout(net2083));
 b15cbf034ar1n64x5 hold328 (.clk(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q),
    .clkout(net2084));
 b15cbf034ar1n64x5 hold329 (.clk(u_gpio_gen_filter_13__u_filter_diff_ctr_q[0]),
    .clkout(net2085));
 b15cbf034ar1n64x5 hold330 (.clk(u_gpio_gen_filter_7__u_filter_filter_synced),
    .clkout(net2086));
 b15cbf034ar1n64x5 hold331 (.clk(net93),
    .clkout(net2087));
 b15cbf034ar1n64x5 hold332 (.clk(u_gpio_gen_filter_29__u_filter_diff_ctr_q[0]),
    .clkout(net2088));
 b15cbf034ar1n64x5 hold333 (.clk(u_gpio_gen_filter_23__u_filter_diff_ctr_q[0]),
    .clkout(net2089));
 b15cbf034ar1n64x5 hold334 (.clk(u_gpio_gen_filter_17__u_filter_diff_ctr_q[3]),
    .clkout(net2090));
 b15cbf034ar1n64x5 hold335 (.clk(u_gpio_gen_filter_17__u_filter_diff_ctr_d[3]),
    .clkout(net2091));
 b15cbf034ar1n64x5 hold336 (.clk(u_gpio_gen_filter_21__u_filter_diff_ctr_q[0]),
    .clkout(net2092));
 b15cbf034ar1n64x5 hold337 (.clk(u_gpio_gen_filter_21__u_filter_diff_ctr_d[0]),
    .clkout(net2093));
 b15cbf034ar1n64x5 hold338 (.clk(u_gpio_gen_filter_6__u_filter_filter_synced),
    .clkout(net2094));
 b15cbf034ar1n64x5 hold339 (.clk(net94),
    .clkout(net2095));
 b15cbf034ar1n64x5 hold340 (.clk(u_gpio_gen_filter_29__u_filter_diff_ctr_q[1]),
    .clkout(net2096));
 b15cbf034ar1n64x5 hold341 (.clk(net106),
    .clkout(net2097));
 b15cbf034ar1n64x5 hold342 (.clk(u_gpio_gen_filter_5__u_filter_diff_ctr_q[2]),
    .clkout(net2098));
 b15cbf034ar1n64x5 hold343 (.clk(u_gpio_gen_filter_5__u_filter_diff_ctr_d[2]),
    .clkout(net2099));
 b15cbf034ar1n64x5 hold344 (.clk(u_gpio_gen_filter_20__u_filter_filter_q),
    .clkout(net2100));
 b15cbf034ar1n64x5 hold345 (.clk(u_gpio_gen_filter_20__u_filter_diff_ctr_d[1]),
    .clkout(net2101));
 b15cbf034ar1n64x5 hold346 (.clk(u_gpio_gen_filter_1__u_filter_diff_ctr_q[3]),
    .clkout(net2102));
 b15cbf034ar1n64x5 hold347 (.clk(net101),
    .clkout(net2103));
 b15cbf034ar1n64x5 hold348 (.clk(u_gpio_data_in_q[8]),
    .clkout(net2104));
 b15cbf034ar1n64x5 hold349 (.clk(u_gpio_gen_filter_14__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2105));
 b15cbf034ar1n64x5 hold350 (.clk(net95),
    .clkout(net2106));
 b15cbf034ar1n64x5 hold351 (.clk(u_gpio_gen_filter_25__u_filter_diff_ctr_q[1]),
    .clkout(net2107));
 b15cbf034ar1n64x5 hold352 (.clk(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_intq_0_),
    .clkout(net2108));
 b15cbf034ar1n64x5 hold353 (.clk(u_gpio_gen_filter_3__u_filter_diff_ctr_q[0]),
    .clkout(net2109));
 b15cbf034ar1n64x5 hold354 (.clk(u_gpio_u_reg_data_in_qs[3]),
    .clkout(net2110));
 b15cbf034ar1n64x5 hold355 (.clk(u_gpio_gen_filter_11__u_filter_diff_ctr_q[0]),
    .clkout(net2111));
 b15cbf034ar1n64x5 hold356 (.clk(u_gpio_gen_filter_31__u_filter_diff_ctr_q[3]),
    .clkout(net2112));
 b15cbf034ar1n64x5 hold357 (.clk(u_gpio_gen_filter_24__u_filter_diff_ctr_q[2]),
    .clkout(net2113));
 b15cbf034ar1n64x5 hold358 (.clk(u_gpio_gen_filter_5__u_filter_diff_ctr_q[3]),
    .clkout(net2114));
 b15cbf034ar1n64x5 hold359 (.clk(u_gpio_data_in_q[20]),
    .clkout(net2115));
 b15cbf034ar1n64x5 hold360 (.clk(n3567),
    .clkout(net2116));
 b15cbf034ar1n64x5 hold361 (.clk(u_gpio_gen_filter_15__u_filter_diff_ctr_q[1]),
    .clkout(net2117));
 b15cbf034ar1n64x5 hold362 (.clk(n2676),
    .clkout(net2118));
 b15cbf034ar1n64x5 hold363 (.clk(u_gpio_gen_filter_22__u_filter_filter_synced),
    .clkout(net2119));
 b15cbf034ar1n64x5 hold364 (.clk(u_gpio_reg2hw[222]),
    .clkout(net2120));
 b15cbf034ar1n64x5 hold365 (.clk(net82),
    .clkout(net2121));
 b15cbf034ar1n64x5 hold366 (.clk(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .clkout(net2122));
 b15cbf034ar1n64x5 hold367 (.clk(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_n5),
    .clkout(net2123));
 b15cbf034ar1n64x5 hold368 (.clk(u_gpio_gen_filter_11__u_filter_stored_value_q),
    .clkout(net2124));
 b15cbf034ar1n64x5 hold369 (.clk(u_gpio_u_reg_masked_oe_upper_data_qs[9]),
    .clkout(net2125));
 b15cbf034ar1n64x5 hold370 (.clk(net89),
    .clkout(net2126));
 b15cbf034ar1n64x5 hold371 (.clk(u_gpio_reg2hw[13]),
    .clkout(net2127));
 b15cbf034ar1n64x5 hold372 (.clk(u_gpio_gen_filter_22__u_filter_diff_ctr_q[1]),
    .clkout(net2128));
 b15cbf034ar1n64x5 hold373 (.clk(u_gpio_gen_filter_4__u_filter_filter_q),
    .clkout(net2129));
 b15cbf034ar1n64x5 hold374 (.clk(u_gpio_gen_filter_15__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2130));
 b15cbf034ar1n64x5 hold375 (.clk(u_gpio_gen_filter_20__u_filter_diff_ctr_q[3]),
    .clkout(net2131));
 b15cbf034ar1n64x5 hold376 (.clk(u_gpio_gen_filter_20__u_filter_diff_ctr_q[0]),
    .clkout(net2132));
 b15cbf034ar1n64x5 hold377 (.clk(u_gpio_gen_filter_16__u_filter_diff_ctr_q[3]),
    .clkout(net2133));
 b15cbf034ar1n64x5 hold378 (.clk(u_gpio_data_in_q[1]),
    .clkout(net2134));
 b15cbf034ar1n64x5 hold379 (.clk(u_gpio_gen_filter_31__u_filter_diff_ctr_q[0]),
    .clkout(net2135));
 b15cbf034ar1n64x5 hold380 (.clk(u_gpio_gen_filter_0__u_filter_diff_ctr_q[1]),
    .clkout(net2136));
 b15cbf034ar1n64x5 hold381 (.clk(u_gpio_data_in_q[19]),
    .clkout(net2137));
 b15cbf034ar1n64x5 hold382 (.clk(u_gpio_gen_filter_30__u_filter_diff_ctr_q[2]),
    .clkout(net2138));
 b15cbf034ar1n64x5 hold383 (.clk(n2770),
    .clkout(net2139));
 b15cbf034ar1n64x5 hold384 (.clk(u_gpio_gen_filter_30__u_filter_diff_ctr_d[1]),
    .clkout(net2140));
 b15cbf034ar1n64x5 hold385 (.clk(u_gpio_reg2hw[1]),
    .clkout(net2141));
 b15cbf034ar1n64x5 hold386 (.clk(u_gpio_gen_filter_0__u_filter_stored_value_q),
    .clkout(net2142));
 b15cbf034ar1n64x5 hold387 (.clk(u_gpio_gen_filter_24__u_filter_diff_ctr_q[0]),
    .clkout(net2143));
 b15cbf034ar1n64x5 hold388 (.clk(u_gpio_gen_filter_24__u_filter_diff_ctr_d[0]),
    .clkout(net2144));
 b15cbf034ar1n64x5 hold389 (.clk(u_gpio_gen_filter_26__u_filter_stored_value_q),
    .clkout(net2145));
 b15cbf034ar1n64x5 hold390 (.clk(u_gpio_u_reg_masked_oe_upper_data_qs[10]),
    .clkout(net2146));
 b15cbf034ar1n64x5 hold391 (.clk(u_xbar_periph_u_s1n_6_num_req_outstanding[8]),
    .clkout(net2147));
 b15cbf034ar1n64x5 hold392 (.clk(u_xbar_periph_u_s1n_6_num_req_outstanding[4]),
    .clkout(net2148));
 b15cbf034ar1n64x5 hold393 (.clk(u_gpio_gen_filter_27__u_filter_stored_value_q),
    .clkout(net2149));
 b15cbf034ar1n64x5 hold394 (.clk(u_gpio_data_in_q[23]),
    .clkout(net2150));
 b15cbf034ar1n64x5 hold395 (.clk(n3574),
    .clkout(net2151));
 b15cbf034ar1n64x5 hold396 (.clk(u_gpio_gen_filter_19__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2152));
 b15cbf034ar1n64x5 hold397 (.clk(u_gpio_reg2hw[198]),
    .clkout(net2153));
 b15cbf034ar1n64x5 hold398 (.clk(u_gpio_u_reg_u_intr_state_wr_data[6]),
    .clkout(net2154));
 b15cbf034ar1n64x5 hold399 (.clk(u_gpio_data_in_q[9]),
    .clkout(net2155));
 b15cbf034ar1n64x5 hold400 (.clk(u_gpio_gen_filter_14__u_filter_filter_synced),
    .clkout(net2156));
 b15cbf034ar1n64x5 hold401 (.clk(u_gpio_gen_filter_30__u_filter_filter_q),
    .clkout(net2157));
 b15cbf034ar1n64x5 hold402 (.clk(net104),
    .clkout(net2158));
 b15cbf034ar1n64x5 hold403 (.clk(u_gpio_gen_filter_30__u_filter_diff_ctr_q[3]),
    .clkout(net2159));
 b15cbf034ar1n64x5 hold404 (.clk(u_xbar_periph_u_s1n_6_num_req_outstanding[2]),
    .clkout(net2160));
 b15cbf034ar1n64x5 hold405 (.clk(u_gpio_u_reg_data_in_qs[26]),
    .clkout(net2161));
 b15cbf034ar1n64x5 hold406 (.clk(u_gpio_gen_filter_23__u_filter_filter_synced),
    .clkout(net2162));
 b15cbf034ar1n64x5 hold407 (.clk(u_gpio_gen_filter_10__u_filter_diff_ctr_q[0]),
    .clkout(net2163));
 b15cbf034ar1n64x5 hold408 (.clk(n2720),
    .clkout(net2164));
 b15cbf034ar1n64x5 hold409 (.clk(u_gpio_gen_filter_10__u_filter_diff_ctr_d[3]),
    .clkout(net2165));
 b15cbf034ar1n64x5 hold410 (.clk(u_gpio_gen_filter_7__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2166));
 b15cbf034ar1n64x5 hold411 (.clk(u_gpio_gen_filter_14__u_filter_filter_q),
    .clkout(net2167));
 b15cbf034ar1n64x5 hold412 (.clk(u_gpio_gen_filter_14__u_filter_diff_ctr_d[3]),
    .clkout(net2168));
 b15cbf034ar1n64x5 hold413 (.clk(u_gpio_gen_filter_2__u_filter_diff_ctr_q[3]),
    .clkout(net2169));
 b15cbf034ar1n64x5 hold414 (.clk(u_gpio_gen_filter_5__u_filter_filter_synced),
    .clkout(net2170));
 b15cbf034ar1n64x5 hold415 (.clk(u_gpio_gen_filter_3__u_filter_diff_ctr_q[1]),
    .clkout(net2171));
 b15cbf034ar1n64x5 hold416 (.clk(n2851),
    .clkout(net2172));
 b15cbf034ar1n64x5 hold417 (.clk(u_gpio_gen_filter_3__u_filter_diff_ctr_d[1]),
    .clkout(net2173));
 b15cbf034ar1n64x5 hold418 (.clk(u_gpio_gen_filter_26__u_filter_diff_ctr_q[2]),
    .clkout(net2174));
 b15cbf034ar1n64x5 hold419 (.clk(u_gpio_gen_filter_26__u_filter_diff_ctr_d[3]),
    .clkout(net2175));
 b15cbf034ar1n64x5 hold420 (.clk(u_gpio_data_in_q[27]),
    .clkout(net2176));
 b15cbf034ar1n64x5 hold421 (.clk(u_gpio_data_in_q[16]),
    .clkout(net2177));
 b15cbf034ar1n64x5 hold422 (.clk(net97),
    .clkout(net2178));
 b15cbf034ar1n64x5 hold423 (.clk(u_gpio_u_reg_data_in_qs[2]),
    .clkout(net2179));
 b15cbf034ar1n64x5 hold424 (.clk(u_gpio_gen_filter_1__u_filter_diff_ctr_q[0]),
    .clkout(net2180));
 b15cbf034ar1n64x5 hold425 (.clk(u_gpio_reg2hw[15]),
    .clkout(net2181));
 b15cbf034ar1n64x5 hold426 (.clk(u_gpio_gen_filter_14__u_filter_diff_ctr_q[3]),
    .clkout(net2182));
 b15cbf034ar1n64x5 hold427 (.clk(n2629),
    .clkout(net2183));
 b15cbf034ar1n64x5 hold428 (.clk(u_gpio_gen_filter_2__u_filter_diff_ctr_q[0]),
    .clkout(net2184));
 b15cbf034ar1n64x5 hold429 (.clk(u_gpio_gen_filter_2__u_filter_diff_ctr_d[1]),
    .clkout(net2185));
 b15cbf034ar1n64x5 hold430 (.clk(u_gpio_gen_filter_14__u_filter_diff_ctr_q[0]),
    .clkout(net2186));
 b15cbf034ar1n64x5 hold431 (.clk(u_gpio_gen_filter_21__u_filter_diff_ctr_q[3]),
    .clkout(net2187));
 b15cbf034ar1n64x5 hold432 (.clk(n2777),
    .clkout(net2188));
 b15cbf034ar1n64x5 hold433 (.clk(u_gpio_gen_filter_14__u_filter_stored_value_q),
    .clkout(net2189));
 b15cbf034ar1n64x5 hold434 (.clk(u_gpio_gen_filter_10__u_filter_diff_ctr_q[2]),
    .clkout(net2190));
 b15cbf034ar1n64x5 hold435 (.clk(u_gpio_gen_filter_10__u_filter_diff_ctr_d[1]),
    .clkout(net2191));
 b15cbf034ar1n64x5 hold436 (.clk(net91),
    .clkout(net2192));
 b15cbf034ar1n64x5 hold437 (.clk(u_gpio_gen_filter_7__u_filter_stored_value_q),
    .clkout(net2193));
 b15cbf034ar1n64x5 hold438 (.clk(u_gpio_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[0]),
    .clkout(net2194));
 b15cbf034ar1n64x5 hold439 (.clk(u_gpio_gen_filter_22__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2195));
 b15cbf034ar1n64x5 hold440 (.clk(u_gpio_gen_filter_2__u_filter_diff_ctr_q[2]),
    .clkout(net2196));
 b15cbf034ar1n64x5 hold441 (.clk(u_gpio_u_reg_masked_oe_upper_data_qs[1]),
    .clkout(net2197));
 b15cbf034ar1n64x5 hold442 (.clk(u_gpio_gen_filter_24__u_filter_diff_ctr_q[3]),
    .clkout(net2198));
 b15cbf034ar1n64x5 hold443 (.clk(u_gpio_gen_filter_31__u_filter_stored_value_q),
    .clkout(net2199));
 b15cbf034ar1n64x5 hold444 (.clk(rst_ni),
    .clkout(net2200));
 b15cbf034ar1n64x5 hold445 (.clk(u_gpio_gen_filter_0__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2201));
 b15cbf034ar1n64x5 hold446 (.clk(u_gpio_gen_filter_3__u_filter_diff_ctr_q[1]),
    .clkout(net2202));
 b15cbf034ar1n64x5 hold447 (.clk(u_gpio_u_reg_data_in_qs[0]),
    .clkout(net2203));
 b15cbf034ar1n64x5 hold448 (.clk(net83),
    .clkout(net2204));
 b15cbf034ar1n64x5 hold449 (.clk(u_gpio_data_in_q[26]),
    .clkout(net2205));
 b15cbf034ar1n64x5 hold450 (.clk(u_gpio_u_reg_data_in_qs[19]),
    .clkout(net2206));
 b15cbf034ar1n64x5 hold451 (.clk(u_gpio_gen_filter_26__u_filter_diff_ctr_q[2]),
    .clkout(net2207));
 b15cbf034ar1n64x5 hold452 (.clk(u_gpio_gen_filter_26__u_filter_diff_ctr_d[0]),
    .clkout(net2208));
 b15cbf034ar1n64x5 hold453 (.clk(u_gpio_u_reg_data_in_qs[29]),
    .clkout(net2209));
 b15cbf034ar1n64x5 hold454 (.clk(u_xbar_periph_u_s1n_6_dev_select_outstanding[2]),
    .clkout(net2210));
 b15cbf034ar1n64x5 hold455 (.clk(u_gpio_reg2hw[1]),
    .clkout(net2211));
 b15cbf034ar1n64x5 hold456 (.clk(u_gpio_reg2hw[15]),
    .clkout(net2212));
 b15cbf034ar1n64x5 hold457 (.clk(u_xbar_periph_u_s1n_6_tl_u_i[17]),
    .clkout(net2213));
 b15cbf034ar1n64x5 hold458 (.clk(u_gpio_gen_filter_26__u_filter_diff_ctr_q[2]),
    .clkout(net2214));
 b15cbf034ar1n64x5 hold459 (.clk(u_gpio_gen_filter_2__u_filter_diff_ctr_q[3]),
    .clkout(net2215));
 b15cbf034ar1n64x5 hold460 (.clk(u_gpio_reg2hw[12]),
    .clkout(net2216));
 b15cbf034ar1n64x5 hold461 (.clk(gpio_2_xbar[18]),
    .clkout(net2217));
 b15cbf034ar1n64x5 hold462 (.clk(u_gpio_gen_filter_3__u_filter_diff_ctr_q[2]),
    .clkout(net2218));
 b15cbf034ar1n64x5 hold463 (.clk(u_gpio_gen_filter_21__u_filter_diff_ctr_q[3]),
    .clkout(net2219));
 b15cbf034ar1n64x5 hold464 (.clk(u_gpio_gen_filter_10__u_filter_diff_ctr_q[2]),
    .clkout(net2220));
 b15cbf034ar1n64x5 hold465 (.clk(u_gpio_gen_filter_11__u_filter_diff_ctr_q[0]),
    .clkout(net2221));
 b15cbf034ar1n64x5 hold466 (.clk(u_xbar_periph_u_s1n_6_dev_select_outstanding[2]),
    .clkout(net2222));
 b15cbf034ar1n64x5 hold467 (.clk(u_xbar_periph_u_s1n_6_dev_select_outstanding[2]),
    .clkout(net2223));
 b15zdnd11an1n64x5 FILLER_0_8 ();
 b15zdnd11an1n64x5 FILLER_0_72 ();
 b15zdnd11an1n64x5 FILLER_0_136 ();
 b15zdnd11an1n64x5 FILLER_0_200 ();
 b15zdnd11an1n64x5 FILLER_0_264 ();
 b15zdnd11an1n64x5 FILLER_0_328 ();
 b15zdnd11an1n64x5 FILLER_0_392 ();
 b15zdnd11an1n64x5 FILLER_0_456 ();
 b15zdnd11an1n64x5 FILLER_0_520 ();
 b15zdnd11an1n64x5 FILLER_0_584 ();
 b15zdnd11an1n64x5 FILLER_0_648 ();
 b15zdnd11an1n04x5 FILLER_0_712 ();
 b15zdnd00an1n02x5 FILLER_0_716 ();
 b15zdnd11an1n64x5 FILLER_0_726 ();
 b15zdnd11an1n64x5 FILLER_0_790 ();
 b15zdnd11an1n64x5 FILLER_0_854 ();
 b15zdnd11an1n64x5 FILLER_0_918 ();
 b15zdnd11an1n32x5 FILLER_0_982 ();
 b15zdnd11an1n16x5 FILLER_0_1014 ();
 b15zdnd11an1n08x5 FILLER_0_1030 ();
 b15zdnd00an1n01x5 FILLER_0_1038 ();
 b15zdnd11an1n08x5 FILLER_0_1043 ();
 b15zdnd11an1n04x5 FILLER_0_1051 ();
 b15zdnd00an1n01x5 FILLER_0_1055 ();
 b15zdnd11an1n16x5 FILLER_0_1060 ();
 b15zdnd11an1n08x5 FILLER_0_1076 ();
 b15zdnd00an1n02x5 FILLER_0_1084 ();
 b15zdnd00an1n01x5 FILLER_0_1086 ();
 b15zdnd11an1n16x5 FILLER_0_1091 ();
 b15zdnd11an1n04x5 FILLER_0_1107 ();
 b15zdnd00an1n02x5 FILLER_0_1111 ();
 b15zdnd00an1n01x5 FILLER_0_1113 ();
 b15zdnd11an1n32x5 FILLER_0_1122 ();
 b15zdnd11an1n04x5 FILLER_0_1154 ();
 b15zdnd00an1n01x5 FILLER_0_1158 ();
 b15zdnd11an1n32x5 FILLER_0_1166 ();
 b15zdnd11an1n16x5 FILLER_0_1198 ();
 b15zdnd00an1n02x5 FILLER_0_1214 ();
 b15zdnd00an1n01x5 FILLER_0_1216 ();
 b15zdnd11an1n64x5 FILLER_0_1221 ();
 b15zdnd11an1n16x5 FILLER_0_1285 ();
 b15zdnd11an1n04x5 FILLER_0_1309 ();
 b15zdnd11an1n08x5 FILLER_0_1320 ();
 b15zdnd11an1n04x5 FILLER_0_1328 ();
 b15zdnd00an1n02x5 FILLER_0_1332 ();
 b15zdnd11an1n32x5 FILLER_0_1342 ();
 b15zdnd11an1n16x5 FILLER_0_1374 ();
 b15zdnd11an1n04x5 FILLER_0_1394 ();
 b15zdnd11an1n32x5 FILLER_0_1402 ();
 b15zdnd00an1n02x5 FILLER_0_1434 ();
 b15zdnd11an1n16x5 FILLER_0_1444 ();
 b15zdnd11an1n04x5 FILLER_0_1460 ();
 b15zdnd00an1n01x5 FILLER_0_1464 ();
 b15zdnd11an1n64x5 FILLER_0_1469 ();
 b15zdnd11an1n64x5 FILLER_0_1533 ();
 b15zdnd11an1n64x5 FILLER_0_1597 ();
 b15zdnd11an1n64x5 FILLER_0_1661 ();
 b15zdnd11an1n64x5 FILLER_0_1725 ();
 b15zdnd11an1n64x5 FILLER_0_1789 ();
 b15zdnd11an1n64x5 FILLER_0_1853 ();
 b15zdnd11an1n64x5 FILLER_0_1917 ();
 b15zdnd11an1n64x5 FILLER_0_1981 ();
 b15zdnd11an1n64x5 FILLER_0_2045 ();
 b15zdnd11an1n32x5 FILLER_0_2109 ();
 b15zdnd11an1n08x5 FILLER_0_2141 ();
 b15zdnd11an1n04x5 FILLER_0_2149 ();
 b15zdnd00an1n01x5 FILLER_0_2153 ();
 b15zdnd11an1n64x5 FILLER_0_2162 ();
 b15zdnd11an1n32x5 FILLER_0_2226 ();
 b15zdnd11an1n16x5 FILLER_0_2258 ();
 b15zdnd00an1n02x5 FILLER_0_2274 ();
 b15zdnd11an1n64x5 FILLER_1_0 ();
 b15zdnd11an1n64x5 FILLER_1_64 ();
 b15zdnd11an1n64x5 FILLER_1_128 ();
 b15zdnd11an1n64x5 FILLER_1_192 ();
 b15zdnd11an1n64x5 FILLER_1_256 ();
 b15zdnd11an1n64x5 FILLER_1_320 ();
 b15zdnd11an1n64x5 FILLER_1_384 ();
 b15zdnd11an1n64x5 FILLER_1_448 ();
 b15zdnd11an1n64x5 FILLER_1_512 ();
 b15zdnd11an1n64x5 FILLER_1_576 ();
 b15zdnd11an1n64x5 FILLER_1_640 ();
 b15zdnd11an1n64x5 FILLER_1_704 ();
 b15zdnd11an1n64x5 FILLER_1_768 ();
 b15zdnd11an1n64x5 FILLER_1_832 ();
 b15zdnd11an1n64x5 FILLER_1_896 ();
 b15zdnd11an1n32x5 FILLER_1_960 ();
 b15zdnd11an1n16x5 FILLER_1_992 ();
 b15zdnd11an1n64x5 FILLER_1_1012 ();
 b15zdnd11an1n32x5 FILLER_1_1076 ();
 b15zdnd11an1n04x5 FILLER_1_1115 ();
 b15zdnd00an1n01x5 FILLER_1_1119 ();
 b15zdnd11an1n64x5 FILLER_1_1131 ();
 b15zdnd11an1n64x5 FILLER_1_1195 ();
 b15zdnd11an1n64x5 FILLER_1_1259 ();
 b15zdnd11an1n08x5 FILLER_1_1323 ();
 b15zdnd11an1n04x5 FILLER_1_1331 ();
 b15zdnd00an1n02x5 FILLER_1_1335 ();
 b15zdnd11an1n64x5 FILLER_1_1345 ();
 b15zdnd11an1n64x5 FILLER_1_1409 ();
 b15zdnd11an1n64x5 FILLER_1_1473 ();
 b15zdnd11an1n64x5 FILLER_1_1537 ();
 b15zdnd11an1n64x5 FILLER_1_1601 ();
 b15zdnd11an1n64x5 FILLER_1_1665 ();
 b15zdnd11an1n64x5 FILLER_1_1729 ();
 b15zdnd11an1n64x5 FILLER_1_1793 ();
 b15zdnd11an1n64x5 FILLER_1_1857 ();
 b15zdnd11an1n64x5 FILLER_1_1921 ();
 b15zdnd11an1n64x5 FILLER_1_1985 ();
 b15zdnd11an1n64x5 FILLER_1_2049 ();
 b15zdnd11an1n64x5 FILLER_1_2113 ();
 b15zdnd11an1n64x5 FILLER_1_2177 ();
 b15zdnd11an1n32x5 FILLER_1_2241 ();
 b15zdnd11an1n08x5 FILLER_1_2273 ();
 b15zdnd00an1n02x5 FILLER_1_2281 ();
 b15zdnd00an1n01x5 FILLER_1_2283 ();
 b15zdnd11an1n64x5 FILLER_2_8 ();
 b15zdnd11an1n64x5 FILLER_2_72 ();
 b15zdnd11an1n64x5 FILLER_2_136 ();
 b15zdnd11an1n64x5 FILLER_2_200 ();
 b15zdnd11an1n64x5 FILLER_2_264 ();
 b15zdnd11an1n64x5 FILLER_2_328 ();
 b15zdnd11an1n64x5 FILLER_2_392 ();
 b15zdnd11an1n64x5 FILLER_2_456 ();
 b15zdnd11an1n64x5 FILLER_2_520 ();
 b15zdnd11an1n64x5 FILLER_2_584 ();
 b15zdnd11an1n64x5 FILLER_2_648 ();
 b15zdnd11an1n04x5 FILLER_2_712 ();
 b15zdnd00an1n02x5 FILLER_2_716 ();
 b15zdnd11an1n64x5 FILLER_2_726 ();
 b15zdnd11an1n64x5 FILLER_2_790 ();
 b15zdnd11an1n64x5 FILLER_2_854 ();
 b15zdnd11an1n64x5 FILLER_2_918 ();
 b15zdnd11an1n64x5 FILLER_2_982 ();
 b15zdnd11an1n64x5 FILLER_2_1046 ();
 b15zdnd11an1n64x5 FILLER_2_1110 ();
 b15zdnd11an1n64x5 FILLER_2_1174 ();
 b15zdnd11an1n64x5 FILLER_2_1238 ();
 b15zdnd11an1n64x5 FILLER_2_1302 ();
 b15zdnd11an1n64x5 FILLER_2_1366 ();
 b15zdnd11an1n64x5 FILLER_2_1430 ();
 b15zdnd11an1n64x5 FILLER_2_1494 ();
 b15zdnd11an1n64x5 FILLER_2_1558 ();
 b15zdnd11an1n64x5 FILLER_2_1622 ();
 b15zdnd11an1n64x5 FILLER_2_1686 ();
 b15zdnd11an1n64x5 FILLER_2_1750 ();
 b15zdnd11an1n64x5 FILLER_2_1814 ();
 b15zdnd11an1n64x5 FILLER_2_1878 ();
 b15zdnd11an1n64x5 FILLER_2_1942 ();
 b15zdnd11an1n64x5 FILLER_2_2006 ();
 b15zdnd11an1n64x5 FILLER_2_2070 ();
 b15zdnd11an1n16x5 FILLER_2_2134 ();
 b15zdnd11an1n04x5 FILLER_2_2150 ();
 b15zdnd11an1n64x5 FILLER_2_2162 ();
 b15zdnd11an1n32x5 FILLER_2_2226 ();
 b15zdnd11an1n16x5 FILLER_2_2258 ();
 b15zdnd00an1n02x5 FILLER_2_2274 ();
 b15zdnd11an1n64x5 FILLER_3_0 ();
 b15zdnd11an1n64x5 FILLER_3_64 ();
 b15zdnd11an1n64x5 FILLER_3_128 ();
 b15zdnd11an1n64x5 FILLER_3_192 ();
 b15zdnd11an1n64x5 FILLER_3_256 ();
 b15zdnd11an1n64x5 FILLER_3_320 ();
 b15zdnd11an1n64x5 FILLER_3_384 ();
 b15zdnd11an1n64x5 FILLER_3_448 ();
 b15zdnd11an1n64x5 FILLER_3_512 ();
 b15zdnd11an1n64x5 FILLER_3_576 ();
 b15zdnd11an1n64x5 FILLER_3_640 ();
 b15zdnd11an1n64x5 FILLER_3_704 ();
 b15zdnd11an1n64x5 FILLER_3_768 ();
 b15zdnd11an1n64x5 FILLER_3_832 ();
 b15zdnd11an1n64x5 FILLER_3_896 ();
 b15zdnd11an1n64x5 FILLER_3_960 ();
 b15zdnd11an1n64x5 FILLER_3_1024 ();
 b15zdnd11an1n64x5 FILLER_3_1088 ();
 b15zdnd11an1n64x5 FILLER_3_1152 ();
 b15zdnd11an1n64x5 FILLER_3_1216 ();
 b15zdnd11an1n64x5 FILLER_3_1280 ();
 b15zdnd11an1n64x5 FILLER_3_1344 ();
 b15zdnd11an1n64x5 FILLER_3_1408 ();
 b15zdnd11an1n64x5 FILLER_3_1472 ();
 b15zdnd11an1n64x5 FILLER_3_1536 ();
 b15zdnd11an1n64x5 FILLER_3_1600 ();
 b15zdnd11an1n64x5 FILLER_3_1664 ();
 b15zdnd11an1n64x5 FILLER_3_1728 ();
 b15zdnd11an1n64x5 FILLER_3_1792 ();
 b15zdnd11an1n64x5 FILLER_3_1856 ();
 b15zdnd11an1n64x5 FILLER_3_1920 ();
 b15zdnd11an1n64x5 FILLER_3_1984 ();
 b15zdnd11an1n64x5 FILLER_3_2048 ();
 b15zdnd11an1n64x5 FILLER_3_2112 ();
 b15zdnd11an1n64x5 FILLER_3_2176 ();
 b15zdnd11an1n32x5 FILLER_3_2240 ();
 b15zdnd11an1n08x5 FILLER_3_2272 ();
 b15zdnd11an1n04x5 FILLER_3_2280 ();
 b15zdnd11an1n64x5 FILLER_4_8 ();
 b15zdnd11an1n64x5 FILLER_4_72 ();
 b15zdnd11an1n64x5 FILLER_4_136 ();
 b15zdnd11an1n64x5 FILLER_4_200 ();
 b15zdnd11an1n64x5 FILLER_4_264 ();
 b15zdnd11an1n64x5 FILLER_4_328 ();
 b15zdnd11an1n64x5 FILLER_4_392 ();
 b15zdnd11an1n64x5 FILLER_4_456 ();
 b15zdnd11an1n64x5 FILLER_4_520 ();
 b15zdnd11an1n64x5 FILLER_4_584 ();
 b15zdnd11an1n64x5 FILLER_4_648 ();
 b15zdnd11an1n04x5 FILLER_4_712 ();
 b15zdnd00an1n02x5 FILLER_4_716 ();
 b15zdnd11an1n64x5 FILLER_4_726 ();
 b15zdnd11an1n64x5 FILLER_4_790 ();
 b15zdnd11an1n64x5 FILLER_4_854 ();
 b15zdnd11an1n64x5 FILLER_4_918 ();
 b15zdnd11an1n64x5 FILLER_4_982 ();
 b15zdnd11an1n64x5 FILLER_4_1046 ();
 b15zdnd11an1n64x5 FILLER_4_1110 ();
 b15zdnd11an1n64x5 FILLER_4_1174 ();
 b15zdnd11an1n64x5 FILLER_4_1238 ();
 b15zdnd11an1n64x5 FILLER_4_1302 ();
 b15zdnd11an1n64x5 FILLER_4_1366 ();
 b15zdnd11an1n64x5 FILLER_4_1430 ();
 b15zdnd11an1n64x5 FILLER_4_1494 ();
 b15zdnd11an1n64x5 FILLER_4_1558 ();
 b15zdnd11an1n64x5 FILLER_4_1622 ();
 b15zdnd11an1n64x5 FILLER_4_1686 ();
 b15zdnd11an1n64x5 FILLER_4_1750 ();
 b15zdnd11an1n64x5 FILLER_4_1814 ();
 b15zdnd11an1n64x5 FILLER_4_1878 ();
 b15zdnd11an1n64x5 FILLER_4_1942 ();
 b15zdnd11an1n64x5 FILLER_4_2006 ();
 b15zdnd11an1n64x5 FILLER_4_2070 ();
 b15zdnd11an1n16x5 FILLER_4_2134 ();
 b15zdnd11an1n04x5 FILLER_4_2150 ();
 b15zdnd11an1n64x5 FILLER_4_2162 ();
 b15zdnd11an1n32x5 FILLER_4_2226 ();
 b15zdnd11an1n16x5 FILLER_4_2258 ();
 b15zdnd00an1n02x5 FILLER_4_2274 ();
 b15zdnd11an1n64x5 FILLER_5_0 ();
 b15zdnd11an1n64x5 FILLER_5_64 ();
 b15zdnd11an1n64x5 FILLER_5_128 ();
 b15zdnd11an1n64x5 FILLER_5_192 ();
 b15zdnd11an1n64x5 FILLER_5_256 ();
 b15zdnd11an1n64x5 FILLER_5_320 ();
 b15zdnd11an1n64x5 FILLER_5_384 ();
 b15zdnd11an1n64x5 FILLER_5_448 ();
 b15zdnd11an1n64x5 FILLER_5_512 ();
 b15zdnd11an1n64x5 FILLER_5_576 ();
 b15zdnd11an1n64x5 FILLER_5_640 ();
 b15zdnd11an1n64x5 FILLER_5_704 ();
 b15zdnd11an1n64x5 FILLER_5_768 ();
 b15zdnd11an1n64x5 FILLER_5_832 ();
 b15zdnd11an1n64x5 FILLER_5_896 ();
 b15zdnd11an1n64x5 FILLER_5_960 ();
 b15zdnd11an1n64x5 FILLER_5_1024 ();
 b15zdnd11an1n64x5 FILLER_5_1088 ();
 b15zdnd11an1n64x5 FILLER_5_1152 ();
 b15zdnd11an1n64x5 FILLER_5_1216 ();
 b15zdnd11an1n64x5 FILLER_5_1280 ();
 b15zdnd11an1n64x5 FILLER_5_1344 ();
 b15zdnd11an1n64x5 FILLER_5_1408 ();
 b15zdnd11an1n64x5 FILLER_5_1472 ();
 b15zdnd11an1n64x5 FILLER_5_1536 ();
 b15zdnd11an1n64x5 FILLER_5_1600 ();
 b15zdnd11an1n64x5 FILLER_5_1664 ();
 b15zdnd11an1n64x5 FILLER_5_1728 ();
 b15zdnd11an1n64x5 FILLER_5_1792 ();
 b15zdnd11an1n64x5 FILLER_5_1856 ();
 b15zdnd11an1n64x5 FILLER_5_1920 ();
 b15zdnd11an1n64x5 FILLER_5_1984 ();
 b15zdnd11an1n64x5 FILLER_5_2048 ();
 b15zdnd11an1n64x5 FILLER_5_2112 ();
 b15zdnd11an1n64x5 FILLER_5_2176 ();
 b15zdnd11an1n32x5 FILLER_5_2240 ();
 b15zdnd11an1n08x5 FILLER_5_2272 ();
 b15zdnd11an1n04x5 FILLER_5_2280 ();
 b15zdnd11an1n64x5 FILLER_6_8 ();
 b15zdnd11an1n64x5 FILLER_6_72 ();
 b15zdnd11an1n64x5 FILLER_6_136 ();
 b15zdnd11an1n64x5 FILLER_6_200 ();
 b15zdnd11an1n64x5 FILLER_6_264 ();
 b15zdnd11an1n64x5 FILLER_6_328 ();
 b15zdnd11an1n64x5 FILLER_6_392 ();
 b15zdnd11an1n64x5 FILLER_6_456 ();
 b15zdnd11an1n64x5 FILLER_6_520 ();
 b15zdnd11an1n64x5 FILLER_6_584 ();
 b15zdnd11an1n64x5 FILLER_6_648 ();
 b15zdnd11an1n04x5 FILLER_6_712 ();
 b15zdnd00an1n02x5 FILLER_6_716 ();
 b15zdnd11an1n64x5 FILLER_6_726 ();
 b15zdnd11an1n64x5 FILLER_6_790 ();
 b15zdnd11an1n64x5 FILLER_6_854 ();
 b15zdnd11an1n64x5 FILLER_6_918 ();
 b15zdnd11an1n64x5 FILLER_6_982 ();
 b15zdnd11an1n64x5 FILLER_6_1046 ();
 b15zdnd11an1n64x5 FILLER_6_1110 ();
 b15zdnd11an1n64x5 FILLER_6_1174 ();
 b15zdnd11an1n64x5 FILLER_6_1238 ();
 b15zdnd11an1n64x5 FILLER_6_1302 ();
 b15zdnd11an1n64x5 FILLER_6_1366 ();
 b15zdnd11an1n64x5 FILLER_6_1430 ();
 b15zdnd11an1n64x5 FILLER_6_1494 ();
 b15zdnd11an1n64x5 FILLER_6_1558 ();
 b15zdnd11an1n64x5 FILLER_6_1622 ();
 b15zdnd11an1n64x5 FILLER_6_1686 ();
 b15zdnd11an1n64x5 FILLER_6_1750 ();
 b15zdnd11an1n64x5 FILLER_6_1814 ();
 b15zdnd11an1n64x5 FILLER_6_1878 ();
 b15zdnd11an1n64x5 FILLER_6_1942 ();
 b15zdnd11an1n64x5 FILLER_6_2006 ();
 b15zdnd11an1n64x5 FILLER_6_2070 ();
 b15zdnd11an1n16x5 FILLER_6_2134 ();
 b15zdnd11an1n04x5 FILLER_6_2150 ();
 b15zdnd11an1n64x5 FILLER_6_2162 ();
 b15zdnd11an1n32x5 FILLER_6_2226 ();
 b15zdnd11an1n16x5 FILLER_6_2258 ();
 b15zdnd00an1n02x5 FILLER_6_2274 ();
 b15zdnd11an1n64x5 FILLER_7_0 ();
 b15zdnd11an1n64x5 FILLER_7_64 ();
 b15zdnd11an1n64x5 FILLER_7_128 ();
 b15zdnd11an1n64x5 FILLER_7_192 ();
 b15zdnd11an1n64x5 FILLER_7_256 ();
 b15zdnd11an1n64x5 FILLER_7_320 ();
 b15zdnd11an1n64x5 FILLER_7_384 ();
 b15zdnd11an1n64x5 FILLER_7_448 ();
 b15zdnd11an1n64x5 FILLER_7_512 ();
 b15zdnd11an1n64x5 FILLER_7_576 ();
 b15zdnd11an1n64x5 FILLER_7_640 ();
 b15zdnd11an1n64x5 FILLER_7_704 ();
 b15zdnd11an1n64x5 FILLER_7_768 ();
 b15zdnd11an1n64x5 FILLER_7_832 ();
 b15zdnd11an1n64x5 FILLER_7_896 ();
 b15zdnd11an1n32x5 FILLER_7_960 ();
 b15zdnd11an1n16x5 FILLER_7_992 ();
 b15zdnd11an1n08x5 FILLER_7_1008 ();
 b15zdnd11an1n04x5 FILLER_7_1058 ();
 b15zdnd00an1n02x5 FILLER_7_1062 ();
 b15zdnd11an1n64x5 FILLER_7_1106 ();
 b15zdnd11an1n64x5 FILLER_7_1170 ();
 b15zdnd11an1n64x5 FILLER_7_1234 ();
 b15zdnd11an1n64x5 FILLER_7_1298 ();
 b15zdnd11an1n16x5 FILLER_7_1362 ();
 b15zdnd11an1n08x5 FILLER_7_1378 ();
 b15zdnd11an1n04x5 FILLER_7_1386 ();
 b15zdnd11an1n32x5 FILLER_7_1399 ();
 b15zdnd11an1n16x5 FILLER_7_1431 ();
 b15zdnd11an1n04x5 FILLER_7_1447 ();
 b15zdnd00an1n01x5 FILLER_7_1451 ();
 b15zdnd11an1n16x5 FILLER_7_1466 ();
 b15zdnd00an1n02x5 FILLER_7_1482 ();
 b15zdnd00an1n01x5 FILLER_7_1484 ();
 b15zdnd11an1n64x5 FILLER_7_1516 ();
 b15zdnd11an1n64x5 FILLER_7_1580 ();
 b15zdnd11an1n64x5 FILLER_7_1644 ();
 b15zdnd11an1n64x5 FILLER_7_1708 ();
 b15zdnd11an1n64x5 FILLER_7_1772 ();
 b15zdnd11an1n64x5 FILLER_7_1836 ();
 b15zdnd11an1n64x5 FILLER_7_1900 ();
 b15zdnd11an1n64x5 FILLER_7_1964 ();
 b15zdnd11an1n64x5 FILLER_7_2028 ();
 b15zdnd11an1n64x5 FILLER_7_2092 ();
 b15zdnd11an1n64x5 FILLER_7_2156 ();
 b15zdnd11an1n64x5 FILLER_7_2220 ();
 b15zdnd11an1n64x5 FILLER_8_8 ();
 b15zdnd11an1n64x5 FILLER_8_72 ();
 b15zdnd11an1n64x5 FILLER_8_136 ();
 b15zdnd11an1n64x5 FILLER_8_200 ();
 b15zdnd11an1n64x5 FILLER_8_264 ();
 b15zdnd11an1n64x5 FILLER_8_328 ();
 b15zdnd11an1n64x5 FILLER_8_392 ();
 b15zdnd11an1n64x5 FILLER_8_456 ();
 b15zdnd11an1n64x5 FILLER_8_520 ();
 b15zdnd11an1n64x5 FILLER_8_584 ();
 b15zdnd11an1n64x5 FILLER_8_648 ();
 b15zdnd11an1n04x5 FILLER_8_712 ();
 b15zdnd00an1n02x5 FILLER_8_716 ();
 b15zdnd11an1n64x5 FILLER_8_726 ();
 b15zdnd11an1n64x5 FILLER_8_790 ();
 b15zdnd11an1n64x5 FILLER_8_854 ();
 b15zdnd11an1n64x5 FILLER_8_918 ();
 b15zdnd11an1n32x5 FILLER_8_982 ();
 b15zdnd11an1n08x5 FILLER_8_1014 ();
 b15zdnd11an1n04x5 FILLER_8_1022 ();
 b15zdnd00an1n02x5 FILLER_8_1026 ();
 b15zdnd00an1n01x5 FILLER_8_1028 ();
 b15zdnd11an1n32x5 FILLER_8_1038 ();
 b15zdnd11an1n04x5 FILLER_8_1070 ();
 b15zdnd11an1n16x5 FILLER_8_1081 ();
 b15zdnd11an1n64x5 FILLER_8_1104 ();
 b15zdnd11an1n32x5 FILLER_8_1168 ();
 b15zdnd11an1n16x5 FILLER_8_1200 ();
 b15zdnd11an1n08x5 FILLER_8_1216 ();
 b15zdnd00an1n02x5 FILLER_8_1224 ();
 b15zdnd11an1n04x5 FILLER_8_1231 ();
 b15zdnd11an1n08x5 FILLER_8_1244 ();
 b15zdnd11an1n04x5 FILLER_8_1252 ();
 b15zdnd00an1n02x5 FILLER_8_1256 ();
 b15zdnd00an1n01x5 FILLER_8_1258 ();
 b15zdnd11an1n32x5 FILLER_8_1266 ();
 b15zdnd11an1n16x5 FILLER_8_1298 ();
 b15zdnd11an1n04x5 FILLER_8_1314 ();
 b15zdnd11an1n08x5 FILLER_8_1332 ();
 b15zdnd00an1n02x5 FILLER_8_1340 ();
 b15zdnd00an1n01x5 FILLER_8_1342 ();
 b15zdnd11an1n32x5 FILLER_8_1353 ();
 b15zdnd11an1n08x5 FILLER_8_1385 ();
 b15zdnd00an1n02x5 FILLER_8_1393 ();
 b15zdnd00an1n01x5 FILLER_8_1395 ();
 b15zdnd11an1n16x5 FILLER_8_1438 ();
 b15zdnd00an1n02x5 FILLER_8_1454 ();
 b15zdnd00an1n01x5 FILLER_8_1456 ();
 b15zdnd11an1n64x5 FILLER_8_1499 ();
 b15zdnd11an1n64x5 FILLER_8_1563 ();
 b15zdnd11an1n64x5 FILLER_8_1627 ();
 b15zdnd11an1n64x5 FILLER_8_1691 ();
 b15zdnd11an1n64x5 FILLER_8_1755 ();
 b15zdnd11an1n64x5 FILLER_8_1819 ();
 b15zdnd11an1n64x5 FILLER_8_1883 ();
 b15zdnd11an1n64x5 FILLER_8_1947 ();
 b15zdnd11an1n64x5 FILLER_8_2011 ();
 b15zdnd11an1n64x5 FILLER_8_2075 ();
 b15zdnd11an1n08x5 FILLER_8_2139 ();
 b15zdnd11an1n04x5 FILLER_8_2147 ();
 b15zdnd00an1n02x5 FILLER_8_2151 ();
 b15zdnd00an1n01x5 FILLER_8_2153 ();
 b15zdnd11an1n64x5 FILLER_8_2162 ();
 b15zdnd11an1n32x5 FILLER_8_2226 ();
 b15zdnd11an1n16x5 FILLER_8_2258 ();
 b15zdnd00an1n02x5 FILLER_8_2274 ();
 b15zdnd11an1n64x5 FILLER_9_0 ();
 b15zdnd11an1n64x5 FILLER_9_64 ();
 b15zdnd11an1n64x5 FILLER_9_128 ();
 b15zdnd11an1n64x5 FILLER_9_192 ();
 b15zdnd11an1n64x5 FILLER_9_256 ();
 b15zdnd11an1n64x5 FILLER_9_320 ();
 b15zdnd11an1n64x5 FILLER_9_384 ();
 b15zdnd11an1n64x5 FILLER_9_448 ();
 b15zdnd11an1n64x5 FILLER_9_512 ();
 b15zdnd11an1n64x5 FILLER_9_576 ();
 b15zdnd11an1n64x5 FILLER_9_640 ();
 b15zdnd11an1n64x5 FILLER_9_704 ();
 b15zdnd11an1n64x5 FILLER_9_768 ();
 b15zdnd11an1n64x5 FILLER_9_832 ();
 b15zdnd11an1n64x5 FILLER_9_896 ();
 b15zdnd11an1n32x5 FILLER_9_960 ();
 b15zdnd11an1n04x5 FILLER_9_992 ();
 b15zdnd11an1n16x5 FILLER_9_1016 ();
 b15zdnd11an1n04x5 FILLER_9_1032 ();
 b15zdnd11an1n04x5 FILLER_9_1067 ();
 b15zdnd11an1n04x5 FILLER_9_1078 ();
 b15zdnd00an1n02x5 FILLER_9_1082 ();
 b15zdnd00an1n01x5 FILLER_9_1084 ();
 b15zdnd11an1n64x5 FILLER_9_1096 ();
 b15zdnd11an1n64x5 FILLER_9_1160 ();
 b15zdnd11an1n32x5 FILLER_9_1224 ();
 b15zdnd00an1n02x5 FILLER_9_1256 ();
 b15zdnd00an1n01x5 FILLER_9_1258 ();
 b15zdnd11an1n32x5 FILLER_9_1266 ();
 b15zdnd11an1n16x5 FILLER_9_1298 ();
 b15zdnd11an1n08x5 FILLER_9_1314 ();
 b15zdnd00an1n02x5 FILLER_9_1322 ();
 b15zdnd00an1n01x5 FILLER_9_1324 ();
 b15zdnd11an1n32x5 FILLER_9_1331 ();
 b15zdnd11an1n16x5 FILLER_9_1363 ();
 b15zdnd11an1n08x5 FILLER_9_1379 ();
 b15zdnd11an1n04x5 FILLER_9_1387 ();
 b15zdnd00an1n01x5 FILLER_9_1391 ();
 b15zdnd11an1n64x5 FILLER_9_1423 ();
 b15zdnd11an1n64x5 FILLER_9_1487 ();
 b15zdnd11an1n64x5 FILLER_9_1551 ();
 b15zdnd11an1n64x5 FILLER_9_1615 ();
 b15zdnd11an1n64x5 FILLER_9_1679 ();
 b15zdnd11an1n64x5 FILLER_9_1743 ();
 b15zdnd11an1n64x5 FILLER_9_1807 ();
 b15zdnd11an1n64x5 FILLER_9_1871 ();
 b15zdnd11an1n64x5 FILLER_9_1935 ();
 b15zdnd11an1n64x5 FILLER_9_1999 ();
 b15zdnd11an1n64x5 FILLER_9_2063 ();
 b15zdnd11an1n64x5 FILLER_9_2127 ();
 b15zdnd11an1n64x5 FILLER_9_2191 ();
 b15zdnd11an1n16x5 FILLER_9_2255 ();
 b15zdnd11an1n08x5 FILLER_9_2271 ();
 b15zdnd11an1n04x5 FILLER_9_2279 ();
 b15zdnd00an1n01x5 FILLER_9_2283 ();
 b15zdnd11an1n64x5 FILLER_10_8 ();
 b15zdnd11an1n64x5 FILLER_10_72 ();
 b15zdnd11an1n64x5 FILLER_10_136 ();
 b15zdnd11an1n64x5 FILLER_10_200 ();
 b15zdnd11an1n64x5 FILLER_10_264 ();
 b15zdnd11an1n64x5 FILLER_10_328 ();
 b15zdnd11an1n64x5 FILLER_10_392 ();
 b15zdnd11an1n64x5 FILLER_10_456 ();
 b15zdnd11an1n64x5 FILLER_10_520 ();
 b15zdnd11an1n64x5 FILLER_10_584 ();
 b15zdnd11an1n64x5 FILLER_10_648 ();
 b15zdnd11an1n04x5 FILLER_10_712 ();
 b15zdnd00an1n02x5 FILLER_10_716 ();
 b15zdnd11an1n64x5 FILLER_10_726 ();
 b15zdnd11an1n64x5 FILLER_10_790 ();
 b15zdnd11an1n64x5 FILLER_10_854 ();
 b15zdnd11an1n64x5 FILLER_10_918 ();
 b15zdnd11an1n64x5 FILLER_10_982 ();
 b15zdnd11an1n16x5 FILLER_10_1046 ();
 b15zdnd11an1n04x5 FILLER_10_1062 ();
 b15zdnd00an1n01x5 FILLER_10_1066 ();
 b15zdnd11an1n64x5 FILLER_10_1078 ();
 b15zdnd11an1n64x5 FILLER_10_1142 ();
 b15zdnd11an1n64x5 FILLER_10_1206 ();
 b15zdnd11an1n64x5 FILLER_10_1270 ();
 b15zdnd11an1n64x5 FILLER_10_1334 ();
 b15zdnd11an1n16x5 FILLER_10_1398 ();
 b15zdnd11an1n08x5 FILLER_10_1414 ();
 b15zdnd11an1n64x5 FILLER_10_1427 ();
 b15zdnd11an1n64x5 FILLER_10_1491 ();
 b15zdnd11an1n64x5 FILLER_10_1555 ();
 b15zdnd11an1n64x5 FILLER_10_1619 ();
 b15zdnd11an1n64x5 FILLER_10_1683 ();
 b15zdnd11an1n64x5 FILLER_10_1747 ();
 b15zdnd11an1n64x5 FILLER_10_1811 ();
 b15zdnd11an1n64x5 FILLER_10_1875 ();
 b15zdnd11an1n64x5 FILLER_10_1939 ();
 b15zdnd11an1n64x5 FILLER_10_2003 ();
 b15zdnd11an1n64x5 FILLER_10_2067 ();
 b15zdnd11an1n16x5 FILLER_10_2131 ();
 b15zdnd11an1n04x5 FILLER_10_2147 ();
 b15zdnd00an1n02x5 FILLER_10_2151 ();
 b15zdnd00an1n01x5 FILLER_10_2153 ();
 b15zdnd11an1n64x5 FILLER_10_2162 ();
 b15zdnd11an1n32x5 FILLER_10_2226 ();
 b15zdnd11an1n16x5 FILLER_10_2258 ();
 b15zdnd00an1n02x5 FILLER_10_2274 ();
 b15zdnd11an1n64x5 FILLER_11_0 ();
 b15zdnd11an1n64x5 FILLER_11_64 ();
 b15zdnd11an1n64x5 FILLER_11_128 ();
 b15zdnd11an1n64x5 FILLER_11_192 ();
 b15zdnd11an1n64x5 FILLER_11_256 ();
 b15zdnd11an1n64x5 FILLER_11_320 ();
 b15zdnd11an1n64x5 FILLER_11_384 ();
 b15zdnd11an1n64x5 FILLER_11_448 ();
 b15zdnd11an1n64x5 FILLER_11_512 ();
 b15zdnd11an1n64x5 FILLER_11_576 ();
 b15zdnd11an1n64x5 FILLER_11_640 ();
 b15zdnd11an1n64x5 FILLER_11_704 ();
 b15zdnd11an1n64x5 FILLER_11_768 ();
 b15zdnd11an1n64x5 FILLER_11_832 ();
 b15zdnd11an1n64x5 FILLER_11_896 ();
 b15zdnd11an1n64x5 FILLER_11_960 ();
 b15zdnd11an1n64x5 FILLER_11_1024 ();
 b15zdnd11an1n64x5 FILLER_11_1088 ();
 b15zdnd11an1n64x5 FILLER_11_1152 ();
 b15zdnd11an1n32x5 FILLER_11_1216 ();
 b15zdnd11an1n16x5 FILLER_11_1248 ();
 b15zdnd11an1n08x5 FILLER_11_1264 ();
 b15zdnd11an1n04x5 FILLER_11_1272 ();
 b15zdnd00an1n01x5 FILLER_11_1276 ();
 b15zdnd11an1n32x5 FILLER_11_1286 ();
 b15zdnd11an1n08x5 FILLER_11_1318 ();
 b15zdnd11an1n04x5 FILLER_11_1326 ();
 b15zdnd11an1n64x5 FILLER_11_1372 ();
 b15zdnd11an1n32x5 FILLER_11_1436 ();
 b15zdnd11an1n04x5 FILLER_11_1468 ();
 b15zdnd00an1n02x5 FILLER_11_1472 ();
 b15zdnd11an1n64x5 FILLER_11_1481 ();
 b15zdnd11an1n64x5 FILLER_11_1545 ();
 b15zdnd11an1n64x5 FILLER_11_1609 ();
 b15zdnd11an1n64x5 FILLER_11_1673 ();
 b15zdnd11an1n64x5 FILLER_11_1737 ();
 b15zdnd11an1n64x5 FILLER_11_1801 ();
 b15zdnd11an1n64x5 FILLER_11_1865 ();
 b15zdnd11an1n64x5 FILLER_11_1929 ();
 b15zdnd11an1n64x5 FILLER_11_1993 ();
 b15zdnd11an1n64x5 FILLER_11_2057 ();
 b15zdnd11an1n64x5 FILLER_11_2121 ();
 b15zdnd11an1n64x5 FILLER_11_2185 ();
 b15zdnd11an1n32x5 FILLER_11_2249 ();
 b15zdnd00an1n02x5 FILLER_11_2281 ();
 b15zdnd00an1n01x5 FILLER_11_2283 ();
 b15zdnd11an1n64x5 FILLER_12_8 ();
 b15zdnd11an1n64x5 FILLER_12_72 ();
 b15zdnd11an1n64x5 FILLER_12_136 ();
 b15zdnd11an1n64x5 FILLER_12_200 ();
 b15zdnd11an1n64x5 FILLER_12_264 ();
 b15zdnd11an1n64x5 FILLER_12_328 ();
 b15zdnd11an1n64x5 FILLER_12_392 ();
 b15zdnd11an1n64x5 FILLER_12_456 ();
 b15zdnd11an1n64x5 FILLER_12_520 ();
 b15zdnd11an1n64x5 FILLER_12_584 ();
 b15zdnd11an1n64x5 FILLER_12_648 ();
 b15zdnd11an1n04x5 FILLER_12_712 ();
 b15zdnd00an1n02x5 FILLER_12_716 ();
 b15zdnd11an1n64x5 FILLER_12_726 ();
 b15zdnd11an1n64x5 FILLER_12_790 ();
 b15zdnd11an1n64x5 FILLER_12_854 ();
 b15zdnd11an1n64x5 FILLER_12_918 ();
 b15zdnd11an1n64x5 FILLER_12_982 ();
 b15zdnd00an1n01x5 FILLER_12_1046 ();
 b15zdnd11an1n08x5 FILLER_12_1050 ();
 b15zdnd11an1n04x5 FILLER_12_1058 ();
 b15zdnd00an1n02x5 FILLER_12_1062 ();
 b15zdnd00an1n01x5 FILLER_12_1064 ();
 b15zdnd11an1n32x5 FILLER_12_1107 ();
 b15zdnd11an1n04x5 FILLER_12_1139 ();
 b15zdnd00an1n01x5 FILLER_12_1143 ();
 b15zdnd11an1n32x5 FILLER_12_1152 ();
 b15zdnd11an1n16x5 FILLER_12_1184 ();
 b15zdnd11an1n08x5 FILLER_12_1200 ();
 b15zdnd00an1n02x5 FILLER_12_1208 ();
 b15zdnd11an1n64x5 FILLER_12_1227 ();
 b15zdnd11an1n08x5 FILLER_12_1291 ();
 b15zdnd00an1n02x5 FILLER_12_1299 ();
 b15zdnd00an1n01x5 FILLER_12_1301 ();
 b15zdnd11an1n64x5 FILLER_12_1316 ();
 b15zdnd11an1n64x5 FILLER_12_1380 ();
 b15zdnd11an1n64x5 FILLER_12_1444 ();
 b15zdnd11an1n64x5 FILLER_12_1508 ();
 b15zdnd11an1n64x5 FILLER_12_1572 ();
 b15zdnd11an1n64x5 FILLER_12_1636 ();
 b15zdnd11an1n64x5 FILLER_12_1700 ();
 b15zdnd11an1n64x5 FILLER_12_1764 ();
 b15zdnd11an1n64x5 FILLER_12_1828 ();
 b15zdnd11an1n64x5 FILLER_12_1892 ();
 b15zdnd11an1n64x5 FILLER_12_1956 ();
 b15zdnd11an1n64x5 FILLER_12_2020 ();
 b15zdnd11an1n64x5 FILLER_12_2084 ();
 b15zdnd11an1n04x5 FILLER_12_2148 ();
 b15zdnd00an1n02x5 FILLER_12_2152 ();
 b15zdnd11an1n64x5 FILLER_12_2162 ();
 b15zdnd11an1n32x5 FILLER_12_2226 ();
 b15zdnd11an1n16x5 FILLER_12_2258 ();
 b15zdnd00an1n02x5 FILLER_12_2274 ();
 b15zdnd11an1n64x5 FILLER_13_0 ();
 b15zdnd11an1n64x5 FILLER_13_64 ();
 b15zdnd11an1n64x5 FILLER_13_128 ();
 b15zdnd11an1n64x5 FILLER_13_192 ();
 b15zdnd11an1n64x5 FILLER_13_256 ();
 b15zdnd11an1n64x5 FILLER_13_320 ();
 b15zdnd11an1n64x5 FILLER_13_384 ();
 b15zdnd11an1n64x5 FILLER_13_448 ();
 b15zdnd11an1n64x5 FILLER_13_512 ();
 b15zdnd11an1n64x5 FILLER_13_576 ();
 b15zdnd11an1n64x5 FILLER_13_640 ();
 b15zdnd11an1n64x5 FILLER_13_704 ();
 b15zdnd11an1n64x5 FILLER_13_768 ();
 b15zdnd11an1n64x5 FILLER_13_832 ();
 b15zdnd11an1n64x5 FILLER_13_896 ();
 b15zdnd11an1n32x5 FILLER_13_960 ();
 b15zdnd11an1n16x5 FILLER_13_992 ();
 b15zdnd11an1n08x5 FILLER_13_1008 ();
 b15zdnd11an1n04x5 FILLER_13_1016 ();
 b15zdnd11an1n32x5 FILLER_13_1072 ();
 b15zdnd11an1n08x5 FILLER_13_1104 ();
 b15zdnd00an1n01x5 FILLER_13_1112 ();
 b15zdnd11an1n64x5 FILLER_13_1155 ();
 b15zdnd11an1n04x5 FILLER_13_1219 ();
 b15zdnd00an1n02x5 FILLER_13_1223 ();
 b15zdnd00an1n01x5 FILLER_13_1225 ();
 b15zdnd11an1n64x5 FILLER_13_1271 ();
 b15zdnd11an1n64x5 FILLER_13_1335 ();
 b15zdnd11an1n16x5 FILLER_13_1399 ();
 b15zdnd11an1n04x5 FILLER_13_1418 ();
 b15zdnd11an1n64x5 FILLER_13_1425 ();
 b15zdnd11an1n64x5 FILLER_13_1489 ();
 b15zdnd11an1n64x5 FILLER_13_1553 ();
 b15zdnd11an1n64x5 FILLER_13_1617 ();
 b15zdnd11an1n64x5 FILLER_13_1681 ();
 b15zdnd11an1n64x5 FILLER_13_1745 ();
 b15zdnd11an1n64x5 FILLER_13_1809 ();
 b15zdnd11an1n64x5 FILLER_13_1873 ();
 b15zdnd11an1n64x5 FILLER_13_1937 ();
 b15zdnd11an1n64x5 FILLER_13_2001 ();
 b15zdnd11an1n64x5 FILLER_13_2065 ();
 b15zdnd11an1n64x5 FILLER_13_2129 ();
 b15zdnd11an1n64x5 FILLER_13_2193 ();
 b15zdnd11an1n16x5 FILLER_13_2257 ();
 b15zdnd11an1n08x5 FILLER_13_2273 ();
 b15zdnd00an1n02x5 FILLER_13_2281 ();
 b15zdnd00an1n01x5 FILLER_13_2283 ();
 b15zdnd11an1n64x5 FILLER_14_8 ();
 b15zdnd11an1n64x5 FILLER_14_72 ();
 b15zdnd11an1n64x5 FILLER_14_136 ();
 b15zdnd11an1n64x5 FILLER_14_200 ();
 b15zdnd11an1n64x5 FILLER_14_264 ();
 b15zdnd11an1n64x5 FILLER_14_328 ();
 b15zdnd11an1n64x5 FILLER_14_392 ();
 b15zdnd11an1n64x5 FILLER_14_456 ();
 b15zdnd11an1n64x5 FILLER_14_520 ();
 b15zdnd11an1n64x5 FILLER_14_584 ();
 b15zdnd11an1n64x5 FILLER_14_648 ();
 b15zdnd11an1n04x5 FILLER_14_712 ();
 b15zdnd00an1n02x5 FILLER_14_716 ();
 b15zdnd11an1n64x5 FILLER_14_726 ();
 b15zdnd11an1n64x5 FILLER_14_790 ();
 b15zdnd11an1n64x5 FILLER_14_854 ();
 b15zdnd11an1n64x5 FILLER_14_918 ();
 b15zdnd11an1n32x5 FILLER_14_982 ();
 b15zdnd11an1n16x5 FILLER_14_1014 ();
 b15zdnd11an1n04x5 FILLER_14_1030 ();
 b15zdnd00an1n02x5 FILLER_14_1034 ();
 b15zdnd00an1n01x5 FILLER_14_1036 ();
 b15zdnd11an1n04x5 FILLER_14_1042 ();
 b15zdnd11an1n64x5 FILLER_14_1049 ();
 b15zdnd11an1n64x5 FILLER_14_1113 ();
 b15zdnd11an1n64x5 FILLER_14_1177 ();
 b15zdnd11an1n64x5 FILLER_14_1241 ();
 b15zdnd11an1n64x5 FILLER_14_1305 ();
 b15zdnd11an1n16x5 FILLER_14_1369 ();
 b15zdnd11an1n08x5 FILLER_14_1385 ();
 b15zdnd11an1n04x5 FILLER_14_1393 ();
 b15zdnd11an1n64x5 FILLER_14_1449 ();
 b15zdnd11an1n16x5 FILLER_14_1513 ();
 b15zdnd11an1n04x5 FILLER_14_1529 ();
 b15zdnd00an1n02x5 FILLER_14_1533 ();
 b15zdnd00an1n01x5 FILLER_14_1535 ();
 b15zdnd11an1n64x5 FILLER_14_1546 ();
 b15zdnd11an1n64x5 FILLER_14_1610 ();
 b15zdnd11an1n64x5 FILLER_14_1674 ();
 b15zdnd11an1n64x5 FILLER_14_1738 ();
 b15zdnd11an1n64x5 FILLER_14_1802 ();
 b15zdnd11an1n64x5 FILLER_14_1866 ();
 b15zdnd11an1n64x5 FILLER_14_1930 ();
 b15zdnd11an1n64x5 FILLER_14_1994 ();
 b15zdnd11an1n64x5 FILLER_14_2058 ();
 b15zdnd11an1n32x5 FILLER_14_2122 ();
 b15zdnd11an1n64x5 FILLER_14_2162 ();
 b15zdnd11an1n32x5 FILLER_14_2226 ();
 b15zdnd11an1n16x5 FILLER_14_2258 ();
 b15zdnd00an1n02x5 FILLER_14_2274 ();
 b15zdnd11an1n64x5 FILLER_15_0 ();
 b15zdnd11an1n64x5 FILLER_15_64 ();
 b15zdnd11an1n64x5 FILLER_15_128 ();
 b15zdnd11an1n64x5 FILLER_15_192 ();
 b15zdnd11an1n64x5 FILLER_15_256 ();
 b15zdnd11an1n64x5 FILLER_15_320 ();
 b15zdnd11an1n64x5 FILLER_15_384 ();
 b15zdnd11an1n64x5 FILLER_15_448 ();
 b15zdnd11an1n64x5 FILLER_15_512 ();
 b15zdnd11an1n64x5 FILLER_15_576 ();
 b15zdnd11an1n64x5 FILLER_15_640 ();
 b15zdnd11an1n64x5 FILLER_15_704 ();
 b15zdnd11an1n64x5 FILLER_15_768 ();
 b15zdnd11an1n64x5 FILLER_15_832 ();
 b15zdnd11an1n64x5 FILLER_15_896 ();
 b15zdnd11an1n64x5 FILLER_15_960 ();
 b15zdnd11an1n16x5 FILLER_15_1024 ();
 b15zdnd11an1n04x5 FILLER_15_1040 ();
 b15zdnd11an1n64x5 FILLER_15_1047 ();
 b15zdnd11an1n64x5 FILLER_15_1111 ();
 b15zdnd11an1n64x5 FILLER_15_1175 ();
 b15zdnd11an1n64x5 FILLER_15_1239 ();
 b15zdnd11an1n64x5 FILLER_15_1303 ();
 b15zdnd11an1n32x5 FILLER_15_1367 ();
 b15zdnd11an1n16x5 FILLER_15_1399 ();
 b15zdnd11an1n04x5 FILLER_15_1415 ();
 b15zdnd00an1n02x5 FILLER_15_1419 ();
 b15zdnd00an1n01x5 FILLER_15_1421 ();
 b15zdnd11an1n64x5 FILLER_15_1425 ();
 b15zdnd11an1n64x5 FILLER_15_1489 ();
 b15zdnd11an1n64x5 FILLER_15_1553 ();
 b15zdnd11an1n08x5 FILLER_15_1617 ();
 b15zdnd11an1n04x5 FILLER_15_1625 ();
 b15zdnd00an1n02x5 FILLER_15_1629 ();
 b15zdnd00an1n01x5 FILLER_15_1631 ();
 b15zdnd11an1n04x5 FILLER_15_1636 ();
 b15zdnd11an1n04x5 FILLER_15_1644 ();
 b15zdnd00an1n02x5 FILLER_15_1648 ();
 b15zdnd11an1n64x5 FILLER_15_1654 ();
 b15zdnd11an1n64x5 FILLER_15_1718 ();
 b15zdnd11an1n64x5 FILLER_15_1782 ();
 b15zdnd11an1n64x5 FILLER_15_1846 ();
 b15zdnd11an1n64x5 FILLER_15_1910 ();
 b15zdnd11an1n64x5 FILLER_15_1974 ();
 b15zdnd11an1n64x5 FILLER_15_2038 ();
 b15zdnd11an1n64x5 FILLER_15_2102 ();
 b15zdnd11an1n64x5 FILLER_15_2166 ();
 b15zdnd11an1n32x5 FILLER_15_2230 ();
 b15zdnd11an1n16x5 FILLER_15_2262 ();
 b15zdnd11an1n04x5 FILLER_15_2278 ();
 b15zdnd00an1n02x5 FILLER_15_2282 ();
 b15zdnd11an1n64x5 FILLER_16_8 ();
 b15zdnd11an1n64x5 FILLER_16_72 ();
 b15zdnd11an1n64x5 FILLER_16_136 ();
 b15zdnd11an1n64x5 FILLER_16_200 ();
 b15zdnd11an1n64x5 FILLER_16_264 ();
 b15zdnd11an1n64x5 FILLER_16_328 ();
 b15zdnd11an1n64x5 FILLER_16_392 ();
 b15zdnd11an1n64x5 FILLER_16_456 ();
 b15zdnd11an1n64x5 FILLER_16_520 ();
 b15zdnd11an1n64x5 FILLER_16_584 ();
 b15zdnd11an1n64x5 FILLER_16_648 ();
 b15zdnd11an1n04x5 FILLER_16_712 ();
 b15zdnd00an1n02x5 FILLER_16_716 ();
 b15zdnd11an1n64x5 FILLER_16_726 ();
 b15zdnd11an1n64x5 FILLER_16_790 ();
 b15zdnd11an1n64x5 FILLER_16_854 ();
 b15zdnd11an1n64x5 FILLER_16_918 ();
 b15zdnd11an1n64x5 FILLER_16_982 ();
 b15zdnd11an1n64x5 FILLER_16_1046 ();
 b15zdnd11an1n64x5 FILLER_16_1110 ();
 b15zdnd11an1n64x5 FILLER_16_1174 ();
 b15zdnd11an1n64x5 FILLER_16_1238 ();
 b15zdnd11an1n64x5 FILLER_16_1302 ();
 b15zdnd11an1n64x5 FILLER_16_1366 ();
 b15zdnd11an1n64x5 FILLER_16_1430 ();
 b15zdnd11an1n64x5 FILLER_16_1494 ();
 b15zdnd11an1n32x5 FILLER_16_1558 ();
 b15zdnd11an1n08x5 FILLER_16_1590 ();
 b15zdnd11an1n04x5 FILLER_16_1598 ();
 b15zdnd00an1n01x5 FILLER_16_1602 ();
 b15zdnd11an1n16x5 FILLER_16_1617 ();
 b15zdnd11an1n08x5 FILLER_16_1633 ();
 b15zdnd00an1n01x5 FILLER_16_1641 ();
 b15zdnd11an1n64x5 FILLER_16_1646 ();
 b15zdnd11an1n64x5 FILLER_16_1710 ();
 b15zdnd11an1n64x5 FILLER_16_1774 ();
 b15zdnd11an1n64x5 FILLER_16_1838 ();
 b15zdnd11an1n64x5 FILLER_16_1902 ();
 b15zdnd11an1n64x5 FILLER_16_1966 ();
 b15zdnd11an1n64x5 FILLER_16_2030 ();
 b15zdnd11an1n32x5 FILLER_16_2094 ();
 b15zdnd11an1n16x5 FILLER_16_2126 ();
 b15zdnd11an1n08x5 FILLER_16_2142 ();
 b15zdnd11an1n04x5 FILLER_16_2150 ();
 b15zdnd11an1n64x5 FILLER_16_2162 ();
 b15zdnd11an1n32x5 FILLER_16_2226 ();
 b15zdnd11an1n16x5 FILLER_16_2258 ();
 b15zdnd00an1n02x5 FILLER_16_2274 ();
 b15zdnd11an1n64x5 FILLER_17_0 ();
 b15zdnd11an1n64x5 FILLER_17_64 ();
 b15zdnd11an1n64x5 FILLER_17_128 ();
 b15zdnd11an1n64x5 FILLER_17_192 ();
 b15zdnd11an1n64x5 FILLER_17_256 ();
 b15zdnd11an1n64x5 FILLER_17_320 ();
 b15zdnd11an1n64x5 FILLER_17_384 ();
 b15zdnd11an1n64x5 FILLER_17_448 ();
 b15zdnd11an1n64x5 FILLER_17_512 ();
 b15zdnd11an1n64x5 FILLER_17_576 ();
 b15zdnd11an1n64x5 FILLER_17_640 ();
 b15zdnd11an1n64x5 FILLER_17_704 ();
 b15zdnd11an1n64x5 FILLER_17_768 ();
 b15zdnd11an1n64x5 FILLER_17_832 ();
 b15zdnd11an1n64x5 FILLER_17_896 ();
 b15zdnd11an1n64x5 FILLER_17_960 ();
 b15zdnd11an1n64x5 FILLER_17_1024 ();
 b15zdnd11an1n64x5 FILLER_17_1088 ();
 b15zdnd11an1n64x5 FILLER_17_1152 ();
 b15zdnd11an1n64x5 FILLER_17_1216 ();
 b15zdnd11an1n64x5 FILLER_17_1280 ();
 b15zdnd11an1n64x5 FILLER_17_1344 ();
 b15zdnd11an1n64x5 FILLER_17_1408 ();
 b15zdnd11an1n64x5 FILLER_17_1472 ();
 b15zdnd11an1n64x5 FILLER_17_1536 ();
 b15zdnd11an1n64x5 FILLER_17_1600 ();
 b15zdnd11an1n64x5 FILLER_17_1664 ();
 b15zdnd11an1n64x5 FILLER_17_1728 ();
 b15zdnd11an1n64x5 FILLER_17_1792 ();
 b15zdnd11an1n64x5 FILLER_17_1856 ();
 b15zdnd11an1n64x5 FILLER_17_1920 ();
 b15zdnd11an1n64x5 FILLER_17_1984 ();
 b15zdnd11an1n64x5 FILLER_17_2048 ();
 b15zdnd11an1n64x5 FILLER_17_2112 ();
 b15zdnd11an1n64x5 FILLER_17_2176 ();
 b15zdnd11an1n32x5 FILLER_17_2240 ();
 b15zdnd11an1n08x5 FILLER_17_2272 ();
 b15zdnd11an1n04x5 FILLER_17_2280 ();
 b15zdnd11an1n64x5 FILLER_18_8 ();
 b15zdnd11an1n64x5 FILLER_18_72 ();
 b15zdnd11an1n64x5 FILLER_18_136 ();
 b15zdnd11an1n64x5 FILLER_18_200 ();
 b15zdnd11an1n64x5 FILLER_18_264 ();
 b15zdnd11an1n64x5 FILLER_18_328 ();
 b15zdnd11an1n64x5 FILLER_18_392 ();
 b15zdnd11an1n64x5 FILLER_18_456 ();
 b15zdnd11an1n64x5 FILLER_18_520 ();
 b15zdnd11an1n64x5 FILLER_18_584 ();
 b15zdnd11an1n64x5 FILLER_18_648 ();
 b15zdnd11an1n04x5 FILLER_18_712 ();
 b15zdnd00an1n02x5 FILLER_18_716 ();
 b15zdnd11an1n64x5 FILLER_18_726 ();
 b15zdnd11an1n64x5 FILLER_18_790 ();
 b15zdnd11an1n64x5 FILLER_18_854 ();
 b15zdnd11an1n64x5 FILLER_18_918 ();
 b15zdnd11an1n16x5 FILLER_18_982 ();
 b15zdnd11an1n08x5 FILLER_18_998 ();
 b15zdnd11an1n04x5 FILLER_18_1006 ();
 b15zdnd11an1n64x5 FILLER_18_1017 ();
 b15zdnd11an1n64x5 FILLER_18_1081 ();
 b15zdnd11an1n64x5 FILLER_18_1145 ();
 b15zdnd11an1n16x5 FILLER_18_1209 ();
 b15zdnd11an1n08x5 FILLER_18_1225 ();
 b15zdnd00an1n02x5 FILLER_18_1233 ();
 b15zdnd11an1n64x5 FILLER_18_1238 ();
 b15zdnd11an1n64x5 FILLER_18_1302 ();
 b15zdnd11an1n64x5 FILLER_18_1366 ();
 b15zdnd11an1n64x5 FILLER_18_1430 ();
 b15zdnd11an1n64x5 FILLER_18_1494 ();
 b15zdnd11an1n64x5 FILLER_18_1558 ();
 b15zdnd11an1n64x5 FILLER_18_1622 ();
 b15zdnd11an1n64x5 FILLER_18_1686 ();
 b15zdnd11an1n64x5 FILLER_18_1750 ();
 b15zdnd11an1n64x5 FILLER_18_1814 ();
 b15zdnd11an1n64x5 FILLER_18_1878 ();
 b15zdnd11an1n64x5 FILLER_18_1942 ();
 b15zdnd11an1n64x5 FILLER_18_2006 ();
 b15zdnd11an1n64x5 FILLER_18_2070 ();
 b15zdnd11an1n16x5 FILLER_18_2134 ();
 b15zdnd11an1n04x5 FILLER_18_2150 ();
 b15zdnd11an1n64x5 FILLER_18_2162 ();
 b15zdnd11an1n32x5 FILLER_18_2226 ();
 b15zdnd11an1n16x5 FILLER_18_2258 ();
 b15zdnd00an1n02x5 FILLER_18_2274 ();
 b15zdnd11an1n64x5 FILLER_19_0 ();
 b15zdnd11an1n64x5 FILLER_19_64 ();
 b15zdnd11an1n64x5 FILLER_19_128 ();
 b15zdnd11an1n64x5 FILLER_19_192 ();
 b15zdnd11an1n64x5 FILLER_19_256 ();
 b15zdnd11an1n64x5 FILLER_19_320 ();
 b15zdnd11an1n64x5 FILLER_19_384 ();
 b15zdnd11an1n64x5 FILLER_19_448 ();
 b15zdnd11an1n64x5 FILLER_19_512 ();
 b15zdnd11an1n64x5 FILLER_19_576 ();
 b15zdnd11an1n64x5 FILLER_19_640 ();
 b15zdnd11an1n64x5 FILLER_19_704 ();
 b15zdnd11an1n64x5 FILLER_19_768 ();
 b15zdnd11an1n64x5 FILLER_19_832 ();
 b15zdnd11an1n64x5 FILLER_19_896 ();
 b15zdnd11an1n64x5 FILLER_19_960 ();
 b15zdnd11an1n64x5 FILLER_19_1024 ();
 b15zdnd11an1n64x5 FILLER_19_1088 ();
 b15zdnd11an1n64x5 FILLER_19_1152 ();
 b15zdnd11an1n16x5 FILLER_19_1216 ();
 b15zdnd00an1n02x5 FILLER_19_1232 ();
 b15zdnd11an1n64x5 FILLER_19_1237 ();
 b15zdnd11an1n64x5 FILLER_19_1301 ();
 b15zdnd11an1n64x5 FILLER_19_1365 ();
 b15zdnd11an1n64x5 FILLER_19_1429 ();
 b15zdnd11an1n64x5 FILLER_19_1493 ();
 b15zdnd11an1n64x5 FILLER_19_1557 ();
 b15zdnd11an1n64x5 FILLER_19_1621 ();
 b15zdnd11an1n64x5 FILLER_19_1685 ();
 b15zdnd11an1n64x5 FILLER_19_1749 ();
 b15zdnd11an1n64x5 FILLER_19_1813 ();
 b15zdnd11an1n64x5 FILLER_19_1877 ();
 b15zdnd11an1n64x5 FILLER_19_1941 ();
 b15zdnd11an1n64x5 FILLER_19_2005 ();
 b15zdnd11an1n64x5 FILLER_19_2069 ();
 b15zdnd11an1n64x5 FILLER_19_2133 ();
 b15zdnd11an1n64x5 FILLER_19_2197 ();
 b15zdnd11an1n16x5 FILLER_19_2261 ();
 b15zdnd11an1n04x5 FILLER_19_2277 ();
 b15zdnd00an1n02x5 FILLER_19_2281 ();
 b15zdnd00an1n01x5 FILLER_19_2283 ();
 b15zdnd11an1n64x5 FILLER_20_8 ();
 b15zdnd11an1n64x5 FILLER_20_72 ();
 b15zdnd11an1n64x5 FILLER_20_136 ();
 b15zdnd11an1n64x5 FILLER_20_200 ();
 b15zdnd11an1n64x5 FILLER_20_264 ();
 b15zdnd11an1n64x5 FILLER_20_328 ();
 b15zdnd11an1n64x5 FILLER_20_392 ();
 b15zdnd11an1n64x5 FILLER_20_456 ();
 b15zdnd11an1n16x5 FILLER_20_520 ();
 b15zdnd00an1n02x5 FILLER_20_536 ();
 b15zdnd11an1n64x5 FILLER_20_542 ();
 b15zdnd11an1n64x5 FILLER_20_606 ();
 b15zdnd11an1n32x5 FILLER_20_670 ();
 b15zdnd11an1n16x5 FILLER_20_702 ();
 b15zdnd11an1n64x5 FILLER_20_726 ();
 b15zdnd11an1n64x5 FILLER_20_790 ();
 b15zdnd11an1n64x5 FILLER_20_854 ();
 b15zdnd11an1n32x5 FILLER_20_918 ();
 b15zdnd11an1n08x5 FILLER_20_950 ();
 b15zdnd11an1n04x5 FILLER_20_958 ();
 b15zdnd00an1n01x5 FILLER_20_962 ();
 b15zdnd11an1n64x5 FILLER_20_969 ();
 b15zdnd11an1n64x5 FILLER_20_1033 ();
 b15zdnd11an1n64x5 FILLER_20_1097 ();
 b15zdnd11an1n32x5 FILLER_20_1161 ();
 b15zdnd11an1n16x5 FILLER_20_1193 ();
 b15zdnd11an1n16x5 FILLER_20_1261 ();
 b15zdnd00an1n02x5 FILLER_20_1277 ();
 b15zdnd11an1n64x5 FILLER_20_1286 ();
 b15zdnd11an1n64x5 FILLER_20_1350 ();
 b15zdnd11an1n64x5 FILLER_20_1414 ();
 b15zdnd11an1n64x5 FILLER_20_1478 ();
 b15zdnd11an1n64x5 FILLER_20_1542 ();
 b15zdnd11an1n64x5 FILLER_20_1606 ();
 b15zdnd11an1n64x5 FILLER_20_1670 ();
 b15zdnd11an1n64x5 FILLER_20_1734 ();
 b15zdnd11an1n64x5 FILLER_20_1798 ();
 b15zdnd11an1n64x5 FILLER_20_1862 ();
 b15zdnd11an1n64x5 FILLER_20_1926 ();
 b15zdnd11an1n64x5 FILLER_20_1990 ();
 b15zdnd11an1n64x5 FILLER_20_2054 ();
 b15zdnd11an1n32x5 FILLER_20_2118 ();
 b15zdnd11an1n04x5 FILLER_20_2150 ();
 b15zdnd11an1n64x5 FILLER_20_2162 ();
 b15zdnd11an1n32x5 FILLER_20_2226 ();
 b15zdnd11an1n16x5 FILLER_20_2258 ();
 b15zdnd00an1n02x5 FILLER_20_2274 ();
 b15zdnd11an1n64x5 FILLER_21_0 ();
 b15zdnd11an1n64x5 FILLER_21_64 ();
 b15zdnd11an1n64x5 FILLER_21_128 ();
 b15zdnd11an1n64x5 FILLER_21_192 ();
 b15zdnd11an1n64x5 FILLER_21_256 ();
 b15zdnd11an1n64x5 FILLER_21_320 ();
 b15zdnd11an1n64x5 FILLER_21_384 ();
 b15zdnd11an1n64x5 FILLER_21_448 ();
 b15zdnd11an1n64x5 FILLER_21_512 ();
 b15zdnd11an1n64x5 FILLER_21_576 ();
 b15zdnd11an1n08x5 FILLER_21_640 ();
 b15zdnd00an1n02x5 FILLER_21_648 ();
 b15zdnd00an1n01x5 FILLER_21_650 ();
 b15zdnd11an1n64x5 FILLER_21_655 ();
 b15zdnd11an1n64x5 FILLER_21_719 ();
 b15zdnd11an1n64x5 FILLER_21_783 ();
 b15zdnd11an1n64x5 FILLER_21_847 ();
 b15zdnd11an1n64x5 FILLER_21_911 ();
 b15zdnd11an1n64x5 FILLER_21_975 ();
 b15zdnd11an1n64x5 FILLER_21_1039 ();
 b15zdnd11an1n64x5 FILLER_21_1103 ();
 b15zdnd11an1n64x5 FILLER_21_1167 ();
 b15zdnd00an1n02x5 FILLER_21_1231 ();
 b15zdnd00an1n01x5 FILLER_21_1233 ();
 b15zdnd11an1n04x5 FILLER_21_1237 ();
 b15zdnd00an1n02x5 FILLER_21_1241 ();
 b15zdnd11an1n64x5 FILLER_21_1250 ();
 b15zdnd11an1n64x5 FILLER_21_1314 ();
 b15zdnd11an1n64x5 FILLER_21_1378 ();
 b15zdnd11an1n64x5 FILLER_21_1442 ();
 b15zdnd11an1n64x5 FILLER_21_1506 ();
 b15zdnd11an1n64x5 FILLER_21_1570 ();
 b15zdnd11an1n64x5 FILLER_21_1634 ();
 b15zdnd11an1n64x5 FILLER_21_1698 ();
 b15zdnd11an1n64x5 FILLER_21_1762 ();
 b15zdnd11an1n64x5 FILLER_21_1826 ();
 b15zdnd11an1n64x5 FILLER_21_1890 ();
 b15zdnd11an1n64x5 FILLER_21_1954 ();
 b15zdnd11an1n64x5 FILLER_21_2018 ();
 b15zdnd11an1n64x5 FILLER_21_2082 ();
 b15zdnd11an1n64x5 FILLER_21_2146 ();
 b15zdnd11an1n64x5 FILLER_21_2210 ();
 b15zdnd11an1n08x5 FILLER_21_2274 ();
 b15zdnd00an1n02x5 FILLER_21_2282 ();
 b15zdnd11an1n64x5 FILLER_22_8 ();
 b15zdnd11an1n64x5 FILLER_22_72 ();
 b15zdnd11an1n64x5 FILLER_22_136 ();
 b15zdnd11an1n64x5 FILLER_22_200 ();
 b15zdnd11an1n64x5 FILLER_22_264 ();
 b15zdnd11an1n64x5 FILLER_22_328 ();
 b15zdnd11an1n64x5 FILLER_22_392 ();
 b15zdnd11an1n64x5 FILLER_22_456 ();
 b15zdnd11an1n16x5 FILLER_22_520 ();
 b15zdnd11an1n08x5 FILLER_22_536 ();
 b15zdnd11an1n64x5 FILLER_22_548 ();
 b15zdnd11an1n32x5 FILLER_22_612 ();
 b15zdnd11an1n16x5 FILLER_22_644 ();
 b15zdnd11an1n04x5 FILLER_22_660 ();
 b15zdnd00an1n01x5 FILLER_22_664 ();
 b15zdnd11an1n32x5 FILLER_22_669 ();
 b15zdnd11an1n16x5 FILLER_22_701 ();
 b15zdnd00an1n01x5 FILLER_22_717 ();
 b15zdnd11an1n64x5 FILLER_22_726 ();
 b15zdnd11an1n64x5 FILLER_22_790 ();
 b15zdnd11an1n64x5 FILLER_22_854 ();
 b15zdnd11an1n64x5 FILLER_22_918 ();
 b15zdnd11an1n64x5 FILLER_22_982 ();
 b15zdnd11an1n64x5 FILLER_22_1046 ();
 b15zdnd11an1n64x5 FILLER_22_1110 ();
 b15zdnd11an1n64x5 FILLER_22_1174 ();
 b15zdnd11an1n64x5 FILLER_22_1238 ();
 b15zdnd11an1n64x5 FILLER_22_1302 ();
 b15zdnd11an1n64x5 FILLER_22_1366 ();
 b15zdnd11an1n64x5 FILLER_22_1430 ();
 b15zdnd11an1n64x5 FILLER_22_1494 ();
 b15zdnd11an1n64x5 FILLER_22_1558 ();
 b15zdnd11an1n64x5 FILLER_22_1622 ();
 b15zdnd11an1n64x5 FILLER_22_1686 ();
 b15zdnd11an1n64x5 FILLER_22_1750 ();
 b15zdnd11an1n64x5 FILLER_22_1814 ();
 b15zdnd11an1n64x5 FILLER_22_1878 ();
 b15zdnd11an1n64x5 FILLER_22_1942 ();
 b15zdnd11an1n64x5 FILLER_22_2006 ();
 b15zdnd11an1n64x5 FILLER_22_2070 ();
 b15zdnd11an1n16x5 FILLER_22_2134 ();
 b15zdnd11an1n04x5 FILLER_22_2150 ();
 b15zdnd11an1n64x5 FILLER_22_2162 ();
 b15zdnd11an1n32x5 FILLER_22_2226 ();
 b15zdnd11an1n16x5 FILLER_22_2258 ();
 b15zdnd00an1n02x5 FILLER_22_2274 ();
 b15zdnd11an1n64x5 FILLER_23_0 ();
 b15zdnd11an1n64x5 FILLER_23_64 ();
 b15zdnd11an1n64x5 FILLER_23_128 ();
 b15zdnd11an1n64x5 FILLER_23_192 ();
 b15zdnd11an1n64x5 FILLER_23_256 ();
 b15zdnd11an1n64x5 FILLER_23_320 ();
 b15zdnd11an1n64x5 FILLER_23_384 ();
 b15zdnd11an1n64x5 FILLER_23_448 ();
 b15zdnd11an1n64x5 FILLER_23_512 ();
 b15zdnd11an1n64x5 FILLER_23_576 ();
 b15zdnd11an1n64x5 FILLER_23_640 ();
 b15zdnd11an1n64x5 FILLER_23_704 ();
 b15zdnd11an1n64x5 FILLER_23_768 ();
 b15zdnd11an1n64x5 FILLER_23_832 ();
 b15zdnd11an1n64x5 FILLER_23_896 ();
 b15zdnd11an1n64x5 FILLER_23_960 ();
 b15zdnd11an1n64x5 FILLER_23_1024 ();
 b15zdnd11an1n16x5 FILLER_23_1088 ();
 b15zdnd11an1n04x5 FILLER_23_1104 ();
 b15zdnd11an1n08x5 FILLER_23_1113 ();
 b15zdnd11an1n64x5 FILLER_23_1124 ();
 b15zdnd11an1n64x5 FILLER_23_1188 ();
 b15zdnd11an1n64x5 FILLER_23_1252 ();
 b15zdnd11an1n64x5 FILLER_23_1316 ();
 b15zdnd11an1n64x5 FILLER_23_1380 ();
 b15zdnd11an1n64x5 FILLER_23_1444 ();
 b15zdnd11an1n64x5 FILLER_23_1508 ();
 b15zdnd11an1n64x5 FILLER_23_1572 ();
 b15zdnd11an1n64x5 FILLER_23_1636 ();
 b15zdnd11an1n64x5 FILLER_23_1700 ();
 b15zdnd11an1n64x5 FILLER_23_1764 ();
 b15zdnd11an1n64x5 FILLER_23_1828 ();
 b15zdnd11an1n64x5 FILLER_23_1892 ();
 b15zdnd11an1n64x5 FILLER_23_1956 ();
 b15zdnd11an1n64x5 FILLER_23_2020 ();
 b15zdnd11an1n64x5 FILLER_23_2084 ();
 b15zdnd11an1n64x5 FILLER_23_2148 ();
 b15zdnd11an1n64x5 FILLER_23_2212 ();
 b15zdnd11an1n08x5 FILLER_23_2276 ();
 b15zdnd11an1n64x5 FILLER_24_8 ();
 b15zdnd11an1n64x5 FILLER_24_72 ();
 b15zdnd11an1n64x5 FILLER_24_136 ();
 b15zdnd11an1n64x5 FILLER_24_200 ();
 b15zdnd11an1n64x5 FILLER_24_264 ();
 b15zdnd11an1n64x5 FILLER_24_328 ();
 b15zdnd11an1n64x5 FILLER_24_392 ();
 b15zdnd11an1n64x5 FILLER_24_456 ();
 b15zdnd11an1n64x5 FILLER_24_520 ();
 b15zdnd11an1n64x5 FILLER_24_584 ();
 b15zdnd11an1n64x5 FILLER_24_648 ();
 b15zdnd11an1n04x5 FILLER_24_712 ();
 b15zdnd00an1n02x5 FILLER_24_716 ();
 b15zdnd11an1n64x5 FILLER_24_726 ();
 b15zdnd11an1n32x5 FILLER_24_790 ();
 b15zdnd11an1n08x5 FILLER_24_822 ();
 b15zdnd11an1n04x5 FILLER_24_830 ();
 b15zdnd00an1n01x5 FILLER_24_834 ();
 b15zdnd11an1n64x5 FILLER_24_839 ();
 b15zdnd11an1n64x5 FILLER_24_903 ();
 b15zdnd11an1n64x5 FILLER_24_967 ();
 b15zdnd11an1n32x5 FILLER_24_1031 ();
 b15zdnd11an1n08x5 FILLER_24_1063 ();
 b15zdnd11an1n04x5 FILLER_24_1071 ();
 b15zdnd00an1n01x5 FILLER_24_1075 ();
 b15zdnd11an1n04x5 FILLER_24_1083 ();
 b15zdnd11an1n64x5 FILLER_24_1139 ();
 b15zdnd11an1n64x5 FILLER_24_1203 ();
 b15zdnd11an1n64x5 FILLER_24_1267 ();
 b15zdnd11an1n64x5 FILLER_24_1331 ();
 b15zdnd11an1n64x5 FILLER_24_1395 ();
 b15zdnd11an1n64x5 FILLER_24_1459 ();
 b15zdnd11an1n64x5 FILLER_24_1523 ();
 b15zdnd11an1n64x5 FILLER_24_1587 ();
 b15zdnd11an1n64x5 FILLER_24_1651 ();
 b15zdnd11an1n64x5 FILLER_24_1715 ();
 b15zdnd11an1n64x5 FILLER_24_1779 ();
 b15zdnd11an1n64x5 FILLER_24_1843 ();
 b15zdnd11an1n64x5 FILLER_24_1907 ();
 b15zdnd11an1n64x5 FILLER_24_1971 ();
 b15zdnd11an1n64x5 FILLER_24_2035 ();
 b15zdnd11an1n32x5 FILLER_24_2099 ();
 b15zdnd11an1n16x5 FILLER_24_2131 ();
 b15zdnd11an1n04x5 FILLER_24_2147 ();
 b15zdnd00an1n02x5 FILLER_24_2151 ();
 b15zdnd00an1n01x5 FILLER_24_2153 ();
 b15zdnd11an1n64x5 FILLER_24_2162 ();
 b15zdnd11an1n32x5 FILLER_24_2226 ();
 b15zdnd11an1n16x5 FILLER_24_2258 ();
 b15zdnd00an1n02x5 FILLER_24_2274 ();
 b15zdnd11an1n64x5 FILLER_25_0 ();
 b15zdnd11an1n64x5 FILLER_25_64 ();
 b15zdnd11an1n64x5 FILLER_25_128 ();
 b15zdnd11an1n64x5 FILLER_25_192 ();
 b15zdnd11an1n64x5 FILLER_25_256 ();
 b15zdnd11an1n64x5 FILLER_25_320 ();
 b15zdnd11an1n64x5 FILLER_25_384 ();
 b15zdnd11an1n64x5 FILLER_25_448 ();
 b15zdnd11an1n64x5 FILLER_25_512 ();
 b15zdnd11an1n64x5 FILLER_25_576 ();
 b15zdnd11an1n64x5 FILLER_25_640 ();
 b15zdnd11an1n64x5 FILLER_25_704 ();
 b15zdnd11an1n32x5 FILLER_25_768 ();
 b15zdnd11an1n04x5 FILLER_25_800 ();
 b15zdnd11an1n04x5 FILLER_25_815 ();
 b15zdnd11an1n64x5 FILLER_25_823 ();
 b15zdnd11an1n64x5 FILLER_25_887 ();
 b15zdnd11an1n64x5 FILLER_25_951 ();
 b15zdnd11an1n64x5 FILLER_25_1015 ();
 b15zdnd11an1n08x5 FILLER_25_1079 ();
 b15zdnd11an1n04x5 FILLER_25_1087 ();
 b15zdnd00an1n02x5 FILLER_25_1091 ();
 b15zdnd00an1n01x5 FILLER_25_1093 ();
 b15zdnd11an1n32x5 FILLER_25_1101 ();
 b15zdnd11an1n08x5 FILLER_25_1133 ();
 b15zdnd11an1n04x5 FILLER_25_1141 ();
 b15zdnd00an1n01x5 FILLER_25_1145 ();
 b15zdnd11an1n04x5 FILLER_25_1154 ();
 b15zdnd11an1n64x5 FILLER_25_1161 ();
 b15zdnd11an1n64x5 FILLER_25_1225 ();
 b15zdnd11an1n64x5 FILLER_25_1289 ();
 b15zdnd11an1n64x5 FILLER_25_1353 ();
 b15zdnd11an1n64x5 FILLER_25_1417 ();
 b15zdnd11an1n64x5 FILLER_25_1481 ();
 b15zdnd11an1n64x5 FILLER_25_1545 ();
 b15zdnd11an1n64x5 FILLER_25_1609 ();
 b15zdnd11an1n64x5 FILLER_25_1673 ();
 b15zdnd11an1n64x5 FILLER_25_1737 ();
 b15zdnd11an1n64x5 FILLER_25_1801 ();
 b15zdnd11an1n64x5 FILLER_25_1865 ();
 b15zdnd11an1n64x5 FILLER_25_1929 ();
 b15zdnd11an1n64x5 FILLER_25_1993 ();
 b15zdnd11an1n64x5 FILLER_25_2057 ();
 b15zdnd11an1n64x5 FILLER_25_2121 ();
 b15zdnd11an1n64x5 FILLER_25_2185 ();
 b15zdnd11an1n32x5 FILLER_25_2249 ();
 b15zdnd00an1n02x5 FILLER_25_2281 ();
 b15zdnd00an1n01x5 FILLER_25_2283 ();
 b15zdnd11an1n64x5 FILLER_26_8 ();
 b15zdnd11an1n64x5 FILLER_26_72 ();
 b15zdnd11an1n64x5 FILLER_26_136 ();
 b15zdnd11an1n64x5 FILLER_26_200 ();
 b15zdnd11an1n64x5 FILLER_26_264 ();
 b15zdnd11an1n64x5 FILLER_26_328 ();
 b15zdnd11an1n64x5 FILLER_26_392 ();
 b15zdnd11an1n64x5 FILLER_26_456 ();
 b15zdnd11an1n64x5 FILLER_26_520 ();
 b15zdnd11an1n64x5 FILLER_26_584 ();
 b15zdnd11an1n64x5 FILLER_26_648 ();
 b15zdnd11an1n04x5 FILLER_26_712 ();
 b15zdnd00an1n02x5 FILLER_26_716 ();
 b15zdnd11an1n64x5 FILLER_26_726 ();
 b15zdnd11an1n64x5 FILLER_26_790 ();
 b15zdnd11an1n64x5 FILLER_26_854 ();
 b15zdnd11an1n64x5 FILLER_26_918 ();
 b15zdnd11an1n64x5 FILLER_26_982 ();
 b15zdnd11an1n32x5 FILLER_26_1046 ();
 b15zdnd11an1n16x5 FILLER_26_1078 ();
 b15zdnd11an1n08x5 FILLER_26_1094 ();
 b15zdnd11an1n16x5 FILLER_26_1107 ();
 b15zdnd11an1n08x5 FILLER_26_1123 ();
 b15zdnd00an1n02x5 FILLER_26_1131 ();
 b15zdnd00an1n01x5 FILLER_26_1133 ();
 b15zdnd11an1n08x5 FILLER_26_1137 ();
 b15zdnd00an1n02x5 FILLER_26_1145 ();
 b15zdnd00an1n01x5 FILLER_26_1147 ();
 b15zdnd11an1n64x5 FILLER_26_1155 ();
 b15zdnd11an1n64x5 FILLER_26_1219 ();
 b15zdnd11an1n64x5 FILLER_26_1283 ();
 b15zdnd11an1n64x5 FILLER_26_1347 ();
 b15zdnd11an1n64x5 FILLER_26_1411 ();
 b15zdnd11an1n64x5 FILLER_26_1475 ();
 b15zdnd11an1n64x5 FILLER_26_1539 ();
 b15zdnd11an1n64x5 FILLER_26_1603 ();
 b15zdnd11an1n64x5 FILLER_26_1667 ();
 b15zdnd11an1n64x5 FILLER_26_1731 ();
 b15zdnd11an1n64x5 FILLER_26_1795 ();
 b15zdnd11an1n64x5 FILLER_26_1859 ();
 b15zdnd11an1n64x5 FILLER_26_1923 ();
 b15zdnd11an1n64x5 FILLER_26_1987 ();
 b15zdnd11an1n64x5 FILLER_26_2051 ();
 b15zdnd11an1n32x5 FILLER_26_2115 ();
 b15zdnd11an1n04x5 FILLER_26_2147 ();
 b15zdnd00an1n02x5 FILLER_26_2151 ();
 b15zdnd00an1n01x5 FILLER_26_2153 ();
 b15zdnd11an1n64x5 FILLER_26_2162 ();
 b15zdnd11an1n32x5 FILLER_26_2226 ();
 b15zdnd11an1n16x5 FILLER_26_2258 ();
 b15zdnd00an1n02x5 FILLER_26_2274 ();
 b15zdnd11an1n64x5 FILLER_27_0 ();
 b15zdnd11an1n64x5 FILLER_27_64 ();
 b15zdnd11an1n64x5 FILLER_27_128 ();
 b15zdnd11an1n64x5 FILLER_27_192 ();
 b15zdnd11an1n64x5 FILLER_27_256 ();
 b15zdnd11an1n64x5 FILLER_27_320 ();
 b15zdnd11an1n64x5 FILLER_27_384 ();
 b15zdnd11an1n64x5 FILLER_27_448 ();
 b15zdnd11an1n16x5 FILLER_27_512 ();
 b15zdnd11an1n04x5 FILLER_27_528 ();
 b15zdnd00an1n01x5 FILLER_27_532 ();
 b15zdnd11an1n04x5 FILLER_27_536 ();
 b15zdnd11an1n64x5 FILLER_27_543 ();
 b15zdnd11an1n32x5 FILLER_27_607 ();
 b15zdnd11an1n16x5 FILLER_27_639 ();
 b15zdnd11an1n04x5 FILLER_27_655 ();
 b15zdnd00an1n02x5 FILLER_27_659 ();
 b15zdnd00an1n01x5 FILLER_27_661 ();
 b15zdnd11an1n64x5 FILLER_27_665 ();
 b15zdnd11an1n64x5 FILLER_27_729 ();
 b15zdnd11an1n64x5 FILLER_27_793 ();
 b15zdnd11an1n64x5 FILLER_27_857 ();
 b15zdnd11an1n64x5 FILLER_27_921 ();
 b15zdnd11an1n16x5 FILLER_27_985 ();
 b15zdnd11an1n04x5 FILLER_27_1001 ();
 b15zdnd00an1n02x5 FILLER_27_1005 ();
 b15zdnd11an1n64x5 FILLER_27_1011 ();
 b15zdnd11an1n64x5 FILLER_27_1075 ();
 b15zdnd11an1n64x5 FILLER_27_1139 ();
 b15zdnd11an1n64x5 FILLER_27_1203 ();
 b15zdnd11an1n64x5 FILLER_27_1267 ();
 b15zdnd11an1n64x5 FILLER_27_1331 ();
 b15zdnd11an1n64x5 FILLER_27_1395 ();
 b15zdnd11an1n32x5 FILLER_27_1459 ();
 b15zdnd11an1n16x5 FILLER_27_1491 ();
 b15zdnd11an1n08x5 FILLER_27_1507 ();
 b15zdnd00an1n02x5 FILLER_27_1515 ();
 b15zdnd00an1n01x5 FILLER_27_1517 ();
 b15zdnd11an1n04x5 FILLER_27_1521 ();
 b15zdnd11an1n64x5 FILLER_27_1528 ();
 b15zdnd11an1n64x5 FILLER_27_1592 ();
 b15zdnd11an1n64x5 FILLER_27_1656 ();
 b15zdnd11an1n64x5 FILLER_27_1720 ();
 b15zdnd11an1n64x5 FILLER_27_1784 ();
 b15zdnd11an1n64x5 FILLER_27_1848 ();
 b15zdnd11an1n64x5 FILLER_27_1912 ();
 b15zdnd11an1n64x5 FILLER_27_1976 ();
 b15zdnd11an1n64x5 FILLER_27_2040 ();
 b15zdnd11an1n64x5 FILLER_27_2104 ();
 b15zdnd11an1n64x5 FILLER_27_2168 ();
 b15zdnd11an1n32x5 FILLER_27_2232 ();
 b15zdnd11an1n16x5 FILLER_27_2264 ();
 b15zdnd11an1n04x5 FILLER_27_2280 ();
 b15zdnd11an1n64x5 FILLER_28_8 ();
 b15zdnd11an1n64x5 FILLER_28_72 ();
 b15zdnd11an1n64x5 FILLER_28_136 ();
 b15zdnd11an1n64x5 FILLER_28_200 ();
 b15zdnd11an1n64x5 FILLER_28_264 ();
 b15zdnd11an1n64x5 FILLER_28_328 ();
 b15zdnd11an1n64x5 FILLER_28_392 ();
 b15zdnd11an1n32x5 FILLER_28_456 ();
 b15zdnd11an1n16x5 FILLER_28_488 ();
 b15zdnd11an1n08x5 FILLER_28_504 ();
 b15zdnd00an1n01x5 FILLER_28_512 ();
 b15zdnd11an1n64x5 FILLER_28_565 ();
 b15zdnd11an1n04x5 FILLER_28_629 ();
 b15zdnd00an1n02x5 FILLER_28_633 ();
 b15zdnd11an1n16x5 FILLER_28_687 ();
 b15zdnd11an1n08x5 FILLER_28_703 ();
 b15zdnd11an1n04x5 FILLER_28_711 ();
 b15zdnd00an1n02x5 FILLER_28_715 ();
 b15zdnd00an1n01x5 FILLER_28_717 ();
 b15zdnd11an1n64x5 FILLER_28_726 ();
 b15zdnd11an1n64x5 FILLER_28_790 ();
 b15zdnd11an1n64x5 FILLER_28_854 ();
 b15zdnd11an1n64x5 FILLER_28_918 ();
 b15zdnd11an1n64x5 FILLER_28_982 ();
 b15zdnd11an1n64x5 FILLER_28_1046 ();
 b15zdnd11an1n64x5 FILLER_28_1110 ();
 b15zdnd11an1n64x5 FILLER_28_1174 ();
 b15zdnd11an1n64x5 FILLER_28_1238 ();
 b15zdnd11an1n16x5 FILLER_28_1302 ();
 b15zdnd11an1n08x5 FILLER_28_1318 ();
 b15zdnd00an1n02x5 FILLER_28_1326 ();
 b15zdnd00an1n01x5 FILLER_28_1328 ();
 b15zdnd11an1n64x5 FILLER_28_1332 ();
 b15zdnd11an1n64x5 FILLER_28_1396 ();
 b15zdnd11an1n32x5 FILLER_28_1460 ();
 b15zdnd11an1n04x5 FILLER_28_1492 ();
 b15zdnd11an1n64x5 FILLER_28_1540 ();
 b15zdnd11an1n64x5 FILLER_28_1604 ();
 b15zdnd11an1n64x5 FILLER_28_1668 ();
 b15zdnd11an1n64x5 FILLER_28_1732 ();
 b15zdnd11an1n64x5 FILLER_28_1796 ();
 b15zdnd11an1n64x5 FILLER_28_1860 ();
 b15zdnd11an1n64x5 FILLER_28_1924 ();
 b15zdnd11an1n64x5 FILLER_28_1988 ();
 b15zdnd11an1n64x5 FILLER_28_2052 ();
 b15zdnd11an1n32x5 FILLER_28_2116 ();
 b15zdnd11an1n04x5 FILLER_28_2148 ();
 b15zdnd00an1n02x5 FILLER_28_2152 ();
 b15zdnd11an1n64x5 FILLER_28_2162 ();
 b15zdnd11an1n32x5 FILLER_28_2226 ();
 b15zdnd11an1n16x5 FILLER_28_2258 ();
 b15zdnd00an1n02x5 FILLER_28_2274 ();
 b15zdnd11an1n64x5 FILLER_29_0 ();
 b15zdnd11an1n64x5 FILLER_29_64 ();
 b15zdnd11an1n64x5 FILLER_29_128 ();
 b15zdnd11an1n64x5 FILLER_29_192 ();
 b15zdnd11an1n64x5 FILLER_29_256 ();
 b15zdnd11an1n64x5 FILLER_29_320 ();
 b15zdnd11an1n64x5 FILLER_29_384 ();
 b15zdnd11an1n64x5 FILLER_29_448 ();
 b15zdnd11an1n16x5 FILLER_29_512 ();
 b15zdnd11an1n08x5 FILLER_29_528 ();
 b15zdnd00an1n02x5 FILLER_29_536 ();
 b15zdnd11an1n08x5 FILLER_29_541 ();
 b15zdnd00an1n01x5 FILLER_29_549 ();
 b15zdnd11an1n04x5 FILLER_29_553 ();
 b15zdnd11an1n64x5 FILLER_29_584 ();
 b15zdnd11an1n04x5 FILLER_29_648 ();
 b15zdnd00an1n01x5 FILLER_29_652 ();
 b15zdnd11an1n04x5 FILLER_29_656 ();
 b15zdnd11an1n64x5 FILLER_29_663 ();
 b15zdnd11an1n64x5 FILLER_29_727 ();
 b15zdnd11an1n64x5 FILLER_29_791 ();
 b15zdnd11an1n64x5 FILLER_29_855 ();
 b15zdnd11an1n64x5 FILLER_29_919 ();
 b15zdnd11an1n64x5 FILLER_29_983 ();
 b15zdnd11an1n64x5 FILLER_29_1047 ();
 b15zdnd11an1n64x5 FILLER_29_1111 ();
 b15zdnd11an1n64x5 FILLER_29_1175 ();
 b15zdnd11an1n64x5 FILLER_29_1239 ();
 b15zdnd11an1n16x5 FILLER_29_1303 ();
 b15zdnd11an1n08x5 FILLER_29_1319 ();
 b15zdnd00an1n02x5 FILLER_29_1327 ();
 b15zdnd00an1n01x5 FILLER_29_1329 ();
 b15zdnd11an1n04x5 FILLER_29_1333 ();
 b15zdnd11an1n64x5 FILLER_29_1340 ();
 b15zdnd11an1n64x5 FILLER_29_1404 ();
 b15zdnd11an1n16x5 FILLER_29_1468 ();
 b15zdnd11an1n08x5 FILLER_29_1484 ();
 b15zdnd00an1n02x5 FILLER_29_1492 ();
 b15zdnd11an1n04x5 FILLER_29_1497 ();
 b15zdnd11an1n08x5 FILLER_29_1504 ();
 b15zdnd11an1n04x5 FILLER_29_1512 ();
 b15zdnd00an1n02x5 FILLER_29_1516 ();
 b15zdnd00an1n01x5 FILLER_29_1518 ();
 b15zdnd11an1n64x5 FILLER_29_1522 ();
 b15zdnd11an1n64x5 FILLER_29_1586 ();
 b15zdnd11an1n64x5 FILLER_29_1650 ();
 b15zdnd11an1n64x5 FILLER_29_1714 ();
 b15zdnd11an1n64x5 FILLER_29_1778 ();
 b15zdnd11an1n64x5 FILLER_29_1842 ();
 b15zdnd11an1n64x5 FILLER_29_1906 ();
 b15zdnd11an1n64x5 FILLER_29_1970 ();
 b15zdnd11an1n64x5 FILLER_29_2034 ();
 b15zdnd11an1n64x5 FILLER_29_2098 ();
 b15zdnd11an1n64x5 FILLER_29_2162 ();
 b15zdnd11an1n32x5 FILLER_29_2226 ();
 b15zdnd11an1n16x5 FILLER_29_2258 ();
 b15zdnd11an1n08x5 FILLER_29_2274 ();
 b15zdnd00an1n02x5 FILLER_29_2282 ();
 b15zdnd11an1n64x5 FILLER_30_8 ();
 b15zdnd11an1n64x5 FILLER_30_72 ();
 b15zdnd11an1n64x5 FILLER_30_136 ();
 b15zdnd11an1n64x5 FILLER_30_200 ();
 b15zdnd11an1n64x5 FILLER_30_264 ();
 b15zdnd11an1n64x5 FILLER_30_328 ();
 b15zdnd11an1n64x5 FILLER_30_392 ();
 b15zdnd11an1n64x5 FILLER_30_456 ();
 b15zdnd11an1n64x5 FILLER_30_520 ();
 b15zdnd11an1n64x5 FILLER_30_584 ();
 b15zdnd11an1n64x5 FILLER_30_648 ();
 b15zdnd11an1n04x5 FILLER_30_712 ();
 b15zdnd00an1n02x5 FILLER_30_716 ();
 b15zdnd11an1n64x5 FILLER_30_726 ();
 b15zdnd11an1n64x5 FILLER_30_790 ();
 b15zdnd11an1n64x5 FILLER_30_854 ();
 b15zdnd11an1n64x5 FILLER_30_918 ();
 b15zdnd11an1n64x5 FILLER_30_982 ();
 b15zdnd11an1n64x5 FILLER_30_1046 ();
 b15zdnd11an1n64x5 FILLER_30_1110 ();
 b15zdnd11an1n64x5 FILLER_30_1174 ();
 b15zdnd11an1n64x5 FILLER_30_1238 ();
 b15zdnd11an1n04x5 FILLER_30_1302 ();
 b15zdnd00an1n02x5 FILLER_30_1306 ();
 b15zdnd00an1n01x5 FILLER_30_1308 ();
 b15zdnd11an1n04x5 FILLER_30_1361 ();
 b15zdnd00an1n01x5 FILLER_30_1365 ();
 b15zdnd11an1n32x5 FILLER_30_1418 ();
 b15zdnd11an1n16x5 FILLER_30_1450 ();
 b15zdnd00an1n02x5 FILLER_30_1466 ();
 b15zdnd00an1n01x5 FILLER_30_1468 ();
 b15zdnd11an1n64x5 FILLER_30_1521 ();
 b15zdnd11an1n64x5 FILLER_30_1585 ();
 b15zdnd11an1n64x5 FILLER_30_1649 ();
 b15zdnd11an1n64x5 FILLER_30_1713 ();
 b15zdnd11an1n64x5 FILLER_30_1777 ();
 b15zdnd11an1n64x5 FILLER_30_1841 ();
 b15zdnd11an1n64x5 FILLER_30_1905 ();
 b15zdnd11an1n64x5 FILLER_30_1969 ();
 b15zdnd11an1n64x5 FILLER_30_2033 ();
 b15zdnd11an1n32x5 FILLER_30_2097 ();
 b15zdnd11an1n16x5 FILLER_30_2129 ();
 b15zdnd11an1n08x5 FILLER_30_2145 ();
 b15zdnd00an1n01x5 FILLER_30_2153 ();
 b15zdnd11an1n64x5 FILLER_30_2162 ();
 b15zdnd11an1n32x5 FILLER_30_2226 ();
 b15zdnd11an1n16x5 FILLER_30_2258 ();
 b15zdnd00an1n02x5 FILLER_30_2274 ();
 b15zdnd11an1n64x5 FILLER_31_0 ();
 b15zdnd11an1n64x5 FILLER_31_64 ();
 b15zdnd11an1n64x5 FILLER_31_128 ();
 b15zdnd11an1n64x5 FILLER_31_192 ();
 b15zdnd11an1n64x5 FILLER_31_256 ();
 b15zdnd11an1n64x5 FILLER_31_320 ();
 b15zdnd11an1n64x5 FILLER_31_384 ();
 b15zdnd11an1n64x5 FILLER_31_448 ();
 b15zdnd11an1n64x5 FILLER_31_512 ();
 b15zdnd11an1n64x5 FILLER_31_576 ();
 b15zdnd11an1n64x5 FILLER_31_640 ();
 b15zdnd11an1n64x5 FILLER_31_704 ();
 b15zdnd11an1n64x5 FILLER_31_768 ();
 b15zdnd11an1n64x5 FILLER_31_832 ();
 b15zdnd11an1n64x5 FILLER_31_896 ();
 b15zdnd11an1n64x5 FILLER_31_960 ();
 b15zdnd11an1n16x5 FILLER_31_1024 ();
 b15zdnd00an1n01x5 FILLER_31_1040 ();
 b15zdnd11an1n64x5 FILLER_31_1045 ();
 b15zdnd11an1n64x5 FILLER_31_1109 ();
 b15zdnd11an1n64x5 FILLER_31_1173 ();
 b15zdnd11an1n64x5 FILLER_31_1237 ();
 b15zdnd11an1n64x5 FILLER_31_1301 ();
 b15zdnd11an1n16x5 FILLER_31_1365 ();
 b15zdnd11an1n04x5 FILLER_31_1381 ();
 b15zdnd11an1n04x5 FILLER_31_1388 ();
 b15zdnd11an1n64x5 FILLER_31_1395 ();
 b15zdnd11an1n32x5 FILLER_31_1459 ();
 b15zdnd00an1n02x5 FILLER_31_1491 ();
 b15zdnd00an1n01x5 FILLER_31_1493 ();
 b15zdnd11an1n64x5 FILLER_31_1497 ();
 b15zdnd11an1n64x5 FILLER_31_1561 ();
 b15zdnd11an1n64x5 FILLER_31_1625 ();
 b15zdnd11an1n64x5 FILLER_31_1689 ();
 b15zdnd11an1n64x5 FILLER_31_1753 ();
 b15zdnd11an1n64x5 FILLER_31_1817 ();
 b15zdnd11an1n64x5 FILLER_31_1881 ();
 b15zdnd11an1n64x5 FILLER_31_1945 ();
 b15zdnd11an1n64x5 FILLER_31_2009 ();
 b15zdnd11an1n64x5 FILLER_31_2073 ();
 b15zdnd11an1n64x5 FILLER_31_2137 ();
 b15zdnd11an1n64x5 FILLER_31_2201 ();
 b15zdnd11an1n16x5 FILLER_31_2265 ();
 b15zdnd00an1n02x5 FILLER_31_2281 ();
 b15zdnd00an1n01x5 FILLER_31_2283 ();
 b15zdnd11an1n64x5 FILLER_32_8 ();
 b15zdnd11an1n64x5 FILLER_32_72 ();
 b15zdnd11an1n64x5 FILLER_32_136 ();
 b15zdnd11an1n64x5 FILLER_32_200 ();
 b15zdnd11an1n64x5 FILLER_32_264 ();
 b15zdnd11an1n64x5 FILLER_32_328 ();
 b15zdnd11an1n64x5 FILLER_32_392 ();
 b15zdnd11an1n64x5 FILLER_32_456 ();
 b15zdnd11an1n64x5 FILLER_32_520 ();
 b15zdnd11an1n64x5 FILLER_32_584 ();
 b15zdnd11an1n64x5 FILLER_32_648 ();
 b15zdnd11an1n04x5 FILLER_32_712 ();
 b15zdnd00an1n02x5 FILLER_32_716 ();
 b15zdnd11an1n64x5 FILLER_32_726 ();
 b15zdnd11an1n64x5 FILLER_32_790 ();
 b15zdnd11an1n64x5 FILLER_32_854 ();
 b15zdnd11an1n64x5 FILLER_32_918 ();
 b15zdnd11an1n64x5 FILLER_32_982 ();
 b15zdnd11an1n64x5 FILLER_32_1046 ();
 b15zdnd11an1n64x5 FILLER_32_1110 ();
 b15zdnd11an1n64x5 FILLER_32_1174 ();
 b15zdnd11an1n64x5 FILLER_32_1238 ();
 b15zdnd11an1n64x5 FILLER_32_1302 ();
 b15zdnd11an1n08x5 FILLER_32_1366 ();
 b15zdnd11an1n04x5 FILLER_32_1374 ();
 b15zdnd11an1n04x5 FILLER_32_1388 ();
 b15zdnd11an1n64x5 FILLER_32_1395 ();
 b15zdnd11an1n64x5 FILLER_32_1459 ();
 b15zdnd11an1n64x5 FILLER_32_1523 ();
 b15zdnd11an1n32x5 FILLER_32_1587 ();
 b15zdnd11an1n16x5 FILLER_32_1619 ();
 b15zdnd11an1n04x5 FILLER_32_1638 ();
 b15zdnd11an1n64x5 FILLER_32_1645 ();
 b15zdnd11an1n64x5 FILLER_32_1709 ();
 b15zdnd11an1n64x5 FILLER_32_1773 ();
 b15zdnd11an1n64x5 FILLER_32_1837 ();
 b15zdnd11an1n64x5 FILLER_32_1901 ();
 b15zdnd11an1n64x5 FILLER_32_1965 ();
 b15zdnd11an1n64x5 FILLER_32_2029 ();
 b15zdnd11an1n32x5 FILLER_32_2093 ();
 b15zdnd11an1n16x5 FILLER_32_2125 ();
 b15zdnd11an1n08x5 FILLER_32_2141 ();
 b15zdnd11an1n04x5 FILLER_32_2149 ();
 b15zdnd00an1n01x5 FILLER_32_2153 ();
 b15zdnd11an1n64x5 FILLER_32_2162 ();
 b15zdnd11an1n32x5 FILLER_32_2226 ();
 b15zdnd11an1n16x5 FILLER_32_2258 ();
 b15zdnd00an1n02x5 FILLER_32_2274 ();
 b15zdnd11an1n64x5 FILLER_33_0 ();
 b15zdnd11an1n64x5 FILLER_33_64 ();
 b15zdnd11an1n64x5 FILLER_33_128 ();
 b15zdnd11an1n64x5 FILLER_33_192 ();
 b15zdnd11an1n64x5 FILLER_33_256 ();
 b15zdnd11an1n64x5 FILLER_33_320 ();
 b15zdnd11an1n64x5 FILLER_33_384 ();
 b15zdnd11an1n64x5 FILLER_33_448 ();
 b15zdnd11an1n64x5 FILLER_33_512 ();
 b15zdnd11an1n64x5 FILLER_33_576 ();
 b15zdnd11an1n64x5 FILLER_33_640 ();
 b15zdnd11an1n64x5 FILLER_33_704 ();
 b15zdnd11an1n64x5 FILLER_33_768 ();
 b15zdnd11an1n64x5 FILLER_33_832 ();
 b15zdnd11an1n64x5 FILLER_33_896 ();
 b15zdnd11an1n64x5 FILLER_33_960 ();
 b15zdnd11an1n64x5 FILLER_33_1024 ();
 b15zdnd11an1n64x5 FILLER_33_1088 ();
 b15zdnd11an1n64x5 FILLER_33_1152 ();
 b15zdnd11an1n64x5 FILLER_33_1216 ();
 b15zdnd11an1n64x5 FILLER_33_1280 ();
 b15zdnd11an1n16x5 FILLER_33_1344 ();
 b15zdnd11an1n08x5 FILLER_33_1360 ();
 b15zdnd11an1n04x5 FILLER_33_1368 ();
 b15zdnd00an1n02x5 FILLER_33_1372 ();
 b15zdnd00an1n01x5 FILLER_33_1374 ();
 b15zdnd11an1n64x5 FILLER_33_1383 ();
 b15zdnd11an1n64x5 FILLER_33_1447 ();
 b15zdnd11an1n64x5 FILLER_33_1511 ();
 b15zdnd11an1n32x5 FILLER_33_1575 ();
 b15zdnd11an1n08x5 FILLER_33_1607 ();
 b15zdnd11an1n04x5 FILLER_33_1667 ();
 b15zdnd11an1n04x5 FILLER_33_1674 ();
 b15zdnd00an1n01x5 FILLER_33_1678 ();
 b15zdnd11an1n04x5 FILLER_33_1682 ();
 b15zdnd00an1n01x5 FILLER_33_1686 ();
 b15zdnd11an1n64x5 FILLER_33_1714 ();
 b15zdnd11an1n64x5 FILLER_33_1778 ();
 b15zdnd11an1n64x5 FILLER_33_1842 ();
 b15zdnd11an1n64x5 FILLER_33_1906 ();
 b15zdnd11an1n64x5 FILLER_33_1970 ();
 b15zdnd11an1n64x5 FILLER_33_2034 ();
 b15zdnd11an1n64x5 FILLER_33_2098 ();
 b15zdnd11an1n64x5 FILLER_33_2162 ();
 b15zdnd11an1n16x5 FILLER_33_2226 ();
 b15zdnd11an1n08x5 FILLER_33_2242 ();
 b15zdnd11an1n04x5 FILLER_33_2250 ();
 b15zdnd00an1n01x5 FILLER_33_2254 ();
 b15zdnd11an1n16x5 FILLER_33_2258 ();
 b15zdnd11an1n08x5 FILLER_33_2274 ();
 b15zdnd00an1n02x5 FILLER_33_2282 ();
 b15zdnd11an1n64x5 FILLER_34_8 ();
 b15zdnd11an1n64x5 FILLER_34_72 ();
 b15zdnd11an1n64x5 FILLER_34_136 ();
 b15zdnd11an1n64x5 FILLER_34_200 ();
 b15zdnd11an1n64x5 FILLER_34_264 ();
 b15zdnd11an1n64x5 FILLER_34_328 ();
 b15zdnd11an1n64x5 FILLER_34_392 ();
 b15zdnd11an1n64x5 FILLER_34_456 ();
 b15zdnd11an1n64x5 FILLER_34_520 ();
 b15zdnd11an1n64x5 FILLER_34_584 ();
 b15zdnd11an1n64x5 FILLER_34_648 ();
 b15zdnd11an1n04x5 FILLER_34_712 ();
 b15zdnd00an1n02x5 FILLER_34_716 ();
 b15zdnd11an1n64x5 FILLER_34_726 ();
 b15zdnd11an1n64x5 FILLER_34_790 ();
 b15zdnd11an1n64x5 FILLER_34_854 ();
 b15zdnd11an1n64x5 FILLER_34_918 ();
 b15zdnd11an1n64x5 FILLER_34_982 ();
 b15zdnd11an1n64x5 FILLER_34_1046 ();
 b15zdnd11an1n16x5 FILLER_34_1110 ();
 b15zdnd11an1n04x5 FILLER_34_1126 ();
 b15zdnd00an1n01x5 FILLER_34_1130 ();
 b15zdnd11an1n64x5 FILLER_34_1183 ();
 b15zdnd11an1n64x5 FILLER_34_1247 ();
 b15zdnd11an1n64x5 FILLER_34_1311 ();
 b15zdnd11an1n64x5 FILLER_34_1375 ();
 b15zdnd11an1n64x5 FILLER_34_1439 ();
 b15zdnd11an1n64x5 FILLER_34_1503 ();
 b15zdnd11an1n32x5 FILLER_34_1567 ();
 b15zdnd11an1n16x5 FILLER_34_1599 ();
 b15zdnd11an1n08x5 FILLER_34_1615 ();
 b15zdnd11an1n04x5 FILLER_34_1675 ();
 b15zdnd00an1n02x5 FILLER_34_1679 ();
 b15zdnd00an1n01x5 FILLER_34_1681 ();
 b15zdnd11an1n04x5 FILLER_34_1685 ();
 b15zdnd00an1n02x5 FILLER_34_1689 ();
 b15zdnd11an1n64x5 FILLER_34_1694 ();
 b15zdnd11an1n08x5 FILLER_34_1758 ();
 b15zdnd11an1n04x5 FILLER_34_1766 ();
 b15zdnd00an1n02x5 FILLER_34_1770 ();
 b15zdnd11an1n64x5 FILLER_34_1824 ();
 b15zdnd11an1n64x5 FILLER_34_1888 ();
 b15zdnd11an1n64x5 FILLER_34_1952 ();
 b15zdnd11an1n64x5 FILLER_34_2016 ();
 b15zdnd11an1n64x5 FILLER_34_2080 ();
 b15zdnd11an1n08x5 FILLER_34_2144 ();
 b15zdnd00an1n02x5 FILLER_34_2152 ();
 b15zdnd11an1n64x5 FILLER_34_2162 ();
 b15zdnd11an1n16x5 FILLER_34_2226 ();
 b15zdnd11an1n08x5 FILLER_34_2242 ();
 b15zdnd11an1n04x5 FILLER_34_2250 ();
 b15zdnd00an1n01x5 FILLER_34_2254 ();
 b15zdnd11an1n16x5 FILLER_34_2258 ();
 b15zdnd00an1n02x5 FILLER_34_2274 ();
 b15zdnd11an1n64x5 FILLER_35_0 ();
 b15zdnd11an1n64x5 FILLER_35_64 ();
 b15zdnd11an1n64x5 FILLER_35_128 ();
 b15zdnd11an1n64x5 FILLER_35_192 ();
 b15zdnd11an1n64x5 FILLER_35_256 ();
 b15zdnd11an1n64x5 FILLER_35_320 ();
 b15zdnd11an1n64x5 FILLER_35_384 ();
 b15zdnd11an1n64x5 FILLER_35_448 ();
 b15zdnd11an1n32x5 FILLER_35_512 ();
 b15zdnd11an1n16x5 FILLER_35_544 ();
 b15zdnd11an1n08x5 FILLER_35_560 ();
 b15zdnd00an1n02x5 FILLER_35_568 ();
 b15zdnd00an1n01x5 FILLER_35_570 ();
 b15zdnd11an1n32x5 FILLER_35_580 ();
 b15zdnd11an1n08x5 FILLER_35_612 ();
 b15zdnd11an1n04x5 FILLER_35_620 ();
 b15zdnd00an1n02x5 FILLER_35_624 ();
 b15zdnd00an1n01x5 FILLER_35_626 ();
 b15zdnd11an1n64x5 FILLER_35_636 ();
 b15zdnd11an1n64x5 FILLER_35_700 ();
 b15zdnd11an1n64x5 FILLER_35_764 ();
 b15zdnd11an1n64x5 FILLER_35_828 ();
 b15zdnd11an1n64x5 FILLER_35_892 ();
 b15zdnd11an1n64x5 FILLER_35_956 ();
 b15zdnd11an1n64x5 FILLER_35_1020 ();
 b15zdnd11an1n64x5 FILLER_35_1084 ();
 b15zdnd00an1n01x5 FILLER_35_1148 ();
 b15zdnd11an1n04x5 FILLER_35_1152 ();
 b15zdnd11an1n04x5 FILLER_35_1159 ();
 b15zdnd11an1n64x5 FILLER_35_1166 ();
 b15zdnd11an1n64x5 FILLER_35_1230 ();
 b15zdnd11an1n32x5 FILLER_35_1294 ();
 b15zdnd11an1n16x5 FILLER_35_1326 ();
 b15zdnd11an1n08x5 FILLER_35_1342 ();
 b15zdnd11an1n04x5 FILLER_35_1350 ();
 b15zdnd00an1n02x5 FILLER_35_1354 ();
 b15zdnd11an1n64x5 FILLER_35_1361 ();
 b15zdnd11an1n64x5 FILLER_35_1425 ();
 b15zdnd11an1n64x5 FILLER_35_1489 ();
 b15zdnd11an1n64x5 FILLER_35_1553 ();
 b15zdnd11an1n08x5 FILLER_35_1617 ();
 b15zdnd11an1n04x5 FILLER_35_1677 ();
 b15zdnd00an1n01x5 FILLER_35_1681 ();
 b15zdnd11an1n32x5 FILLER_35_1691 ();
 b15zdnd11an1n08x5 FILLER_35_1723 ();
 b15zdnd11an1n04x5 FILLER_35_1731 ();
 b15zdnd00an1n02x5 FILLER_35_1735 ();
 b15zdnd00an1n01x5 FILLER_35_1737 ();
 b15zdnd11an1n16x5 FILLER_35_1747 ();
 b15zdnd11an1n08x5 FILLER_35_1763 ();
 b15zdnd11an1n04x5 FILLER_35_1771 ();
 b15zdnd11an1n64x5 FILLER_35_1827 ();
 b15zdnd11an1n64x5 FILLER_35_1891 ();
 b15zdnd11an1n64x5 FILLER_35_1955 ();
 b15zdnd11an1n64x5 FILLER_35_2019 ();
 b15zdnd11an1n64x5 FILLER_35_2083 ();
 b15zdnd11an1n64x5 FILLER_35_2147 ();
 b15zdnd11an1n64x5 FILLER_35_2211 ();
 b15zdnd11an1n08x5 FILLER_35_2275 ();
 b15zdnd00an1n01x5 FILLER_35_2283 ();
 b15zdnd11an1n64x5 FILLER_36_8 ();
 b15zdnd11an1n64x5 FILLER_36_72 ();
 b15zdnd11an1n64x5 FILLER_36_136 ();
 b15zdnd11an1n64x5 FILLER_36_200 ();
 b15zdnd11an1n64x5 FILLER_36_264 ();
 b15zdnd11an1n64x5 FILLER_36_328 ();
 b15zdnd11an1n64x5 FILLER_36_392 ();
 b15zdnd11an1n64x5 FILLER_36_456 ();
 b15zdnd11an1n64x5 FILLER_36_520 ();
 b15zdnd11an1n64x5 FILLER_36_584 ();
 b15zdnd11an1n64x5 FILLER_36_648 ();
 b15zdnd11an1n04x5 FILLER_36_712 ();
 b15zdnd00an1n02x5 FILLER_36_716 ();
 b15zdnd11an1n64x5 FILLER_36_726 ();
 b15zdnd11an1n64x5 FILLER_36_790 ();
 b15zdnd11an1n64x5 FILLER_36_854 ();
 b15zdnd11an1n64x5 FILLER_36_918 ();
 b15zdnd11an1n64x5 FILLER_36_982 ();
 b15zdnd11an1n64x5 FILLER_36_1046 ();
 b15zdnd11an1n64x5 FILLER_36_1110 ();
 b15zdnd11an1n64x5 FILLER_36_1174 ();
 b15zdnd11an1n64x5 FILLER_36_1238 ();
 b15zdnd11an1n32x5 FILLER_36_1302 ();
 b15zdnd11an1n08x5 FILLER_36_1334 ();
 b15zdnd11an1n04x5 FILLER_36_1342 ();
 b15zdnd00an1n01x5 FILLER_36_1346 ();
 b15zdnd11an1n64x5 FILLER_36_1361 ();
 b15zdnd11an1n64x5 FILLER_36_1425 ();
 b15zdnd11an1n64x5 FILLER_36_1489 ();
 b15zdnd11an1n64x5 FILLER_36_1553 ();
 b15zdnd11an1n08x5 FILLER_36_1617 ();
 b15zdnd11an1n32x5 FILLER_36_1677 ();
 b15zdnd11an1n16x5 FILLER_36_1709 ();
 b15zdnd00an1n02x5 FILLER_36_1725 ();
 b15zdnd11an1n32x5 FILLER_36_1736 ();
 b15zdnd00an1n02x5 FILLER_36_1768 ();
 b15zdnd11an1n04x5 FILLER_36_1822 ();
 b15zdnd11an1n64x5 FILLER_36_1829 ();
 b15zdnd11an1n64x5 FILLER_36_1893 ();
 b15zdnd11an1n64x5 FILLER_36_1957 ();
 b15zdnd11an1n64x5 FILLER_36_2021 ();
 b15zdnd11an1n64x5 FILLER_36_2085 ();
 b15zdnd11an1n04x5 FILLER_36_2149 ();
 b15zdnd00an1n01x5 FILLER_36_2153 ();
 b15zdnd11an1n64x5 FILLER_36_2162 ();
 b15zdnd11an1n32x5 FILLER_36_2226 ();
 b15zdnd11an1n16x5 FILLER_36_2258 ();
 b15zdnd00an1n02x5 FILLER_36_2274 ();
 b15zdnd11an1n64x5 FILLER_37_0 ();
 b15zdnd11an1n64x5 FILLER_37_64 ();
 b15zdnd11an1n64x5 FILLER_37_128 ();
 b15zdnd11an1n64x5 FILLER_37_192 ();
 b15zdnd11an1n64x5 FILLER_37_256 ();
 b15zdnd11an1n64x5 FILLER_37_320 ();
 b15zdnd11an1n64x5 FILLER_37_384 ();
 b15zdnd11an1n64x5 FILLER_37_448 ();
 b15zdnd11an1n64x5 FILLER_37_512 ();
 b15zdnd11an1n32x5 FILLER_37_576 ();
 b15zdnd00an1n02x5 FILLER_37_608 ();
 b15zdnd11an1n64x5 FILLER_37_619 ();
 b15zdnd11an1n64x5 FILLER_37_683 ();
 b15zdnd11an1n64x5 FILLER_37_747 ();
 b15zdnd11an1n16x5 FILLER_37_811 ();
 b15zdnd00an1n01x5 FILLER_37_827 ();
 b15zdnd11an1n64x5 FILLER_37_831 ();
 b15zdnd11an1n64x5 FILLER_37_895 ();
 b15zdnd11an1n64x5 FILLER_37_959 ();
 b15zdnd11an1n64x5 FILLER_37_1023 ();
 b15zdnd11an1n32x5 FILLER_37_1087 ();
 b15zdnd11an1n16x5 FILLER_37_1119 ();
 b15zdnd00an1n02x5 FILLER_37_1135 ();
 b15zdnd11an1n64x5 FILLER_37_1151 ();
 b15zdnd11an1n64x5 FILLER_37_1215 ();
 b15zdnd11an1n64x5 FILLER_37_1279 ();
 b15zdnd11an1n64x5 FILLER_37_1343 ();
 b15zdnd11an1n64x5 FILLER_37_1407 ();
 b15zdnd11an1n64x5 FILLER_37_1471 ();
 b15zdnd11an1n64x5 FILLER_37_1535 ();
 b15zdnd11an1n32x5 FILLER_37_1599 ();
 b15zdnd11an1n08x5 FILLER_37_1631 ();
 b15zdnd11an1n04x5 FILLER_37_1639 ();
 b15zdnd11an1n04x5 FILLER_37_1646 ();
 b15zdnd11an1n04x5 FILLER_37_1653 ();
 b15zdnd11an1n04x5 FILLER_37_1660 ();
 b15zdnd11an1n64x5 FILLER_37_1667 ();
 b15zdnd11an1n32x5 FILLER_37_1731 ();
 b15zdnd11an1n08x5 FILLER_37_1763 ();
 b15zdnd11an1n64x5 FILLER_37_1823 ();
 b15zdnd11an1n64x5 FILLER_37_1887 ();
 b15zdnd11an1n64x5 FILLER_37_1951 ();
 b15zdnd11an1n64x5 FILLER_37_2015 ();
 b15zdnd11an1n64x5 FILLER_37_2079 ();
 b15zdnd11an1n64x5 FILLER_37_2143 ();
 b15zdnd11an1n64x5 FILLER_37_2207 ();
 b15zdnd11an1n08x5 FILLER_37_2271 ();
 b15zdnd11an1n04x5 FILLER_37_2279 ();
 b15zdnd00an1n01x5 FILLER_37_2283 ();
 b15zdnd11an1n64x5 FILLER_38_8 ();
 b15zdnd11an1n64x5 FILLER_38_72 ();
 b15zdnd11an1n64x5 FILLER_38_136 ();
 b15zdnd11an1n64x5 FILLER_38_200 ();
 b15zdnd11an1n64x5 FILLER_38_264 ();
 b15zdnd11an1n64x5 FILLER_38_328 ();
 b15zdnd11an1n64x5 FILLER_38_392 ();
 b15zdnd11an1n64x5 FILLER_38_456 ();
 b15zdnd11an1n64x5 FILLER_38_520 ();
 b15zdnd11an1n64x5 FILLER_38_584 ();
 b15zdnd11an1n08x5 FILLER_38_648 ();
 b15zdnd11an1n04x5 FILLER_38_656 ();
 b15zdnd00an1n02x5 FILLER_38_660 ();
 b15zdnd00an1n01x5 FILLER_38_662 ();
 b15zdnd11an1n32x5 FILLER_38_666 ();
 b15zdnd11an1n16x5 FILLER_38_698 ();
 b15zdnd11an1n04x5 FILLER_38_714 ();
 b15zdnd11an1n64x5 FILLER_38_726 ();
 b15zdnd11an1n08x5 FILLER_38_790 ();
 b15zdnd00an1n02x5 FILLER_38_798 ();
 b15zdnd00an1n01x5 FILLER_38_800 ();
 b15zdnd11an1n64x5 FILLER_38_853 ();
 b15zdnd11an1n64x5 FILLER_38_917 ();
 b15zdnd11an1n08x5 FILLER_38_981 ();
 b15zdnd11an1n04x5 FILLER_38_989 ();
 b15zdnd00an1n01x5 FILLER_38_993 ();
 b15zdnd11an1n04x5 FILLER_38_997 ();
 b15zdnd11an1n64x5 FILLER_38_1004 ();
 b15zdnd11an1n64x5 FILLER_38_1068 ();
 b15zdnd11an1n64x5 FILLER_38_1132 ();
 b15zdnd11an1n64x5 FILLER_38_1196 ();
 b15zdnd11an1n64x5 FILLER_38_1260 ();
 b15zdnd11an1n64x5 FILLER_38_1324 ();
 b15zdnd11an1n64x5 FILLER_38_1388 ();
 b15zdnd11an1n64x5 FILLER_38_1452 ();
 b15zdnd11an1n64x5 FILLER_38_1516 ();
 b15zdnd11an1n32x5 FILLER_38_1580 ();
 b15zdnd11an1n16x5 FILLER_38_1612 ();
 b15zdnd11an1n08x5 FILLER_38_1628 ();
 b15zdnd11an1n04x5 FILLER_38_1636 ();
 b15zdnd00an1n02x5 FILLER_38_1640 ();
 b15zdnd00an1n01x5 FILLER_38_1642 ();
 b15zdnd11an1n04x5 FILLER_38_1646 ();
 b15zdnd11an1n64x5 FILLER_38_1653 ();
 b15zdnd11an1n64x5 FILLER_38_1717 ();
 b15zdnd11an1n04x5 FILLER_38_1784 ();
 b15zdnd11an1n04x5 FILLER_38_1791 ();
 b15zdnd11an1n04x5 FILLER_38_1798 ();
 b15zdnd11an1n04x5 FILLER_38_1805 ();
 b15zdnd11an1n04x5 FILLER_38_1812 ();
 b15zdnd11an1n64x5 FILLER_38_1819 ();
 b15zdnd11an1n64x5 FILLER_38_1883 ();
 b15zdnd11an1n64x5 FILLER_38_1947 ();
 b15zdnd11an1n64x5 FILLER_38_2011 ();
 b15zdnd11an1n64x5 FILLER_38_2075 ();
 b15zdnd11an1n08x5 FILLER_38_2139 ();
 b15zdnd11an1n04x5 FILLER_38_2147 ();
 b15zdnd00an1n02x5 FILLER_38_2151 ();
 b15zdnd00an1n01x5 FILLER_38_2153 ();
 b15zdnd11an1n64x5 FILLER_38_2162 ();
 b15zdnd11an1n32x5 FILLER_38_2226 ();
 b15zdnd11an1n16x5 FILLER_38_2258 ();
 b15zdnd00an1n02x5 FILLER_38_2274 ();
 b15zdnd11an1n64x5 FILLER_39_0 ();
 b15zdnd11an1n64x5 FILLER_39_64 ();
 b15zdnd11an1n64x5 FILLER_39_128 ();
 b15zdnd11an1n64x5 FILLER_39_192 ();
 b15zdnd11an1n64x5 FILLER_39_256 ();
 b15zdnd11an1n64x5 FILLER_39_320 ();
 b15zdnd11an1n64x5 FILLER_39_384 ();
 b15zdnd11an1n64x5 FILLER_39_448 ();
 b15zdnd11an1n64x5 FILLER_39_512 ();
 b15zdnd11an1n64x5 FILLER_39_576 ();
 b15zdnd11an1n16x5 FILLER_39_640 ();
 b15zdnd11an1n04x5 FILLER_39_656 ();
 b15zdnd00an1n02x5 FILLER_39_660 ();
 b15zdnd11an1n04x5 FILLER_39_665 ();
 b15zdnd11an1n64x5 FILLER_39_672 ();
 b15zdnd11an1n64x5 FILLER_39_736 ();
 b15zdnd11an1n16x5 FILLER_39_800 ();
 b15zdnd00an1n02x5 FILLER_39_816 ();
 b15zdnd00an1n01x5 FILLER_39_818 ();
 b15zdnd11an1n04x5 FILLER_39_822 ();
 b15zdnd11an1n64x5 FILLER_39_829 ();
 b15zdnd11an1n64x5 FILLER_39_893 ();
 b15zdnd11an1n16x5 FILLER_39_957 ();
 b15zdnd11an1n08x5 FILLER_39_973 ();
 b15zdnd11an1n04x5 FILLER_39_981 ();
 b15zdnd00an1n02x5 FILLER_39_985 ();
 b15zdnd00an1n01x5 FILLER_39_987 ();
 b15zdnd11an1n64x5 FILLER_39_1040 ();
 b15zdnd11an1n64x5 FILLER_39_1104 ();
 b15zdnd00an1n02x5 FILLER_39_1168 ();
 b15zdnd00an1n01x5 FILLER_39_1170 ();
 b15zdnd11an1n32x5 FILLER_39_1176 ();
 b15zdnd11an1n16x5 FILLER_39_1208 ();
 b15zdnd11an1n64x5 FILLER_39_1230 ();
 b15zdnd11an1n64x5 FILLER_39_1294 ();
 b15zdnd11an1n64x5 FILLER_39_1358 ();
 b15zdnd11an1n64x5 FILLER_39_1422 ();
 b15zdnd11an1n64x5 FILLER_39_1486 ();
 b15zdnd11an1n64x5 FILLER_39_1550 ();
 b15zdnd11an1n32x5 FILLER_39_1614 ();
 b15zdnd00an1n02x5 FILLER_39_1646 ();
 b15zdnd11an1n64x5 FILLER_39_1651 ();
 b15zdnd11an1n64x5 FILLER_39_1715 ();
 b15zdnd11an1n08x5 FILLER_39_1779 ();
 b15zdnd00an1n02x5 FILLER_39_1787 ();
 b15zdnd11an1n04x5 FILLER_39_1792 ();
 b15zdnd11an1n04x5 FILLER_39_1799 ();
 b15zdnd11an1n64x5 FILLER_39_1806 ();
 b15zdnd11an1n64x5 FILLER_39_1870 ();
 b15zdnd11an1n64x5 FILLER_39_1934 ();
 b15zdnd11an1n64x5 FILLER_39_1998 ();
 b15zdnd11an1n64x5 FILLER_39_2062 ();
 b15zdnd11an1n64x5 FILLER_39_2126 ();
 b15zdnd11an1n64x5 FILLER_39_2190 ();
 b15zdnd11an1n16x5 FILLER_39_2254 ();
 b15zdnd11an1n08x5 FILLER_39_2270 ();
 b15zdnd11an1n04x5 FILLER_39_2278 ();
 b15zdnd00an1n02x5 FILLER_39_2282 ();
 b15zdnd11an1n64x5 FILLER_40_8 ();
 b15zdnd11an1n64x5 FILLER_40_72 ();
 b15zdnd11an1n64x5 FILLER_40_136 ();
 b15zdnd11an1n64x5 FILLER_40_200 ();
 b15zdnd11an1n64x5 FILLER_40_264 ();
 b15zdnd11an1n64x5 FILLER_40_328 ();
 b15zdnd11an1n64x5 FILLER_40_392 ();
 b15zdnd11an1n64x5 FILLER_40_456 ();
 b15zdnd11an1n16x5 FILLER_40_520 ();
 b15zdnd11an1n64x5 FILLER_40_539 ();
 b15zdnd11an1n32x5 FILLER_40_603 ();
 b15zdnd11an1n04x5 FILLER_40_635 ();
 b15zdnd00an1n02x5 FILLER_40_639 ();
 b15zdnd00an1n01x5 FILLER_40_641 ();
 b15zdnd11an1n16x5 FILLER_40_694 ();
 b15zdnd11an1n08x5 FILLER_40_710 ();
 b15zdnd11an1n64x5 FILLER_40_726 ();
 b15zdnd11an1n64x5 FILLER_40_790 ();
 b15zdnd11an1n16x5 FILLER_40_854 ();
 b15zdnd11an1n04x5 FILLER_40_870 ();
 b15zdnd00an1n02x5 FILLER_40_874 ();
 b15zdnd00an1n01x5 FILLER_40_876 ();
 b15zdnd11an1n32x5 FILLER_40_886 ();
 b15zdnd11an1n08x5 FILLER_40_918 ();
 b15zdnd11an1n04x5 FILLER_40_926 ();
 b15zdnd00an1n02x5 FILLER_40_930 ();
 b15zdnd11an1n32x5 FILLER_40_941 ();
 b15zdnd11an1n16x5 FILLER_40_973 ();
 b15zdnd11an1n08x5 FILLER_40_989 ();
 b15zdnd00an1n01x5 FILLER_40_997 ();
 b15zdnd11an1n64x5 FILLER_40_1001 ();
 b15zdnd11an1n64x5 FILLER_40_1065 ();
 b15zdnd11an1n64x5 FILLER_40_1129 ();
 b15zdnd11an1n64x5 FILLER_40_1193 ();
 b15zdnd11an1n64x5 FILLER_40_1257 ();
 b15zdnd11an1n64x5 FILLER_40_1321 ();
 b15zdnd11an1n64x5 FILLER_40_1385 ();
 b15zdnd11an1n32x5 FILLER_40_1449 ();
 b15zdnd11an1n16x5 FILLER_40_1481 ();
 b15zdnd00an1n01x5 FILLER_40_1497 ();
 b15zdnd11an1n64x5 FILLER_40_1540 ();
 b15zdnd11an1n64x5 FILLER_40_1604 ();
 b15zdnd11an1n64x5 FILLER_40_1668 ();
 b15zdnd11an1n64x5 FILLER_40_1732 ();
 b15zdnd00an1n01x5 FILLER_40_1796 ();
 b15zdnd11an1n04x5 FILLER_40_1800 ();
 b15zdnd11an1n64x5 FILLER_40_1807 ();
 b15zdnd11an1n32x5 FILLER_40_1871 ();
 b15zdnd11an1n16x5 FILLER_40_1903 ();
 b15zdnd11an1n08x5 FILLER_40_1919 ();
 b15zdnd00an1n01x5 FILLER_40_1927 ();
 b15zdnd11an1n04x5 FILLER_40_1932 ();
 b15zdnd11an1n64x5 FILLER_40_1940 ();
 b15zdnd11an1n64x5 FILLER_40_2004 ();
 b15zdnd11an1n64x5 FILLER_40_2068 ();
 b15zdnd11an1n16x5 FILLER_40_2132 ();
 b15zdnd11an1n04x5 FILLER_40_2148 ();
 b15zdnd00an1n02x5 FILLER_40_2152 ();
 b15zdnd11an1n64x5 FILLER_40_2162 ();
 b15zdnd11an1n32x5 FILLER_40_2226 ();
 b15zdnd11an1n16x5 FILLER_40_2258 ();
 b15zdnd00an1n02x5 FILLER_40_2274 ();
 b15zdnd11an1n64x5 FILLER_41_0 ();
 b15zdnd11an1n64x5 FILLER_41_64 ();
 b15zdnd11an1n64x5 FILLER_41_128 ();
 b15zdnd11an1n64x5 FILLER_41_192 ();
 b15zdnd11an1n64x5 FILLER_41_256 ();
 b15zdnd11an1n64x5 FILLER_41_320 ();
 b15zdnd11an1n64x5 FILLER_41_384 ();
 b15zdnd11an1n64x5 FILLER_41_448 ();
 b15zdnd11an1n16x5 FILLER_41_512 ();
 b15zdnd00an1n02x5 FILLER_41_528 ();
 b15zdnd00an1n01x5 FILLER_41_530 ();
 b15zdnd11an1n04x5 FILLER_41_534 ();
 b15zdnd11an1n64x5 FILLER_41_541 ();
 b15zdnd11an1n32x5 FILLER_41_605 ();
 b15zdnd11an1n04x5 FILLER_41_637 ();
 b15zdnd00an1n02x5 FILLER_41_641 ();
 b15zdnd11an1n64x5 FILLER_41_695 ();
 b15zdnd11an1n64x5 FILLER_41_759 ();
 b15zdnd11an1n64x5 FILLER_41_823 ();
 b15zdnd11an1n16x5 FILLER_41_887 ();
 b15zdnd11an1n04x5 FILLER_41_903 ();
 b15zdnd00an1n02x5 FILLER_41_907 ();
 b15zdnd00an1n01x5 FILLER_41_909 ();
 b15zdnd11an1n04x5 FILLER_41_937 ();
 b15zdnd00an1n01x5 FILLER_41_941 ();
 b15zdnd11an1n64x5 FILLER_41_994 ();
 b15zdnd11an1n64x5 FILLER_41_1058 ();
 b15zdnd11an1n64x5 FILLER_41_1122 ();
 b15zdnd11an1n64x5 FILLER_41_1186 ();
 b15zdnd11an1n64x5 FILLER_41_1250 ();
 b15zdnd11an1n64x5 FILLER_41_1314 ();
 b15zdnd11an1n16x5 FILLER_41_1378 ();
 b15zdnd11an1n08x5 FILLER_41_1394 ();
 b15zdnd11an1n04x5 FILLER_41_1402 ();
 b15zdnd11an1n64x5 FILLER_41_1409 ();
 b15zdnd11an1n64x5 FILLER_41_1473 ();
 b15zdnd11an1n64x5 FILLER_41_1537 ();
 b15zdnd11an1n64x5 FILLER_41_1601 ();
 b15zdnd11an1n64x5 FILLER_41_1665 ();
 b15zdnd11an1n64x5 FILLER_41_1729 ();
 b15zdnd11an1n64x5 FILLER_41_1793 ();
 b15zdnd11an1n64x5 FILLER_41_1857 ();
 b15zdnd11an1n04x5 FILLER_41_1921 ();
 b15zdnd11an1n04x5 FILLER_41_1929 ();
 b15zdnd00an1n02x5 FILLER_41_1933 ();
 b15zdnd11an1n64x5 FILLER_41_1939 ();
 b15zdnd11an1n64x5 FILLER_41_2003 ();
 b15zdnd11an1n64x5 FILLER_41_2067 ();
 b15zdnd11an1n64x5 FILLER_41_2131 ();
 b15zdnd11an1n64x5 FILLER_41_2195 ();
 b15zdnd11an1n16x5 FILLER_41_2259 ();
 b15zdnd11an1n08x5 FILLER_41_2275 ();
 b15zdnd00an1n01x5 FILLER_41_2283 ();
 b15zdnd11an1n64x5 FILLER_42_8 ();
 b15zdnd11an1n64x5 FILLER_42_72 ();
 b15zdnd11an1n64x5 FILLER_42_136 ();
 b15zdnd11an1n64x5 FILLER_42_200 ();
 b15zdnd11an1n64x5 FILLER_42_264 ();
 b15zdnd11an1n64x5 FILLER_42_328 ();
 b15zdnd11an1n64x5 FILLER_42_392 ();
 b15zdnd11an1n32x5 FILLER_42_456 ();
 b15zdnd11an1n16x5 FILLER_42_488 ();
 b15zdnd11an1n04x5 FILLER_42_504 ();
 b15zdnd00an1n02x5 FILLER_42_508 ();
 b15zdnd00an1n01x5 FILLER_42_510 ();
 b15zdnd11an1n64x5 FILLER_42_563 ();
 b15zdnd11an1n16x5 FILLER_42_627 ();
 b15zdnd00an1n01x5 FILLER_42_643 ();
 b15zdnd11an1n16x5 FILLER_42_696 ();
 b15zdnd11an1n04x5 FILLER_42_712 ();
 b15zdnd00an1n02x5 FILLER_42_716 ();
 b15zdnd11an1n64x5 FILLER_42_726 ();
 b15zdnd11an1n16x5 FILLER_42_790 ();
 b15zdnd11an1n08x5 FILLER_42_806 ();
 b15zdnd11an1n04x5 FILLER_42_814 ();
 b15zdnd11an1n04x5 FILLER_42_821 ();
 b15zdnd11an1n04x5 FILLER_42_828 ();
 b15zdnd11an1n64x5 FILLER_42_835 ();
 b15zdnd11an1n08x5 FILLER_42_899 ();
 b15zdnd00an1n02x5 FILLER_42_907 ();
 b15zdnd00an1n01x5 FILLER_42_909 ();
 b15zdnd11an1n04x5 FILLER_42_913 ();
 b15zdnd00an1n02x5 FILLER_42_917 ();
 b15zdnd11an1n08x5 FILLER_42_928 ();
 b15zdnd11an1n04x5 FILLER_42_936 ();
 b15zdnd00an1n02x5 FILLER_42_940 ();
 b15zdnd00an1n01x5 FILLER_42_942 ();
 b15zdnd11an1n08x5 FILLER_42_951 ();
 b15zdnd00an1n02x5 FILLER_42_959 ();
 b15zdnd00an1n01x5 FILLER_42_961 ();
 b15zdnd11an1n04x5 FILLER_42_965 ();
 b15zdnd11an1n64x5 FILLER_42_972 ();
 b15zdnd11an1n64x5 FILLER_42_1036 ();
 b15zdnd11an1n64x5 FILLER_42_1100 ();
 b15zdnd11an1n64x5 FILLER_42_1164 ();
 b15zdnd11an1n64x5 FILLER_42_1228 ();
 b15zdnd00an1n02x5 FILLER_42_1292 ();
 b15zdnd11an1n64x5 FILLER_42_1312 ();
 b15zdnd11an1n16x5 FILLER_42_1376 ();
 b15zdnd11an1n08x5 FILLER_42_1392 ();
 b15zdnd11an1n04x5 FILLER_42_1400 ();
 b15zdnd00an1n01x5 FILLER_42_1404 ();
 b15zdnd11an1n64x5 FILLER_42_1408 ();
 b15zdnd11an1n16x5 FILLER_42_1472 ();
 b15zdnd11an1n08x5 FILLER_42_1488 ();
 b15zdnd00an1n01x5 FILLER_42_1496 ();
 b15zdnd11an1n64x5 FILLER_42_1500 ();
 b15zdnd11an1n64x5 FILLER_42_1564 ();
 b15zdnd11an1n64x5 FILLER_42_1628 ();
 b15zdnd11an1n64x5 FILLER_42_1692 ();
 b15zdnd11an1n64x5 FILLER_42_1756 ();
 b15zdnd11an1n64x5 FILLER_42_1820 ();
 b15zdnd11an1n16x5 FILLER_42_1884 ();
 b15zdnd11an1n08x5 FILLER_42_1900 ();
 b15zdnd00an1n02x5 FILLER_42_1908 ();
 b15zdnd11an1n64x5 FILLER_42_1918 ();
 b15zdnd11an1n64x5 FILLER_42_1982 ();
 b15zdnd11an1n64x5 FILLER_42_2046 ();
 b15zdnd11an1n32x5 FILLER_42_2110 ();
 b15zdnd11an1n08x5 FILLER_42_2142 ();
 b15zdnd11an1n04x5 FILLER_42_2150 ();
 b15zdnd11an1n64x5 FILLER_42_2162 ();
 b15zdnd11an1n32x5 FILLER_42_2226 ();
 b15zdnd11an1n16x5 FILLER_42_2258 ();
 b15zdnd00an1n02x5 FILLER_42_2274 ();
 b15zdnd11an1n64x5 FILLER_43_0 ();
 b15zdnd11an1n64x5 FILLER_43_64 ();
 b15zdnd11an1n64x5 FILLER_43_128 ();
 b15zdnd11an1n64x5 FILLER_43_192 ();
 b15zdnd11an1n64x5 FILLER_43_256 ();
 b15zdnd11an1n64x5 FILLER_43_320 ();
 b15zdnd11an1n64x5 FILLER_43_384 ();
 b15zdnd11an1n64x5 FILLER_43_448 ();
 b15zdnd00an1n01x5 FILLER_43_512 ();
 b15zdnd11an1n64x5 FILLER_43_565 ();
 b15zdnd11an1n32x5 FILLER_43_629 ();
 b15zdnd00an1n02x5 FILLER_43_661 ();
 b15zdnd00an1n01x5 FILLER_43_663 ();
 b15zdnd11an1n04x5 FILLER_43_667 ();
 b15zdnd11an1n04x5 FILLER_43_674 ();
 b15zdnd11an1n04x5 FILLER_43_681 ();
 b15zdnd11an1n64x5 FILLER_43_688 ();
 b15zdnd11an1n32x5 FILLER_43_752 ();
 b15zdnd11an1n08x5 FILLER_43_784 ();
 b15zdnd11an1n04x5 FILLER_43_792 ();
 b15zdnd00an1n02x5 FILLER_43_796 ();
 b15zdnd11an1n64x5 FILLER_43_850 ();
 b15zdnd11an1n32x5 FILLER_43_914 ();
 b15zdnd11an1n16x5 FILLER_43_946 ();
 b15zdnd00an1n01x5 FILLER_43_962 ();
 b15zdnd11an1n04x5 FILLER_43_966 ();
 b15zdnd11an1n08x5 FILLER_43_973 ();
 b15zdnd11an1n16x5 FILLER_43_988 ();
 b15zdnd11an1n08x5 FILLER_43_1004 ();
 b15zdnd11an1n64x5 FILLER_43_1019 ();
 b15zdnd11an1n64x5 FILLER_43_1083 ();
 b15zdnd11an1n64x5 FILLER_43_1147 ();
 b15zdnd11an1n32x5 FILLER_43_1211 ();
 b15zdnd11an1n16x5 FILLER_43_1243 ();
 b15zdnd11an1n04x5 FILLER_43_1259 ();
 b15zdnd00an1n02x5 FILLER_43_1263 ();
 b15zdnd00an1n01x5 FILLER_43_1265 ();
 b15zdnd11an1n64x5 FILLER_43_1269 ();
 b15zdnd11an1n32x5 FILLER_43_1333 ();
 b15zdnd11an1n16x5 FILLER_43_1365 ();
 b15zdnd00an1n02x5 FILLER_43_1381 ();
 b15zdnd11an1n64x5 FILLER_43_1427 ();
 b15zdnd11an1n64x5 FILLER_43_1491 ();
 b15zdnd11an1n64x5 FILLER_43_1555 ();
 b15zdnd11an1n64x5 FILLER_43_1619 ();
 b15zdnd11an1n64x5 FILLER_43_1683 ();
 b15zdnd11an1n64x5 FILLER_43_1747 ();
 b15zdnd11an1n64x5 FILLER_43_1811 ();
 b15zdnd11an1n64x5 FILLER_43_1875 ();
 b15zdnd11an1n64x5 FILLER_43_1939 ();
 b15zdnd11an1n64x5 FILLER_43_2003 ();
 b15zdnd11an1n64x5 FILLER_43_2067 ();
 b15zdnd11an1n64x5 FILLER_43_2131 ();
 b15zdnd11an1n64x5 FILLER_43_2195 ();
 b15zdnd11an1n16x5 FILLER_43_2259 ();
 b15zdnd11an1n08x5 FILLER_43_2275 ();
 b15zdnd00an1n01x5 FILLER_43_2283 ();
 b15zdnd11an1n64x5 FILLER_44_8 ();
 b15zdnd11an1n64x5 FILLER_44_72 ();
 b15zdnd11an1n64x5 FILLER_44_136 ();
 b15zdnd11an1n64x5 FILLER_44_200 ();
 b15zdnd11an1n64x5 FILLER_44_264 ();
 b15zdnd11an1n64x5 FILLER_44_328 ();
 b15zdnd11an1n64x5 FILLER_44_392 ();
 b15zdnd11an1n64x5 FILLER_44_456 ();
 b15zdnd11an1n08x5 FILLER_44_520 ();
 b15zdnd11an1n04x5 FILLER_44_531 ();
 b15zdnd11an1n04x5 FILLER_44_538 ();
 b15zdnd11an1n04x5 FILLER_44_545 ();
 b15zdnd11an1n64x5 FILLER_44_552 ();
 b15zdnd11an1n32x5 FILLER_44_616 ();
 b15zdnd11an1n08x5 FILLER_44_648 ();
 b15zdnd11an1n04x5 FILLER_44_656 ();
 b15zdnd00an1n02x5 FILLER_44_660 ();
 b15zdnd00an1n01x5 FILLER_44_662 ();
 b15zdnd11an1n04x5 FILLER_44_666 ();
 b15zdnd11an1n32x5 FILLER_44_673 ();
 b15zdnd11an1n08x5 FILLER_44_705 ();
 b15zdnd11an1n04x5 FILLER_44_713 ();
 b15zdnd00an1n01x5 FILLER_44_717 ();
 b15zdnd11an1n64x5 FILLER_44_726 ();
 b15zdnd11an1n04x5 FILLER_44_790 ();
 b15zdnd00an1n02x5 FILLER_44_794 ();
 b15zdnd00an1n01x5 FILLER_44_796 ();
 b15zdnd11an1n64x5 FILLER_44_849 ();
 b15zdnd11an1n16x5 FILLER_44_913 ();
 b15zdnd11an1n08x5 FILLER_44_929 ();
 b15zdnd11an1n04x5 FILLER_44_937 ();
 b15zdnd00an1n02x5 FILLER_44_941 ();
 b15zdnd00an1n01x5 FILLER_44_943 ();
 b15zdnd11an1n64x5 FILLER_44_996 ();
 b15zdnd11an1n64x5 FILLER_44_1060 ();
 b15zdnd11an1n64x5 FILLER_44_1124 ();
 b15zdnd11an1n32x5 FILLER_44_1188 ();
 b15zdnd11an1n16x5 FILLER_44_1220 ();
 b15zdnd11an1n04x5 FILLER_44_1236 ();
 b15zdnd11an1n08x5 FILLER_44_1292 ();
 b15zdnd00an1n02x5 FILLER_44_1300 ();
 b15zdnd11an1n04x5 FILLER_44_1305 ();
 b15zdnd11an1n64x5 FILLER_44_1312 ();
 b15zdnd11an1n16x5 FILLER_44_1376 ();
 b15zdnd11an1n08x5 FILLER_44_1392 ();
 b15zdnd11an1n04x5 FILLER_44_1400 ();
 b15zdnd00an1n02x5 FILLER_44_1404 ();
 b15zdnd11an1n64x5 FILLER_44_1409 ();
 b15zdnd11an1n64x5 FILLER_44_1473 ();
 b15zdnd11an1n64x5 FILLER_44_1537 ();
 b15zdnd11an1n64x5 FILLER_44_1601 ();
 b15zdnd11an1n64x5 FILLER_44_1665 ();
 b15zdnd11an1n64x5 FILLER_44_1729 ();
 b15zdnd11an1n64x5 FILLER_44_1793 ();
 b15zdnd11an1n64x5 FILLER_44_1857 ();
 b15zdnd11an1n64x5 FILLER_44_1921 ();
 b15zdnd11an1n64x5 FILLER_44_1985 ();
 b15zdnd11an1n64x5 FILLER_44_2049 ();
 b15zdnd11an1n32x5 FILLER_44_2113 ();
 b15zdnd11an1n08x5 FILLER_44_2145 ();
 b15zdnd00an1n01x5 FILLER_44_2153 ();
 b15zdnd11an1n64x5 FILLER_44_2162 ();
 b15zdnd11an1n32x5 FILLER_44_2226 ();
 b15zdnd11an1n16x5 FILLER_44_2258 ();
 b15zdnd00an1n02x5 FILLER_44_2274 ();
 b15zdnd11an1n64x5 FILLER_45_0 ();
 b15zdnd11an1n64x5 FILLER_45_64 ();
 b15zdnd11an1n64x5 FILLER_45_128 ();
 b15zdnd11an1n64x5 FILLER_45_192 ();
 b15zdnd11an1n64x5 FILLER_45_256 ();
 b15zdnd11an1n64x5 FILLER_45_320 ();
 b15zdnd11an1n64x5 FILLER_45_384 ();
 b15zdnd11an1n64x5 FILLER_45_448 ();
 b15zdnd00an1n02x5 FILLER_45_512 ();
 b15zdnd00an1n01x5 FILLER_45_514 ();
 b15zdnd11an1n64x5 FILLER_45_567 ();
 b15zdnd11an1n64x5 FILLER_45_631 ();
 b15zdnd11an1n64x5 FILLER_45_695 ();
 b15zdnd11an1n32x5 FILLER_45_759 ();
 b15zdnd11an1n08x5 FILLER_45_791 ();
 b15zdnd00an1n02x5 FILLER_45_799 ();
 b15zdnd00an1n01x5 FILLER_45_801 ();
 b15zdnd11an1n64x5 FILLER_45_854 ();
 b15zdnd11an1n32x5 FILLER_45_918 ();
 b15zdnd11an1n08x5 FILLER_45_950 ();
 b15zdnd11an1n64x5 FILLER_45_1010 ();
 b15zdnd11an1n32x5 FILLER_45_1074 ();
 b15zdnd11an1n16x5 FILLER_45_1106 ();
 b15zdnd11an1n08x5 FILLER_45_1122 ();
 b15zdnd11an1n64x5 FILLER_45_1133 ();
 b15zdnd11an1n32x5 FILLER_45_1197 ();
 b15zdnd11an1n16x5 FILLER_45_1229 ();
 b15zdnd11an1n08x5 FILLER_45_1245 ();
 b15zdnd11an1n04x5 FILLER_45_1253 ();
 b15zdnd00an1n01x5 FILLER_45_1257 ();
 b15zdnd11an1n04x5 FILLER_45_1261 ();
 b15zdnd11an1n16x5 FILLER_45_1268 ();
 b15zdnd11an1n64x5 FILLER_45_1336 ();
 b15zdnd11an1n32x5 FILLER_45_1400 ();
 b15zdnd11an1n08x5 FILLER_45_1432 ();
 b15zdnd11an1n64x5 FILLER_45_1443 ();
 b15zdnd11an1n64x5 FILLER_45_1507 ();
 b15zdnd11an1n64x5 FILLER_45_1571 ();
 b15zdnd11an1n64x5 FILLER_45_1635 ();
 b15zdnd11an1n64x5 FILLER_45_1699 ();
 b15zdnd11an1n64x5 FILLER_45_1763 ();
 b15zdnd11an1n64x5 FILLER_45_1827 ();
 b15zdnd11an1n64x5 FILLER_45_1891 ();
 b15zdnd11an1n64x5 FILLER_45_1955 ();
 b15zdnd11an1n64x5 FILLER_45_2019 ();
 b15zdnd11an1n64x5 FILLER_45_2083 ();
 b15zdnd11an1n64x5 FILLER_45_2147 ();
 b15zdnd11an1n32x5 FILLER_45_2211 ();
 b15zdnd11an1n08x5 FILLER_45_2243 ();
 b15zdnd11an1n16x5 FILLER_45_2254 ();
 b15zdnd11an1n08x5 FILLER_45_2270 ();
 b15zdnd11an1n04x5 FILLER_45_2278 ();
 b15zdnd00an1n02x5 FILLER_45_2282 ();
 b15zdnd11an1n64x5 FILLER_46_8 ();
 b15zdnd11an1n64x5 FILLER_46_72 ();
 b15zdnd11an1n64x5 FILLER_46_136 ();
 b15zdnd11an1n64x5 FILLER_46_200 ();
 b15zdnd11an1n64x5 FILLER_46_264 ();
 b15zdnd11an1n64x5 FILLER_46_328 ();
 b15zdnd11an1n64x5 FILLER_46_392 ();
 b15zdnd11an1n64x5 FILLER_46_456 ();
 b15zdnd11an1n08x5 FILLER_46_520 ();
 b15zdnd11an1n04x5 FILLER_46_528 ();
 b15zdnd00an1n02x5 FILLER_46_532 ();
 b15zdnd11an1n04x5 FILLER_46_537 ();
 b15zdnd11an1n64x5 FILLER_46_544 ();
 b15zdnd11an1n64x5 FILLER_46_608 ();
 b15zdnd11an1n32x5 FILLER_46_672 ();
 b15zdnd11an1n08x5 FILLER_46_704 ();
 b15zdnd11an1n04x5 FILLER_46_712 ();
 b15zdnd00an1n02x5 FILLER_46_716 ();
 b15zdnd11an1n64x5 FILLER_46_726 ();
 b15zdnd11an1n16x5 FILLER_46_790 ();
 b15zdnd11an1n08x5 FILLER_46_806 ();
 b15zdnd00an1n01x5 FILLER_46_814 ();
 b15zdnd11an1n04x5 FILLER_46_818 ();
 b15zdnd11an1n04x5 FILLER_46_825 ();
 b15zdnd11an1n04x5 FILLER_46_832 ();
 b15zdnd11an1n64x5 FILLER_46_839 ();
 b15zdnd11an1n32x5 FILLER_46_903 ();
 b15zdnd11an1n16x5 FILLER_46_935 ();
 b15zdnd11an1n08x5 FILLER_46_951 ();
 b15zdnd11an1n04x5 FILLER_46_959 ();
 b15zdnd00an1n01x5 FILLER_46_963 ();
 b15zdnd11an1n04x5 FILLER_46_967 ();
 b15zdnd11an1n04x5 FILLER_46_974 ();
 b15zdnd11an1n04x5 FILLER_46_981 ();
 b15zdnd11an1n16x5 FILLER_46_988 ();
 b15zdnd11an1n04x5 FILLER_46_1004 ();
 b15zdnd00an1n02x5 FILLER_46_1008 ();
 b15zdnd00an1n01x5 FILLER_46_1010 ();
 b15zdnd11an1n64x5 FILLER_46_1019 ();
 b15zdnd11an1n16x5 FILLER_46_1083 ();
 b15zdnd11an1n04x5 FILLER_46_1099 ();
 b15zdnd00an1n02x5 FILLER_46_1103 ();
 b15zdnd00an1n01x5 FILLER_46_1105 ();
 b15zdnd11an1n64x5 FILLER_46_1150 ();
 b15zdnd11an1n64x5 FILLER_46_1214 ();
 b15zdnd11an1n16x5 FILLER_46_1278 ();
 b15zdnd11an1n08x5 FILLER_46_1294 ();
 b15zdnd11an1n04x5 FILLER_46_1302 ();
 b15zdnd00an1n02x5 FILLER_46_1306 ();
 b15zdnd00an1n01x5 FILLER_46_1308 ();
 b15zdnd11an1n64x5 FILLER_46_1312 ();
 b15zdnd11an1n32x5 FILLER_46_1376 ();
 b15zdnd11an1n16x5 FILLER_46_1408 ();
 b15zdnd11an1n08x5 FILLER_46_1424 ();
 b15zdnd00an1n01x5 FILLER_46_1432 ();
 b15zdnd11an1n64x5 FILLER_46_1475 ();
 b15zdnd11an1n64x5 FILLER_46_1539 ();
 b15zdnd11an1n64x5 FILLER_46_1603 ();
 b15zdnd11an1n64x5 FILLER_46_1667 ();
 b15zdnd11an1n64x5 FILLER_46_1731 ();
 b15zdnd11an1n64x5 FILLER_46_1795 ();
 b15zdnd11an1n64x5 FILLER_46_1859 ();
 b15zdnd11an1n64x5 FILLER_46_1923 ();
 b15zdnd11an1n64x5 FILLER_46_1987 ();
 b15zdnd11an1n64x5 FILLER_46_2051 ();
 b15zdnd11an1n32x5 FILLER_46_2115 ();
 b15zdnd11an1n04x5 FILLER_46_2147 ();
 b15zdnd00an1n02x5 FILLER_46_2151 ();
 b15zdnd00an1n01x5 FILLER_46_2153 ();
 b15zdnd11an1n64x5 FILLER_46_2162 ();
 b15zdnd11an1n16x5 FILLER_46_2226 ();
 b15zdnd11an1n08x5 FILLER_46_2242 ();
 b15zdnd00an1n02x5 FILLER_46_2250 ();
 b15zdnd00an1n01x5 FILLER_46_2252 ();
 b15zdnd11an1n16x5 FILLER_46_2256 ();
 b15zdnd11an1n04x5 FILLER_46_2272 ();
 b15zdnd11an1n64x5 FILLER_47_0 ();
 b15zdnd11an1n64x5 FILLER_47_64 ();
 b15zdnd11an1n64x5 FILLER_47_128 ();
 b15zdnd11an1n64x5 FILLER_47_192 ();
 b15zdnd11an1n64x5 FILLER_47_256 ();
 b15zdnd11an1n64x5 FILLER_47_320 ();
 b15zdnd11an1n64x5 FILLER_47_384 ();
 b15zdnd11an1n64x5 FILLER_47_448 ();
 b15zdnd11an1n64x5 FILLER_47_512 ();
 b15zdnd11an1n64x5 FILLER_47_576 ();
 b15zdnd11an1n64x5 FILLER_47_640 ();
 b15zdnd11an1n64x5 FILLER_47_704 ();
 b15zdnd11an1n32x5 FILLER_47_768 ();
 b15zdnd11an1n16x5 FILLER_47_800 ();
 b15zdnd00an1n01x5 FILLER_47_816 ();
 b15zdnd11an1n08x5 FILLER_47_820 ();
 b15zdnd00an1n02x5 FILLER_47_828 ();
 b15zdnd00an1n01x5 FILLER_47_830 ();
 b15zdnd11an1n64x5 FILLER_47_834 ();
 b15zdnd11an1n64x5 FILLER_47_898 ();
 b15zdnd11an1n16x5 FILLER_47_962 ();
 b15zdnd11an1n04x5 FILLER_47_978 ();
 b15zdnd00an1n01x5 FILLER_47_982 ();
 b15zdnd11an1n64x5 FILLER_47_986 ();
 b15zdnd11an1n64x5 FILLER_47_1050 ();
 b15zdnd11an1n08x5 FILLER_47_1114 ();
 b15zdnd11an1n04x5 FILLER_47_1125 ();
 b15zdnd11an1n64x5 FILLER_47_1132 ();
 b15zdnd11an1n32x5 FILLER_47_1196 ();
 b15zdnd11an1n08x5 FILLER_47_1228 ();
 b15zdnd00an1n02x5 FILLER_47_1236 ();
 b15zdnd11an1n64x5 FILLER_47_1249 ();
 b15zdnd11an1n32x5 FILLER_47_1313 ();
 b15zdnd11an1n16x5 FILLER_47_1345 ();
 b15zdnd11an1n04x5 FILLER_47_1361 ();
 b15zdnd00an1n02x5 FILLER_47_1365 ();
 b15zdnd00an1n01x5 FILLER_47_1367 ();
 b15zdnd11an1n64x5 FILLER_47_1410 ();
 b15zdnd11an1n04x5 FILLER_47_1474 ();
 b15zdnd11an1n04x5 FILLER_47_1481 ();
 b15zdnd11an1n16x5 FILLER_47_1488 ();
 b15zdnd11an1n08x5 FILLER_47_1504 ();
 b15zdnd11an1n08x5 FILLER_47_1515 ();
 b15zdnd11an1n04x5 FILLER_47_1523 ();
 b15zdnd11an1n64x5 FILLER_47_1530 ();
 b15zdnd11an1n64x5 FILLER_47_1594 ();
 b15zdnd11an1n64x5 FILLER_47_1658 ();
 b15zdnd11an1n64x5 FILLER_47_1722 ();
 b15zdnd11an1n64x5 FILLER_47_1786 ();
 b15zdnd11an1n64x5 FILLER_47_1850 ();
 b15zdnd11an1n64x5 FILLER_47_1914 ();
 b15zdnd11an1n64x5 FILLER_47_1978 ();
 b15zdnd11an1n64x5 FILLER_47_2042 ();
 b15zdnd11an1n64x5 FILLER_47_2106 ();
 b15zdnd11an1n64x5 FILLER_47_2170 ();
 b15zdnd11an1n32x5 FILLER_47_2234 ();
 b15zdnd11an1n16x5 FILLER_47_2266 ();
 b15zdnd00an1n02x5 FILLER_47_2282 ();
 b15zdnd11an1n64x5 FILLER_48_8 ();
 b15zdnd11an1n64x5 FILLER_48_72 ();
 b15zdnd11an1n64x5 FILLER_48_136 ();
 b15zdnd11an1n64x5 FILLER_48_200 ();
 b15zdnd11an1n64x5 FILLER_48_264 ();
 b15zdnd11an1n64x5 FILLER_48_328 ();
 b15zdnd11an1n64x5 FILLER_48_392 ();
 b15zdnd11an1n64x5 FILLER_48_456 ();
 b15zdnd11an1n64x5 FILLER_48_520 ();
 b15zdnd11an1n64x5 FILLER_48_584 ();
 b15zdnd11an1n64x5 FILLER_48_648 ();
 b15zdnd11an1n04x5 FILLER_48_712 ();
 b15zdnd00an1n02x5 FILLER_48_716 ();
 b15zdnd11an1n64x5 FILLER_48_726 ();
 b15zdnd11an1n64x5 FILLER_48_790 ();
 b15zdnd11an1n64x5 FILLER_48_854 ();
 b15zdnd11an1n64x5 FILLER_48_918 ();
 b15zdnd11an1n64x5 FILLER_48_982 ();
 b15zdnd11an1n32x5 FILLER_48_1046 ();
 b15zdnd11an1n04x5 FILLER_48_1078 ();
 b15zdnd00an1n02x5 FILLER_48_1082 ();
 b15zdnd11an1n64x5 FILLER_48_1098 ();
 b15zdnd11an1n32x5 FILLER_48_1162 ();
 b15zdnd11an1n08x5 FILLER_48_1194 ();
 b15zdnd00an1n01x5 FILLER_48_1202 ();
 b15zdnd11an1n08x5 FILLER_48_1245 ();
 b15zdnd11an1n64x5 FILLER_48_1261 ();
 b15zdnd11an1n64x5 FILLER_48_1325 ();
 b15zdnd11an1n64x5 FILLER_48_1389 ();
 b15zdnd11an1n08x5 FILLER_48_1453 ();
 b15zdnd00an1n02x5 FILLER_48_1461 ();
 b15zdnd11an1n64x5 FILLER_48_1507 ();
 b15zdnd11an1n64x5 FILLER_48_1571 ();
 b15zdnd11an1n64x5 FILLER_48_1635 ();
 b15zdnd11an1n64x5 FILLER_48_1699 ();
 b15zdnd11an1n64x5 FILLER_48_1763 ();
 b15zdnd11an1n64x5 FILLER_48_1827 ();
 b15zdnd11an1n64x5 FILLER_48_1891 ();
 b15zdnd11an1n64x5 FILLER_48_1955 ();
 b15zdnd11an1n64x5 FILLER_48_2019 ();
 b15zdnd11an1n64x5 FILLER_48_2083 ();
 b15zdnd11an1n04x5 FILLER_48_2147 ();
 b15zdnd00an1n02x5 FILLER_48_2151 ();
 b15zdnd00an1n01x5 FILLER_48_2153 ();
 b15zdnd11an1n64x5 FILLER_48_2162 ();
 b15zdnd11an1n32x5 FILLER_48_2226 ();
 b15zdnd11an1n16x5 FILLER_48_2258 ();
 b15zdnd00an1n02x5 FILLER_48_2274 ();
 b15zdnd11an1n64x5 FILLER_49_0 ();
 b15zdnd11an1n64x5 FILLER_49_64 ();
 b15zdnd11an1n64x5 FILLER_49_128 ();
 b15zdnd11an1n64x5 FILLER_49_192 ();
 b15zdnd11an1n64x5 FILLER_49_256 ();
 b15zdnd11an1n64x5 FILLER_49_320 ();
 b15zdnd11an1n64x5 FILLER_49_384 ();
 b15zdnd11an1n64x5 FILLER_49_448 ();
 b15zdnd11an1n64x5 FILLER_49_512 ();
 b15zdnd11an1n64x5 FILLER_49_576 ();
 b15zdnd11an1n64x5 FILLER_49_640 ();
 b15zdnd11an1n64x5 FILLER_49_704 ();
 b15zdnd11an1n64x5 FILLER_49_768 ();
 b15zdnd11an1n64x5 FILLER_49_832 ();
 b15zdnd11an1n64x5 FILLER_49_896 ();
 b15zdnd11an1n64x5 FILLER_49_960 ();
 b15zdnd11an1n64x5 FILLER_49_1024 ();
 b15zdnd11an1n64x5 FILLER_49_1088 ();
 b15zdnd11an1n64x5 FILLER_49_1152 ();
 b15zdnd11an1n04x5 FILLER_49_1216 ();
 b15zdnd00an1n02x5 FILLER_49_1220 ();
 b15zdnd11an1n64x5 FILLER_49_1233 ();
 b15zdnd11an1n64x5 FILLER_49_1297 ();
 b15zdnd11an1n16x5 FILLER_49_1361 ();
 b15zdnd11an1n04x5 FILLER_49_1377 ();
 b15zdnd00an1n02x5 FILLER_49_1381 ();
 b15zdnd00an1n01x5 FILLER_49_1383 ();
 b15zdnd11an1n04x5 FILLER_49_1426 ();
 b15zdnd11an1n04x5 FILLER_49_1434 ();
 b15zdnd11an1n32x5 FILLER_49_1452 ();
 b15zdnd00an1n02x5 FILLER_49_1484 ();
 b15zdnd11an1n32x5 FILLER_49_1489 ();
 b15zdnd11an1n04x5 FILLER_49_1521 ();
 b15zdnd00an1n02x5 FILLER_49_1525 ();
 b15zdnd11an1n64x5 FILLER_49_1530 ();
 b15zdnd11an1n64x5 FILLER_49_1594 ();
 b15zdnd11an1n64x5 FILLER_49_1658 ();
 b15zdnd11an1n64x5 FILLER_49_1722 ();
 b15zdnd11an1n64x5 FILLER_49_1786 ();
 b15zdnd11an1n64x5 FILLER_49_1850 ();
 b15zdnd11an1n64x5 FILLER_49_1914 ();
 b15zdnd11an1n64x5 FILLER_49_1978 ();
 b15zdnd11an1n64x5 FILLER_49_2042 ();
 b15zdnd11an1n64x5 FILLER_49_2106 ();
 b15zdnd11an1n64x5 FILLER_49_2170 ();
 b15zdnd11an1n32x5 FILLER_49_2234 ();
 b15zdnd11an1n16x5 FILLER_49_2266 ();
 b15zdnd00an1n02x5 FILLER_49_2282 ();
 b15zdnd11an1n64x5 FILLER_50_8 ();
 b15zdnd11an1n64x5 FILLER_50_72 ();
 b15zdnd11an1n64x5 FILLER_50_136 ();
 b15zdnd11an1n64x5 FILLER_50_200 ();
 b15zdnd11an1n64x5 FILLER_50_264 ();
 b15zdnd11an1n64x5 FILLER_50_328 ();
 b15zdnd11an1n64x5 FILLER_50_392 ();
 b15zdnd11an1n64x5 FILLER_50_456 ();
 b15zdnd11an1n64x5 FILLER_50_520 ();
 b15zdnd11an1n64x5 FILLER_50_584 ();
 b15zdnd11an1n64x5 FILLER_50_648 ();
 b15zdnd11an1n04x5 FILLER_50_712 ();
 b15zdnd00an1n02x5 FILLER_50_716 ();
 b15zdnd11an1n64x5 FILLER_50_726 ();
 b15zdnd11an1n64x5 FILLER_50_790 ();
 b15zdnd11an1n64x5 FILLER_50_854 ();
 b15zdnd11an1n64x5 FILLER_50_918 ();
 b15zdnd11an1n64x5 FILLER_50_982 ();
 b15zdnd11an1n64x5 FILLER_50_1046 ();
 b15zdnd11an1n64x5 FILLER_50_1110 ();
 b15zdnd11an1n32x5 FILLER_50_1174 ();
 b15zdnd11an1n64x5 FILLER_50_1216 ();
 b15zdnd11an1n64x5 FILLER_50_1280 ();
 b15zdnd11an1n64x5 FILLER_50_1344 ();
 b15zdnd11an1n64x5 FILLER_50_1408 ();
 b15zdnd11an1n16x5 FILLER_50_1472 ();
 b15zdnd11an1n08x5 FILLER_50_1488 ();
 b15zdnd00an1n01x5 FILLER_50_1496 ();
 b15zdnd11an1n04x5 FILLER_50_1511 ();
 b15zdnd11an1n64x5 FILLER_50_1557 ();
 b15zdnd11an1n64x5 FILLER_50_1621 ();
 b15zdnd11an1n64x5 FILLER_50_1685 ();
 b15zdnd11an1n64x5 FILLER_50_1749 ();
 b15zdnd11an1n64x5 FILLER_50_1813 ();
 b15zdnd11an1n64x5 FILLER_50_1877 ();
 b15zdnd11an1n64x5 FILLER_50_1941 ();
 b15zdnd11an1n64x5 FILLER_50_2005 ();
 b15zdnd11an1n64x5 FILLER_50_2069 ();
 b15zdnd11an1n16x5 FILLER_50_2133 ();
 b15zdnd11an1n04x5 FILLER_50_2149 ();
 b15zdnd00an1n01x5 FILLER_50_2153 ();
 b15zdnd11an1n64x5 FILLER_50_2162 ();
 b15zdnd11an1n32x5 FILLER_50_2226 ();
 b15zdnd11an1n16x5 FILLER_50_2258 ();
 b15zdnd00an1n02x5 FILLER_50_2274 ();
 b15zdnd11an1n64x5 FILLER_51_0 ();
 b15zdnd11an1n64x5 FILLER_51_64 ();
 b15zdnd11an1n64x5 FILLER_51_128 ();
 b15zdnd11an1n64x5 FILLER_51_192 ();
 b15zdnd11an1n64x5 FILLER_51_256 ();
 b15zdnd11an1n64x5 FILLER_51_320 ();
 b15zdnd11an1n64x5 FILLER_51_384 ();
 b15zdnd11an1n64x5 FILLER_51_448 ();
 b15zdnd11an1n64x5 FILLER_51_512 ();
 b15zdnd11an1n64x5 FILLER_51_576 ();
 b15zdnd11an1n64x5 FILLER_51_640 ();
 b15zdnd11an1n64x5 FILLER_51_704 ();
 b15zdnd11an1n64x5 FILLER_51_768 ();
 b15zdnd11an1n64x5 FILLER_51_832 ();
 b15zdnd11an1n64x5 FILLER_51_896 ();
 b15zdnd11an1n64x5 FILLER_51_960 ();
 b15zdnd11an1n64x5 FILLER_51_1024 ();
 b15zdnd11an1n16x5 FILLER_51_1088 ();
 b15zdnd11an1n08x5 FILLER_51_1104 ();
 b15zdnd00an1n02x5 FILLER_51_1112 ();
 b15zdnd00an1n01x5 FILLER_51_1114 ();
 b15zdnd11an1n64x5 FILLER_51_1122 ();
 b15zdnd11an1n64x5 FILLER_51_1186 ();
 b15zdnd11an1n64x5 FILLER_51_1250 ();
 b15zdnd11an1n64x5 FILLER_51_1314 ();
 b15zdnd11an1n64x5 FILLER_51_1378 ();
 b15zdnd11an1n64x5 FILLER_51_1442 ();
 b15zdnd11an1n16x5 FILLER_51_1506 ();
 b15zdnd11an1n64x5 FILLER_51_1536 ();
 b15zdnd11an1n64x5 FILLER_51_1600 ();
 b15zdnd11an1n64x5 FILLER_51_1664 ();
 b15zdnd11an1n32x5 FILLER_51_1728 ();
 b15zdnd00an1n01x5 FILLER_51_1760 ();
 b15zdnd11an1n64x5 FILLER_51_1769 ();
 b15zdnd11an1n64x5 FILLER_51_1833 ();
 b15zdnd11an1n64x5 FILLER_51_1897 ();
 b15zdnd11an1n64x5 FILLER_51_1961 ();
 b15zdnd11an1n64x5 FILLER_51_2025 ();
 b15zdnd11an1n64x5 FILLER_51_2089 ();
 b15zdnd11an1n64x5 FILLER_51_2153 ();
 b15zdnd11an1n64x5 FILLER_51_2217 ();
 b15zdnd00an1n02x5 FILLER_51_2281 ();
 b15zdnd00an1n01x5 FILLER_51_2283 ();
 b15zdnd11an1n64x5 FILLER_52_8 ();
 b15zdnd11an1n64x5 FILLER_52_72 ();
 b15zdnd11an1n64x5 FILLER_52_136 ();
 b15zdnd11an1n64x5 FILLER_52_200 ();
 b15zdnd11an1n64x5 FILLER_52_264 ();
 b15zdnd11an1n64x5 FILLER_52_328 ();
 b15zdnd11an1n16x5 FILLER_52_392 ();
 b15zdnd11an1n08x5 FILLER_52_408 ();
 b15zdnd00an1n01x5 FILLER_52_416 ();
 b15zdnd11an1n64x5 FILLER_52_420 ();
 b15zdnd11an1n64x5 FILLER_52_484 ();
 b15zdnd11an1n64x5 FILLER_52_548 ();
 b15zdnd11an1n64x5 FILLER_52_612 ();
 b15zdnd11an1n32x5 FILLER_52_676 ();
 b15zdnd11an1n08x5 FILLER_52_708 ();
 b15zdnd00an1n02x5 FILLER_52_716 ();
 b15zdnd11an1n64x5 FILLER_52_726 ();
 b15zdnd11an1n64x5 FILLER_52_790 ();
 b15zdnd11an1n64x5 FILLER_52_854 ();
 b15zdnd11an1n64x5 FILLER_52_918 ();
 b15zdnd11an1n64x5 FILLER_52_982 ();
 b15zdnd11an1n32x5 FILLER_52_1046 ();
 b15zdnd11an1n08x5 FILLER_52_1078 ();
 b15zdnd00an1n02x5 FILLER_52_1086 ();
 b15zdnd11an1n16x5 FILLER_52_1100 ();
 b15zdnd11an1n64x5 FILLER_52_1158 ();
 b15zdnd11an1n64x5 FILLER_52_1222 ();
 b15zdnd11an1n64x5 FILLER_52_1286 ();
 b15zdnd11an1n08x5 FILLER_52_1350 ();
 b15zdnd11an1n04x5 FILLER_52_1358 ();
 b15zdnd00an1n02x5 FILLER_52_1362 ();
 b15zdnd00an1n01x5 FILLER_52_1364 ();
 b15zdnd11an1n64x5 FILLER_52_1368 ();
 b15zdnd11an1n64x5 FILLER_52_1432 ();
 b15zdnd11an1n64x5 FILLER_52_1496 ();
 b15zdnd11an1n64x5 FILLER_52_1560 ();
 b15zdnd11an1n64x5 FILLER_52_1624 ();
 b15zdnd11an1n64x5 FILLER_52_1688 ();
 b15zdnd11an1n64x5 FILLER_52_1752 ();
 b15zdnd11an1n64x5 FILLER_52_1816 ();
 b15zdnd11an1n32x5 FILLER_52_1880 ();
 b15zdnd11an1n08x5 FILLER_52_1912 ();
 b15zdnd11an1n04x5 FILLER_52_1920 ();
 b15zdnd00an1n02x5 FILLER_52_1924 ();
 b15zdnd11an1n04x5 FILLER_52_1929 ();
 b15zdnd11an1n64x5 FILLER_52_1936 ();
 b15zdnd11an1n64x5 FILLER_52_2000 ();
 b15zdnd11an1n64x5 FILLER_52_2064 ();
 b15zdnd11an1n16x5 FILLER_52_2128 ();
 b15zdnd11an1n08x5 FILLER_52_2144 ();
 b15zdnd00an1n02x5 FILLER_52_2152 ();
 b15zdnd11an1n64x5 FILLER_52_2162 ();
 b15zdnd11an1n32x5 FILLER_52_2226 ();
 b15zdnd11an1n16x5 FILLER_52_2258 ();
 b15zdnd00an1n02x5 FILLER_52_2274 ();
 b15zdnd11an1n64x5 FILLER_53_0 ();
 b15zdnd11an1n64x5 FILLER_53_64 ();
 b15zdnd11an1n64x5 FILLER_53_128 ();
 b15zdnd11an1n64x5 FILLER_53_192 ();
 b15zdnd11an1n64x5 FILLER_53_256 ();
 b15zdnd11an1n64x5 FILLER_53_320 ();
 b15zdnd11an1n16x5 FILLER_53_384 ();
 b15zdnd11an1n04x5 FILLER_53_400 ();
 b15zdnd00an1n02x5 FILLER_53_404 ();
 b15zdnd00an1n01x5 FILLER_53_406 ();
 b15zdnd11an1n64x5 FILLER_53_459 ();
 b15zdnd11an1n64x5 FILLER_53_523 ();
 b15zdnd11an1n64x5 FILLER_53_587 ();
 b15zdnd11an1n16x5 FILLER_53_651 ();
 b15zdnd11an1n04x5 FILLER_53_667 ();
 b15zdnd11an1n64x5 FILLER_53_675 ();
 b15zdnd11an1n64x5 FILLER_53_739 ();
 b15zdnd11an1n64x5 FILLER_53_803 ();
 b15zdnd11an1n64x5 FILLER_53_867 ();
 b15zdnd11an1n64x5 FILLER_53_931 ();
 b15zdnd11an1n64x5 FILLER_53_995 ();
 b15zdnd11an1n32x5 FILLER_53_1059 ();
 b15zdnd11an1n64x5 FILLER_53_1108 ();
 b15zdnd11an1n64x5 FILLER_53_1172 ();
 b15zdnd11an1n64x5 FILLER_53_1236 ();
 b15zdnd11an1n64x5 FILLER_53_1300 ();
 b15zdnd11an1n64x5 FILLER_53_1364 ();
 b15zdnd11an1n64x5 FILLER_53_1428 ();
 b15zdnd11an1n64x5 FILLER_53_1492 ();
 b15zdnd11an1n64x5 FILLER_53_1556 ();
 b15zdnd11an1n64x5 FILLER_53_1620 ();
 b15zdnd11an1n64x5 FILLER_53_1684 ();
 b15zdnd11an1n64x5 FILLER_53_1748 ();
 b15zdnd11an1n64x5 FILLER_53_1812 ();
 b15zdnd11an1n32x5 FILLER_53_1876 ();
 b15zdnd11an1n64x5 FILLER_53_1960 ();
 b15zdnd11an1n64x5 FILLER_53_2024 ();
 b15zdnd11an1n64x5 FILLER_53_2088 ();
 b15zdnd11an1n64x5 FILLER_53_2152 ();
 b15zdnd11an1n64x5 FILLER_53_2216 ();
 b15zdnd11an1n04x5 FILLER_53_2280 ();
 b15zdnd11an1n64x5 FILLER_54_8 ();
 b15zdnd11an1n64x5 FILLER_54_72 ();
 b15zdnd11an1n64x5 FILLER_54_136 ();
 b15zdnd11an1n64x5 FILLER_54_200 ();
 b15zdnd11an1n64x5 FILLER_54_264 ();
 b15zdnd11an1n64x5 FILLER_54_328 ();
 b15zdnd11an1n16x5 FILLER_54_392 ();
 b15zdnd11an1n08x5 FILLER_54_408 ();
 b15zdnd11an1n04x5 FILLER_54_416 ();
 b15zdnd00an1n02x5 FILLER_54_420 ();
 b15zdnd00an1n01x5 FILLER_54_422 ();
 b15zdnd11an1n04x5 FILLER_54_426 ();
 b15zdnd11an1n64x5 FILLER_54_433 ();
 b15zdnd11an1n64x5 FILLER_54_497 ();
 b15zdnd11an1n64x5 FILLER_54_561 ();
 b15zdnd11an1n32x5 FILLER_54_625 ();
 b15zdnd11an1n04x5 FILLER_54_657 ();
 b15zdnd00an1n01x5 FILLER_54_661 ();
 b15zdnd11an1n04x5 FILLER_54_666 ();
 b15zdnd00an1n01x5 FILLER_54_670 ();
 b15zdnd11an1n08x5 FILLER_54_675 ();
 b15zdnd11an1n04x5 FILLER_54_683 ();
 b15zdnd11an1n16x5 FILLER_54_691 ();
 b15zdnd11an1n08x5 FILLER_54_707 ();
 b15zdnd00an1n02x5 FILLER_54_715 ();
 b15zdnd00an1n01x5 FILLER_54_717 ();
 b15zdnd11an1n64x5 FILLER_54_726 ();
 b15zdnd11an1n64x5 FILLER_54_790 ();
 b15zdnd11an1n64x5 FILLER_54_854 ();
 b15zdnd11an1n64x5 FILLER_54_918 ();
 b15zdnd11an1n64x5 FILLER_54_982 ();
 b15zdnd11an1n64x5 FILLER_54_1046 ();
 b15zdnd11an1n64x5 FILLER_54_1110 ();
 b15zdnd11an1n64x5 FILLER_54_1174 ();
 b15zdnd11an1n64x5 FILLER_54_1238 ();
 b15zdnd11an1n64x5 FILLER_54_1302 ();
 b15zdnd11an1n08x5 FILLER_54_1366 ();
 b15zdnd11an1n04x5 FILLER_54_1374 ();
 b15zdnd00an1n02x5 FILLER_54_1378 ();
 b15zdnd00an1n01x5 FILLER_54_1380 ();
 b15zdnd11an1n32x5 FILLER_54_1384 ();
 b15zdnd11an1n16x5 FILLER_54_1416 ();
 b15zdnd11an1n08x5 FILLER_54_1432 ();
 b15zdnd00an1n02x5 FILLER_54_1440 ();
 b15zdnd00an1n01x5 FILLER_54_1442 ();
 b15zdnd11an1n64x5 FILLER_54_1452 ();
 b15zdnd11an1n32x5 FILLER_54_1516 ();
 b15zdnd11an1n16x5 FILLER_54_1548 ();
 b15zdnd11an1n04x5 FILLER_54_1564 ();
 b15zdnd00an1n01x5 FILLER_54_1568 ();
 b15zdnd11an1n64x5 FILLER_54_1613 ();
 b15zdnd11an1n64x5 FILLER_54_1677 ();
 b15zdnd11an1n64x5 FILLER_54_1741 ();
 b15zdnd11an1n64x5 FILLER_54_1805 ();
 b15zdnd11an1n32x5 FILLER_54_1869 ();
 b15zdnd11an1n04x5 FILLER_54_1901 ();
 b15zdnd00an1n02x5 FILLER_54_1905 ();
 b15zdnd11an1n64x5 FILLER_54_1959 ();
 b15zdnd11an1n64x5 FILLER_54_2023 ();
 b15zdnd11an1n64x5 FILLER_54_2087 ();
 b15zdnd00an1n02x5 FILLER_54_2151 ();
 b15zdnd00an1n01x5 FILLER_54_2153 ();
 b15zdnd11an1n64x5 FILLER_54_2162 ();
 b15zdnd11an1n32x5 FILLER_54_2226 ();
 b15zdnd11an1n16x5 FILLER_54_2258 ();
 b15zdnd00an1n02x5 FILLER_54_2274 ();
 b15zdnd11an1n64x5 FILLER_55_0 ();
 b15zdnd11an1n64x5 FILLER_55_64 ();
 b15zdnd11an1n64x5 FILLER_55_128 ();
 b15zdnd11an1n64x5 FILLER_55_192 ();
 b15zdnd11an1n64x5 FILLER_55_256 ();
 b15zdnd11an1n64x5 FILLER_55_320 ();
 b15zdnd11an1n64x5 FILLER_55_384 ();
 b15zdnd11an1n04x5 FILLER_55_448 ();
 b15zdnd00an1n01x5 FILLER_55_452 ();
 b15zdnd11an1n64x5 FILLER_55_459 ();
 b15zdnd11an1n64x5 FILLER_55_523 ();
 b15zdnd11an1n64x5 FILLER_55_587 ();
 b15zdnd11an1n04x5 FILLER_55_651 ();
 b15zdnd00an1n02x5 FILLER_55_655 ();
 b15zdnd00an1n01x5 FILLER_55_657 ();
 b15zdnd11an1n32x5 FILLER_55_662 ();
 b15zdnd11an1n08x5 FILLER_55_694 ();
 b15zdnd11an1n64x5 FILLER_55_710 ();
 b15zdnd11an1n64x5 FILLER_55_774 ();
 b15zdnd11an1n64x5 FILLER_55_838 ();
 b15zdnd11an1n64x5 FILLER_55_902 ();
 b15zdnd11an1n64x5 FILLER_55_966 ();
 b15zdnd11an1n64x5 FILLER_55_1030 ();
 b15zdnd11an1n64x5 FILLER_55_1094 ();
 b15zdnd11an1n64x5 FILLER_55_1158 ();
 b15zdnd11an1n64x5 FILLER_55_1222 ();
 b15zdnd11an1n32x5 FILLER_55_1286 ();
 b15zdnd11an1n16x5 FILLER_55_1318 ();
 b15zdnd11an1n32x5 FILLER_55_1346 ();
 b15zdnd11an1n04x5 FILLER_55_1378 ();
 b15zdnd11an1n64x5 FILLER_55_1395 ();
 b15zdnd11an1n64x5 FILLER_55_1459 ();
 b15zdnd11an1n64x5 FILLER_55_1523 ();
 b15zdnd11an1n04x5 FILLER_55_1587 ();
 b15zdnd11an1n04x5 FILLER_55_1594 ();
 b15zdnd11an1n32x5 FILLER_55_1601 ();
 b15zdnd11an1n16x5 FILLER_55_1633 ();
 b15zdnd00an1n02x5 FILLER_55_1649 ();
 b15zdnd00an1n01x5 FILLER_55_1651 ();
 b15zdnd11an1n64x5 FILLER_55_1656 ();
 b15zdnd11an1n64x5 FILLER_55_1720 ();
 b15zdnd11an1n64x5 FILLER_55_1784 ();
 b15zdnd11an1n64x5 FILLER_55_1848 ();
 b15zdnd11an1n08x5 FILLER_55_1912 ();
 b15zdnd11an1n04x5 FILLER_55_1920 ();
 b15zdnd00an1n01x5 FILLER_55_1924 ();
 b15zdnd11an1n04x5 FILLER_55_1928 ();
 b15zdnd11an1n04x5 FILLER_55_1935 ();
 b15zdnd11an1n32x5 FILLER_55_1942 ();
 b15zdnd11an1n16x5 FILLER_55_1974 ();
 b15zdnd11an1n08x5 FILLER_55_1990 ();
 b15zdnd11an1n04x5 FILLER_55_1998 ();
 b15zdnd00an1n02x5 FILLER_55_2002 ();
 b15zdnd11an1n64x5 FILLER_55_2007 ();
 b15zdnd11an1n64x5 FILLER_55_2071 ();
 b15zdnd11an1n64x5 FILLER_55_2135 ();
 b15zdnd11an1n64x5 FILLER_55_2199 ();
 b15zdnd11an1n16x5 FILLER_55_2263 ();
 b15zdnd11an1n04x5 FILLER_55_2279 ();
 b15zdnd00an1n01x5 FILLER_55_2283 ();
 b15zdnd11an1n64x5 FILLER_56_8 ();
 b15zdnd11an1n64x5 FILLER_56_72 ();
 b15zdnd11an1n64x5 FILLER_56_136 ();
 b15zdnd11an1n64x5 FILLER_56_200 ();
 b15zdnd11an1n64x5 FILLER_56_264 ();
 b15zdnd11an1n64x5 FILLER_56_328 ();
 b15zdnd11an1n32x5 FILLER_56_392 ();
 b15zdnd11an1n16x5 FILLER_56_424 ();
 b15zdnd11an1n08x5 FILLER_56_440 ();
 b15zdnd11an1n04x5 FILLER_56_448 ();
 b15zdnd00an1n01x5 FILLER_56_452 ();
 b15zdnd11an1n64x5 FILLER_56_457 ();
 b15zdnd11an1n64x5 FILLER_56_521 ();
 b15zdnd11an1n64x5 FILLER_56_585 ();
 b15zdnd11an1n08x5 FILLER_56_649 ();
 b15zdnd00an1n02x5 FILLER_56_657 ();
 b15zdnd00an1n01x5 FILLER_56_659 ();
 b15zdnd11an1n32x5 FILLER_56_664 ();
 b15zdnd11an1n16x5 FILLER_56_696 ();
 b15zdnd11an1n04x5 FILLER_56_712 ();
 b15zdnd00an1n02x5 FILLER_56_716 ();
 b15zdnd11an1n64x5 FILLER_56_726 ();
 b15zdnd11an1n64x5 FILLER_56_790 ();
 b15zdnd11an1n64x5 FILLER_56_854 ();
 b15zdnd11an1n64x5 FILLER_56_918 ();
 b15zdnd11an1n64x5 FILLER_56_982 ();
 b15zdnd11an1n64x5 FILLER_56_1046 ();
 b15zdnd11an1n64x5 FILLER_56_1110 ();
 b15zdnd11an1n64x5 FILLER_56_1174 ();
 b15zdnd11an1n64x5 FILLER_56_1238 ();
 b15zdnd11an1n64x5 FILLER_56_1302 ();
 b15zdnd11an1n64x5 FILLER_56_1366 ();
 b15zdnd11an1n64x5 FILLER_56_1430 ();
 b15zdnd11an1n64x5 FILLER_56_1494 ();
 b15zdnd11an1n32x5 FILLER_56_1558 ();
 b15zdnd00an1n01x5 FILLER_56_1590 ();
 b15zdnd11an1n32x5 FILLER_56_1594 ();
 b15zdnd11an1n16x5 FILLER_56_1626 ();
 b15zdnd11an1n04x5 FILLER_56_1648 ();
 b15zdnd11an1n64x5 FILLER_56_1656 ();
 b15zdnd11an1n16x5 FILLER_56_1720 ();
 b15zdnd11an1n08x5 FILLER_56_1736 ();
 b15zdnd11an1n04x5 FILLER_56_1744 ();
 b15zdnd00an1n02x5 FILLER_56_1748 ();
 b15zdnd00an1n01x5 FILLER_56_1750 ();
 b15zdnd11an1n64x5 FILLER_56_1759 ();
 b15zdnd11an1n64x5 FILLER_56_1823 ();
 b15zdnd11an1n32x5 FILLER_56_1887 ();
 b15zdnd11an1n08x5 FILLER_56_1919 ();
 b15zdnd11an1n04x5 FILLER_56_1927 ();
 b15zdnd00an1n02x5 FILLER_56_1931 ();
 b15zdnd11an1n64x5 FILLER_56_1936 ();
 b15zdnd11an1n04x5 FILLER_56_2000 ();
 b15zdnd11an1n64x5 FILLER_56_2031 ();
 b15zdnd11an1n32x5 FILLER_56_2095 ();
 b15zdnd11an1n16x5 FILLER_56_2127 ();
 b15zdnd11an1n08x5 FILLER_56_2143 ();
 b15zdnd00an1n02x5 FILLER_56_2151 ();
 b15zdnd00an1n01x5 FILLER_56_2153 ();
 b15zdnd11an1n64x5 FILLER_56_2162 ();
 b15zdnd11an1n32x5 FILLER_56_2226 ();
 b15zdnd11an1n16x5 FILLER_56_2258 ();
 b15zdnd00an1n02x5 FILLER_56_2274 ();
 b15zdnd11an1n64x5 FILLER_57_0 ();
 b15zdnd11an1n64x5 FILLER_57_64 ();
 b15zdnd11an1n64x5 FILLER_57_128 ();
 b15zdnd11an1n64x5 FILLER_57_192 ();
 b15zdnd11an1n64x5 FILLER_57_256 ();
 b15zdnd11an1n64x5 FILLER_57_320 ();
 b15zdnd11an1n64x5 FILLER_57_384 ();
 b15zdnd11an1n64x5 FILLER_57_448 ();
 b15zdnd11an1n16x5 FILLER_57_512 ();
 b15zdnd11an1n08x5 FILLER_57_528 ();
 b15zdnd11an1n64x5 FILLER_57_540 ();
 b15zdnd11an1n64x5 FILLER_57_604 ();
 b15zdnd11an1n64x5 FILLER_57_668 ();
 b15zdnd11an1n64x5 FILLER_57_732 ();
 b15zdnd11an1n64x5 FILLER_57_796 ();
 b15zdnd11an1n64x5 FILLER_57_860 ();
 b15zdnd11an1n32x5 FILLER_57_924 ();
 b15zdnd11an1n08x5 FILLER_57_956 ();
 b15zdnd11an1n04x5 FILLER_57_964 ();
 b15zdnd00an1n02x5 FILLER_57_968 ();
 b15zdnd00an1n01x5 FILLER_57_970 ();
 b15zdnd11an1n64x5 FILLER_57_975 ();
 b15zdnd11an1n64x5 FILLER_57_1039 ();
 b15zdnd11an1n16x5 FILLER_57_1103 ();
 b15zdnd11an1n04x5 FILLER_57_1119 ();
 b15zdnd00an1n01x5 FILLER_57_1123 ();
 b15zdnd11an1n64x5 FILLER_57_1138 ();
 b15zdnd11an1n32x5 FILLER_57_1202 ();
 b15zdnd11an1n16x5 FILLER_57_1234 ();
 b15zdnd11an1n08x5 FILLER_57_1250 ();
 b15zdnd11an1n04x5 FILLER_57_1258 ();
 b15zdnd00an1n02x5 FILLER_57_1262 ();
 b15zdnd11an1n64x5 FILLER_57_1271 ();
 b15zdnd11an1n64x5 FILLER_57_1335 ();
 b15zdnd11an1n64x5 FILLER_57_1399 ();
 b15zdnd11an1n64x5 FILLER_57_1463 ();
 b15zdnd11an1n64x5 FILLER_57_1527 ();
 b15zdnd11an1n32x5 FILLER_57_1591 ();
 b15zdnd11an1n16x5 FILLER_57_1623 ();
 b15zdnd11an1n04x5 FILLER_57_1639 ();
 b15zdnd11an1n64x5 FILLER_57_1647 ();
 b15zdnd11an1n64x5 FILLER_57_1711 ();
 b15zdnd11an1n08x5 FILLER_57_1775 ();
 b15zdnd11an1n04x5 FILLER_57_1783 ();
 b15zdnd00an1n02x5 FILLER_57_1787 ();
 b15zdnd11an1n64x5 FILLER_57_1793 ();
 b15zdnd11an1n64x5 FILLER_57_1857 ();
 b15zdnd11an1n64x5 FILLER_57_1921 ();
 b15zdnd11an1n64x5 FILLER_57_1985 ();
 b15zdnd11an1n64x5 FILLER_57_2049 ();
 b15zdnd11an1n64x5 FILLER_57_2113 ();
 b15zdnd11an1n64x5 FILLER_57_2177 ();
 b15zdnd11an1n32x5 FILLER_57_2241 ();
 b15zdnd11an1n08x5 FILLER_57_2273 ();
 b15zdnd00an1n02x5 FILLER_57_2281 ();
 b15zdnd00an1n01x5 FILLER_57_2283 ();
 b15zdnd11an1n64x5 FILLER_58_8 ();
 b15zdnd11an1n64x5 FILLER_58_72 ();
 b15zdnd11an1n64x5 FILLER_58_136 ();
 b15zdnd11an1n64x5 FILLER_58_200 ();
 b15zdnd11an1n64x5 FILLER_58_264 ();
 b15zdnd11an1n64x5 FILLER_58_328 ();
 b15zdnd11an1n64x5 FILLER_58_392 ();
 b15zdnd11an1n64x5 FILLER_58_456 ();
 b15zdnd11an1n08x5 FILLER_58_520 ();
 b15zdnd11an1n04x5 FILLER_58_528 ();
 b15zdnd11an1n04x5 FILLER_58_538 ();
 b15zdnd11an1n64x5 FILLER_58_546 ();
 b15zdnd11an1n64x5 FILLER_58_610 ();
 b15zdnd11an1n32x5 FILLER_58_674 ();
 b15zdnd11an1n08x5 FILLER_58_706 ();
 b15zdnd11an1n04x5 FILLER_58_714 ();
 b15zdnd11an1n64x5 FILLER_58_726 ();
 b15zdnd11an1n64x5 FILLER_58_790 ();
 b15zdnd11an1n64x5 FILLER_58_854 ();
 b15zdnd11an1n32x5 FILLER_58_918 ();
 b15zdnd11an1n08x5 FILLER_58_950 ();
 b15zdnd11an1n04x5 FILLER_58_958 ();
 b15zdnd11an1n32x5 FILLER_58_966 ();
 b15zdnd11an1n16x5 FILLER_58_998 ();
 b15zdnd11an1n04x5 FILLER_58_1014 ();
 b15zdnd00an1n02x5 FILLER_58_1018 ();
 b15zdnd00an1n01x5 FILLER_58_1020 ();
 b15zdnd11an1n64x5 FILLER_58_1029 ();
 b15zdnd11an1n64x5 FILLER_58_1093 ();
 b15zdnd11an1n64x5 FILLER_58_1157 ();
 b15zdnd11an1n32x5 FILLER_58_1221 ();
 b15zdnd11an1n04x5 FILLER_58_1253 ();
 b15zdnd00an1n01x5 FILLER_58_1257 ();
 b15zdnd11an1n32x5 FILLER_58_1275 ();
 b15zdnd11an1n08x5 FILLER_58_1307 ();
 b15zdnd00an1n01x5 FILLER_58_1315 ();
 b15zdnd11an1n64x5 FILLER_58_1327 ();
 b15zdnd11an1n64x5 FILLER_58_1391 ();
 b15zdnd11an1n32x5 FILLER_58_1455 ();
 b15zdnd11an1n16x5 FILLER_58_1487 ();
 b15zdnd11an1n08x5 FILLER_58_1503 ();
 b15zdnd11an1n16x5 FILLER_58_1528 ();
 b15zdnd11an1n08x5 FILLER_58_1544 ();
 b15zdnd00an1n02x5 FILLER_58_1552 ();
 b15zdnd00an1n01x5 FILLER_58_1554 ();
 b15zdnd11an1n64x5 FILLER_58_1586 ();
 b15zdnd11an1n64x5 FILLER_58_1650 ();
 b15zdnd11an1n64x5 FILLER_58_1714 ();
 b15zdnd11an1n08x5 FILLER_58_1778 ();
 b15zdnd00an1n02x5 FILLER_58_1786 ();
 b15zdnd00an1n01x5 FILLER_58_1788 ();
 b15zdnd11an1n04x5 FILLER_58_1793 ();
 b15zdnd00an1n02x5 FILLER_58_1797 ();
 b15zdnd00an1n01x5 FILLER_58_1799 ();
 b15zdnd11an1n64x5 FILLER_58_1806 ();
 b15zdnd11an1n64x5 FILLER_58_1870 ();
 b15zdnd11an1n64x5 FILLER_58_1934 ();
 b15zdnd11an1n64x5 FILLER_58_1998 ();
 b15zdnd11an1n64x5 FILLER_58_2062 ();
 b15zdnd11an1n16x5 FILLER_58_2126 ();
 b15zdnd11an1n08x5 FILLER_58_2142 ();
 b15zdnd11an1n04x5 FILLER_58_2150 ();
 b15zdnd11an1n64x5 FILLER_58_2162 ();
 b15zdnd11an1n32x5 FILLER_58_2226 ();
 b15zdnd11an1n16x5 FILLER_58_2258 ();
 b15zdnd00an1n02x5 FILLER_58_2274 ();
 b15zdnd11an1n64x5 FILLER_59_0 ();
 b15zdnd11an1n64x5 FILLER_59_64 ();
 b15zdnd11an1n64x5 FILLER_59_128 ();
 b15zdnd11an1n64x5 FILLER_59_192 ();
 b15zdnd11an1n64x5 FILLER_59_256 ();
 b15zdnd11an1n64x5 FILLER_59_320 ();
 b15zdnd11an1n64x5 FILLER_59_384 ();
 b15zdnd11an1n64x5 FILLER_59_448 ();
 b15zdnd11an1n16x5 FILLER_59_512 ();
 b15zdnd00an1n02x5 FILLER_59_528 ();
 b15zdnd11an1n64x5 FILLER_59_534 ();
 b15zdnd11an1n64x5 FILLER_59_598 ();
 b15zdnd11an1n64x5 FILLER_59_662 ();
 b15zdnd11an1n64x5 FILLER_59_726 ();
 b15zdnd11an1n64x5 FILLER_59_790 ();
 b15zdnd11an1n64x5 FILLER_59_854 ();
 b15zdnd11an1n32x5 FILLER_59_918 ();
 b15zdnd11an1n16x5 FILLER_59_950 ();
 b15zdnd11an1n04x5 FILLER_59_972 ();
 b15zdnd11an1n64x5 FILLER_59_980 ();
 b15zdnd11an1n64x5 FILLER_59_1044 ();
 b15zdnd11an1n32x5 FILLER_59_1108 ();
 b15zdnd00an1n02x5 FILLER_59_1140 ();
 b15zdnd11an1n64x5 FILLER_59_1145 ();
 b15zdnd11an1n64x5 FILLER_59_1209 ();
 b15zdnd11an1n64x5 FILLER_59_1273 ();
 b15zdnd11an1n64x5 FILLER_59_1337 ();
 b15zdnd11an1n64x5 FILLER_59_1401 ();
 b15zdnd11an1n64x5 FILLER_59_1465 ();
 b15zdnd11an1n16x5 FILLER_59_1529 ();
 b15zdnd11an1n04x5 FILLER_59_1545 ();
 b15zdnd00an1n01x5 FILLER_59_1549 ();
 b15zdnd11an1n08x5 FILLER_59_1592 ();
 b15zdnd11an1n04x5 FILLER_59_1600 ();
 b15zdnd11an1n64x5 FILLER_59_1646 ();
 b15zdnd11an1n64x5 FILLER_59_1710 ();
 b15zdnd11an1n16x5 FILLER_59_1774 ();
 b15zdnd00an1n02x5 FILLER_59_1790 ();
 b15zdnd00an1n01x5 FILLER_59_1792 ();
 b15zdnd11an1n04x5 FILLER_59_1797 ();
 b15zdnd11an1n64x5 FILLER_59_1805 ();
 b15zdnd11an1n64x5 FILLER_59_1869 ();
 b15zdnd11an1n16x5 FILLER_59_1933 ();
 b15zdnd11an1n08x5 FILLER_59_1949 ();
 b15zdnd00an1n02x5 FILLER_59_1957 ();
 b15zdnd00an1n01x5 FILLER_59_1959 ();
 b15zdnd11an1n16x5 FILLER_59_1969 ();
 b15zdnd00an1n02x5 FILLER_59_1985 ();
 b15zdnd00an1n01x5 FILLER_59_1987 ();
 b15zdnd11an1n64x5 FILLER_59_1997 ();
 b15zdnd11an1n64x5 FILLER_59_2061 ();
 b15zdnd11an1n64x5 FILLER_59_2125 ();
 b15zdnd11an1n64x5 FILLER_59_2189 ();
 b15zdnd11an1n16x5 FILLER_59_2253 ();
 b15zdnd11an1n08x5 FILLER_59_2269 ();
 b15zdnd11an1n04x5 FILLER_59_2277 ();
 b15zdnd00an1n02x5 FILLER_59_2281 ();
 b15zdnd00an1n01x5 FILLER_59_2283 ();
 b15zdnd11an1n64x5 FILLER_60_8 ();
 b15zdnd11an1n64x5 FILLER_60_72 ();
 b15zdnd11an1n64x5 FILLER_60_136 ();
 b15zdnd11an1n64x5 FILLER_60_200 ();
 b15zdnd11an1n64x5 FILLER_60_264 ();
 b15zdnd11an1n64x5 FILLER_60_328 ();
 b15zdnd11an1n64x5 FILLER_60_392 ();
 b15zdnd11an1n64x5 FILLER_60_456 ();
 b15zdnd11an1n64x5 FILLER_60_520 ();
 b15zdnd11an1n64x5 FILLER_60_584 ();
 b15zdnd11an1n32x5 FILLER_60_648 ();
 b15zdnd00an1n02x5 FILLER_60_680 ();
 b15zdnd00an1n01x5 FILLER_60_682 ();
 b15zdnd11an1n16x5 FILLER_60_687 ();
 b15zdnd11an1n08x5 FILLER_60_703 ();
 b15zdnd11an1n04x5 FILLER_60_711 ();
 b15zdnd00an1n02x5 FILLER_60_715 ();
 b15zdnd00an1n01x5 FILLER_60_717 ();
 b15zdnd11an1n64x5 FILLER_60_726 ();
 b15zdnd11an1n16x5 FILLER_60_790 ();
 b15zdnd11an1n08x5 FILLER_60_806 ();
 b15zdnd11an1n04x5 FILLER_60_814 ();
 b15zdnd00an1n02x5 FILLER_60_818 ();
 b15zdnd11an1n04x5 FILLER_60_824 ();
 b15zdnd11an1n08x5 FILLER_60_832 ();
 b15zdnd11an1n04x5 FILLER_60_840 ();
 b15zdnd00an1n01x5 FILLER_60_844 ();
 b15zdnd11an1n64x5 FILLER_60_849 ();
 b15zdnd11an1n32x5 FILLER_60_913 ();
 b15zdnd11an1n08x5 FILLER_60_945 ();
 b15zdnd11an1n04x5 FILLER_60_953 ();
 b15zdnd00an1n02x5 FILLER_60_957 ();
 b15zdnd11an1n16x5 FILLER_60_963 ();
 b15zdnd11an1n04x5 FILLER_60_979 ();
 b15zdnd00an1n02x5 FILLER_60_983 ();
 b15zdnd11an1n64x5 FILLER_60_989 ();
 b15zdnd11an1n64x5 FILLER_60_1053 ();
 b15zdnd11an1n08x5 FILLER_60_1117 ();
 b15zdnd00an1n01x5 FILLER_60_1125 ();
 b15zdnd11an1n64x5 FILLER_60_1138 ();
 b15zdnd11an1n64x5 FILLER_60_1202 ();
 b15zdnd11an1n64x5 FILLER_60_1266 ();
 b15zdnd11an1n64x5 FILLER_60_1330 ();
 b15zdnd11an1n32x5 FILLER_60_1394 ();
 b15zdnd11an1n16x5 FILLER_60_1426 ();
 b15zdnd11an1n08x5 FILLER_60_1442 ();
 b15zdnd11an1n04x5 FILLER_60_1450 ();
 b15zdnd00an1n02x5 FILLER_60_1454 ();
 b15zdnd11an1n08x5 FILLER_60_1470 ();
 b15zdnd00an1n02x5 FILLER_60_1478 ();
 b15zdnd00an1n01x5 FILLER_60_1480 ();
 b15zdnd11an1n64x5 FILLER_60_1495 ();
 b15zdnd11an1n64x5 FILLER_60_1559 ();
 b15zdnd11an1n64x5 FILLER_60_1623 ();
 b15zdnd11an1n64x5 FILLER_60_1687 ();
 b15zdnd11an1n32x5 FILLER_60_1751 ();
 b15zdnd11an1n16x5 FILLER_60_1783 ();
 b15zdnd00an1n02x5 FILLER_60_1799 ();
 b15zdnd11an1n64x5 FILLER_60_1805 ();
 b15zdnd11an1n32x5 FILLER_60_1869 ();
 b15zdnd11an1n16x5 FILLER_60_1901 ();
 b15zdnd11an1n04x5 FILLER_60_1917 ();
 b15zdnd00an1n01x5 FILLER_60_1921 ();
 b15zdnd11an1n64x5 FILLER_60_1925 ();
 b15zdnd11an1n64x5 FILLER_60_1989 ();
 b15zdnd11an1n64x5 FILLER_60_2053 ();
 b15zdnd11an1n32x5 FILLER_60_2117 ();
 b15zdnd11an1n04x5 FILLER_60_2149 ();
 b15zdnd00an1n01x5 FILLER_60_2153 ();
 b15zdnd11an1n64x5 FILLER_60_2162 ();
 b15zdnd11an1n32x5 FILLER_60_2226 ();
 b15zdnd11an1n16x5 FILLER_60_2258 ();
 b15zdnd00an1n02x5 FILLER_60_2274 ();
 b15zdnd11an1n64x5 FILLER_61_0 ();
 b15zdnd11an1n64x5 FILLER_61_64 ();
 b15zdnd11an1n32x5 FILLER_61_128 ();
 b15zdnd11an1n08x5 FILLER_61_160 ();
 b15zdnd11an1n04x5 FILLER_61_168 ();
 b15zdnd00an1n02x5 FILLER_61_172 ();
 b15zdnd11an1n64x5 FILLER_61_177 ();
 b15zdnd11an1n64x5 FILLER_61_241 ();
 b15zdnd11an1n64x5 FILLER_61_305 ();
 b15zdnd11an1n64x5 FILLER_61_369 ();
 b15zdnd11an1n64x5 FILLER_61_433 ();
 b15zdnd11an1n64x5 FILLER_61_497 ();
 b15zdnd11an1n64x5 FILLER_61_561 ();
 b15zdnd11an1n64x5 FILLER_61_625 ();
 b15zdnd11an1n64x5 FILLER_61_689 ();
 b15zdnd11an1n32x5 FILLER_61_753 ();
 b15zdnd11an1n16x5 FILLER_61_785 ();
 b15zdnd11an1n08x5 FILLER_61_801 ();
 b15zdnd11an1n04x5 FILLER_61_809 ();
 b15zdnd00an1n01x5 FILLER_61_813 ();
 b15zdnd11an1n64x5 FILLER_61_818 ();
 b15zdnd11an1n64x5 FILLER_61_882 ();
 b15zdnd11an1n64x5 FILLER_61_946 ();
 b15zdnd11an1n64x5 FILLER_61_1010 ();
 b15zdnd11an1n32x5 FILLER_61_1074 ();
 b15zdnd11an1n08x5 FILLER_61_1106 ();
 b15zdnd00an1n02x5 FILLER_61_1114 ();
 b15zdnd00an1n01x5 FILLER_61_1116 ();
 b15zdnd11an1n64x5 FILLER_61_1120 ();
 b15zdnd11an1n16x5 FILLER_61_1184 ();
 b15zdnd11an1n08x5 FILLER_61_1200 ();
 b15zdnd00an1n02x5 FILLER_61_1208 ();
 b15zdnd11an1n64x5 FILLER_61_1222 ();
 b15zdnd11an1n08x5 FILLER_61_1286 ();
 b15zdnd00an1n02x5 FILLER_61_1294 ();
 b15zdnd00an1n01x5 FILLER_61_1296 ();
 b15zdnd11an1n64x5 FILLER_61_1304 ();
 b15zdnd11an1n64x5 FILLER_61_1368 ();
 b15zdnd11an1n32x5 FILLER_61_1432 ();
 b15zdnd00an1n01x5 FILLER_61_1464 ();
 b15zdnd11an1n32x5 FILLER_61_1507 ();
 b15zdnd00an1n01x5 FILLER_61_1539 ();
 b15zdnd11an1n32x5 FILLER_61_1543 ();
 b15zdnd11an1n16x5 FILLER_61_1575 ();
 b15zdnd11an1n04x5 FILLER_61_1591 ();
 b15zdnd11an1n32x5 FILLER_61_1598 ();
 b15zdnd11an1n16x5 FILLER_61_1630 ();
 b15zdnd11an1n08x5 FILLER_61_1646 ();
 b15zdnd11an1n04x5 FILLER_61_1654 ();
 b15zdnd00an1n02x5 FILLER_61_1658 ();
 b15zdnd11an1n08x5 FILLER_61_1666 ();
 b15zdnd00an1n01x5 FILLER_61_1674 ();
 b15zdnd11an1n64x5 FILLER_61_1681 ();
 b15zdnd11an1n32x5 FILLER_61_1745 ();
 b15zdnd11an1n08x5 FILLER_61_1777 ();
 b15zdnd11an1n04x5 FILLER_61_1785 ();
 b15zdnd11an1n04x5 FILLER_61_1793 ();
 b15zdnd00an1n02x5 FILLER_61_1797 ();
 b15zdnd00an1n01x5 FILLER_61_1799 ();
 b15zdnd11an1n64x5 FILLER_61_1804 ();
 b15zdnd11an1n16x5 FILLER_61_1868 ();
 b15zdnd11an1n08x5 FILLER_61_1884 ();
 b15zdnd11an1n04x5 FILLER_61_1892 ();
 b15zdnd11an1n64x5 FILLER_61_1948 ();
 b15zdnd11an1n64x5 FILLER_61_2012 ();
 b15zdnd11an1n64x5 FILLER_61_2076 ();
 b15zdnd11an1n64x5 FILLER_61_2140 ();
 b15zdnd11an1n64x5 FILLER_61_2204 ();
 b15zdnd11an1n16x5 FILLER_61_2268 ();
 b15zdnd11an1n64x5 FILLER_62_8 ();
 b15zdnd11an1n64x5 FILLER_62_72 ();
 b15zdnd11an1n08x5 FILLER_62_136 ();
 b15zdnd00an1n02x5 FILLER_62_144 ();
 b15zdnd00an1n01x5 FILLER_62_146 ();
 b15zdnd11an1n64x5 FILLER_62_199 ();
 b15zdnd11an1n64x5 FILLER_62_263 ();
 b15zdnd11an1n64x5 FILLER_62_327 ();
 b15zdnd11an1n64x5 FILLER_62_391 ();
 b15zdnd11an1n64x5 FILLER_62_455 ();
 b15zdnd11an1n64x5 FILLER_62_519 ();
 b15zdnd11an1n64x5 FILLER_62_583 ();
 b15zdnd11an1n64x5 FILLER_62_647 ();
 b15zdnd11an1n04x5 FILLER_62_711 ();
 b15zdnd00an1n02x5 FILLER_62_715 ();
 b15zdnd00an1n01x5 FILLER_62_717 ();
 b15zdnd11an1n64x5 FILLER_62_726 ();
 b15zdnd11an1n32x5 FILLER_62_790 ();
 b15zdnd00an1n02x5 FILLER_62_822 ();
 b15zdnd00an1n01x5 FILLER_62_824 ();
 b15zdnd11an1n04x5 FILLER_62_829 ();
 b15zdnd00an1n02x5 FILLER_62_833 ();
 b15zdnd11an1n64x5 FILLER_62_839 ();
 b15zdnd11an1n64x5 FILLER_62_903 ();
 b15zdnd11an1n64x5 FILLER_62_967 ();
 b15zdnd11an1n64x5 FILLER_62_1031 ();
 b15zdnd11an1n08x5 FILLER_62_1095 ();
 b15zdnd11an1n04x5 FILLER_62_1103 ();
 b15zdnd00an1n02x5 FILLER_62_1107 ();
 b15zdnd11an1n64x5 FILLER_62_1123 ();
 b15zdnd11an1n16x5 FILLER_62_1193 ();
 b15zdnd11an1n08x5 FILLER_62_1209 ();
 b15zdnd11an1n04x5 FILLER_62_1217 ();
 b15zdnd11an1n64x5 FILLER_62_1229 ();
 b15zdnd11an1n64x5 FILLER_62_1293 ();
 b15zdnd11an1n64x5 FILLER_62_1357 ();
 b15zdnd11an1n64x5 FILLER_62_1442 ();
 b15zdnd11an1n08x5 FILLER_62_1506 ();
 b15zdnd11an1n04x5 FILLER_62_1514 ();
 b15zdnd11an1n04x5 FILLER_62_1525 ();
 b15zdnd11an1n32x5 FILLER_62_1543 ();
 b15zdnd11an1n16x5 FILLER_62_1575 ();
 b15zdnd11an1n04x5 FILLER_62_1591 ();
 b15zdnd11an1n16x5 FILLER_62_1609 ();
 b15zdnd11an1n04x5 FILLER_62_1625 ();
 b15zdnd00an1n02x5 FILLER_62_1629 ();
 b15zdnd11an1n08x5 FILLER_62_1662 ();
 b15zdnd11an1n04x5 FILLER_62_1670 ();
 b15zdnd00an1n02x5 FILLER_62_1674 ();
 b15zdnd11an1n04x5 FILLER_62_1683 ();
 b15zdnd11an1n64x5 FILLER_62_1694 ();
 b15zdnd11an1n64x5 FILLER_62_1758 ();
 b15zdnd11an1n64x5 FILLER_62_1822 ();
 b15zdnd11an1n16x5 FILLER_62_1886 ();
 b15zdnd11an1n08x5 FILLER_62_1902 ();
 b15zdnd11an1n04x5 FILLER_62_1910 ();
 b15zdnd11an1n04x5 FILLER_62_1917 ();
 b15zdnd11an1n64x5 FILLER_62_1924 ();
 b15zdnd11an1n08x5 FILLER_62_1988 ();
 b15zdnd11an1n04x5 FILLER_62_1996 ();
 b15zdnd11an1n64x5 FILLER_62_2009 ();
 b15zdnd11an1n64x5 FILLER_62_2073 ();
 b15zdnd11an1n16x5 FILLER_62_2137 ();
 b15zdnd00an1n01x5 FILLER_62_2153 ();
 b15zdnd11an1n64x5 FILLER_62_2162 ();
 b15zdnd11an1n32x5 FILLER_62_2226 ();
 b15zdnd11an1n16x5 FILLER_62_2258 ();
 b15zdnd00an1n02x5 FILLER_62_2274 ();
 b15zdnd11an1n64x5 FILLER_63_0 ();
 b15zdnd11an1n64x5 FILLER_63_64 ();
 b15zdnd11an1n32x5 FILLER_63_128 ();
 b15zdnd11an1n04x5 FILLER_63_160 ();
 b15zdnd00an1n01x5 FILLER_63_164 ();
 b15zdnd11an1n04x5 FILLER_63_168 ();
 b15zdnd11an1n16x5 FILLER_63_175 ();
 b15zdnd11an1n04x5 FILLER_63_191 ();
 b15zdnd00an1n02x5 FILLER_63_195 ();
 b15zdnd11an1n64x5 FILLER_63_239 ();
 b15zdnd11an1n64x5 FILLER_63_303 ();
 b15zdnd11an1n64x5 FILLER_63_367 ();
 b15zdnd11an1n64x5 FILLER_63_431 ();
 b15zdnd11an1n64x5 FILLER_63_495 ();
 b15zdnd11an1n32x5 FILLER_63_559 ();
 b15zdnd11an1n16x5 FILLER_63_591 ();
 b15zdnd11an1n08x5 FILLER_63_607 ();
 b15zdnd00an1n02x5 FILLER_63_615 ();
 b15zdnd00an1n01x5 FILLER_63_617 ();
 b15zdnd11an1n64x5 FILLER_63_622 ();
 b15zdnd11an1n64x5 FILLER_63_686 ();
 b15zdnd11an1n64x5 FILLER_63_750 ();
 b15zdnd11an1n64x5 FILLER_63_814 ();
 b15zdnd11an1n64x5 FILLER_63_878 ();
 b15zdnd11an1n64x5 FILLER_63_942 ();
 b15zdnd11an1n64x5 FILLER_63_1006 ();
 b15zdnd11an1n64x5 FILLER_63_1070 ();
 b15zdnd00an1n02x5 FILLER_63_1134 ();
 b15zdnd00an1n01x5 FILLER_63_1136 ();
 b15zdnd11an1n64x5 FILLER_63_1142 ();
 b15zdnd11an1n16x5 FILLER_63_1206 ();
 b15zdnd00an1n02x5 FILLER_63_1222 ();
 b15zdnd11an1n32x5 FILLER_63_1238 ();
 b15zdnd11an1n16x5 FILLER_63_1270 ();
 b15zdnd11an1n08x5 FILLER_63_1286 ();
 b15zdnd00an1n02x5 FILLER_63_1294 ();
 b15zdnd00an1n01x5 FILLER_63_1296 ();
 b15zdnd11an1n64x5 FILLER_63_1303 ();
 b15zdnd11an1n08x5 FILLER_63_1367 ();
 b15zdnd11an1n04x5 FILLER_63_1375 ();
 b15zdnd00an1n02x5 FILLER_63_1379 ();
 b15zdnd00an1n01x5 FILLER_63_1381 ();
 b15zdnd11an1n32x5 FILLER_63_1392 ();
 b15zdnd11an1n08x5 FILLER_63_1424 ();
 b15zdnd00an1n01x5 FILLER_63_1432 ();
 b15zdnd11an1n32x5 FILLER_63_1440 ();
 b15zdnd11an1n08x5 FILLER_63_1472 ();
 b15zdnd00an1n02x5 FILLER_63_1480 ();
 b15zdnd11an1n64x5 FILLER_63_1502 ();
 b15zdnd11an1n64x5 FILLER_63_1566 ();
 b15zdnd11an1n32x5 FILLER_63_1630 ();
 b15zdnd11an1n08x5 FILLER_63_1662 ();
 b15zdnd11an1n04x5 FILLER_63_1670 ();
 b15zdnd00an1n01x5 FILLER_63_1674 ();
 b15zdnd11an1n64x5 FILLER_63_1679 ();
 b15zdnd11an1n64x5 FILLER_63_1743 ();
 b15zdnd11an1n64x5 FILLER_63_1807 ();
 b15zdnd11an1n64x5 FILLER_63_1871 ();
 b15zdnd11an1n64x5 FILLER_63_1935 ();
 b15zdnd11an1n32x5 FILLER_63_1999 ();
 b15zdnd11an1n16x5 FILLER_63_2031 ();
 b15zdnd11an1n04x5 FILLER_63_2047 ();
 b15zdnd00an1n01x5 FILLER_63_2051 ();
 b15zdnd11an1n64x5 FILLER_63_2055 ();
 b15zdnd11an1n64x5 FILLER_63_2119 ();
 b15zdnd11an1n32x5 FILLER_63_2183 ();
 b15zdnd11an1n16x5 FILLER_63_2215 ();
 b15zdnd11an1n08x5 FILLER_63_2231 ();
 b15zdnd00an1n02x5 FILLER_63_2239 ();
 b15zdnd11an1n04x5 FILLER_63_2244 ();
 b15zdnd11an1n08x5 FILLER_63_2251 ();
 b15zdnd00an1n01x5 FILLER_63_2259 ();
 b15zdnd11an1n16x5 FILLER_63_2263 ();
 b15zdnd11an1n04x5 FILLER_63_2279 ();
 b15zdnd00an1n01x5 FILLER_63_2283 ();
 b15zdnd11an1n64x5 FILLER_64_8 ();
 b15zdnd11an1n64x5 FILLER_64_72 ();
 b15zdnd11an1n16x5 FILLER_64_136 ();
 b15zdnd11an1n04x5 FILLER_64_152 ();
 b15zdnd00an1n02x5 FILLER_64_156 ();
 b15zdnd00an1n01x5 FILLER_64_158 ();
 b15zdnd11an1n64x5 FILLER_64_201 ();
 b15zdnd11an1n64x5 FILLER_64_265 ();
 b15zdnd11an1n64x5 FILLER_64_329 ();
 b15zdnd11an1n64x5 FILLER_64_393 ();
 b15zdnd11an1n64x5 FILLER_64_457 ();
 b15zdnd11an1n32x5 FILLER_64_521 ();
 b15zdnd11an1n08x5 FILLER_64_553 ();
 b15zdnd11an1n04x5 FILLER_64_561 ();
 b15zdnd00an1n02x5 FILLER_64_565 ();
 b15zdnd11an1n64x5 FILLER_64_571 ();
 b15zdnd11an1n32x5 FILLER_64_635 ();
 b15zdnd00an1n02x5 FILLER_64_667 ();
 b15zdnd00an1n01x5 FILLER_64_669 ();
 b15zdnd11an1n32x5 FILLER_64_674 ();
 b15zdnd11an1n08x5 FILLER_64_706 ();
 b15zdnd11an1n04x5 FILLER_64_714 ();
 b15zdnd11an1n64x5 FILLER_64_726 ();
 b15zdnd11an1n32x5 FILLER_64_790 ();
 b15zdnd00an1n01x5 FILLER_64_822 ();
 b15zdnd11an1n64x5 FILLER_64_830 ();
 b15zdnd11an1n64x5 FILLER_64_894 ();
 b15zdnd11an1n64x5 FILLER_64_958 ();
 b15zdnd11an1n64x5 FILLER_64_1022 ();
 b15zdnd11an1n08x5 FILLER_64_1086 ();
 b15zdnd00an1n01x5 FILLER_64_1094 ();
 b15zdnd11an1n64x5 FILLER_64_1109 ();
 b15zdnd11an1n08x5 FILLER_64_1173 ();
 b15zdnd00an1n01x5 FILLER_64_1181 ();
 b15zdnd11an1n64x5 FILLER_64_1189 ();
 b15zdnd11an1n08x5 FILLER_64_1253 ();
 b15zdnd11an1n04x5 FILLER_64_1261 ();
 b15zdnd00an1n02x5 FILLER_64_1265 ();
 b15zdnd11an1n64x5 FILLER_64_1284 ();
 b15zdnd11an1n08x5 FILLER_64_1354 ();
 b15zdnd11an1n04x5 FILLER_64_1362 ();
 b15zdnd00an1n01x5 FILLER_64_1366 ();
 b15zdnd11an1n16x5 FILLER_64_1374 ();
 b15zdnd00an1n02x5 FILLER_64_1390 ();
 b15zdnd11an1n16x5 FILLER_64_1416 ();
 b15zdnd11an1n08x5 FILLER_64_1432 ();
 b15zdnd00an1n02x5 FILLER_64_1440 ();
 b15zdnd11an1n64x5 FILLER_64_1462 ();
 b15zdnd11an1n64x5 FILLER_64_1526 ();
 b15zdnd11an1n64x5 FILLER_64_1590 ();
 b15zdnd11an1n64x5 FILLER_64_1654 ();
 b15zdnd00an1n01x5 FILLER_64_1718 ();
 b15zdnd11an1n64x5 FILLER_64_1725 ();
 b15zdnd11an1n64x5 FILLER_64_1789 ();
 b15zdnd11an1n64x5 FILLER_64_1853 ();
 b15zdnd11an1n64x5 FILLER_64_1917 ();
 b15zdnd11an1n64x5 FILLER_64_1981 ();
 b15zdnd11an1n04x5 FILLER_64_2045 ();
 b15zdnd00an1n02x5 FILLER_64_2049 ();
 b15zdnd11an1n04x5 FILLER_64_2054 ();
 b15zdnd11an1n64x5 FILLER_64_2061 ();
 b15zdnd11an1n16x5 FILLER_64_2125 ();
 b15zdnd11an1n08x5 FILLER_64_2141 ();
 b15zdnd11an1n04x5 FILLER_64_2149 ();
 b15zdnd00an1n01x5 FILLER_64_2153 ();
 b15zdnd11an1n64x5 FILLER_64_2162 ();
 b15zdnd11an1n16x5 FILLER_64_2226 ();
 b15zdnd11an1n08x5 FILLER_64_2242 ();
 b15zdnd00an1n02x5 FILLER_64_2250 ();
 b15zdnd11an1n16x5 FILLER_64_2255 ();
 b15zdnd11an1n04x5 FILLER_64_2271 ();
 b15zdnd00an1n01x5 FILLER_64_2275 ();
 b15zdnd11an1n64x5 FILLER_65_0 ();
 b15zdnd11an1n64x5 FILLER_65_64 ();
 b15zdnd11an1n32x5 FILLER_65_128 ();
 b15zdnd11an1n04x5 FILLER_65_160 ();
 b15zdnd00an1n02x5 FILLER_65_164 ();
 b15zdnd00an1n01x5 FILLER_65_166 ();
 b15zdnd11an1n16x5 FILLER_65_172 ();
 b15zdnd11an1n04x5 FILLER_65_188 ();
 b15zdnd00an1n01x5 FILLER_65_192 ();
 b15zdnd11an1n64x5 FILLER_65_224 ();
 b15zdnd11an1n64x5 FILLER_65_288 ();
 b15zdnd11an1n64x5 FILLER_65_352 ();
 b15zdnd11an1n64x5 FILLER_65_416 ();
 b15zdnd11an1n64x5 FILLER_65_480 ();
 b15zdnd11an1n32x5 FILLER_65_544 ();
 b15zdnd00an1n01x5 FILLER_65_576 ();
 b15zdnd11an1n64x5 FILLER_65_581 ();
 b15zdnd11an1n16x5 FILLER_65_645 ();
 b15zdnd11an1n08x5 FILLER_65_661 ();
 b15zdnd00an1n01x5 FILLER_65_669 ();
 b15zdnd11an1n64x5 FILLER_65_674 ();
 b15zdnd11an1n32x5 FILLER_65_738 ();
 b15zdnd11an1n16x5 FILLER_65_770 ();
 b15zdnd11an1n04x5 FILLER_65_786 ();
 b15zdnd00an1n02x5 FILLER_65_790 ();
 b15zdnd00an1n01x5 FILLER_65_792 ();
 b15zdnd11an1n64x5 FILLER_65_807 ();
 b15zdnd11an1n64x5 FILLER_65_871 ();
 b15zdnd11an1n32x5 FILLER_65_935 ();
 b15zdnd11an1n08x5 FILLER_65_967 ();
 b15zdnd11an1n64x5 FILLER_65_999 ();
 b15zdnd11an1n64x5 FILLER_65_1063 ();
 b15zdnd11an1n64x5 FILLER_65_1127 ();
 b15zdnd11an1n64x5 FILLER_65_1191 ();
 b15zdnd11an1n64x5 FILLER_65_1255 ();
 b15zdnd11an1n08x5 FILLER_65_1319 ();
 b15zdnd11an1n04x5 FILLER_65_1327 ();
 b15zdnd00an1n02x5 FILLER_65_1331 ();
 b15zdnd11an1n64x5 FILLER_65_1354 ();
 b15zdnd11an1n64x5 FILLER_65_1418 ();
 b15zdnd11an1n64x5 FILLER_65_1482 ();
 b15zdnd11an1n64x5 FILLER_65_1546 ();
 b15zdnd11an1n64x5 FILLER_65_1610 ();
 b15zdnd11an1n64x5 FILLER_65_1674 ();
 b15zdnd11an1n32x5 FILLER_65_1738 ();
 b15zdnd00an1n01x5 FILLER_65_1770 ();
 b15zdnd11an1n64x5 FILLER_65_1775 ();
 b15zdnd11an1n64x5 FILLER_65_1839 ();
 b15zdnd11an1n64x5 FILLER_65_1903 ();
 b15zdnd11an1n64x5 FILLER_65_1967 ();
 b15zdnd00an1n01x5 FILLER_65_2031 ();
 b15zdnd11an1n64x5 FILLER_65_2084 ();
 b15zdnd11an1n64x5 FILLER_65_2148 ();
 b15zdnd11an1n64x5 FILLER_65_2212 ();
 b15zdnd11an1n08x5 FILLER_65_2276 ();
 b15zdnd11an1n64x5 FILLER_66_8 ();
 b15zdnd11an1n64x5 FILLER_66_72 ();
 b15zdnd11an1n64x5 FILLER_66_136 ();
 b15zdnd11an1n32x5 FILLER_66_200 ();
 b15zdnd11an1n16x5 FILLER_66_232 ();
 b15zdnd11an1n08x5 FILLER_66_248 ();
 b15zdnd11an1n04x5 FILLER_66_296 ();
 b15zdnd11an1n64x5 FILLER_66_303 ();
 b15zdnd11an1n64x5 FILLER_66_367 ();
 b15zdnd11an1n64x5 FILLER_66_431 ();
 b15zdnd11an1n64x5 FILLER_66_495 ();
 b15zdnd11an1n64x5 FILLER_66_559 ();
 b15zdnd11an1n64x5 FILLER_66_623 ();
 b15zdnd11an1n16x5 FILLER_66_687 ();
 b15zdnd11an1n08x5 FILLER_66_703 ();
 b15zdnd11an1n04x5 FILLER_66_711 ();
 b15zdnd00an1n02x5 FILLER_66_715 ();
 b15zdnd00an1n01x5 FILLER_66_717 ();
 b15zdnd11an1n16x5 FILLER_66_726 ();
 b15zdnd00an1n01x5 FILLER_66_742 ();
 b15zdnd11an1n32x5 FILLER_66_751 ();
 b15zdnd11an1n04x5 FILLER_66_783 ();
 b15zdnd11an1n04x5 FILLER_66_801 ();
 b15zdnd00an1n01x5 FILLER_66_805 ();
 b15zdnd11an1n64x5 FILLER_66_809 ();
 b15zdnd11an1n64x5 FILLER_66_873 ();
 b15zdnd11an1n32x5 FILLER_66_937 ();
 b15zdnd11an1n16x5 FILLER_66_969 ();
 b15zdnd11an1n08x5 FILLER_66_985 ();
 b15zdnd11an1n04x5 FILLER_66_993 ();
 b15zdnd00an1n02x5 FILLER_66_997 ();
 b15zdnd00an1n01x5 FILLER_66_999 ();
 b15zdnd11an1n64x5 FILLER_66_1008 ();
 b15zdnd11an1n64x5 FILLER_66_1072 ();
 b15zdnd11an1n08x5 FILLER_66_1136 ();
 b15zdnd11an1n04x5 FILLER_66_1144 ();
 b15zdnd11an1n64x5 FILLER_66_1162 ();
 b15zdnd11an1n64x5 FILLER_66_1226 ();
 b15zdnd11an1n64x5 FILLER_66_1290 ();
 b15zdnd11an1n16x5 FILLER_66_1354 ();
 b15zdnd11an1n08x5 FILLER_66_1370 ();
 b15zdnd11an1n64x5 FILLER_66_1409 ();
 b15zdnd11an1n32x5 FILLER_66_1473 ();
 b15zdnd11an1n16x5 FILLER_66_1505 ();
 b15zdnd11an1n08x5 FILLER_66_1521 ();
 b15zdnd00an1n02x5 FILLER_66_1529 ();
 b15zdnd00an1n01x5 FILLER_66_1531 ();
 b15zdnd11an1n32x5 FILLER_66_1535 ();
 b15zdnd11an1n08x5 FILLER_66_1567 ();
 b15zdnd11an1n04x5 FILLER_66_1575 ();
 b15zdnd00an1n02x5 FILLER_66_1579 ();
 b15zdnd00an1n01x5 FILLER_66_1581 ();
 b15zdnd11an1n64x5 FILLER_66_1585 ();
 b15zdnd11an1n64x5 FILLER_66_1649 ();
 b15zdnd11an1n16x5 FILLER_66_1713 ();
 b15zdnd11an1n08x5 FILLER_66_1729 ();
 b15zdnd11an1n04x5 FILLER_66_1737 ();
 b15zdnd00an1n02x5 FILLER_66_1741 ();
 b15zdnd11an1n16x5 FILLER_66_1747 ();
 b15zdnd11an1n08x5 FILLER_66_1763 ();
 b15zdnd00an1n02x5 FILLER_66_1771 ();
 b15zdnd11an1n64x5 FILLER_66_1779 ();
 b15zdnd11an1n64x5 FILLER_66_1843 ();
 b15zdnd11an1n08x5 FILLER_66_1907 ();
 b15zdnd11an1n04x5 FILLER_66_1915 ();
 b15zdnd11an1n64x5 FILLER_66_1922 ();
 b15zdnd11an1n32x5 FILLER_66_1986 ();
 b15zdnd11an1n08x5 FILLER_66_2018 ();
 b15zdnd11an1n04x5 FILLER_66_2026 ();
 b15zdnd11an1n16x5 FILLER_66_2082 ();
 b15zdnd11an1n04x5 FILLER_66_2098 ();
 b15zdnd11an1n32x5 FILLER_66_2106 ();
 b15zdnd11an1n16x5 FILLER_66_2138 ();
 b15zdnd11an1n64x5 FILLER_66_2162 ();
 b15zdnd11an1n32x5 FILLER_66_2226 ();
 b15zdnd11an1n16x5 FILLER_66_2258 ();
 b15zdnd00an1n02x5 FILLER_66_2274 ();
 b15zdnd11an1n64x5 FILLER_67_0 ();
 b15zdnd11an1n64x5 FILLER_67_64 ();
 b15zdnd11an1n64x5 FILLER_67_128 ();
 b15zdnd11an1n64x5 FILLER_67_192 ();
 b15zdnd11an1n08x5 FILLER_67_256 ();
 b15zdnd11an1n04x5 FILLER_67_264 ();
 b15zdnd11an1n16x5 FILLER_67_272 ();
 b15zdnd11an1n04x5 FILLER_67_288 ();
 b15zdnd11an1n64x5 FILLER_67_295 ();
 b15zdnd11an1n64x5 FILLER_67_359 ();
 b15zdnd11an1n64x5 FILLER_67_423 ();
 b15zdnd11an1n64x5 FILLER_67_487 ();
 b15zdnd11an1n64x5 FILLER_67_551 ();
 b15zdnd11an1n64x5 FILLER_67_615 ();
 b15zdnd11an1n64x5 FILLER_67_679 ();
 b15zdnd11an1n64x5 FILLER_67_743 ();
 b15zdnd11an1n64x5 FILLER_67_807 ();
 b15zdnd11an1n64x5 FILLER_67_871 ();
 b15zdnd11an1n16x5 FILLER_67_935 ();
 b15zdnd00an1n01x5 FILLER_67_951 ();
 b15zdnd11an1n64x5 FILLER_67_955 ();
 b15zdnd11an1n32x5 FILLER_67_1019 ();
 b15zdnd11an1n16x5 FILLER_67_1051 ();
 b15zdnd11an1n08x5 FILLER_67_1067 ();
 b15zdnd11an1n64x5 FILLER_67_1082 ();
 b15zdnd11an1n64x5 FILLER_67_1146 ();
 b15zdnd11an1n64x5 FILLER_67_1210 ();
 b15zdnd11an1n64x5 FILLER_67_1274 ();
 b15zdnd11an1n64x5 FILLER_67_1338 ();
 b15zdnd11an1n64x5 FILLER_67_1402 ();
 b15zdnd11an1n64x5 FILLER_67_1466 ();
 b15zdnd11an1n64x5 FILLER_67_1530 ();
 b15zdnd11an1n64x5 FILLER_67_1594 ();
 b15zdnd11an1n64x5 FILLER_67_1658 ();
 b15zdnd11an1n32x5 FILLER_67_1722 ();
 b15zdnd11an1n16x5 FILLER_67_1754 ();
 b15zdnd11an1n04x5 FILLER_67_1770 ();
 b15zdnd11an1n64x5 FILLER_67_1778 ();
 b15zdnd11an1n64x5 FILLER_67_1842 ();
 b15zdnd11an1n08x5 FILLER_67_1906 ();
 b15zdnd11an1n04x5 FILLER_67_1914 ();
 b15zdnd11an1n04x5 FILLER_67_1921 ();
 b15zdnd11an1n64x5 FILLER_67_1928 ();
 b15zdnd11an1n32x5 FILLER_67_1992 ();
 b15zdnd11an1n08x5 FILLER_67_2024 ();
 b15zdnd11an1n04x5 FILLER_67_2032 ();
 b15zdnd00an1n02x5 FILLER_67_2036 ();
 b15zdnd00an1n01x5 FILLER_67_2038 ();
 b15zdnd11an1n04x5 FILLER_67_2091 ();
 b15zdnd11an1n64x5 FILLER_67_2099 ();
 b15zdnd11an1n64x5 FILLER_67_2163 ();
 b15zdnd11an1n32x5 FILLER_67_2227 ();
 b15zdnd11an1n16x5 FILLER_67_2259 ();
 b15zdnd11an1n08x5 FILLER_67_2275 ();
 b15zdnd00an1n01x5 FILLER_67_2283 ();
 b15zdnd11an1n64x5 FILLER_68_8 ();
 b15zdnd11an1n64x5 FILLER_68_72 ();
 b15zdnd11an1n64x5 FILLER_68_136 ();
 b15zdnd11an1n64x5 FILLER_68_200 ();
 b15zdnd11an1n64x5 FILLER_68_264 ();
 b15zdnd11an1n08x5 FILLER_68_328 ();
 b15zdnd11an1n04x5 FILLER_68_336 ();
 b15zdnd00an1n01x5 FILLER_68_340 ();
 b15zdnd11an1n64x5 FILLER_68_383 ();
 b15zdnd11an1n32x5 FILLER_68_447 ();
 b15zdnd11an1n04x5 FILLER_68_483 ();
 b15zdnd11an1n64x5 FILLER_68_491 ();
 b15zdnd11an1n64x5 FILLER_68_555 ();
 b15zdnd11an1n64x5 FILLER_68_619 ();
 b15zdnd11an1n32x5 FILLER_68_683 ();
 b15zdnd00an1n02x5 FILLER_68_715 ();
 b15zdnd00an1n01x5 FILLER_68_717 ();
 b15zdnd11an1n64x5 FILLER_68_726 ();
 b15zdnd11an1n64x5 FILLER_68_790 ();
 b15zdnd11an1n32x5 FILLER_68_854 ();
 b15zdnd11an1n16x5 FILLER_68_886 ();
 b15zdnd11an1n08x5 FILLER_68_902 ();
 b15zdnd11an1n04x5 FILLER_68_910 ();
 b15zdnd00an1n02x5 FILLER_68_914 ();
 b15zdnd00an1n01x5 FILLER_68_916 ();
 b15zdnd11an1n04x5 FILLER_68_924 ();
 b15zdnd11an1n04x5 FILLER_68_972 ();
 b15zdnd00an1n02x5 FILLER_68_976 ();
 b15zdnd11an1n64x5 FILLER_68_992 ();
 b15zdnd11an1n64x5 FILLER_68_1056 ();
 b15zdnd11an1n08x5 FILLER_68_1120 ();
 b15zdnd11an1n64x5 FILLER_68_1131 ();
 b15zdnd11an1n64x5 FILLER_68_1195 ();
 b15zdnd11an1n32x5 FILLER_68_1259 ();
 b15zdnd11an1n08x5 FILLER_68_1291 ();
 b15zdnd11an1n04x5 FILLER_68_1299 ();
 b15zdnd00an1n02x5 FILLER_68_1303 ();
 b15zdnd11an1n32x5 FILLER_68_1313 ();
 b15zdnd11an1n08x5 FILLER_68_1345 ();
 b15zdnd00an1n02x5 FILLER_68_1353 ();
 b15zdnd00an1n01x5 FILLER_68_1355 ();
 b15zdnd11an1n04x5 FILLER_68_1370 ();
 b15zdnd11an1n32x5 FILLER_68_1390 ();
 b15zdnd11an1n04x5 FILLER_68_1422 ();
 b15zdnd00an1n01x5 FILLER_68_1426 ();
 b15zdnd11an1n32x5 FILLER_68_1435 ();
 b15zdnd11an1n16x5 FILLER_68_1467 ();
 b15zdnd11an1n08x5 FILLER_68_1483 ();
 b15zdnd11an1n04x5 FILLER_68_1491 ();
 b15zdnd00an1n02x5 FILLER_68_1495 ();
 b15zdnd11an1n64x5 FILLER_68_1510 ();
 b15zdnd11an1n64x5 FILLER_68_1574 ();
 b15zdnd11an1n64x5 FILLER_68_1638 ();
 b15zdnd11an1n64x5 FILLER_68_1702 ();
 b15zdnd11an1n64x5 FILLER_68_1766 ();
 b15zdnd11an1n64x5 FILLER_68_1830 ();
 b15zdnd11an1n04x5 FILLER_68_1894 ();
 b15zdnd00an1n01x5 FILLER_68_1898 ();
 b15zdnd11an1n64x5 FILLER_68_1951 ();
 b15zdnd11an1n32x5 FILLER_68_2015 ();
 b15zdnd00an1n01x5 FILLER_68_2047 ();
 b15zdnd11an1n04x5 FILLER_68_2051 ();
 b15zdnd11an1n04x5 FILLER_68_2058 ();
 b15zdnd11an1n04x5 FILLER_68_2065 ();
 b15zdnd11an1n08x5 FILLER_68_2072 ();
 b15zdnd11an1n04x5 FILLER_68_2080 ();
 b15zdnd00an1n01x5 FILLER_68_2084 ();
 b15zdnd11an1n08x5 FILLER_68_2093 ();
 b15zdnd11an1n32x5 FILLER_68_2105 ();
 b15zdnd11an1n16x5 FILLER_68_2137 ();
 b15zdnd00an1n01x5 FILLER_68_2153 ();
 b15zdnd11an1n64x5 FILLER_68_2162 ();
 b15zdnd11an1n32x5 FILLER_68_2226 ();
 b15zdnd11an1n16x5 FILLER_68_2258 ();
 b15zdnd00an1n02x5 FILLER_68_2274 ();
 b15zdnd11an1n64x5 FILLER_69_0 ();
 b15zdnd11an1n64x5 FILLER_69_64 ();
 b15zdnd11an1n64x5 FILLER_69_128 ();
 b15zdnd11an1n64x5 FILLER_69_192 ();
 b15zdnd11an1n64x5 FILLER_69_256 ();
 b15zdnd11an1n64x5 FILLER_69_320 ();
 b15zdnd11an1n64x5 FILLER_69_384 ();
 b15zdnd11an1n64x5 FILLER_69_448 ();
 b15zdnd11an1n64x5 FILLER_69_512 ();
 b15zdnd11an1n64x5 FILLER_69_579 ();
 b15zdnd11an1n64x5 FILLER_69_643 ();
 b15zdnd11an1n64x5 FILLER_69_707 ();
 b15zdnd11an1n16x5 FILLER_69_771 ();
 b15zdnd00an1n02x5 FILLER_69_787 ();
 b15zdnd11an1n64x5 FILLER_69_792 ();
 b15zdnd11an1n64x5 FILLER_69_856 ();
 b15zdnd11an1n16x5 FILLER_69_920 ();
 b15zdnd11an1n08x5 FILLER_69_936 ();
 b15zdnd11an1n04x5 FILLER_69_947 ();
 b15zdnd11an1n16x5 FILLER_69_954 ();
 b15zdnd11an1n04x5 FILLER_69_970 ();
 b15zdnd00an1n01x5 FILLER_69_974 ();
 b15zdnd11an1n64x5 FILLER_69_1017 ();
 b15zdnd11an1n64x5 FILLER_69_1081 ();
 b15zdnd11an1n32x5 FILLER_69_1145 ();
 b15zdnd11an1n16x5 FILLER_69_1177 ();
 b15zdnd11an1n08x5 FILLER_69_1193 ();
 b15zdnd00an1n02x5 FILLER_69_1201 ();
 b15zdnd00an1n01x5 FILLER_69_1203 ();
 b15zdnd11an1n64x5 FILLER_69_1211 ();
 b15zdnd11an1n16x5 FILLER_69_1275 ();
 b15zdnd00an1n02x5 FILLER_69_1291 ();
 b15zdnd00an1n01x5 FILLER_69_1293 ();
 b15zdnd11an1n16x5 FILLER_69_1306 ();
 b15zdnd11an1n08x5 FILLER_69_1322 ();
 b15zdnd00an1n01x5 FILLER_69_1330 ();
 b15zdnd11an1n64x5 FILLER_69_1338 ();
 b15zdnd11an1n64x5 FILLER_69_1402 ();
 b15zdnd11an1n64x5 FILLER_69_1466 ();
 b15zdnd11an1n64x5 FILLER_69_1530 ();
 b15zdnd11an1n64x5 FILLER_69_1594 ();
 b15zdnd11an1n64x5 FILLER_69_1658 ();
 b15zdnd11an1n64x5 FILLER_69_1722 ();
 b15zdnd11an1n64x5 FILLER_69_1786 ();
 b15zdnd11an1n32x5 FILLER_69_1850 ();
 b15zdnd11an1n16x5 FILLER_69_1882 ();
 b15zdnd00an1n02x5 FILLER_69_1898 ();
 b15zdnd00an1n01x5 FILLER_69_1900 ();
 b15zdnd11an1n64x5 FILLER_69_1953 ();
 b15zdnd11an1n32x5 FILLER_69_2017 ();
 b15zdnd00an1n01x5 FILLER_69_2049 ();
 b15zdnd11an1n04x5 FILLER_69_2053 ();
 b15zdnd11an1n16x5 FILLER_69_2060 ();
 b15zdnd11an1n08x5 FILLER_69_2076 ();
 b15zdnd11an1n04x5 FILLER_69_2084 ();
 b15zdnd00an1n01x5 FILLER_69_2088 ();
 b15zdnd11an1n04x5 FILLER_69_2093 ();
 b15zdnd00an1n02x5 FILLER_69_2097 ();
 b15zdnd11an1n64x5 FILLER_69_2103 ();
 b15zdnd11an1n64x5 FILLER_69_2167 ();
 b15zdnd11an1n32x5 FILLER_69_2231 ();
 b15zdnd11an1n16x5 FILLER_69_2263 ();
 b15zdnd11an1n04x5 FILLER_69_2279 ();
 b15zdnd00an1n01x5 FILLER_69_2283 ();
 b15zdnd11an1n64x5 FILLER_70_8 ();
 b15zdnd11an1n64x5 FILLER_70_72 ();
 b15zdnd11an1n64x5 FILLER_70_136 ();
 b15zdnd11an1n64x5 FILLER_70_200 ();
 b15zdnd11an1n64x5 FILLER_70_264 ();
 b15zdnd11an1n64x5 FILLER_70_328 ();
 b15zdnd11an1n16x5 FILLER_70_392 ();
 b15zdnd11an1n08x5 FILLER_70_408 ();
 b15zdnd00an1n02x5 FILLER_70_416 ();
 b15zdnd11an1n64x5 FILLER_70_424 ();
 b15zdnd11an1n32x5 FILLER_70_488 ();
 b15zdnd11an1n16x5 FILLER_70_520 ();
 b15zdnd11an1n08x5 FILLER_70_536 ();
 b15zdnd11an1n04x5 FILLER_70_544 ();
 b15zdnd00an1n01x5 FILLER_70_548 ();
 b15zdnd11an1n64x5 FILLER_70_601 ();
 b15zdnd11an1n08x5 FILLER_70_665 ();
 b15zdnd11an1n04x5 FILLER_70_673 ();
 b15zdnd00an1n02x5 FILLER_70_677 ();
 b15zdnd11an1n32x5 FILLER_70_682 ();
 b15zdnd11an1n04x5 FILLER_70_714 ();
 b15zdnd11an1n64x5 FILLER_70_726 ();
 b15zdnd11an1n16x5 FILLER_70_790 ();
 b15zdnd11an1n08x5 FILLER_70_806 ();
 b15zdnd11an1n64x5 FILLER_70_831 ();
 b15zdnd11an1n64x5 FILLER_70_895 ();
 b15zdnd11an1n16x5 FILLER_70_959 ();
 b15zdnd11an1n08x5 FILLER_70_975 ();
 b15zdnd11an1n04x5 FILLER_70_983 ();
 b15zdnd11an1n64x5 FILLER_70_990 ();
 b15zdnd11an1n64x5 FILLER_70_1054 ();
 b15zdnd00an1n01x5 FILLER_70_1118 ();
 b15zdnd11an1n64x5 FILLER_70_1126 ();
 b15zdnd11an1n08x5 FILLER_70_1190 ();
 b15zdnd11an1n04x5 FILLER_70_1198 ();
 b15zdnd00an1n02x5 FILLER_70_1202 ();
 b15zdnd00an1n01x5 FILLER_70_1204 ();
 b15zdnd11an1n64x5 FILLER_70_1217 ();
 b15zdnd11an1n16x5 FILLER_70_1281 ();
 b15zdnd11an1n64x5 FILLER_70_1303 ();
 b15zdnd11an1n64x5 FILLER_70_1367 ();
 b15zdnd11an1n64x5 FILLER_70_1431 ();
 b15zdnd00an1n01x5 FILLER_70_1495 ();
 b15zdnd11an1n08x5 FILLER_70_1512 ();
 b15zdnd00an1n01x5 FILLER_70_1520 ();
 b15zdnd11an1n04x5 FILLER_70_1538 ();
 b15zdnd11an1n64x5 FILLER_70_1551 ();
 b15zdnd11an1n64x5 FILLER_70_1615 ();
 b15zdnd11an1n64x5 FILLER_70_1679 ();
 b15zdnd11an1n64x5 FILLER_70_1743 ();
 b15zdnd11an1n64x5 FILLER_70_1807 ();
 b15zdnd11an1n32x5 FILLER_70_1871 ();
 b15zdnd11an1n16x5 FILLER_70_1903 ();
 b15zdnd11an1n04x5 FILLER_70_1922 ();
 b15zdnd11an1n04x5 FILLER_70_1929 ();
 b15zdnd11an1n64x5 FILLER_70_1936 ();
 b15zdnd11an1n64x5 FILLER_70_2000 ();
 b15zdnd11an1n64x5 FILLER_70_2064 ();
 b15zdnd11an1n16x5 FILLER_70_2128 ();
 b15zdnd11an1n08x5 FILLER_70_2144 ();
 b15zdnd00an1n02x5 FILLER_70_2152 ();
 b15zdnd11an1n64x5 FILLER_70_2162 ();
 b15zdnd11an1n32x5 FILLER_70_2226 ();
 b15zdnd11an1n16x5 FILLER_70_2258 ();
 b15zdnd00an1n02x5 FILLER_70_2274 ();
 b15zdnd11an1n64x5 FILLER_71_0 ();
 b15zdnd11an1n64x5 FILLER_71_64 ();
 b15zdnd11an1n64x5 FILLER_71_128 ();
 b15zdnd11an1n16x5 FILLER_71_192 ();
 b15zdnd11an1n64x5 FILLER_71_213 ();
 b15zdnd11an1n64x5 FILLER_71_277 ();
 b15zdnd11an1n64x5 FILLER_71_341 ();
 b15zdnd11an1n64x5 FILLER_71_449 ();
 b15zdnd11an1n32x5 FILLER_71_513 ();
 b15zdnd00an1n02x5 FILLER_71_545 ();
 b15zdnd00an1n01x5 FILLER_71_547 ();
 b15zdnd11an1n32x5 FILLER_71_600 ();
 b15zdnd11an1n16x5 FILLER_71_632 ();
 b15zdnd11an1n04x5 FILLER_71_648 ();
 b15zdnd11an1n64x5 FILLER_71_704 ();
 b15zdnd11an1n32x5 FILLER_71_768 ();
 b15zdnd11an1n16x5 FILLER_71_800 ();
 b15zdnd11an1n04x5 FILLER_71_816 ();
 b15zdnd00an1n01x5 FILLER_71_820 ();
 b15zdnd11an1n64x5 FILLER_71_828 ();
 b15zdnd11an1n64x5 FILLER_71_892 ();
 b15zdnd11an1n64x5 FILLER_71_956 ();
 b15zdnd11an1n08x5 FILLER_71_1020 ();
 b15zdnd11an1n04x5 FILLER_71_1028 ();
 b15zdnd00an1n02x5 FILLER_71_1032 ();
 b15zdnd11an1n16x5 FILLER_71_1050 ();
 b15zdnd11an1n08x5 FILLER_71_1066 ();
 b15zdnd11an1n16x5 FILLER_71_1081 ();
 b15zdnd11an1n08x5 FILLER_71_1097 ();
 b15zdnd00an1n02x5 FILLER_71_1105 ();
 b15zdnd00an1n01x5 FILLER_71_1107 ();
 b15zdnd11an1n64x5 FILLER_71_1111 ();
 b15zdnd11an1n64x5 FILLER_71_1175 ();
 b15zdnd11an1n16x5 FILLER_71_1239 ();
 b15zdnd11an1n64x5 FILLER_71_1266 ();
 b15zdnd11an1n64x5 FILLER_71_1330 ();
 b15zdnd11an1n64x5 FILLER_71_1394 ();
 b15zdnd11an1n64x5 FILLER_71_1458 ();
 b15zdnd11an1n64x5 FILLER_71_1522 ();
 b15zdnd11an1n64x5 FILLER_71_1586 ();
 b15zdnd11an1n64x5 FILLER_71_1650 ();
 b15zdnd11an1n64x5 FILLER_71_1714 ();
 b15zdnd11an1n64x5 FILLER_71_1778 ();
 b15zdnd11an1n64x5 FILLER_71_1842 ();
 b15zdnd11an1n64x5 FILLER_71_1906 ();
 b15zdnd11an1n64x5 FILLER_71_1970 ();
 b15zdnd11an1n64x5 FILLER_71_2034 ();
 b15zdnd11an1n64x5 FILLER_71_2098 ();
 b15zdnd11an1n64x5 FILLER_71_2162 ();
 b15zdnd11an1n32x5 FILLER_71_2226 ();
 b15zdnd11an1n16x5 FILLER_71_2258 ();
 b15zdnd11an1n08x5 FILLER_71_2274 ();
 b15zdnd00an1n02x5 FILLER_71_2282 ();
 b15zdnd11an1n64x5 FILLER_72_8 ();
 b15zdnd11an1n64x5 FILLER_72_72 ();
 b15zdnd11an1n64x5 FILLER_72_136 ();
 b15zdnd11an1n64x5 FILLER_72_200 ();
 b15zdnd11an1n64x5 FILLER_72_264 ();
 b15zdnd11an1n08x5 FILLER_72_328 ();
 b15zdnd00an1n02x5 FILLER_72_336 ();
 b15zdnd00an1n01x5 FILLER_72_338 ();
 b15zdnd11an1n64x5 FILLER_72_343 ();
 b15zdnd11an1n16x5 FILLER_72_407 ();
 b15zdnd00an1n01x5 FILLER_72_423 ();
 b15zdnd11an1n64x5 FILLER_72_466 ();
 b15zdnd11an1n32x5 FILLER_72_530 ();
 b15zdnd11an1n04x5 FILLER_72_562 ();
 b15zdnd00an1n02x5 FILLER_72_566 ();
 b15zdnd11an1n04x5 FILLER_72_571 ();
 b15zdnd11an1n04x5 FILLER_72_578 ();
 b15zdnd11an1n08x5 FILLER_72_585 ();
 b15zdnd11an1n04x5 FILLER_72_593 ();
 b15zdnd00an1n01x5 FILLER_72_597 ();
 b15zdnd11an1n32x5 FILLER_72_605 ();
 b15zdnd11an1n16x5 FILLER_72_637 ();
 b15zdnd11an1n08x5 FILLER_72_705 ();
 b15zdnd11an1n04x5 FILLER_72_713 ();
 b15zdnd00an1n01x5 FILLER_72_717 ();
 b15zdnd11an1n64x5 FILLER_72_726 ();
 b15zdnd11an1n64x5 FILLER_72_790 ();
 b15zdnd11an1n64x5 FILLER_72_854 ();
 b15zdnd11an1n64x5 FILLER_72_918 ();
 b15zdnd11an1n64x5 FILLER_72_982 ();
 b15zdnd11an1n64x5 FILLER_72_1046 ();
 b15zdnd11an1n64x5 FILLER_72_1110 ();
 b15zdnd11an1n64x5 FILLER_72_1174 ();
 b15zdnd11an1n64x5 FILLER_72_1238 ();
 b15zdnd11an1n64x5 FILLER_72_1302 ();
 b15zdnd11an1n64x5 FILLER_72_1366 ();
 b15zdnd11an1n32x5 FILLER_72_1430 ();
 b15zdnd11an1n08x5 FILLER_72_1462 ();
 b15zdnd11an1n04x5 FILLER_72_1470 ();
 b15zdnd00an1n01x5 FILLER_72_1474 ();
 b15zdnd11an1n64x5 FILLER_72_1478 ();
 b15zdnd11an1n64x5 FILLER_72_1542 ();
 b15zdnd11an1n64x5 FILLER_72_1606 ();
 b15zdnd11an1n64x5 FILLER_72_1670 ();
 b15zdnd11an1n64x5 FILLER_72_1734 ();
 b15zdnd11an1n64x5 FILLER_72_1798 ();
 b15zdnd11an1n64x5 FILLER_72_1862 ();
 b15zdnd11an1n64x5 FILLER_72_1926 ();
 b15zdnd11an1n64x5 FILLER_72_1990 ();
 b15zdnd00an1n02x5 FILLER_72_2054 ();
 b15zdnd00an1n01x5 FILLER_72_2056 ();
 b15zdnd11an1n64x5 FILLER_72_2061 ();
 b15zdnd11an1n16x5 FILLER_72_2125 ();
 b15zdnd11an1n08x5 FILLER_72_2141 ();
 b15zdnd11an1n04x5 FILLER_72_2149 ();
 b15zdnd00an1n01x5 FILLER_72_2153 ();
 b15zdnd11an1n32x5 FILLER_72_2162 ();
 b15zdnd11an1n08x5 FILLER_72_2194 ();
 b15zdnd00an1n02x5 FILLER_72_2202 ();
 b15zdnd00an1n01x5 FILLER_72_2204 ();
 b15zdnd11an1n64x5 FILLER_72_2208 ();
 b15zdnd11an1n04x5 FILLER_72_2272 ();
 b15zdnd11an1n64x5 FILLER_73_0 ();
 b15zdnd11an1n64x5 FILLER_73_64 ();
 b15zdnd11an1n64x5 FILLER_73_128 ();
 b15zdnd11an1n64x5 FILLER_73_192 ();
 b15zdnd11an1n64x5 FILLER_73_256 ();
 b15zdnd11an1n64x5 FILLER_73_320 ();
 b15zdnd11an1n16x5 FILLER_73_384 ();
 b15zdnd11an1n08x5 FILLER_73_400 ();
 b15zdnd11an1n04x5 FILLER_73_429 ();
 b15zdnd11an1n04x5 FILLER_73_436 ();
 b15zdnd11an1n04x5 FILLER_73_443 ();
 b15zdnd00an1n02x5 FILLER_73_447 ();
 b15zdnd00an1n01x5 FILLER_73_449 ();
 b15zdnd11an1n16x5 FILLER_73_459 ();
 b15zdnd11an1n04x5 FILLER_73_475 ();
 b15zdnd00an1n02x5 FILLER_73_479 ();
 b15zdnd00an1n01x5 FILLER_73_481 ();
 b15zdnd11an1n08x5 FILLER_73_488 ();
 b15zdnd11an1n04x5 FILLER_73_496 ();
 b15zdnd00an1n02x5 FILLER_73_500 ();
 b15zdnd11an1n32x5 FILLER_73_508 ();
 b15zdnd11an1n16x5 FILLER_73_540 ();
 b15zdnd11an1n08x5 FILLER_73_556 ();
 b15zdnd11an1n04x5 FILLER_73_564 ();
 b15zdnd11an1n04x5 FILLER_73_571 ();
 b15zdnd11an1n32x5 FILLER_73_578 ();
 b15zdnd11an1n04x5 FILLER_73_610 ();
 b15zdnd00an1n02x5 FILLER_73_614 ();
 b15zdnd11an1n32x5 FILLER_73_623 ();
 b15zdnd11an1n08x5 FILLER_73_655 ();
 b15zdnd00an1n02x5 FILLER_73_663 ();
 b15zdnd00an1n01x5 FILLER_73_665 ();
 b15zdnd11an1n04x5 FILLER_73_669 ();
 b15zdnd11an1n04x5 FILLER_73_676 ();
 b15zdnd11an1n04x5 FILLER_73_683 ();
 b15zdnd11an1n64x5 FILLER_73_690 ();
 b15zdnd11an1n32x5 FILLER_73_754 ();
 b15zdnd11an1n16x5 FILLER_73_786 ();
 b15zdnd00an1n02x5 FILLER_73_802 ();
 b15zdnd00an1n01x5 FILLER_73_804 ();
 b15zdnd11an1n64x5 FILLER_73_819 ();
 b15zdnd11an1n16x5 FILLER_73_883 ();
 b15zdnd11an1n04x5 FILLER_73_899 ();
 b15zdnd00an1n02x5 FILLER_73_903 ();
 b15zdnd11an1n64x5 FILLER_73_912 ();
 b15zdnd11an1n64x5 FILLER_73_976 ();
 b15zdnd11an1n32x5 FILLER_73_1040 ();
 b15zdnd00an1n02x5 FILLER_73_1072 ();
 b15zdnd00an1n01x5 FILLER_73_1074 ();
 b15zdnd11an1n04x5 FILLER_73_1078 ();
 b15zdnd11an1n64x5 FILLER_73_1094 ();
 b15zdnd11an1n64x5 FILLER_73_1158 ();
 b15zdnd11an1n16x5 FILLER_73_1222 ();
 b15zdnd11an1n04x5 FILLER_73_1238 ();
 b15zdnd00an1n02x5 FILLER_73_1242 ();
 b15zdnd00an1n01x5 FILLER_73_1244 ();
 b15zdnd11an1n64x5 FILLER_73_1249 ();
 b15zdnd11an1n64x5 FILLER_73_1313 ();
 b15zdnd11an1n16x5 FILLER_73_1377 ();
 b15zdnd11an1n04x5 FILLER_73_1393 ();
 b15zdnd00an1n01x5 FILLER_73_1397 ();
 b15zdnd11an1n32x5 FILLER_73_1410 ();
 b15zdnd11an1n16x5 FILLER_73_1442 ();
 b15zdnd11an1n04x5 FILLER_73_1458 ();
 b15zdnd00an1n02x5 FILLER_73_1462 ();
 b15zdnd11an1n16x5 FILLER_73_1478 ();
 b15zdnd00an1n01x5 FILLER_73_1494 ();
 b15zdnd11an1n32x5 FILLER_73_1506 ();
 b15zdnd11an1n16x5 FILLER_73_1538 ();
 b15zdnd00an1n02x5 FILLER_73_1554 ();
 b15zdnd00an1n01x5 FILLER_73_1556 ();
 b15zdnd11an1n64x5 FILLER_73_1566 ();
 b15zdnd11an1n64x5 FILLER_73_1630 ();
 b15zdnd11an1n64x5 FILLER_73_1694 ();
 b15zdnd11an1n64x5 FILLER_73_1758 ();
 b15zdnd11an1n64x5 FILLER_73_1822 ();
 b15zdnd11an1n64x5 FILLER_73_1886 ();
 b15zdnd11an1n64x5 FILLER_73_1950 ();
 b15zdnd11an1n64x5 FILLER_73_2014 ();
 b15zdnd11an1n64x5 FILLER_73_2078 ();
 b15zdnd11an1n32x5 FILLER_73_2142 ();
 b15zdnd11an1n04x5 FILLER_73_2174 ();
 b15zdnd00an1n01x5 FILLER_73_2178 ();
 b15zdnd11an1n32x5 FILLER_73_2231 ();
 b15zdnd11an1n16x5 FILLER_73_2263 ();
 b15zdnd11an1n04x5 FILLER_73_2279 ();
 b15zdnd00an1n01x5 FILLER_73_2283 ();
 b15zdnd11an1n64x5 FILLER_74_8 ();
 b15zdnd11an1n64x5 FILLER_74_72 ();
 b15zdnd11an1n64x5 FILLER_74_136 ();
 b15zdnd11an1n64x5 FILLER_74_200 ();
 b15zdnd11an1n64x5 FILLER_74_264 ();
 b15zdnd11an1n64x5 FILLER_74_328 ();
 b15zdnd11an1n16x5 FILLER_74_392 ();
 b15zdnd11an1n08x5 FILLER_74_408 ();
 b15zdnd11an1n04x5 FILLER_74_416 ();
 b15zdnd00an1n02x5 FILLER_74_420 ();
 b15zdnd11an1n32x5 FILLER_74_425 ();
 b15zdnd11an1n16x5 FILLER_74_457 ();
 b15zdnd11an1n04x5 FILLER_74_473 ();
 b15zdnd00an1n02x5 FILLER_74_477 ();
 b15zdnd00an1n01x5 FILLER_74_479 ();
 b15zdnd11an1n04x5 FILLER_74_486 ();
 b15zdnd11an1n64x5 FILLER_74_496 ();
 b15zdnd11an1n64x5 FILLER_74_560 ();
 b15zdnd11an1n32x5 FILLER_74_624 ();
 b15zdnd11an1n16x5 FILLER_74_656 ();
 b15zdnd11an1n04x5 FILLER_74_672 ();
 b15zdnd00an1n02x5 FILLER_74_676 ();
 b15zdnd11an1n32x5 FILLER_74_681 ();
 b15zdnd11an1n04x5 FILLER_74_713 ();
 b15zdnd00an1n01x5 FILLER_74_717 ();
 b15zdnd11an1n32x5 FILLER_74_726 ();
 b15zdnd11an1n08x5 FILLER_74_758 ();
 b15zdnd00an1n01x5 FILLER_74_766 ();
 b15zdnd11an1n08x5 FILLER_74_774 ();
 b15zdnd11an1n04x5 FILLER_74_782 ();
 b15zdnd00an1n02x5 FILLER_74_786 ();
 b15zdnd11an1n08x5 FILLER_74_805 ();
 b15zdnd11an1n04x5 FILLER_74_813 ();
 b15zdnd11an1n64x5 FILLER_74_820 ();
 b15zdnd11an1n16x5 FILLER_74_884 ();
 b15zdnd00an1n02x5 FILLER_74_900 ();
 b15zdnd11an1n64x5 FILLER_74_908 ();
 b15zdnd11an1n32x5 FILLER_74_972 ();
 b15zdnd11an1n16x5 FILLER_74_1004 ();
 b15zdnd11an1n04x5 FILLER_74_1020 ();
 b15zdnd00an1n02x5 FILLER_74_1024 ();
 b15zdnd00an1n01x5 FILLER_74_1026 ();
 b15zdnd11an1n16x5 FILLER_74_1039 ();
 b15zdnd11an1n08x5 FILLER_74_1055 ();
 b15zdnd00an1n01x5 FILLER_74_1063 ();
 b15zdnd11an1n08x5 FILLER_74_1106 ();
 b15zdnd11an1n04x5 FILLER_74_1114 ();
 b15zdnd00an1n02x5 FILLER_74_1118 ();
 b15zdnd11an1n64x5 FILLER_74_1136 ();
 b15zdnd11an1n64x5 FILLER_74_1200 ();
 b15zdnd11an1n64x5 FILLER_74_1264 ();
 b15zdnd11an1n64x5 FILLER_74_1328 ();
 b15zdnd11an1n08x5 FILLER_74_1392 ();
 b15zdnd00an1n02x5 FILLER_74_1400 ();
 b15zdnd00an1n01x5 FILLER_74_1402 ();
 b15zdnd11an1n16x5 FILLER_74_1411 ();
 b15zdnd00an1n02x5 FILLER_74_1427 ();
 b15zdnd00an1n01x5 FILLER_74_1429 ();
 b15zdnd11an1n64x5 FILLER_74_1443 ();
 b15zdnd11an1n32x5 FILLER_74_1507 ();
 b15zdnd11an1n04x5 FILLER_74_1539 ();
 b15zdnd00an1n02x5 FILLER_74_1543 ();
 b15zdnd11an1n64x5 FILLER_74_1562 ();
 b15zdnd11an1n16x5 FILLER_74_1626 ();
 b15zdnd11an1n08x5 FILLER_74_1642 ();
 b15zdnd00an1n02x5 FILLER_74_1650 ();
 b15zdnd00an1n01x5 FILLER_74_1652 ();
 b15zdnd11an1n64x5 FILLER_74_1656 ();
 b15zdnd11an1n64x5 FILLER_74_1720 ();
 b15zdnd11an1n64x5 FILLER_74_1784 ();
 b15zdnd11an1n64x5 FILLER_74_1848 ();
 b15zdnd11an1n08x5 FILLER_74_1912 ();
 b15zdnd00an1n02x5 FILLER_74_1920 ();
 b15zdnd11an1n64x5 FILLER_74_1936 ();
 b15zdnd11an1n64x5 FILLER_74_2000 ();
 b15zdnd11an1n64x5 FILLER_74_2064 ();
 b15zdnd11an1n16x5 FILLER_74_2128 ();
 b15zdnd11an1n08x5 FILLER_74_2144 ();
 b15zdnd00an1n02x5 FILLER_74_2152 ();
 b15zdnd11an1n32x5 FILLER_74_2162 ();
 b15zdnd11an1n08x5 FILLER_74_2194 ();
 b15zdnd00an1n02x5 FILLER_74_2202 ();
 b15zdnd11an1n04x5 FILLER_74_2207 ();
 b15zdnd11an1n32x5 FILLER_74_2214 ();
 b15zdnd11an1n16x5 FILLER_74_2246 ();
 b15zdnd11an1n08x5 FILLER_74_2262 ();
 b15zdnd11an1n04x5 FILLER_74_2270 ();
 b15zdnd00an1n02x5 FILLER_74_2274 ();
 b15zdnd11an1n64x5 FILLER_75_0 ();
 b15zdnd11an1n64x5 FILLER_75_64 ();
 b15zdnd11an1n64x5 FILLER_75_128 ();
 b15zdnd11an1n64x5 FILLER_75_192 ();
 b15zdnd11an1n64x5 FILLER_75_256 ();
 b15zdnd11an1n64x5 FILLER_75_320 ();
 b15zdnd11an1n64x5 FILLER_75_384 ();
 b15zdnd11an1n64x5 FILLER_75_448 ();
 b15zdnd11an1n64x5 FILLER_75_512 ();
 b15zdnd11an1n64x5 FILLER_75_576 ();
 b15zdnd11an1n64x5 FILLER_75_640 ();
 b15zdnd11an1n64x5 FILLER_75_704 ();
 b15zdnd11an1n16x5 FILLER_75_768 ();
 b15zdnd11an1n04x5 FILLER_75_784 ();
 b15zdnd00an1n02x5 FILLER_75_788 ();
 b15zdnd11an1n64x5 FILLER_75_804 ();
 b15zdnd11an1n08x5 FILLER_75_868 ();
 b15zdnd11an1n04x5 FILLER_75_876 ();
 b15zdnd00an1n02x5 FILLER_75_880 ();
 b15zdnd00an1n01x5 FILLER_75_882 ();
 b15zdnd11an1n64x5 FILLER_75_899 ();
 b15zdnd11an1n64x5 FILLER_75_963 ();
 b15zdnd11an1n16x5 FILLER_75_1027 ();
 b15zdnd11an1n08x5 FILLER_75_1043 ();
 b15zdnd11an1n64x5 FILLER_75_1103 ();
 b15zdnd11an1n64x5 FILLER_75_1167 ();
 b15zdnd11an1n64x5 FILLER_75_1231 ();
 b15zdnd11an1n64x5 FILLER_75_1295 ();
 b15zdnd11an1n64x5 FILLER_75_1359 ();
 b15zdnd11an1n64x5 FILLER_75_1423 ();
 b15zdnd11an1n64x5 FILLER_75_1487 ();
 b15zdnd11an1n32x5 FILLER_75_1551 ();
 b15zdnd11an1n16x5 FILLER_75_1583 ();
 b15zdnd11an1n32x5 FILLER_75_1603 ();
 b15zdnd11an1n08x5 FILLER_75_1635 ();
 b15zdnd11an1n04x5 FILLER_75_1643 ();
 b15zdnd00an1n02x5 FILLER_75_1647 ();
 b15zdnd11an1n32x5 FILLER_75_1701 ();
 b15zdnd11an1n16x5 FILLER_75_1733 ();
 b15zdnd11an1n04x5 FILLER_75_1749 ();
 b15zdnd11an1n64x5 FILLER_75_1805 ();
 b15zdnd11an1n64x5 FILLER_75_1869 ();
 b15zdnd11an1n64x5 FILLER_75_1933 ();
 b15zdnd11an1n64x5 FILLER_75_1997 ();
 b15zdnd11an1n64x5 FILLER_75_2061 ();
 b15zdnd11an1n64x5 FILLER_75_2125 ();
 b15zdnd11an1n64x5 FILLER_75_2189 ();
 b15zdnd11an1n16x5 FILLER_75_2253 ();
 b15zdnd11an1n08x5 FILLER_75_2269 ();
 b15zdnd11an1n04x5 FILLER_75_2277 ();
 b15zdnd00an1n02x5 FILLER_75_2281 ();
 b15zdnd00an1n01x5 FILLER_75_2283 ();
 b15zdnd11an1n64x5 FILLER_76_8 ();
 b15zdnd11an1n64x5 FILLER_76_72 ();
 b15zdnd11an1n64x5 FILLER_76_136 ();
 b15zdnd11an1n64x5 FILLER_76_200 ();
 b15zdnd11an1n64x5 FILLER_76_264 ();
 b15zdnd11an1n64x5 FILLER_76_328 ();
 b15zdnd11an1n64x5 FILLER_76_392 ();
 b15zdnd11an1n64x5 FILLER_76_456 ();
 b15zdnd11an1n64x5 FILLER_76_520 ();
 b15zdnd11an1n64x5 FILLER_76_584 ();
 b15zdnd11an1n64x5 FILLER_76_648 ();
 b15zdnd11an1n04x5 FILLER_76_712 ();
 b15zdnd00an1n02x5 FILLER_76_716 ();
 b15zdnd11an1n64x5 FILLER_76_726 ();
 b15zdnd11an1n64x5 FILLER_76_790 ();
 b15zdnd11an1n16x5 FILLER_76_854 ();
 b15zdnd11an1n08x5 FILLER_76_870 ();
 b15zdnd11an1n32x5 FILLER_76_892 ();
 b15zdnd11an1n04x5 FILLER_76_924 ();
 b15zdnd00an1n01x5 FILLER_76_928 ();
 b15zdnd11an1n64x5 FILLER_76_971 ();
 b15zdnd11an1n32x5 FILLER_76_1035 ();
 b15zdnd11an1n04x5 FILLER_76_1067 ();
 b15zdnd11an1n04x5 FILLER_76_1074 ();
 b15zdnd11an1n64x5 FILLER_76_1081 ();
 b15zdnd11an1n64x5 FILLER_76_1145 ();
 b15zdnd11an1n64x5 FILLER_76_1209 ();
 b15zdnd11an1n64x5 FILLER_76_1273 ();
 b15zdnd11an1n64x5 FILLER_76_1337 ();
 b15zdnd11an1n16x5 FILLER_76_1401 ();
 b15zdnd11an1n08x5 FILLER_76_1417 ();
 b15zdnd11an1n04x5 FILLER_76_1425 ();
 b15zdnd00an1n02x5 FILLER_76_1429 ();
 b15zdnd00an1n01x5 FILLER_76_1431 ();
 b15zdnd11an1n64x5 FILLER_76_1448 ();
 b15zdnd11an1n04x5 FILLER_76_1512 ();
 b15zdnd00an1n01x5 FILLER_76_1516 ();
 b15zdnd11an1n64x5 FILLER_76_1533 ();
 b15zdnd11an1n16x5 FILLER_76_1597 ();
 b15zdnd11an1n08x5 FILLER_76_1613 ();
 b15zdnd11an1n04x5 FILLER_76_1621 ();
 b15zdnd00an1n01x5 FILLER_76_1625 ();
 b15zdnd11an1n04x5 FILLER_76_1678 ();
 b15zdnd11an1n64x5 FILLER_76_1685 ();
 b15zdnd11an1n16x5 FILLER_76_1749 ();
 b15zdnd11an1n04x5 FILLER_76_1765 ();
 b15zdnd00an1n02x5 FILLER_76_1769 ();
 b15zdnd00an1n01x5 FILLER_76_1771 ();
 b15zdnd11an1n04x5 FILLER_76_1775 ();
 b15zdnd11an1n64x5 FILLER_76_1782 ();
 b15zdnd11an1n64x5 FILLER_76_1846 ();
 b15zdnd11an1n64x5 FILLER_76_1910 ();
 b15zdnd11an1n64x5 FILLER_76_1974 ();
 b15zdnd11an1n64x5 FILLER_76_2038 ();
 b15zdnd11an1n32x5 FILLER_76_2102 ();
 b15zdnd11an1n16x5 FILLER_76_2134 ();
 b15zdnd11an1n04x5 FILLER_76_2150 ();
 b15zdnd11an1n64x5 FILLER_76_2162 ();
 b15zdnd11an1n32x5 FILLER_76_2226 ();
 b15zdnd11an1n16x5 FILLER_76_2258 ();
 b15zdnd00an1n02x5 FILLER_76_2274 ();
 b15zdnd11an1n64x5 FILLER_77_0 ();
 b15zdnd11an1n64x5 FILLER_77_64 ();
 b15zdnd11an1n64x5 FILLER_77_128 ();
 b15zdnd11an1n64x5 FILLER_77_192 ();
 b15zdnd11an1n64x5 FILLER_77_256 ();
 b15zdnd11an1n64x5 FILLER_77_320 ();
 b15zdnd11an1n64x5 FILLER_77_384 ();
 b15zdnd11an1n64x5 FILLER_77_448 ();
 b15zdnd11an1n64x5 FILLER_77_512 ();
 b15zdnd11an1n64x5 FILLER_77_576 ();
 b15zdnd11an1n64x5 FILLER_77_640 ();
 b15zdnd11an1n64x5 FILLER_77_704 ();
 b15zdnd11an1n16x5 FILLER_77_768 ();
 b15zdnd11an1n04x5 FILLER_77_784 ();
 b15zdnd00an1n01x5 FILLER_77_788 ();
 b15zdnd11an1n64x5 FILLER_77_795 ();
 b15zdnd11an1n64x5 FILLER_77_859 ();
 b15zdnd11an1n64x5 FILLER_77_923 ();
 b15zdnd11an1n64x5 FILLER_77_987 ();
 b15zdnd11an1n32x5 FILLER_77_1051 ();
 b15zdnd11an1n16x5 FILLER_77_1083 ();
 b15zdnd11an1n08x5 FILLER_77_1099 ();
 b15zdnd00an1n02x5 FILLER_77_1107 ();
 b15zdnd11an1n64x5 FILLER_77_1122 ();
 b15zdnd11an1n64x5 FILLER_77_1186 ();
 b15zdnd11an1n64x5 FILLER_77_1250 ();
 b15zdnd11an1n64x5 FILLER_77_1314 ();
 b15zdnd11an1n64x5 FILLER_77_1378 ();
 b15zdnd11an1n64x5 FILLER_77_1442 ();
 b15zdnd11an1n32x5 FILLER_77_1506 ();
 b15zdnd11an1n08x5 FILLER_77_1538 ();
 b15zdnd11an1n08x5 FILLER_77_1562 ();
 b15zdnd00an1n01x5 FILLER_77_1570 ();
 b15zdnd11an1n64x5 FILLER_77_1581 ();
 b15zdnd11an1n04x5 FILLER_77_1648 ();
 b15zdnd11an1n16x5 FILLER_77_1655 ();
 b15zdnd00an1n02x5 FILLER_77_1671 ();
 b15zdnd00an1n01x5 FILLER_77_1673 ();
 b15zdnd11an1n64x5 FILLER_77_1677 ();
 b15zdnd11an1n32x5 FILLER_77_1741 ();
 b15zdnd11an1n04x5 FILLER_77_1773 ();
 b15zdnd11an1n64x5 FILLER_77_1780 ();
 b15zdnd11an1n64x5 FILLER_77_1844 ();
 b15zdnd11an1n64x5 FILLER_77_1908 ();
 b15zdnd11an1n64x5 FILLER_77_1972 ();
 b15zdnd11an1n64x5 FILLER_77_2036 ();
 b15zdnd11an1n64x5 FILLER_77_2100 ();
 b15zdnd11an1n64x5 FILLER_77_2164 ();
 b15zdnd11an1n32x5 FILLER_77_2228 ();
 b15zdnd11an1n16x5 FILLER_77_2260 ();
 b15zdnd11an1n08x5 FILLER_77_2276 ();
 b15zdnd11an1n64x5 FILLER_78_8 ();
 b15zdnd11an1n64x5 FILLER_78_72 ();
 b15zdnd11an1n64x5 FILLER_78_136 ();
 b15zdnd11an1n64x5 FILLER_78_200 ();
 b15zdnd11an1n64x5 FILLER_78_264 ();
 b15zdnd11an1n64x5 FILLER_78_328 ();
 b15zdnd11an1n64x5 FILLER_78_392 ();
 b15zdnd11an1n64x5 FILLER_78_456 ();
 b15zdnd11an1n64x5 FILLER_78_520 ();
 b15zdnd11an1n08x5 FILLER_78_584 ();
 b15zdnd11an1n04x5 FILLER_78_592 ();
 b15zdnd00an1n02x5 FILLER_78_596 ();
 b15zdnd00an1n01x5 FILLER_78_598 ();
 b15zdnd11an1n32x5 FILLER_78_608 ();
 b15zdnd11an1n08x5 FILLER_78_640 ();
 b15zdnd11an1n04x5 FILLER_78_648 ();
 b15zdnd00an1n02x5 FILLER_78_652 ();
 b15zdnd00an1n01x5 FILLER_78_654 ();
 b15zdnd11an1n32x5 FILLER_78_664 ();
 b15zdnd11an1n16x5 FILLER_78_696 ();
 b15zdnd11an1n04x5 FILLER_78_712 ();
 b15zdnd00an1n02x5 FILLER_78_716 ();
 b15zdnd11an1n64x5 FILLER_78_726 ();
 b15zdnd11an1n16x5 FILLER_78_790 ();
 b15zdnd00an1n01x5 FILLER_78_806 ();
 b15zdnd11an1n08x5 FILLER_78_810 ();
 b15zdnd11an1n04x5 FILLER_78_818 ();
 b15zdnd11an1n64x5 FILLER_78_835 ();
 b15zdnd11an1n64x5 FILLER_78_899 ();
 b15zdnd11an1n64x5 FILLER_78_963 ();
 b15zdnd11an1n64x5 FILLER_78_1027 ();
 b15zdnd11an1n64x5 FILLER_78_1091 ();
 b15zdnd11an1n64x5 FILLER_78_1155 ();
 b15zdnd11an1n64x5 FILLER_78_1219 ();
 b15zdnd11an1n64x5 FILLER_78_1283 ();
 b15zdnd11an1n64x5 FILLER_78_1347 ();
 b15zdnd11an1n32x5 FILLER_78_1411 ();
 b15zdnd11an1n04x5 FILLER_78_1443 ();
 b15zdnd00an1n01x5 FILLER_78_1447 ();
 b15zdnd11an1n64x5 FILLER_78_1454 ();
 b15zdnd11an1n64x5 FILLER_78_1518 ();
 b15zdnd11an1n64x5 FILLER_78_1582 ();
 b15zdnd11an1n16x5 FILLER_78_1646 ();
 b15zdnd11an1n08x5 FILLER_78_1662 ();
 b15zdnd11an1n04x5 FILLER_78_1670 ();
 b15zdnd11an1n64x5 FILLER_78_1677 ();
 b15zdnd11an1n64x5 FILLER_78_1741 ();
 b15zdnd11an1n64x5 FILLER_78_1805 ();
 b15zdnd11an1n32x5 FILLER_78_1869 ();
 b15zdnd11an1n08x5 FILLER_78_1901 ();
 b15zdnd11an1n04x5 FILLER_78_1909 ();
 b15zdnd00an1n01x5 FILLER_78_1913 ();
 b15zdnd11an1n64x5 FILLER_78_1918 ();
 b15zdnd11an1n64x5 FILLER_78_1982 ();
 b15zdnd11an1n64x5 FILLER_78_2046 ();
 b15zdnd11an1n32x5 FILLER_78_2110 ();
 b15zdnd11an1n08x5 FILLER_78_2142 ();
 b15zdnd11an1n04x5 FILLER_78_2150 ();
 b15zdnd11an1n64x5 FILLER_78_2162 ();
 b15zdnd11an1n32x5 FILLER_78_2226 ();
 b15zdnd11an1n16x5 FILLER_78_2258 ();
 b15zdnd00an1n02x5 FILLER_78_2274 ();
 b15zdnd11an1n64x5 FILLER_79_0 ();
 b15zdnd11an1n64x5 FILLER_79_64 ();
 b15zdnd11an1n64x5 FILLER_79_128 ();
 b15zdnd11an1n64x5 FILLER_79_192 ();
 b15zdnd11an1n64x5 FILLER_79_256 ();
 b15zdnd11an1n64x5 FILLER_79_320 ();
 b15zdnd11an1n64x5 FILLER_79_384 ();
 b15zdnd11an1n64x5 FILLER_79_448 ();
 b15zdnd11an1n64x5 FILLER_79_512 ();
 b15zdnd11an1n64x5 FILLER_79_576 ();
 b15zdnd11an1n64x5 FILLER_79_640 ();
 b15zdnd11an1n64x5 FILLER_79_704 ();
 b15zdnd11an1n16x5 FILLER_79_768 ();
 b15zdnd11an1n04x5 FILLER_79_784 ();
 b15zdnd00an1n01x5 FILLER_79_788 ();
 b15zdnd11an1n64x5 FILLER_79_805 ();
 b15zdnd11an1n64x5 FILLER_79_869 ();
 b15zdnd11an1n64x5 FILLER_79_933 ();
 b15zdnd11an1n64x5 FILLER_79_997 ();
 b15zdnd11an1n16x5 FILLER_79_1061 ();
 b15zdnd00an1n02x5 FILLER_79_1077 ();
 b15zdnd11an1n64x5 FILLER_79_1090 ();
 b15zdnd11an1n64x5 FILLER_79_1154 ();
 b15zdnd11an1n64x5 FILLER_79_1218 ();
 b15zdnd11an1n64x5 FILLER_79_1282 ();
 b15zdnd11an1n32x5 FILLER_79_1346 ();
 b15zdnd11an1n16x5 FILLER_79_1378 ();
 b15zdnd11an1n08x5 FILLER_79_1394 ();
 b15zdnd11an1n04x5 FILLER_79_1402 ();
 b15zdnd00an1n01x5 FILLER_79_1406 ();
 b15zdnd11an1n16x5 FILLER_79_1410 ();
 b15zdnd11an1n04x5 FILLER_79_1426 ();
 b15zdnd00an1n02x5 FILLER_79_1430 ();
 b15zdnd11an1n04x5 FILLER_79_1442 ();
 b15zdnd11an1n32x5 FILLER_79_1461 ();
 b15zdnd11an1n16x5 FILLER_79_1493 ();
 b15zdnd11an1n04x5 FILLER_79_1509 ();
 b15zdnd11an1n16x5 FILLER_79_1526 ();
 b15zdnd11an1n08x5 FILLER_79_1542 ();
 b15zdnd00an1n01x5 FILLER_79_1550 ();
 b15zdnd11an1n64x5 FILLER_79_1561 ();
 b15zdnd11an1n64x5 FILLER_79_1625 ();
 b15zdnd11an1n64x5 FILLER_79_1689 ();
 b15zdnd11an1n64x5 FILLER_79_1753 ();
 b15zdnd11an1n64x5 FILLER_79_1817 ();
 b15zdnd11an1n32x5 FILLER_79_1881 ();
 b15zdnd11an1n04x5 FILLER_79_1913 ();
 b15zdnd00an1n02x5 FILLER_79_1917 ();
 b15zdnd11an1n04x5 FILLER_79_1923 ();
 b15zdnd00an1n02x5 FILLER_79_1927 ();
 b15zdnd11an1n64x5 FILLER_79_1933 ();
 b15zdnd11an1n64x5 FILLER_79_1997 ();
 b15zdnd11an1n64x5 FILLER_79_2061 ();
 b15zdnd11an1n64x5 FILLER_79_2125 ();
 b15zdnd11an1n64x5 FILLER_79_2189 ();
 b15zdnd11an1n16x5 FILLER_79_2253 ();
 b15zdnd11an1n08x5 FILLER_79_2269 ();
 b15zdnd11an1n04x5 FILLER_79_2277 ();
 b15zdnd00an1n02x5 FILLER_79_2281 ();
 b15zdnd00an1n01x5 FILLER_79_2283 ();
 b15zdnd11an1n64x5 FILLER_80_8 ();
 b15zdnd11an1n64x5 FILLER_80_72 ();
 b15zdnd11an1n64x5 FILLER_80_136 ();
 b15zdnd11an1n32x5 FILLER_80_200 ();
 b15zdnd11an1n16x5 FILLER_80_232 ();
 b15zdnd11an1n08x5 FILLER_80_248 ();
 b15zdnd00an1n01x5 FILLER_80_256 ();
 b15zdnd11an1n64x5 FILLER_80_270 ();
 b15zdnd11an1n64x5 FILLER_80_334 ();
 b15zdnd11an1n16x5 FILLER_80_398 ();
 b15zdnd00an1n02x5 FILLER_80_414 ();
 b15zdnd00an1n01x5 FILLER_80_416 ();
 b15zdnd11an1n64x5 FILLER_80_421 ();
 b15zdnd11an1n64x5 FILLER_80_485 ();
 b15zdnd11an1n64x5 FILLER_80_549 ();
 b15zdnd11an1n64x5 FILLER_80_613 ();
 b15zdnd11an1n32x5 FILLER_80_677 ();
 b15zdnd11an1n08x5 FILLER_80_709 ();
 b15zdnd00an1n01x5 FILLER_80_717 ();
 b15zdnd11an1n64x5 FILLER_80_726 ();
 b15zdnd11an1n64x5 FILLER_80_790 ();
 b15zdnd11an1n64x5 FILLER_80_854 ();
 b15zdnd11an1n64x5 FILLER_80_918 ();
 b15zdnd11an1n32x5 FILLER_80_982 ();
 b15zdnd11an1n08x5 FILLER_80_1014 ();
 b15zdnd00an1n02x5 FILLER_80_1022 ();
 b15zdnd11an1n64x5 FILLER_80_1036 ();
 b15zdnd11an1n64x5 FILLER_80_1100 ();
 b15zdnd11an1n64x5 FILLER_80_1164 ();
 b15zdnd11an1n64x5 FILLER_80_1228 ();
 b15zdnd11an1n64x5 FILLER_80_1292 ();
 b15zdnd11an1n64x5 FILLER_80_1356 ();
 b15zdnd11an1n64x5 FILLER_80_1420 ();
 b15zdnd11an1n64x5 FILLER_80_1484 ();
 b15zdnd11an1n64x5 FILLER_80_1548 ();
 b15zdnd11an1n64x5 FILLER_80_1612 ();
 b15zdnd11an1n64x5 FILLER_80_1676 ();
 b15zdnd11an1n64x5 FILLER_80_1740 ();
 b15zdnd11an1n64x5 FILLER_80_1804 ();
 b15zdnd11an1n32x5 FILLER_80_1868 ();
 b15zdnd11an1n16x5 FILLER_80_1900 ();
 b15zdnd11an1n04x5 FILLER_80_1920 ();
 b15zdnd11an1n04x5 FILLER_80_1930 ();
 b15zdnd11an1n64x5 FILLER_80_1938 ();
 b15zdnd11an1n64x5 FILLER_80_2002 ();
 b15zdnd11an1n64x5 FILLER_80_2066 ();
 b15zdnd11an1n16x5 FILLER_80_2130 ();
 b15zdnd11an1n08x5 FILLER_80_2146 ();
 b15zdnd11an1n64x5 FILLER_80_2162 ();
 b15zdnd11an1n32x5 FILLER_80_2226 ();
 b15zdnd11an1n16x5 FILLER_80_2258 ();
 b15zdnd00an1n02x5 FILLER_80_2274 ();
 b15zdnd11an1n64x5 FILLER_81_0 ();
 b15zdnd11an1n64x5 FILLER_81_64 ();
 b15zdnd11an1n64x5 FILLER_81_128 ();
 b15zdnd11an1n16x5 FILLER_81_192 ();
 b15zdnd11an1n08x5 FILLER_81_208 ();
 b15zdnd11an1n04x5 FILLER_81_216 ();
 b15zdnd00an1n02x5 FILLER_81_220 ();
 b15zdnd11an1n16x5 FILLER_81_225 ();
 b15zdnd11an1n08x5 FILLER_81_241 ();
 b15zdnd00an1n02x5 FILLER_81_249 ();
 b15zdnd11an1n04x5 FILLER_81_258 ();
 b15zdnd11an1n64x5 FILLER_81_278 ();
 b15zdnd11an1n64x5 FILLER_81_342 ();
 b15zdnd11an1n64x5 FILLER_81_406 ();
 b15zdnd11an1n64x5 FILLER_81_470 ();
 b15zdnd11an1n64x5 FILLER_81_534 ();
 b15zdnd11an1n32x5 FILLER_81_598 ();
 b15zdnd11an1n08x5 FILLER_81_630 ();
 b15zdnd11an1n04x5 FILLER_81_638 ();
 b15zdnd00an1n02x5 FILLER_81_642 ();
 b15zdnd00an1n01x5 FILLER_81_644 ();
 b15zdnd11an1n64x5 FILLER_81_654 ();
 b15zdnd11an1n16x5 FILLER_81_718 ();
 b15zdnd11an1n04x5 FILLER_81_734 ();
 b15zdnd00an1n01x5 FILLER_81_738 ();
 b15zdnd11an1n64x5 FILLER_81_749 ();
 b15zdnd11an1n08x5 FILLER_81_813 ();
 b15zdnd11an1n04x5 FILLER_81_821 ();
 b15zdnd00an1n01x5 FILLER_81_825 ();
 b15zdnd11an1n64x5 FILLER_81_842 ();
 b15zdnd11an1n16x5 FILLER_81_906 ();
 b15zdnd11an1n08x5 FILLER_81_922 ();
 b15zdnd11an1n04x5 FILLER_81_930 ();
 b15zdnd00an1n02x5 FILLER_81_934 ();
 b15zdnd00an1n01x5 FILLER_81_936 ();
 b15zdnd11an1n16x5 FILLER_81_940 ();
 b15zdnd11an1n04x5 FILLER_81_956 ();
 b15zdnd00an1n02x5 FILLER_81_960 ();
 b15zdnd11an1n04x5 FILLER_81_976 ();
 b15zdnd11an1n64x5 FILLER_81_983 ();
 b15zdnd11an1n64x5 FILLER_81_1047 ();
 b15zdnd11an1n64x5 FILLER_81_1111 ();
 b15zdnd11an1n64x5 FILLER_81_1175 ();
 b15zdnd11an1n64x5 FILLER_81_1239 ();
 b15zdnd11an1n64x5 FILLER_81_1303 ();
 b15zdnd11an1n64x5 FILLER_81_1367 ();
 b15zdnd11an1n64x5 FILLER_81_1431 ();
 b15zdnd11an1n64x5 FILLER_81_1495 ();
 b15zdnd11an1n64x5 FILLER_81_1559 ();
 b15zdnd11an1n64x5 FILLER_81_1623 ();
 b15zdnd11an1n64x5 FILLER_81_1687 ();
 b15zdnd11an1n64x5 FILLER_81_1751 ();
 b15zdnd11an1n64x5 FILLER_81_1815 ();
 b15zdnd11an1n64x5 FILLER_81_1879 ();
 b15zdnd11an1n64x5 FILLER_81_1943 ();
 b15zdnd11an1n64x5 FILLER_81_2007 ();
 b15zdnd11an1n64x5 FILLER_81_2071 ();
 b15zdnd11an1n32x5 FILLER_81_2135 ();
 b15zdnd11an1n08x5 FILLER_81_2167 ();
 b15zdnd11an1n64x5 FILLER_81_2196 ();
 b15zdnd11an1n16x5 FILLER_81_2260 ();
 b15zdnd11an1n08x5 FILLER_81_2276 ();
 b15zdnd11an1n64x5 FILLER_82_8 ();
 b15zdnd11an1n64x5 FILLER_82_72 ();
 b15zdnd11an1n64x5 FILLER_82_136 ();
 b15zdnd11an1n64x5 FILLER_82_200 ();
 b15zdnd00an1n02x5 FILLER_82_264 ();
 b15zdnd11an1n64x5 FILLER_82_276 ();
 b15zdnd11an1n64x5 FILLER_82_340 ();
 b15zdnd11an1n08x5 FILLER_82_404 ();
 b15zdnd11an1n04x5 FILLER_82_412 ();
 b15zdnd00an1n01x5 FILLER_82_416 ();
 b15zdnd11an1n64x5 FILLER_82_421 ();
 b15zdnd11an1n64x5 FILLER_82_485 ();
 b15zdnd11an1n16x5 FILLER_82_549 ();
 b15zdnd11an1n08x5 FILLER_82_565 ();
 b15zdnd11an1n04x5 FILLER_82_573 ();
 b15zdnd00an1n02x5 FILLER_82_577 ();
 b15zdnd11an1n08x5 FILLER_82_582 ();
 b15zdnd11an1n04x5 FILLER_82_590 ();
 b15zdnd00an1n01x5 FILLER_82_594 ();
 b15zdnd11an1n64x5 FILLER_82_622 ();
 b15zdnd11an1n32x5 FILLER_82_686 ();
 b15zdnd11an1n64x5 FILLER_82_726 ();
 b15zdnd11an1n16x5 FILLER_82_790 ();
 b15zdnd11an1n64x5 FILLER_82_820 ();
 b15zdnd11an1n32x5 FILLER_82_884 ();
 b15zdnd11an1n08x5 FILLER_82_916 ();
 b15zdnd11an1n04x5 FILLER_82_924 ();
 b15zdnd11an1n64x5 FILLER_82_941 ();
 b15zdnd11an1n64x5 FILLER_82_1005 ();
 b15zdnd11an1n64x5 FILLER_82_1069 ();
 b15zdnd11an1n64x5 FILLER_82_1133 ();
 b15zdnd11an1n64x5 FILLER_82_1197 ();
 b15zdnd11an1n64x5 FILLER_82_1261 ();
 b15zdnd11an1n64x5 FILLER_82_1325 ();
 b15zdnd11an1n64x5 FILLER_82_1389 ();
 b15zdnd11an1n08x5 FILLER_82_1453 ();
 b15zdnd11an1n04x5 FILLER_82_1461 ();
 b15zdnd00an1n02x5 FILLER_82_1465 ();
 b15zdnd11an1n64x5 FILLER_82_1470 ();
 b15zdnd11an1n64x5 FILLER_82_1534 ();
 b15zdnd11an1n64x5 FILLER_82_1598 ();
 b15zdnd11an1n64x5 FILLER_82_1662 ();
 b15zdnd11an1n64x5 FILLER_82_1726 ();
 b15zdnd11an1n64x5 FILLER_82_1790 ();
 b15zdnd11an1n64x5 FILLER_82_1854 ();
 b15zdnd11an1n64x5 FILLER_82_1918 ();
 b15zdnd11an1n64x5 FILLER_82_1982 ();
 b15zdnd11an1n64x5 FILLER_82_2046 ();
 b15zdnd11an1n32x5 FILLER_82_2110 ();
 b15zdnd11an1n08x5 FILLER_82_2142 ();
 b15zdnd11an1n04x5 FILLER_82_2150 ();
 b15zdnd11an1n64x5 FILLER_82_2162 ();
 b15zdnd11an1n32x5 FILLER_82_2226 ();
 b15zdnd11an1n16x5 FILLER_82_2258 ();
 b15zdnd00an1n02x5 FILLER_82_2274 ();
 b15zdnd11an1n64x5 FILLER_83_0 ();
 b15zdnd11an1n64x5 FILLER_83_64 ();
 b15zdnd11an1n64x5 FILLER_83_128 ();
 b15zdnd11an1n64x5 FILLER_83_192 ();
 b15zdnd00an1n02x5 FILLER_83_256 ();
 b15zdnd11an1n64x5 FILLER_83_263 ();
 b15zdnd11an1n64x5 FILLER_83_327 ();
 b15zdnd11an1n64x5 FILLER_83_391 ();
 b15zdnd11an1n64x5 FILLER_83_455 ();
 b15zdnd11an1n64x5 FILLER_83_519 ();
 b15zdnd11an1n64x5 FILLER_83_583 ();
 b15zdnd11an1n64x5 FILLER_83_647 ();
 b15zdnd11an1n32x5 FILLER_83_711 ();
 b15zdnd00an1n02x5 FILLER_83_743 ();
 b15zdnd11an1n04x5 FILLER_83_753 ();
 b15zdnd11an1n64x5 FILLER_83_765 ();
 b15zdnd11an1n64x5 FILLER_83_829 ();
 b15zdnd11an1n32x5 FILLER_83_893 ();
 b15zdnd11an1n64x5 FILLER_83_928 ();
 b15zdnd11an1n64x5 FILLER_83_992 ();
 b15zdnd11an1n64x5 FILLER_83_1056 ();
 b15zdnd11an1n16x5 FILLER_83_1120 ();
 b15zdnd11an1n04x5 FILLER_83_1136 ();
 b15zdnd00an1n02x5 FILLER_83_1140 ();
 b15zdnd11an1n64x5 FILLER_83_1162 ();
 b15zdnd11an1n64x5 FILLER_83_1226 ();
 b15zdnd11an1n64x5 FILLER_83_1290 ();
 b15zdnd11an1n64x5 FILLER_83_1354 ();
 b15zdnd11an1n64x5 FILLER_83_1418 ();
 b15zdnd11an1n64x5 FILLER_83_1482 ();
 b15zdnd11an1n64x5 FILLER_83_1546 ();
 b15zdnd11an1n64x5 FILLER_83_1610 ();
 b15zdnd11an1n08x5 FILLER_83_1674 ();
 b15zdnd11an1n32x5 FILLER_83_1691 ();
 b15zdnd11an1n08x5 FILLER_83_1723 ();
 b15zdnd11an1n04x5 FILLER_83_1731 ();
 b15zdnd00an1n02x5 FILLER_83_1735 ();
 b15zdnd00an1n01x5 FILLER_83_1737 ();
 b15zdnd11an1n64x5 FILLER_83_1747 ();
 b15zdnd11an1n64x5 FILLER_83_1811 ();
 b15zdnd11an1n64x5 FILLER_83_1875 ();
 b15zdnd11an1n64x5 FILLER_83_1939 ();
 b15zdnd11an1n64x5 FILLER_83_2003 ();
 b15zdnd11an1n64x5 FILLER_83_2067 ();
 b15zdnd11an1n64x5 FILLER_83_2131 ();
 b15zdnd11an1n64x5 FILLER_83_2195 ();
 b15zdnd11an1n16x5 FILLER_83_2259 ();
 b15zdnd11an1n08x5 FILLER_83_2275 ();
 b15zdnd00an1n01x5 FILLER_83_2283 ();
 b15zdnd11an1n64x5 FILLER_84_8 ();
 b15zdnd11an1n64x5 FILLER_84_72 ();
 b15zdnd11an1n64x5 FILLER_84_136 ();
 b15zdnd11an1n32x5 FILLER_84_200 ();
 b15zdnd11an1n16x5 FILLER_84_232 ();
 b15zdnd11an1n08x5 FILLER_84_248 ();
 b15zdnd11an1n04x5 FILLER_84_256 ();
 b15zdnd00an1n01x5 FILLER_84_260 ();
 b15zdnd11an1n64x5 FILLER_84_272 ();
 b15zdnd11an1n64x5 FILLER_84_336 ();
 b15zdnd11an1n64x5 FILLER_84_400 ();
 b15zdnd11an1n64x5 FILLER_84_464 ();
 b15zdnd11an1n64x5 FILLER_84_528 ();
 b15zdnd11an1n64x5 FILLER_84_592 ();
 b15zdnd11an1n32x5 FILLER_84_656 ();
 b15zdnd11an1n16x5 FILLER_84_688 ();
 b15zdnd11an1n08x5 FILLER_84_704 ();
 b15zdnd11an1n04x5 FILLER_84_712 ();
 b15zdnd00an1n02x5 FILLER_84_716 ();
 b15zdnd11an1n64x5 FILLER_84_726 ();
 b15zdnd11an1n16x5 FILLER_84_790 ();
 b15zdnd11an1n04x5 FILLER_84_806 ();
 b15zdnd00an1n02x5 FILLER_84_810 ();
 b15zdnd00an1n01x5 FILLER_84_812 ();
 b15zdnd11an1n64x5 FILLER_84_827 ();
 b15zdnd11an1n64x5 FILLER_84_891 ();
 b15zdnd11an1n64x5 FILLER_84_955 ();
 b15zdnd11an1n64x5 FILLER_84_1019 ();
 b15zdnd11an1n32x5 FILLER_84_1083 ();
 b15zdnd11an1n16x5 FILLER_84_1115 ();
 b15zdnd11an1n08x5 FILLER_84_1131 ();
 b15zdnd11an1n32x5 FILLER_84_1155 ();
 b15zdnd11an1n16x5 FILLER_84_1187 ();
 b15zdnd11an1n04x5 FILLER_84_1203 ();
 b15zdnd11an1n04x5 FILLER_84_1210 ();
 b15zdnd11an1n64x5 FILLER_84_1217 ();
 b15zdnd11an1n64x5 FILLER_84_1281 ();
 b15zdnd11an1n64x5 FILLER_84_1345 ();
 b15zdnd11an1n64x5 FILLER_84_1409 ();
 b15zdnd11an1n64x5 FILLER_84_1473 ();
 b15zdnd11an1n64x5 FILLER_84_1537 ();
 b15zdnd11an1n16x5 FILLER_84_1601 ();
 b15zdnd11an1n04x5 FILLER_84_1617 ();
 b15zdnd00an1n02x5 FILLER_84_1621 ();
 b15zdnd00an1n01x5 FILLER_84_1623 ();
 b15zdnd11an1n64x5 FILLER_84_1651 ();
 b15zdnd00an1n02x5 FILLER_84_1715 ();
 b15zdnd11an1n64x5 FILLER_84_1726 ();
 b15zdnd11an1n64x5 FILLER_84_1790 ();
 b15zdnd11an1n64x5 FILLER_84_1854 ();
 b15zdnd11an1n64x5 FILLER_84_1918 ();
 b15zdnd11an1n64x5 FILLER_84_1982 ();
 b15zdnd11an1n64x5 FILLER_84_2046 ();
 b15zdnd11an1n32x5 FILLER_84_2110 ();
 b15zdnd11an1n08x5 FILLER_84_2142 ();
 b15zdnd11an1n04x5 FILLER_84_2150 ();
 b15zdnd11an1n64x5 FILLER_84_2162 ();
 b15zdnd11an1n32x5 FILLER_84_2226 ();
 b15zdnd11an1n16x5 FILLER_84_2258 ();
 b15zdnd00an1n02x5 FILLER_84_2274 ();
 b15zdnd11an1n64x5 FILLER_85_0 ();
 b15zdnd11an1n64x5 FILLER_85_64 ();
 b15zdnd11an1n64x5 FILLER_85_128 ();
 b15zdnd11an1n32x5 FILLER_85_192 ();
 b15zdnd11an1n16x5 FILLER_85_224 ();
 b15zdnd11an1n08x5 FILLER_85_240 ();
 b15zdnd11an1n04x5 FILLER_85_248 ();
 b15zdnd00an1n02x5 FILLER_85_252 ();
 b15zdnd11an1n04x5 FILLER_85_259 ();
 b15zdnd11an1n64x5 FILLER_85_305 ();
 b15zdnd11an1n64x5 FILLER_85_369 ();
 b15zdnd11an1n64x5 FILLER_85_433 ();
 b15zdnd11an1n64x5 FILLER_85_497 ();
 b15zdnd11an1n64x5 FILLER_85_561 ();
 b15zdnd11an1n64x5 FILLER_85_625 ();
 b15zdnd11an1n64x5 FILLER_85_689 ();
 b15zdnd11an1n64x5 FILLER_85_753 ();
 b15zdnd11an1n64x5 FILLER_85_817 ();
 b15zdnd11an1n64x5 FILLER_85_881 ();
 b15zdnd11an1n64x5 FILLER_85_945 ();
 b15zdnd11an1n64x5 FILLER_85_1009 ();
 b15zdnd11an1n64x5 FILLER_85_1073 ();
 b15zdnd11an1n64x5 FILLER_85_1137 ();
 b15zdnd11an1n04x5 FILLER_85_1201 ();
 b15zdnd00an1n02x5 FILLER_85_1205 ();
 b15zdnd11an1n04x5 FILLER_85_1210 ();
 b15zdnd11an1n16x5 FILLER_85_1217 ();
 b15zdnd11an1n08x5 FILLER_85_1233 ();
 b15zdnd11an1n04x5 FILLER_85_1241 ();
 b15zdnd00an1n02x5 FILLER_85_1245 ();
 b15zdnd00an1n01x5 FILLER_85_1247 ();
 b15zdnd11an1n32x5 FILLER_85_1251 ();
 b15zdnd11an1n16x5 FILLER_85_1283 ();
 b15zdnd11an1n04x5 FILLER_85_1299 ();
 b15zdnd00an1n02x5 FILLER_85_1303 ();
 b15zdnd11an1n32x5 FILLER_85_1308 ();
 b15zdnd11an1n08x5 FILLER_85_1347 ();
 b15zdnd11an1n04x5 FILLER_85_1355 ();
 b15zdnd00an1n02x5 FILLER_85_1359 ();
 b15zdnd11an1n04x5 FILLER_85_1364 ();
 b15zdnd11an1n64x5 FILLER_85_1371 ();
 b15zdnd11an1n64x5 FILLER_85_1435 ();
 b15zdnd11an1n64x5 FILLER_85_1499 ();
 b15zdnd11an1n32x5 FILLER_85_1563 ();
 b15zdnd11an1n16x5 FILLER_85_1595 ();
 b15zdnd11an1n08x5 FILLER_85_1611 ();
 b15zdnd11an1n04x5 FILLER_85_1619 ();
 b15zdnd00an1n01x5 FILLER_85_1623 ();
 b15zdnd11an1n64x5 FILLER_85_1627 ();
 b15zdnd11an1n64x5 FILLER_85_1691 ();
 b15zdnd11an1n16x5 FILLER_85_1755 ();
 b15zdnd00an1n02x5 FILLER_85_1771 ();
 b15zdnd00an1n01x5 FILLER_85_1773 ();
 b15zdnd11an1n04x5 FILLER_85_1777 ();
 b15zdnd11an1n64x5 FILLER_85_1784 ();
 b15zdnd11an1n64x5 FILLER_85_1848 ();
 b15zdnd11an1n64x5 FILLER_85_1912 ();
 b15zdnd11an1n64x5 FILLER_85_1976 ();
 b15zdnd11an1n64x5 FILLER_85_2040 ();
 b15zdnd11an1n64x5 FILLER_85_2104 ();
 b15zdnd11an1n64x5 FILLER_85_2168 ();
 b15zdnd11an1n32x5 FILLER_85_2232 ();
 b15zdnd11an1n16x5 FILLER_85_2264 ();
 b15zdnd11an1n04x5 FILLER_85_2280 ();
 b15zdnd11an1n64x5 FILLER_86_8 ();
 b15zdnd11an1n64x5 FILLER_86_72 ();
 b15zdnd11an1n64x5 FILLER_86_136 ();
 b15zdnd11an1n32x5 FILLER_86_200 ();
 b15zdnd11an1n16x5 FILLER_86_232 ();
 b15zdnd11an1n08x5 FILLER_86_248 ();
 b15zdnd11an1n04x5 FILLER_86_256 ();
 b15zdnd00an1n02x5 FILLER_86_260 ();
 b15zdnd11an1n64x5 FILLER_86_266 ();
 b15zdnd11an1n64x5 FILLER_86_330 ();
 b15zdnd11an1n64x5 FILLER_86_394 ();
 b15zdnd11an1n64x5 FILLER_86_458 ();
 b15zdnd11an1n64x5 FILLER_86_522 ();
 b15zdnd11an1n64x5 FILLER_86_586 ();
 b15zdnd11an1n64x5 FILLER_86_650 ();
 b15zdnd11an1n04x5 FILLER_86_714 ();
 b15zdnd11an1n64x5 FILLER_86_726 ();
 b15zdnd11an1n64x5 FILLER_86_790 ();
 b15zdnd11an1n64x5 FILLER_86_854 ();
 b15zdnd11an1n64x5 FILLER_86_918 ();
 b15zdnd11an1n64x5 FILLER_86_982 ();
 b15zdnd11an1n08x5 FILLER_86_1046 ();
 b15zdnd11an1n04x5 FILLER_86_1054 ();
 b15zdnd00an1n01x5 FILLER_86_1058 ();
 b15zdnd11an1n32x5 FILLER_86_1066 ();
 b15zdnd11an1n16x5 FILLER_86_1098 ();
 b15zdnd00an1n02x5 FILLER_86_1114 ();
 b15zdnd11an1n32x5 FILLER_86_1128 ();
 b15zdnd11an1n16x5 FILLER_86_1160 ();
 b15zdnd11an1n08x5 FILLER_86_1176 ();
 b15zdnd00an1n02x5 FILLER_86_1184 ();
 b15zdnd00an1n01x5 FILLER_86_1186 ();
 b15zdnd11an1n04x5 FILLER_86_1239 ();
 b15zdnd00an1n02x5 FILLER_86_1243 ();
 b15zdnd00an1n01x5 FILLER_86_1245 ();
 b15zdnd11an1n04x5 FILLER_86_1273 ();
 b15zdnd00an1n02x5 FILLER_86_1277 ();
 b15zdnd11an1n08x5 FILLER_86_1331 ();
 b15zdnd11an1n04x5 FILLER_86_1339 ();
 b15zdnd11an1n64x5 FILLER_86_1395 ();
 b15zdnd11an1n64x5 FILLER_86_1459 ();
 b15zdnd11an1n16x5 FILLER_86_1523 ();
 b15zdnd11an1n04x5 FILLER_86_1539 ();
 b15zdnd00an1n01x5 FILLER_86_1543 ();
 b15zdnd11an1n64x5 FILLER_86_1556 ();
 b15zdnd11an1n64x5 FILLER_86_1620 ();
 b15zdnd11an1n64x5 FILLER_86_1684 ();
 b15zdnd11an1n08x5 FILLER_86_1748 ();
 b15zdnd11an1n64x5 FILLER_86_1808 ();
 b15zdnd11an1n64x5 FILLER_86_1872 ();
 b15zdnd11an1n64x5 FILLER_86_1936 ();
 b15zdnd11an1n64x5 FILLER_86_2000 ();
 b15zdnd11an1n64x5 FILLER_86_2064 ();
 b15zdnd11an1n16x5 FILLER_86_2128 ();
 b15zdnd11an1n08x5 FILLER_86_2144 ();
 b15zdnd00an1n02x5 FILLER_86_2152 ();
 b15zdnd11an1n64x5 FILLER_86_2162 ();
 b15zdnd11an1n32x5 FILLER_86_2226 ();
 b15zdnd11an1n16x5 FILLER_86_2258 ();
 b15zdnd00an1n02x5 FILLER_86_2274 ();
 b15zdnd11an1n64x5 FILLER_87_0 ();
 b15zdnd11an1n64x5 FILLER_87_64 ();
 b15zdnd11an1n64x5 FILLER_87_128 ();
 b15zdnd11an1n64x5 FILLER_87_192 ();
 b15zdnd11an1n08x5 FILLER_87_256 ();
 b15zdnd11an1n04x5 FILLER_87_264 ();
 b15zdnd00an1n02x5 FILLER_87_268 ();
 b15zdnd00an1n01x5 FILLER_87_270 ();
 b15zdnd11an1n64x5 FILLER_87_274 ();
 b15zdnd11an1n64x5 FILLER_87_338 ();
 b15zdnd11an1n64x5 FILLER_87_402 ();
 b15zdnd11an1n64x5 FILLER_87_466 ();
 b15zdnd11an1n64x5 FILLER_87_530 ();
 b15zdnd11an1n64x5 FILLER_87_594 ();
 b15zdnd11an1n64x5 FILLER_87_658 ();
 b15zdnd11an1n64x5 FILLER_87_722 ();
 b15zdnd11an1n64x5 FILLER_87_786 ();
 b15zdnd11an1n32x5 FILLER_87_850 ();
 b15zdnd11an1n08x5 FILLER_87_882 ();
 b15zdnd11an1n04x5 FILLER_87_890 ();
 b15zdnd00an1n01x5 FILLER_87_894 ();
 b15zdnd11an1n04x5 FILLER_87_919 ();
 b15zdnd11an1n04x5 FILLER_87_936 ();
 b15zdnd00an1n01x5 FILLER_87_940 ();
 b15zdnd11an1n64x5 FILLER_87_972 ();
 b15zdnd11an1n64x5 FILLER_87_1036 ();
 b15zdnd11an1n08x5 FILLER_87_1100 ();
 b15zdnd00an1n01x5 FILLER_87_1108 ();
 b15zdnd11an1n64x5 FILLER_87_1125 ();
 b15zdnd11an1n32x5 FILLER_87_1241 ();
 b15zdnd11an1n16x5 FILLER_87_1273 ();
 b15zdnd11an1n08x5 FILLER_87_1289 ();
 b15zdnd11an1n04x5 FILLER_87_1300 ();
 b15zdnd11an1n32x5 FILLER_87_1307 ();
 b15zdnd11an1n16x5 FILLER_87_1339 ();
 b15zdnd11an1n08x5 FILLER_87_1355 ();
 b15zdnd11an1n04x5 FILLER_87_1363 ();
 b15zdnd00an1n01x5 FILLER_87_1367 ();
 b15zdnd11an1n32x5 FILLER_87_1371 ();
 b15zdnd11an1n08x5 FILLER_87_1403 ();
 b15zdnd00an1n02x5 FILLER_87_1411 ();
 b15zdnd11an1n64x5 FILLER_87_1420 ();
 b15zdnd11an1n64x5 FILLER_87_1484 ();
 b15zdnd11an1n64x5 FILLER_87_1548 ();
 b15zdnd11an1n64x5 FILLER_87_1612 ();
 b15zdnd11an1n64x5 FILLER_87_1676 ();
 b15zdnd11an1n32x5 FILLER_87_1740 ();
 b15zdnd11an1n08x5 FILLER_87_1772 ();
 b15zdnd00an1n01x5 FILLER_87_1780 ();
 b15zdnd11an1n64x5 FILLER_87_1784 ();
 b15zdnd11an1n16x5 FILLER_87_1848 ();
 b15zdnd11an1n08x5 FILLER_87_1864 ();
 b15zdnd00an1n02x5 FILLER_87_1872 ();
 b15zdnd11an1n64x5 FILLER_87_1878 ();
 b15zdnd11an1n64x5 FILLER_87_1942 ();
 b15zdnd11an1n64x5 FILLER_87_2006 ();
 b15zdnd11an1n64x5 FILLER_87_2070 ();
 b15zdnd11an1n64x5 FILLER_87_2134 ();
 b15zdnd11an1n64x5 FILLER_87_2198 ();
 b15zdnd11an1n16x5 FILLER_87_2262 ();
 b15zdnd11an1n04x5 FILLER_87_2278 ();
 b15zdnd00an1n02x5 FILLER_87_2282 ();
 b15zdnd11an1n64x5 FILLER_88_8 ();
 b15zdnd11an1n64x5 FILLER_88_72 ();
 b15zdnd11an1n64x5 FILLER_88_136 ();
 b15zdnd11an1n32x5 FILLER_88_200 ();
 b15zdnd11an1n08x5 FILLER_88_232 ();
 b15zdnd11an1n04x5 FILLER_88_240 ();
 b15zdnd11an1n64x5 FILLER_88_296 ();
 b15zdnd11an1n64x5 FILLER_88_360 ();
 b15zdnd11an1n64x5 FILLER_88_424 ();
 b15zdnd11an1n64x5 FILLER_88_488 ();
 b15zdnd11an1n16x5 FILLER_88_552 ();
 b15zdnd11an1n04x5 FILLER_88_568 ();
 b15zdnd00an1n02x5 FILLER_88_572 ();
 b15zdnd00an1n01x5 FILLER_88_574 ();
 b15zdnd11an1n64x5 FILLER_88_578 ();
 b15zdnd11an1n64x5 FILLER_88_642 ();
 b15zdnd11an1n08x5 FILLER_88_706 ();
 b15zdnd11an1n04x5 FILLER_88_714 ();
 b15zdnd11an1n64x5 FILLER_88_726 ();
 b15zdnd11an1n64x5 FILLER_88_790 ();
 b15zdnd11an1n64x5 FILLER_88_854 ();
 b15zdnd11an1n04x5 FILLER_88_918 ();
 b15zdnd00an1n02x5 FILLER_88_922 ();
 b15zdnd11an1n64x5 FILLER_88_940 ();
 b15zdnd11an1n64x5 FILLER_88_1004 ();
 b15zdnd11an1n64x5 FILLER_88_1068 ();
 b15zdnd00an1n02x5 FILLER_88_1132 ();
 b15zdnd00an1n01x5 FILLER_88_1134 ();
 b15zdnd11an1n32x5 FILLER_88_1146 ();
 b15zdnd11an1n16x5 FILLER_88_1178 ();
 b15zdnd11an1n08x5 FILLER_88_1194 ();
 b15zdnd11an1n04x5 FILLER_88_1202 ();
 b15zdnd00an1n02x5 FILLER_88_1206 ();
 b15zdnd11an1n04x5 FILLER_88_1211 ();
 b15zdnd11an1n04x5 FILLER_88_1235 ();
 b15zdnd00an1n02x5 FILLER_88_1239 ();
 b15zdnd00an1n01x5 FILLER_88_1241 ();
 b15zdnd11an1n64x5 FILLER_88_1284 ();
 b15zdnd11an1n64x5 FILLER_88_1348 ();
 b15zdnd11an1n16x5 FILLER_88_1412 ();
 b15zdnd11an1n08x5 FILLER_88_1428 ();
 b15zdnd00an1n02x5 FILLER_88_1436 ();
 b15zdnd11an1n64x5 FILLER_88_1452 ();
 b15zdnd11an1n64x5 FILLER_88_1516 ();
 b15zdnd11an1n64x5 FILLER_88_1580 ();
 b15zdnd11an1n64x5 FILLER_88_1644 ();
 b15zdnd11an1n64x5 FILLER_88_1708 ();
 b15zdnd11an1n04x5 FILLER_88_1772 ();
 b15zdnd11an1n64x5 FILLER_88_1779 ();
 b15zdnd11an1n32x5 FILLER_88_1843 ();
 b15zdnd11an1n08x5 FILLER_88_1875 ();
 b15zdnd11an1n04x5 FILLER_88_1883 ();
 b15zdnd00an1n02x5 FILLER_88_1887 ();
 b15zdnd11an1n64x5 FILLER_88_1895 ();
 b15zdnd11an1n64x5 FILLER_88_1959 ();
 b15zdnd11an1n64x5 FILLER_88_2023 ();
 b15zdnd11an1n64x5 FILLER_88_2087 ();
 b15zdnd00an1n02x5 FILLER_88_2151 ();
 b15zdnd00an1n01x5 FILLER_88_2153 ();
 b15zdnd11an1n64x5 FILLER_88_2162 ();
 b15zdnd11an1n32x5 FILLER_88_2226 ();
 b15zdnd11an1n16x5 FILLER_88_2258 ();
 b15zdnd00an1n02x5 FILLER_88_2274 ();
 b15zdnd11an1n64x5 FILLER_89_0 ();
 b15zdnd11an1n64x5 FILLER_89_64 ();
 b15zdnd11an1n64x5 FILLER_89_128 ();
 b15zdnd11an1n64x5 FILLER_89_192 ();
 b15zdnd11an1n04x5 FILLER_89_256 ();
 b15zdnd00an1n02x5 FILLER_89_260 ();
 b15zdnd11an1n04x5 FILLER_89_265 ();
 b15zdnd11an1n64x5 FILLER_89_272 ();
 b15zdnd11an1n64x5 FILLER_89_336 ();
 b15zdnd11an1n64x5 FILLER_89_400 ();
 b15zdnd11an1n64x5 FILLER_89_464 ();
 b15zdnd11an1n16x5 FILLER_89_528 ();
 b15zdnd11an1n04x5 FILLER_89_544 ();
 b15zdnd11an1n64x5 FILLER_89_600 ();
 b15zdnd11an1n08x5 FILLER_89_664 ();
 b15zdnd11an1n04x5 FILLER_89_672 ();
 b15zdnd00an1n02x5 FILLER_89_676 ();
 b15zdnd11an1n08x5 FILLER_89_681 ();
 b15zdnd11an1n04x5 FILLER_89_689 ();
 b15zdnd00an1n02x5 FILLER_89_693 ();
 b15zdnd11an1n04x5 FILLER_89_698 ();
 b15zdnd11an1n64x5 FILLER_89_705 ();
 b15zdnd11an1n64x5 FILLER_89_769 ();
 b15zdnd11an1n64x5 FILLER_89_833 ();
 b15zdnd11an1n64x5 FILLER_89_897 ();
 b15zdnd11an1n64x5 FILLER_89_961 ();
 b15zdnd11an1n64x5 FILLER_89_1025 ();
 b15zdnd11an1n64x5 FILLER_89_1089 ();
 b15zdnd11an1n16x5 FILLER_89_1153 ();
 b15zdnd11an1n08x5 FILLER_89_1169 ();
 b15zdnd00an1n02x5 FILLER_89_1177 ();
 b15zdnd00an1n01x5 FILLER_89_1179 ();
 b15zdnd11an1n16x5 FILLER_89_1188 ();
 b15zdnd11an1n08x5 FILLER_89_1204 ();
 b15zdnd00an1n02x5 FILLER_89_1212 ();
 b15zdnd11an1n16x5 FILLER_89_1217 ();
 b15zdnd11an1n08x5 FILLER_89_1233 ();
 b15zdnd00an1n02x5 FILLER_89_1241 ();
 b15zdnd00an1n01x5 FILLER_89_1243 ();
 b15zdnd11an1n64x5 FILLER_89_1251 ();
 b15zdnd11an1n64x5 FILLER_89_1315 ();
 b15zdnd11an1n64x5 FILLER_89_1379 ();
 b15zdnd11an1n32x5 FILLER_89_1443 ();
 b15zdnd11an1n04x5 FILLER_89_1475 ();
 b15zdnd00an1n01x5 FILLER_89_1479 ();
 b15zdnd11an1n16x5 FILLER_89_1488 ();
 b15zdnd00an1n01x5 FILLER_89_1504 ();
 b15zdnd11an1n64x5 FILLER_89_1547 ();
 b15zdnd11an1n32x5 FILLER_89_1611 ();
 b15zdnd00an1n02x5 FILLER_89_1643 ();
 b15zdnd00an1n01x5 FILLER_89_1645 ();
 b15zdnd11an1n64x5 FILLER_89_1649 ();
 b15zdnd11an1n32x5 FILLER_89_1713 ();
 b15zdnd11an1n16x5 FILLER_89_1745 ();
 b15zdnd11an1n08x5 FILLER_89_1761 ();
 b15zdnd11an1n04x5 FILLER_89_1769 ();
 b15zdnd00an1n02x5 FILLER_89_1773 ();
 b15zdnd11an1n04x5 FILLER_89_1778 ();
 b15zdnd11an1n64x5 FILLER_89_1785 ();
 b15zdnd11an1n64x5 FILLER_89_1849 ();
 b15zdnd11an1n64x5 FILLER_89_1913 ();
 b15zdnd11an1n64x5 FILLER_89_1977 ();
 b15zdnd11an1n64x5 FILLER_89_2041 ();
 b15zdnd11an1n64x5 FILLER_89_2105 ();
 b15zdnd11an1n64x5 FILLER_89_2169 ();
 b15zdnd11an1n32x5 FILLER_89_2233 ();
 b15zdnd11an1n16x5 FILLER_89_2265 ();
 b15zdnd00an1n02x5 FILLER_89_2281 ();
 b15zdnd00an1n01x5 FILLER_89_2283 ();
 b15zdnd11an1n64x5 FILLER_90_8 ();
 b15zdnd11an1n64x5 FILLER_90_72 ();
 b15zdnd11an1n64x5 FILLER_90_136 ();
 b15zdnd11an1n64x5 FILLER_90_200 ();
 b15zdnd11an1n64x5 FILLER_90_264 ();
 b15zdnd11an1n64x5 FILLER_90_328 ();
 b15zdnd11an1n64x5 FILLER_90_392 ();
 b15zdnd11an1n64x5 FILLER_90_456 ();
 b15zdnd11an1n16x5 FILLER_90_520 ();
 b15zdnd11an1n08x5 FILLER_90_536 ();
 b15zdnd11an1n04x5 FILLER_90_544 ();
 b15zdnd00an1n02x5 FILLER_90_548 ();
 b15zdnd11an1n32x5 FILLER_90_602 ();
 b15zdnd11an1n16x5 FILLER_90_634 ();
 b15zdnd11an1n08x5 FILLER_90_650 ();
 b15zdnd11an1n08x5 FILLER_90_710 ();
 b15zdnd11an1n08x5 FILLER_90_726 ();
 b15zdnd11an1n04x5 FILLER_90_734 ();
 b15zdnd00an1n01x5 FILLER_90_738 ();
 b15zdnd11an1n64x5 FILLER_90_747 ();
 b15zdnd11an1n64x5 FILLER_90_811 ();
 b15zdnd11an1n64x5 FILLER_90_875 ();
 b15zdnd11an1n64x5 FILLER_90_939 ();
 b15zdnd00an1n02x5 FILLER_90_1003 ();
 b15zdnd00an1n01x5 FILLER_90_1005 ();
 b15zdnd11an1n04x5 FILLER_90_1019 ();
 b15zdnd11an1n64x5 FILLER_90_1039 ();
 b15zdnd11an1n64x5 FILLER_90_1103 ();
 b15zdnd11an1n64x5 FILLER_90_1167 ();
 b15zdnd11an1n64x5 FILLER_90_1231 ();
 b15zdnd11an1n64x5 FILLER_90_1295 ();
 b15zdnd11an1n64x5 FILLER_90_1359 ();
 b15zdnd11an1n32x5 FILLER_90_1423 ();
 b15zdnd11an1n16x5 FILLER_90_1455 ();
 b15zdnd11an1n08x5 FILLER_90_1471 ();
 b15zdnd11an1n04x5 FILLER_90_1479 ();
 b15zdnd00an1n02x5 FILLER_90_1483 ();
 b15zdnd11an1n64x5 FILLER_90_1493 ();
 b15zdnd00an1n01x5 FILLER_90_1557 ();
 b15zdnd11an1n64x5 FILLER_90_1578 ();
 b15zdnd00an1n02x5 FILLER_90_1642 ();
 b15zdnd00an1n01x5 FILLER_90_1644 ();
 b15zdnd11an1n64x5 FILLER_90_1648 ();
 b15zdnd11an1n32x5 FILLER_90_1712 ();
 b15zdnd11an1n08x5 FILLER_90_1744 ();
 b15zdnd11an1n04x5 FILLER_90_1752 ();
 b15zdnd11an1n64x5 FILLER_90_1808 ();
 b15zdnd00an1n02x5 FILLER_90_1872 ();
 b15zdnd00an1n01x5 FILLER_90_1874 ();
 b15zdnd11an1n64x5 FILLER_90_1881 ();
 b15zdnd11an1n64x5 FILLER_90_1945 ();
 b15zdnd11an1n32x5 FILLER_90_2009 ();
 b15zdnd11an1n08x5 FILLER_90_2041 ();
 b15zdnd11an1n04x5 FILLER_90_2049 ();
 b15zdnd00an1n01x5 FILLER_90_2053 ();
 b15zdnd11an1n04x5 FILLER_90_2057 ();
 b15zdnd11an1n64x5 FILLER_90_2064 ();
 b15zdnd11an1n16x5 FILLER_90_2128 ();
 b15zdnd11an1n08x5 FILLER_90_2144 ();
 b15zdnd00an1n02x5 FILLER_90_2152 ();
 b15zdnd11an1n64x5 FILLER_90_2162 ();
 b15zdnd11an1n32x5 FILLER_90_2226 ();
 b15zdnd11an1n16x5 FILLER_90_2258 ();
 b15zdnd00an1n02x5 FILLER_90_2274 ();
 b15zdnd11an1n64x5 FILLER_91_0 ();
 b15zdnd11an1n64x5 FILLER_91_64 ();
 b15zdnd11an1n64x5 FILLER_91_128 ();
 b15zdnd11an1n64x5 FILLER_91_192 ();
 b15zdnd11an1n64x5 FILLER_91_256 ();
 b15zdnd11an1n64x5 FILLER_91_320 ();
 b15zdnd11an1n64x5 FILLER_91_384 ();
 b15zdnd11an1n64x5 FILLER_91_448 ();
 b15zdnd11an1n32x5 FILLER_91_512 ();
 b15zdnd11an1n16x5 FILLER_91_544 ();
 b15zdnd00an1n02x5 FILLER_91_560 ();
 b15zdnd00an1n01x5 FILLER_91_562 ();
 b15zdnd11an1n04x5 FILLER_91_566 ();
 b15zdnd11an1n04x5 FILLER_91_573 ();
 b15zdnd11an1n04x5 FILLER_91_580 ();
 b15zdnd11an1n64x5 FILLER_91_587 ();
 b15zdnd11an1n16x5 FILLER_91_651 ();
 b15zdnd11an1n08x5 FILLER_91_667 ();
 b15zdnd00an1n02x5 FILLER_91_675 ();
 b15zdnd11an1n32x5 FILLER_91_729 ();
 b15zdnd11an1n16x5 FILLER_91_761 ();
 b15zdnd11an1n08x5 FILLER_91_777 ();
 b15zdnd00an1n02x5 FILLER_91_785 ();
 b15zdnd00an1n01x5 FILLER_91_787 ();
 b15zdnd11an1n32x5 FILLER_91_792 ();
 b15zdnd11an1n16x5 FILLER_91_824 ();
 b15zdnd11an1n04x5 FILLER_91_840 ();
 b15zdnd00an1n01x5 FILLER_91_844 ();
 b15zdnd11an1n64x5 FILLER_91_865 ();
 b15zdnd11an1n64x5 FILLER_91_929 ();
 b15zdnd11an1n64x5 FILLER_91_993 ();
 b15zdnd11an1n64x5 FILLER_91_1057 ();
 b15zdnd11an1n64x5 FILLER_91_1121 ();
 b15zdnd11an1n64x5 FILLER_91_1185 ();
 b15zdnd11an1n64x5 FILLER_91_1249 ();
 b15zdnd11an1n64x5 FILLER_91_1313 ();
 b15zdnd11an1n64x5 FILLER_91_1377 ();
 b15zdnd11an1n64x5 FILLER_91_1441 ();
 b15zdnd11an1n64x5 FILLER_91_1505 ();
 b15zdnd11an1n32x5 FILLER_91_1569 ();
 b15zdnd11an1n16x5 FILLER_91_1601 ();
 b15zdnd00an1n02x5 FILLER_91_1617 ();
 b15zdnd00an1n01x5 FILLER_91_1619 ();
 b15zdnd11an1n64x5 FILLER_91_1672 ();
 b15zdnd11an1n16x5 FILLER_91_1736 ();
 b15zdnd11an1n04x5 FILLER_91_1752 ();
 b15zdnd11an1n64x5 FILLER_91_1808 ();
 b15zdnd11an1n64x5 FILLER_91_1872 ();
 b15zdnd11an1n64x5 FILLER_91_1936 ();
 b15zdnd11an1n32x5 FILLER_91_2000 ();
 b15zdnd11an1n04x5 FILLER_91_2032 ();
 b15zdnd11an1n04x5 FILLER_91_2088 ();
 b15zdnd11an1n64x5 FILLER_91_2095 ();
 b15zdnd11an1n64x5 FILLER_91_2159 ();
 b15zdnd11an1n32x5 FILLER_91_2223 ();
 b15zdnd11an1n16x5 FILLER_91_2255 ();
 b15zdnd11an1n08x5 FILLER_91_2271 ();
 b15zdnd11an1n04x5 FILLER_91_2279 ();
 b15zdnd00an1n01x5 FILLER_91_2283 ();
 b15zdnd11an1n64x5 FILLER_92_8 ();
 b15zdnd11an1n64x5 FILLER_92_72 ();
 b15zdnd11an1n64x5 FILLER_92_136 ();
 b15zdnd11an1n64x5 FILLER_92_200 ();
 b15zdnd11an1n64x5 FILLER_92_264 ();
 b15zdnd11an1n64x5 FILLER_92_328 ();
 b15zdnd11an1n08x5 FILLER_92_392 ();
 b15zdnd11an1n04x5 FILLER_92_400 ();
 b15zdnd00an1n02x5 FILLER_92_404 ();
 b15zdnd11an1n04x5 FILLER_92_409 ();
 b15zdnd11an1n64x5 FILLER_92_416 ();
 b15zdnd11an1n64x5 FILLER_92_480 ();
 b15zdnd11an1n16x5 FILLER_92_544 ();
 b15zdnd11an1n08x5 FILLER_92_560 ();
 b15zdnd11an1n04x5 FILLER_92_568 ();
 b15zdnd00an1n01x5 FILLER_92_572 ();
 b15zdnd11an1n64x5 FILLER_92_576 ();
 b15zdnd11an1n32x5 FILLER_92_640 ();
 b15zdnd11an1n08x5 FILLER_92_672 ();
 b15zdnd11an1n04x5 FILLER_92_683 ();
 b15zdnd11an1n04x5 FILLER_92_690 ();
 b15zdnd00an1n02x5 FILLER_92_694 ();
 b15zdnd00an1n01x5 FILLER_92_696 ();
 b15zdnd11an1n16x5 FILLER_92_700 ();
 b15zdnd00an1n02x5 FILLER_92_716 ();
 b15zdnd11an1n32x5 FILLER_92_726 ();
 b15zdnd11an1n16x5 FILLER_92_758 ();
 b15zdnd00an1n02x5 FILLER_92_774 ();
 b15zdnd11an1n16x5 FILLER_92_782 ();
 b15zdnd11an1n64x5 FILLER_92_809 ();
 b15zdnd11an1n32x5 FILLER_92_873 ();
 b15zdnd00an1n02x5 FILLER_92_905 ();
 b15zdnd11an1n64x5 FILLER_92_923 ();
 b15zdnd11an1n64x5 FILLER_92_987 ();
 b15zdnd11an1n64x5 FILLER_92_1051 ();
 b15zdnd11an1n64x5 FILLER_92_1115 ();
 b15zdnd11an1n32x5 FILLER_92_1179 ();
 b15zdnd11an1n16x5 FILLER_92_1211 ();
 b15zdnd11an1n08x5 FILLER_92_1227 ();
 b15zdnd00an1n02x5 FILLER_92_1235 ();
 b15zdnd00an1n01x5 FILLER_92_1237 ();
 b15zdnd11an1n64x5 FILLER_92_1247 ();
 b15zdnd11an1n64x5 FILLER_92_1311 ();
 b15zdnd11an1n64x5 FILLER_92_1375 ();
 b15zdnd11an1n64x5 FILLER_92_1439 ();
 b15zdnd11an1n32x5 FILLER_92_1503 ();
 b15zdnd11an1n16x5 FILLER_92_1535 ();
 b15zdnd00an1n01x5 FILLER_92_1551 ();
 b15zdnd11an1n32x5 FILLER_92_1568 ();
 b15zdnd11an1n16x5 FILLER_92_1600 ();
 b15zdnd11an1n04x5 FILLER_92_1616 ();
 b15zdnd11an1n64x5 FILLER_92_1672 ();
 b15zdnd11an1n32x5 FILLER_92_1736 ();
 b15zdnd11an1n04x5 FILLER_92_1768 ();
 b15zdnd00an1n02x5 FILLER_92_1772 ();
 b15zdnd00an1n01x5 FILLER_92_1774 ();
 b15zdnd11an1n04x5 FILLER_92_1778 ();
 b15zdnd11an1n16x5 FILLER_92_1785 ();
 b15zdnd11an1n08x5 FILLER_92_1801 ();
 b15zdnd11an1n32x5 FILLER_92_1829 ();
 b15zdnd11an1n16x5 FILLER_92_1861 ();
 b15zdnd11an1n08x5 FILLER_92_1877 ();
 b15zdnd00an1n02x5 FILLER_92_1885 ();
 b15zdnd11an1n04x5 FILLER_92_1891 ();
 b15zdnd11an1n32x5 FILLER_92_1899 ();
 b15zdnd00an1n01x5 FILLER_92_1931 ();
 b15zdnd11an1n04x5 FILLER_92_1936 ();
 b15zdnd11an1n04x5 FILLER_92_1944 ();
 b15zdnd00an1n02x5 FILLER_92_1948 ();
 b15zdnd11an1n08x5 FILLER_92_1954 ();
 b15zdnd00an1n02x5 FILLER_92_1962 ();
 b15zdnd11an1n32x5 FILLER_92_1968 ();
 b15zdnd11an1n08x5 FILLER_92_2000 ();
 b15zdnd11an1n04x5 FILLER_92_2008 ();
 b15zdnd11an1n16x5 FILLER_92_2020 ();
 b15zdnd11an1n04x5 FILLER_92_2088 ();
 b15zdnd11an1n32x5 FILLER_92_2095 ();
 b15zdnd11an1n16x5 FILLER_92_2127 ();
 b15zdnd11an1n08x5 FILLER_92_2143 ();
 b15zdnd00an1n02x5 FILLER_92_2151 ();
 b15zdnd00an1n01x5 FILLER_92_2153 ();
 b15zdnd11an1n64x5 FILLER_92_2162 ();
 b15zdnd11an1n32x5 FILLER_92_2226 ();
 b15zdnd11an1n16x5 FILLER_92_2258 ();
 b15zdnd00an1n02x5 FILLER_92_2274 ();
 b15zdnd11an1n64x5 FILLER_93_0 ();
 b15zdnd11an1n64x5 FILLER_93_64 ();
 b15zdnd11an1n64x5 FILLER_93_128 ();
 b15zdnd11an1n64x5 FILLER_93_192 ();
 b15zdnd11an1n64x5 FILLER_93_256 ();
 b15zdnd11an1n64x5 FILLER_93_320 ();
 b15zdnd00an1n02x5 FILLER_93_384 ();
 b15zdnd11an1n64x5 FILLER_93_438 ();
 b15zdnd11an1n64x5 FILLER_93_502 ();
 b15zdnd11an1n64x5 FILLER_93_566 ();
 b15zdnd11an1n16x5 FILLER_93_630 ();
 b15zdnd11an1n08x5 FILLER_93_646 ();
 b15zdnd11an1n04x5 FILLER_93_654 ();
 b15zdnd00an1n02x5 FILLER_93_658 ();
 b15zdnd11an1n64x5 FILLER_93_686 ();
 b15zdnd11an1n64x5 FILLER_93_750 ();
 b15zdnd11an1n64x5 FILLER_93_814 ();
 b15zdnd11an1n64x5 FILLER_93_878 ();
 b15zdnd11an1n64x5 FILLER_93_942 ();
 b15zdnd11an1n32x5 FILLER_93_1006 ();
 b15zdnd11an1n16x5 FILLER_93_1038 ();
 b15zdnd11an1n08x5 FILLER_93_1054 ();
 b15zdnd00an1n01x5 FILLER_93_1062 ();
 b15zdnd11an1n64x5 FILLER_93_1072 ();
 b15zdnd11an1n64x5 FILLER_93_1136 ();
 b15zdnd11an1n64x5 FILLER_93_1200 ();
 b15zdnd11an1n64x5 FILLER_93_1264 ();
 b15zdnd11an1n64x5 FILLER_93_1328 ();
 b15zdnd11an1n64x5 FILLER_93_1392 ();
 b15zdnd11an1n04x5 FILLER_93_1456 ();
 b15zdnd11an1n64x5 FILLER_93_1476 ();
 b15zdnd11an1n64x5 FILLER_93_1540 ();
 b15zdnd11an1n32x5 FILLER_93_1604 ();
 b15zdnd00an1n02x5 FILLER_93_1636 ();
 b15zdnd11an1n04x5 FILLER_93_1641 ();
 b15zdnd11an1n04x5 FILLER_93_1648 ();
 b15zdnd11an1n64x5 FILLER_93_1655 ();
 b15zdnd11an1n32x5 FILLER_93_1719 ();
 b15zdnd11an1n16x5 FILLER_93_1751 ();
 b15zdnd11an1n08x5 FILLER_93_1767 ();
 b15zdnd11an1n04x5 FILLER_93_1775 ();
 b15zdnd00an1n02x5 FILLER_93_1779 ();
 b15zdnd11an1n64x5 FILLER_93_1784 ();
 b15zdnd11an1n64x5 FILLER_93_1848 ();
 b15zdnd11an1n16x5 FILLER_93_1912 ();
 b15zdnd11an1n16x5 FILLER_93_1932 ();
 b15zdnd00an1n02x5 FILLER_93_1948 ();
 b15zdnd11an1n64x5 FILLER_93_1954 ();
 b15zdnd11an1n16x5 FILLER_93_2018 ();
 b15zdnd00an1n01x5 FILLER_93_2034 ();
 b15zdnd11an1n04x5 FILLER_93_2087 ();
 b15zdnd11an1n64x5 FILLER_93_2094 ();
 b15zdnd11an1n64x5 FILLER_93_2158 ();
 b15zdnd11an1n32x5 FILLER_93_2222 ();
 b15zdnd11an1n16x5 FILLER_93_2254 ();
 b15zdnd11an1n08x5 FILLER_93_2270 ();
 b15zdnd11an1n04x5 FILLER_93_2278 ();
 b15zdnd00an1n02x5 FILLER_93_2282 ();
 b15zdnd11an1n64x5 FILLER_94_8 ();
 b15zdnd11an1n64x5 FILLER_94_72 ();
 b15zdnd11an1n64x5 FILLER_94_136 ();
 b15zdnd11an1n64x5 FILLER_94_200 ();
 b15zdnd11an1n64x5 FILLER_94_264 ();
 b15zdnd11an1n64x5 FILLER_94_328 ();
 b15zdnd11an1n08x5 FILLER_94_392 ();
 b15zdnd00an1n01x5 FILLER_94_400 ();
 b15zdnd11an1n04x5 FILLER_94_404 ();
 b15zdnd00an1n01x5 FILLER_94_408 ();
 b15zdnd11an1n64x5 FILLER_94_461 ();
 b15zdnd11an1n64x5 FILLER_94_525 ();
 b15zdnd11an1n64x5 FILLER_94_589 ();
 b15zdnd11an1n64x5 FILLER_94_653 ();
 b15zdnd00an1n01x5 FILLER_94_717 ();
 b15zdnd11an1n64x5 FILLER_94_726 ();
 b15zdnd11an1n64x5 FILLER_94_790 ();
 b15zdnd11an1n64x5 FILLER_94_854 ();
 b15zdnd11an1n16x5 FILLER_94_918 ();
 b15zdnd00an1n02x5 FILLER_94_934 ();
 b15zdnd00an1n01x5 FILLER_94_936 ();
 b15zdnd11an1n64x5 FILLER_94_957 ();
 b15zdnd11an1n64x5 FILLER_94_1021 ();
 b15zdnd11an1n64x5 FILLER_94_1085 ();
 b15zdnd11an1n64x5 FILLER_94_1149 ();
 b15zdnd11an1n64x5 FILLER_94_1213 ();
 b15zdnd11an1n64x5 FILLER_94_1277 ();
 b15zdnd11an1n64x5 FILLER_94_1341 ();
 b15zdnd11an1n16x5 FILLER_94_1405 ();
 b15zdnd11an1n08x5 FILLER_94_1421 ();
 b15zdnd11an1n04x5 FILLER_94_1429 ();
 b15zdnd00an1n02x5 FILLER_94_1433 ();
 b15zdnd11an1n04x5 FILLER_94_1441 ();
 b15zdnd11an1n04x5 FILLER_94_1466 ();
 b15zdnd11an1n64x5 FILLER_94_1483 ();
 b15zdnd11an1n64x5 FILLER_94_1547 ();
 b15zdnd11an1n16x5 FILLER_94_1611 ();
 b15zdnd11an1n08x5 FILLER_94_1627 ();
 b15zdnd11an1n04x5 FILLER_94_1635 ();
 b15zdnd00an1n01x5 FILLER_94_1639 ();
 b15zdnd11an1n64x5 FILLER_94_1643 ();
 b15zdnd11an1n64x5 FILLER_94_1707 ();
 b15zdnd11an1n64x5 FILLER_94_1771 ();
 b15zdnd11an1n64x5 FILLER_94_1835 ();
 b15zdnd11an1n16x5 FILLER_94_1899 ();
 b15zdnd11an1n08x5 FILLER_94_1915 ();
 b15zdnd11an1n16x5 FILLER_94_1927 ();
 b15zdnd11an1n08x5 FILLER_94_1943 ();
 b15zdnd00an1n01x5 FILLER_94_1951 ();
 b15zdnd11an1n64x5 FILLER_94_1956 ();
 b15zdnd11an1n08x5 FILLER_94_2026 ();
 b15zdnd00an1n02x5 FILLER_94_2034 ();
 b15zdnd11an1n64x5 FILLER_94_2088 ();
 b15zdnd00an1n02x5 FILLER_94_2152 ();
 b15zdnd11an1n64x5 FILLER_94_2162 ();
 b15zdnd11an1n32x5 FILLER_94_2226 ();
 b15zdnd11an1n16x5 FILLER_94_2258 ();
 b15zdnd00an1n02x5 FILLER_94_2274 ();
 b15zdnd11an1n64x5 FILLER_95_0 ();
 b15zdnd11an1n64x5 FILLER_95_64 ();
 b15zdnd11an1n64x5 FILLER_95_128 ();
 b15zdnd11an1n64x5 FILLER_95_192 ();
 b15zdnd11an1n64x5 FILLER_95_256 ();
 b15zdnd11an1n64x5 FILLER_95_320 ();
 b15zdnd11an1n04x5 FILLER_95_384 ();
 b15zdnd00an1n02x5 FILLER_95_388 ();
 b15zdnd00an1n01x5 FILLER_95_390 ();
 b15zdnd11an1n04x5 FILLER_95_443 ();
 b15zdnd11an1n16x5 FILLER_95_455 ();
 b15zdnd11an1n04x5 FILLER_95_471 ();
 b15zdnd00an1n02x5 FILLER_95_475 ();
 b15zdnd11an1n32x5 FILLER_95_481 ();
 b15zdnd11an1n16x5 FILLER_95_513 ();
 b15zdnd11an1n04x5 FILLER_95_529 ();
 b15zdnd11an1n64x5 FILLER_95_541 ();
 b15zdnd11an1n64x5 FILLER_95_605 ();
 b15zdnd11an1n64x5 FILLER_95_669 ();
 b15zdnd11an1n64x5 FILLER_95_733 ();
 b15zdnd11an1n64x5 FILLER_95_797 ();
 b15zdnd11an1n32x5 FILLER_95_861 ();
 b15zdnd11an1n16x5 FILLER_95_893 ();
 b15zdnd11an1n08x5 FILLER_95_909 ();
 b15zdnd00an1n02x5 FILLER_95_917 ();
 b15zdnd11an1n64x5 FILLER_95_935 ();
 b15zdnd11an1n64x5 FILLER_95_999 ();
 b15zdnd11an1n64x5 FILLER_95_1063 ();
 b15zdnd11an1n64x5 FILLER_95_1127 ();
 b15zdnd11an1n64x5 FILLER_95_1191 ();
 b15zdnd11an1n64x5 FILLER_95_1255 ();
 b15zdnd11an1n64x5 FILLER_95_1319 ();
 b15zdnd11an1n64x5 FILLER_95_1383 ();
 b15zdnd11an1n64x5 FILLER_95_1447 ();
 b15zdnd11an1n08x5 FILLER_95_1511 ();
 b15zdnd11an1n04x5 FILLER_95_1519 ();
 b15zdnd00an1n02x5 FILLER_95_1523 ();
 b15zdnd11an1n64x5 FILLER_95_1541 ();
 b15zdnd11an1n64x5 FILLER_95_1605 ();
 b15zdnd11an1n64x5 FILLER_95_1669 ();
 b15zdnd11an1n64x5 FILLER_95_1733 ();
 b15zdnd11an1n64x5 FILLER_95_1797 ();
 b15zdnd11an1n64x5 FILLER_95_1861 ();
 b15zdnd11an1n64x5 FILLER_95_1925 ();
 b15zdnd11an1n64x5 FILLER_95_1989 ();
 b15zdnd11an1n04x5 FILLER_95_2056 ();
 b15zdnd11an1n04x5 FILLER_95_2063 ();
 b15zdnd11an1n04x5 FILLER_95_2070 ();
 b15zdnd11an1n64x5 FILLER_95_2077 ();
 b15zdnd11an1n64x5 FILLER_95_2141 ();
 b15zdnd11an1n64x5 FILLER_95_2205 ();
 b15zdnd11an1n08x5 FILLER_95_2269 ();
 b15zdnd11an1n04x5 FILLER_95_2277 ();
 b15zdnd00an1n02x5 FILLER_95_2281 ();
 b15zdnd00an1n01x5 FILLER_95_2283 ();
 b15zdnd11an1n64x5 FILLER_96_8 ();
 b15zdnd11an1n64x5 FILLER_96_72 ();
 b15zdnd11an1n64x5 FILLER_96_136 ();
 b15zdnd11an1n64x5 FILLER_96_200 ();
 b15zdnd11an1n64x5 FILLER_96_264 ();
 b15zdnd11an1n64x5 FILLER_96_328 ();
 b15zdnd00an1n01x5 FILLER_96_392 ();
 b15zdnd11an1n04x5 FILLER_96_420 ();
 b15zdnd11an1n04x5 FILLER_96_427 ();
 b15zdnd11an1n04x5 FILLER_96_434 ();
 b15zdnd11an1n64x5 FILLER_96_441 ();
 b15zdnd11an1n64x5 FILLER_96_505 ();
 b15zdnd11an1n64x5 FILLER_96_569 ();
 b15zdnd11an1n64x5 FILLER_96_633 ();
 b15zdnd00an1n02x5 FILLER_96_697 ();
 b15zdnd00an1n01x5 FILLER_96_699 ();
 b15zdnd11an1n08x5 FILLER_96_704 ();
 b15zdnd11an1n04x5 FILLER_96_712 ();
 b15zdnd00an1n02x5 FILLER_96_716 ();
 b15zdnd11an1n64x5 FILLER_96_726 ();
 b15zdnd11an1n64x5 FILLER_96_790 ();
 b15zdnd11an1n64x5 FILLER_96_854 ();
 b15zdnd11an1n64x5 FILLER_96_918 ();
 b15zdnd11an1n64x5 FILLER_96_982 ();
 b15zdnd11an1n64x5 FILLER_96_1046 ();
 b15zdnd11an1n64x5 FILLER_96_1110 ();
 b15zdnd11an1n64x5 FILLER_96_1174 ();
 b15zdnd11an1n64x5 FILLER_96_1238 ();
 b15zdnd11an1n32x5 FILLER_96_1302 ();
 b15zdnd00an1n01x5 FILLER_96_1334 ();
 b15zdnd11an1n64x5 FILLER_96_1343 ();
 b15zdnd11an1n64x5 FILLER_96_1407 ();
 b15zdnd11an1n04x5 FILLER_96_1471 ();
 b15zdnd11an1n16x5 FILLER_96_1489 ();
 b15zdnd00an1n02x5 FILLER_96_1505 ();
 b15zdnd00an1n01x5 FILLER_96_1507 ();
 b15zdnd11an1n16x5 FILLER_96_1514 ();
 b15zdnd00an1n02x5 FILLER_96_1530 ();
 b15zdnd00an1n01x5 FILLER_96_1532 ();
 b15zdnd11an1n16x5 FILLER_96_1543 ();
 b15zdnd11an1n08x5 FILLER_96_1559 ();
 b15zdnd00an1n01x5 FILLER_96_1567 ();
 b15zdnd11an1n64x5 FILLER_96_1585 ();
 b15zdnd11an1n64x5 FILLER_96_1649 ();
 b15zdnd11an1n08x5 FILLER_96_1713 ();
 b15zdnd00an1n01x5 FILLER_96_1721 ();
 b15zdnd11an1n64x5 FILLER_96_1730 ();
 b15zdnd11an1n64x5 FILLER_96_1794 ();
 b15zdnd11an1n64x5 FILLER_96_1858 ();
 b15zdnd11an1n64x5 FILLER_96_1930 ();
 b15zdnd11an1n32x5 FILLER_96_1994 ();
 b15zdnd11an1n16x5 FILLER_96_2026 ();
 b15zdnd00an1n02x5 FILLER_96_2042 ();
 b15zdnd11an1n04x5 FILLER_96_2053 ();
 b15zdnd11an1n04x5 FILLER_96_2060 ();
 b15zdnd11an1n04x5 FILLER_96_2067 ();
 b15zdnd11an1n64x5 FILLER_96_2074 ();
 b15zdnd11an1n16x5 FILLER_96_2138 ();
 b15zdnd11an1n64x5 FILLER_96_2162 ();
 b15zdnd11an1n32x5 FILLER_96_2226 ();
 b15zdnd11an1n16x5 FILLER_96_2258 ();
 b15zdnd00an1n02x5 FILLER_96_2274 ();
 b15zdnd11an1n64x5 FILLER_97_0 ();
 b15zdnd11an1n64x5 FILLER_97_64 ();
 b15zdnd11an1n64x5 FILLER_97_128 ();
 b15zdnd11an1n64x5 FILLER_97_192 ();
 b15zdnd11an1n64x5 FILLER_97_256 ();
 b15zdnd11an1n64x5 FILLER_97_320 ();
 b15zdnd11an1n08x5 FILLER_97_384 ();
 b15zdnd00an1n01x5 FILLER_97_392 ();
 b15zdnd11an1n08x5 FILLER_97_396 ();
 b15zdnd11an1n04x5 FILLER_97_404 ();
 b15zdnd00an1n02x5 FILLER_97_408 ();
 b15zdnd00an1n01x5 FILLER_97_410 ();
 b15zdnd11an1n04x5 FILLER_97_414 ();
 b15zdnd11an1n08x5 FILLER_97_421 ();
 b15zdnd00an1n02x5 FILLER_97_429 ();
 b15zdnd11an1n64x5 FILLER_97_434 ();
 b15zdnd11an1n64x5 FILLER_97_498 ();
 b15zdnd11an1n64x5 FILLER_97_562 ();
 b15zdnd11an1n32x5 FILLER_97_626 ();
 b15zdnd11an1n16x5 FILLER_97_658 ();
 b15zdnd11an1n04x5 FILLER_97_674 ();
 b15zdnd00an1n02x5 FILLER_97_678 ();
 b15zdnd11an1n64x5 FILLER_97_684 ();
 b15zdnd11an1n64x5 FILLER_97_748 ();
 b15zdnd11an1n64x5 FILLER_97_812 ();
 b15zdnd11an1n64x5 FILLER_97_876 ();
 b15zdnd11an1n64x5 FILLER_97_940 ();
 b15zdnd11an1n32x5 FILLER_97_1004 ();
 b15zdnd11an1n08x5 FILLER_97_1036 ();
 b15zdnd11an1n04x5 FILLER_97_1044 ();
 b15zdnd11an1n64x5 FILLER_97_1100 ();
 b15zdnd11an1n64x5 FILLER_97_1164 ();
 b15zdnd11an1n32x5 FILLER_97_1228 ();
 b15zdnd11an1n04x5 FILLER_97_1260 ();
 b15zdnd00an1n02x5 FILLER_97_1264 ();
 b15zdnd11an1n04x5 FILLER_97_1275 ();
 b15zdnd11an1n64x5 FILLER_97_1288 ();
 b15zdnd11an1n64x5 FILLER_97_1352 ();
 b15zdnd11an1n64x5 FILLER_97_1416 ();
 b15zdnd11an1n16x5 FILLER_97_1480 ();
 b15zdnd11an1n04x5 FILLER_97_1496 ();
 b15zdnd00an1n02x5 FILLER_97_1500 ();
 b15zdnd11an1n64x5 FILLER_97_1509 ();
 b15zdnd11an1n64x5 FILLER_97_1573 ();
 b15zdnd11an1n64x5 FILLER_97_1637 ();
 b15zdnd11an1n64x5 FILLER_97_1701 ();
 b15zdnd11an1n64x5 FILLER_97_1765 ();
 b15zdnd11an1n64x5 FILLER_97_1829 ();
 b15zdnd11an1n64x5 FILLER_97_1893 ();
 b15zdnd11an1n64x5 FILLER_97_1957 ();
 b15zdnd11an1n08x5 FILLER_97_2021 ();
 b15zdnd00an1n01x5 FILLER_97_2029 ();
 b15zdnd11an1n64x5 FILLER_97_2057 ();
 b15zdnd11an1n64x5 FILLER_97_2121 ();
 b15zdnd11an1n64x5 FILLER_97_2185 ();
 b15zdnd11an1n32x5 FILLER_97_2249 ();
 b15zdnd00an1n02x5 FILLER_97_2281 ();
 b15zdnd00an1n01x5 FILLER_97_2283 ();
 b15zdnd11an1n64x5 FILLER_98_8 ();
 b15zdnd11an1n64x5 FILLER_98_72 ();
 b15zdnd11an1n64x5 FILLER_98_136 ();
 b15zdnd11an1n64x5 FILLER_98_200 ();
 b15zdnd11an1n64x5 FILLER_98_264 ();
 b15zdnd11an1n64x5 FILLER_98_328 ();
 b15zdnd11an1n64x5 FILLER_98_392 ();
 b15zdnd11an1n32x5 FILLER_98_456 ();
 b15zdnd11an1n08x5 FILLER_98_488 ();
 b15zdnd00an1n02x5 FILLER_98_496 ();
 b15zdnd11an1n08x5 FILLER_98_502 ();
 b15zdnd11an1n04x5 FILLER_98_510 ();
 b15zdnd11an1n04x5 FILLER_98_518 ();
 b15zdnd11an1n64x5 FILLER_98_526 ();
 b15zdnd11an1n64x5 FILLER_98_590 ();
 b15zdnd11an1n64x5 FILLER_98_654 ();
 b15zdnd11an1n16x5 FILLER_98_726 ();
 b15zdnd11an1n08x5 FILLER_98_742 ();
 b15zdnd11an1n04x5 FILLER_98_750 ();
 b15zdnd00an1n01x5 FILLER_98_754 ();
 b15zdnd11an1n16x5 FILLER_98_766 ();
 b15zdnd00an1n02x5 FILLER_98_782 ();
 b15zdnd11an1n64x5 FILLER_98_794 ();
 b15zdnd11an1n32x5 FILLER_98_858 ();
 b15zdnd00an1n02x5 FILLER_98_890 ();
 b15zdnd11an1n64x5 FILLER_98_909 ();
 b15zdnd11an1n32x5 FILLER_98_973 ();
 b15zdnd11an1n16x5 FILLER_98_1005 ();
 b15zdnd11an1n08x5 FILLER_98_1021 ();
 b15zdnd11an1n04x5 FILLER_98_1081 ();
 b15zdnd11an1n64x5 FILLER_98_1088 ();
 b15zdnd11an1n64x5 FILLER_98_1152 ();
 b15zdnd11an1n64x5 FILLER_98_1216 ();
 b15zdnd11an1n64x5 FILLER_98_1280 ();
 b15zdnd11an1n64x5 FILLER_98_1344 ();
 b15zdnd11an1n64x5 FILLER_98_1408 ();
 b15zdnd11an1n16x5 FILLER_98_1472 ();
 b15zdnd00an1n02x5 FILLER_98_1488 ();
 b15zdnd00an1n01x5 FILLER_98_1490 ();
 b15zdnd11an1n64x5 FILLER_98_1512 ();
 b15zdnd11an1n64x5 FILLER_98_1576 ();
 b15zdnd11an1n64x5 FILLER_98_1640 ();
 b15zdnd11an1n64x5 FILLER_98_1704 ();
 b15zdnd11an1n64x5 FILLER_98_1768 ();
 b15zdnd11an1n64x5 FILLER_98_1832 ();
 b15zdnd11an1n64x5 FILLER_98_1896 ();
 b15zdnd11an1n64x5 FILLER_98_1960 ();
 b15zdnd11an1n04x5 FILLER_98_2024 ();
 b15zdnd00an1n02x5 FILLER_98_2028 ();
 b15zdnd11an1n64x5 FILLER_98_2033 ();
 b15zdnd11an1n32x5 FILLER_98_2097 ();
 b15zdnd11an1n16x5 FILLER_98_2129 ();
 b15zdnd11an1n08x5 FILLER_98_2145 ();
 b15zdnd00an1n01x5 FILLER_98_2153 ();
 b15zdnd11an1n64x5 FILLER_98_2162 ();
 b15zdnd11an1n32x5 FILLER_98_2226 ();
 b15zdnd11an1n16x5 FILLER_98_2258 ();
 b15zdnd00an1n02x5 FILLER_98_2274 ();
 b15zdnd11an1n64x5 FILLER_99_0 ();
 b15zdnd11an1n64x5 FILLER_99_64 ();
 b15zdnd11an1n64x5 FILLER_99_128 ();
 b15zdnd11an1n64x5 FILLER_99_192 ();
 b15zdnd11an1n64x5 FILLER_99_256 ();
 b15zdnd11an1n64x5 FILLER_99_320 ();
 b15zdnd11an1n64x5 FILLER_99_384 ();
 b15zdnd11an1n64x5 FILLER_99_448 ();
 b15zdnd11an1n64x5 FILLER_99_512 ();
 b15zdnd11an1n64x5 FILLER_99_576 ();
 b15zdnd11an1n64x5 FILLER_99_640 ();
 b15zdnd11an1n64x5 FILLER_99_704 ();
 b15zdnd11an1n32x5 FILLER_99_768 ();
 b15zdnd11an1n08x5 FILLER_99_800 ();
 b15zdnd11an1n04x5 FILLER_99_808 ();
 b15zdnd00an1n02x5 FILLER_99_812 ();
 b15zdnd11an1n64x5 FILLER_99_817 ();
 b15zdnd11an1n32x5 FILLER_99_881 ();
 b15zdnd11an1n04x5 FILLER_99_913 ();
 b15zdnd00an1n01x5 FILLER_99_917 ();
 b15zdnd11an1n04x5 FILLER_99_921 ();
 b15zdnd11an1n64x5 FILLER_99_928 ();
 b15zdnd11an1n32x5 FILLER_99_992 ();
 b15zdnd11an1n16x5 FILLER_99_1024 ();
 b15zdnd11an1n08x5 FILLER_99_1040 ();
 b15zdnd00an1n01x5 FILLER_99_1048 ();
 b15zdnd11an1n04x5 FILLER_99_1052 ();
 b15zdnd11an1n04x5 FILLER_99_1059 ();
 b15zdnd00an1n02x5 FILLER_99_1063 ();
 b15zdnd00an1n01x5 FILLER_99_1065 ();
 b15zdnd11an1n04x5 FILLER_99_1069 ();
 b15zdnd11an1n64x5 FILLER_99_1076 ();
 b15zdnd11an1n64x5 FILLER_99_1140 ();
 b15zdnd11an1n64x5 FILLER_99_1204 ();
 b15zdnd11an1n64x5 FILLER_99_1268 ();
 b15zdnd11an1n64x5 FILLER_99_1332 ();
 b15zdnd11an1n64x5 FILLER_99_1396 ();
 b15zdnd11an1n64x5 FILLER_99_1460 ();
 b15zdnd11an1n64x5 FILLER_99_1524 ();
 b15zdnd11an1n64x5 FILLER_99_1588 ();
 b15zdnd11an1n64x5 FILLER_99_1652 ();
 b15zdnd11an1n64x5 FILLER_99_1716 ();
 b15zdnd11an1n64x5 FILLER_99_1780 ();
 b15zdnd11an1n64x5 FILLER_99_1844 ();
 b15zdnd11an1n64x5 FILLER_99_1908 ();
 b15zdnd11an1n64x5 FILLER_99_1972 ();
 b15zdnd11an1n64x5 FILLER_99_2036 ();
 b15zdnd11an1n64x5 FILLER_99_2100 ();
 b15zdnd11an1n64x5 FILLER_99_2164 ();
 b15zdnd11an1n32x5 FILLER_99_2228 ();
 b15zdnd11an1n16x5 FILLER_99_2260 ();
 b15zdnd11an1n08x5 FILLER_99_2276 ();
 b15zdnd11an1n64x5 FILLER_100_8 ();
 b15zdnd11an1n64x5 FILLER_100_72 ();
 b15zdnd11an1n64x5 FILLER_100_136 ();
 b15zdnd11an1n64x5 FILLER_100_200 ();
 b15zdnd11an1n64x5 FILLER_100_264 ();
 b15zdnd11an1n64x5 FILLER_100_328 ();
 b15zdnd11an1n64x5 FILLER_100_392 ();
 b15zdnd11an1n64x5 FILLER_100_456 ();
 b15zdnd11an1n64x5 FILLER_100_520 ();
 b15zdnd11an1n64x5 FILLER_100_584 ();
 b15zdnd11an1n64x5 FILLER_100_648 ();
 b15zdnd11an1n04x5 FILLER_100_712 ();
 b15zdnd00an1n02x5 FILLER_100_716 ();
 b15zdnd11an1n32x5 FILLER_100_726 ();
 b15zdnd11an1n16x5 FILLER_100_758 ();
 b15zdnd11an1n08x5 FILLER_100_774 ();
 b15zdnd11an1n04x5 FILLER_100_782 ();
 b15zdnd00an1n01x5 FILLER_100_786 ();
 b15zdnd11an1n16x5 FILLER_100_839 ();
 b15zdnd11an1n04x5 FILLER_100_855 ();
 b15zdnd00an1n02x5 FILLER_100_859 ();
 b15zdnd11an1n16x5 FILLER_100_867 ();
 b15zdnd11an1n08x5 FILLER_100_883 ();
 b15zdnd11an1n64x5 FILLER_100_943 ();
 b15zdnd11an1n32x5 FILLER_100_1007 ();
 b15zdnd11an1n08x5 FILLER_100_1039 ();
 b15zdnd00an1n01x5 FILLER_100_1047 ();
 b15zdnd11an1n64x5 FILLER_100_1051 ();
 b15zdnd11an1n64x5 FILLER_100_1115 ();
 b15zdnd11an1n64x5 FILLER_100_1179 ();
 b15zdnd11an1n64x5 FILLER_100_1243 ();
 b15zdnd11an1n64x5 FILLER_100_1307 ();
 b15zdnd11an1n64x5 FILLER_100_1371 ();
 b15zdnd11an1n64x5 FILLER_100_1435 ();
 b15zdnd11an1n64x5 FILLER_100_1499 ();
 b15zdnd11an1n64x5 FILLER_100_1563 ();
 b15zdnd11an1n64x5 FILLER_100_1627 ();
 b15zdnd11an1n64x5 FILLER_100_1691 ();
 b15zdnd11an1n64x5 FILLER_100_1755 ();
 b15zdnd11an1n64x5 FILLER_100_1819 ();
 b15zdnd11an1n64x5 FILLER_100_1883 ();
 b15zdnd11an1n64x5 FILLER_100_1947 ();
 b15zdnd11an1n64x5 FILLER_100_2011 ();
 b15zdnd11an1n64x5 FILLER_100_2075 ();
 b15zdnd11an1n08x5 FILLER_100_2139 ();
 b15zdnd11an1n04x5 FILLER_100_2147 ();
 b15zdnd00an1n02x5 FILLER_100_2151 ();
 b15zdnd00an1n01x5 FILLER_100_2153 ();
 b15zdnd11an1n64x5 FILLER_100_2162 ();
 b15zdnd11an1n32x5 FILLER_100_2226 ();
 b15zdnd11an1n16x5 FILLER_100_2258 ();
 b15zdnd00an1n02x5 FILLER_100_2274 ();
 b15zdnd11an1n64x5 FILLER_101_0 ();
 b15zdnd11an1n64x5 FILLER_101_64 ();
 b15zdnd11an1n64x5 FILLER_101_128 ();
 b15zdnd11an1n64x5 FILLER_101_192 ();
 b15zdnd11an1n16x5 FILLER_101_256 ();
 b15zdnd11an1n08x5 FILLER_101_272 ();
 b15zdnd00an1n01x5 FILLER_101_280 ();
 b15zdnd11an1n64x5 FILLER_101_284 ();
 b15zdnd11an1n64x5 FILLER_101_348 ();
 b15zdnd11an1n64x5 FILLER_101_412 ();
 b15zdnd11an1n64x5 FILLER_101_476 ();
 b15zdnd11an1n64x5 FILLER_101_540 ();
 b15zdnd11an1n64x5 FILLER_101_604 ();
 b15zdnd11an1n64x5 FILLER_101_668 ();
 b15zdnd11an1n64x5 FILLER_101_732 ();
 b15zdnd11an1n08x5 FILLER_101_796 ();
 b15zdnd00an1n02x5 FILLER_101_804 ();
 b15zdnd11an1n04x5 FILLER_101_809 ();
 b15zdnd11an1n16x5 FILLER_101_816 ();
 b15zdnd11an1n08x5 FILLER_101_832 ();
 b15zdnd00an1n02x5 FILLER_101_840 ();
 b15zdnd00an1n01x5 FILLER_101_842 ();
 b15zdnd11an1n64x5 FILLER_101_857 ();
 b15zdnd11an1n08x5 FILLER_101_921 ();
 b15zdnd11an1n04x5 FILLER_101_929 ();
 b15zdnd11an1n64x5 FILLER_101_936 ();
 b15zdnd11an1n64x5 FILLER_101_1000 ();
 b15zdnd11an1n64x5 FILLER_101_1064 ();
 b15zdnd11an1n64x5 FILLER_101_1128 ();
 b15zdnd11an1n64x5 FILLER_101_1192 ();
 b15zdnd11an1n64x5 FILLER_101_1256 ();
 b15zdnd11an1n64x5 FILLER_101_1320 ();
 b15zdnd11an1n64x5 FILLER_101_1384 ();
 b15zdnd11an1n64x5 FILLER_101_1448 ();
 b15zdnd11an1n08x5 FILLER_101_1512 ();
 b15zdnd00an1n02x5 FILLER_101_1520 ();
 b15zdnd11an1n64x5 FILLER_101_1564 ();
 b15zdnd11an1n64x5 FILLER_101_1628 ();
 b15zdnd11an1n64x5 FILLER_101_1692 ();
 b15zdnd11an1n64x5 FILLER_101_1756 ();
 b15zdnd11an1n64x5 FILLER_101_1820 ();
 b15zdnd11an1n64x5 FILLER_101_1884 ();
 b15zdnd11an1n64x5 FILLER_101_1948 ();
 b15zdnd11an1n64x5 FILLER_101_2012 ();
 b15zdnd11an1n64x5 FILLER_101_2076 ();
 b15zdnd11an1n64x5 FILLER_101_2140 ();
 b15zdnd11an1n64x5 FILLER_101_2204 ();
 b15zdnd11an1n16x5 FILLER_101_2268 ();
 b15zdnd11an1n64x5 FILLER_102_8 ();
 b15zdnd11an1n64x5 FILLER_102_72 ();
 b15zdnd11an1n64x5 FILLER_102_136 ();
 b15zdnd11an1n32x5 FILLER_102_200 ();
 b15zdnd11an1n16x5 FILLER_102_232 ();
 b15zdnd11an1n04x5 FILLER_102_248 ();
 b15zdnd00an1n02x5 FILLER_102_252 ();
 b15zdnd11an1n64x5 FILLER_102_306 ();
 b15zdnd11an1n32x5 FILLER_102_370 ();
 b15zdnd00an1n02x5 FILLER_102_402 ();
 b15zdnd00an1n01x5 FILLER_102_404 ();
 b15zdnd11an1n64x5 FILLER_102_414 ();
 b15zdnd11an1n64x5 FILLER_102_478 ();
 b15zdnd11an1n64x5 FILLER_102_542 ();
 b15zdnd11an1n64x5 FILLER_102_606 ();
 b15zdnd11an1n32x5 FILLER_102_670 ();
 b15zdnd11an1n16x5 FILLER_102_702 ();
 b15zdnd00an1n02x5 FILLER_102_726 ();
 b15zdnd11an1n32x5 FILLER_102_759 ();
 b15zdnd00an1n02x5 FILLER_102_791 ();
 b15zdnd00an1n01x5 FILLER_102_793 ();
 b15zdnd11an1n32x5 FILLER_102_802 ();
 b15zdnd11an1n08x5 FILLER_102_834 ();
 b15zdnd11an1n04x5 FILLER_102_842 ();
 b15zdnd00an1n02x5 FILLER_102_846 ();
 b15zdnd00an1n01x5 FILLER_102_848 ();
 b15zdnd11an1n32x5 FILLER_102_855 ();
 b15zdnd11an1n16x5 FILLER_102_887 ();
 b15zdnd00an1n02x5 FILLER_102_903 ();
 b15zdnd00an1n01x5 FILLER_102_905 ();
 b15zdnd11an1n32x5 FILLER_102_914 ();
 b15zdnd11an1n08x5 FILLER_102_946 ();
 b15zdnd11an1n04x5 FILLER_102_954 ();
 b15zdnd00an1n02x5 FILLER_102_958 ();
 b15zdnd11an1n64x5 FILLER_102_969 ();
 b15zdnd11an1n64x5 FILLER_102_1033 ();
 b15zdnd11an1n64x5 FILLER_102_1097 ();
 b15zdnd11an1n32x5 FILLER_102_1161 ();
 b15zdnd11an1n04x5 FILLER_102_1193 ();
 b15zdnd11an1n04x5 FILLER_102_1200 ();
 b15zdnd11an1n64x5 FILLER_102_1207 ();
 b15zdnd11an1n64x5 FILLER_102_1271 ();
 b15zdnd11an1n64x5 FILLER_102_1335 ();
 b15zdnd11an1n64x5 FILLER_102_1399 ();
 b15zdnd11an1n64x5 FILLER_102_1463 ();
 b15zdnd11an1n64x5 FILLER_102_1527 ();
 b15zdnd11an1n64x5 FILLER_102_1591 ();
 b15zdnd11an1n64x5 FILLER_102_1655 ();
 b15zdnd11an1n64x5 FILLER_102_1719 ();
 b15zdnd11an1n64x5 FILLER_102_1783 ();
 b15zdnd11an1n64x5 FILLER_102_1847 ();
 b15zdnd11an1n64x5 FILLER_102_1911 ();
 b15zdnd11an1n64x5 FILLER_102_1975 ();
 b15zdnd11an1n64x5 FILLER_102_2039 ();
 b15zdnd11an1n32x5 FILLER_102_2103 ();
 b15zdnd11an1n16x5 FILLER_102_2135 ();
 b15zdnd00an1n02x5 FILLER_102_2151 ();
 b15zdnd00an1n01x5 FILLER_102_2153 ();
 b15zdnd11an1n64x5 FILLER_102_2162 ();
 b15zdnd11an1n32x5 FILLER_102_2226 ();
 b15zdnd11an1n16x5 FILLER_102_2258 ();
 b15zdnd00an1n02x5 FILLER_102_2274 ();
 b15zdnd11an1n64x5 FILLER_103_0 ();
 b15zdnd11an1n64x5 FILLER_103_64 ();
 b15zdnd11an1n64x5 FILLER_103_128 ();
 b15zdnd11an1n64x5 FILLER_103_192 ();
 b15zdnd11an1n16x5 FILLER_103_256 ();
 b15zdnd00an1n01x5 FILLER_103_272 ();
 b15zdnd11an1n04x5 FILLER_103_276 ();
 b15zdnd11an1n64x5 FILLER_103_283 ();
 b15zdnd11an1n64x5 FILLER_103_347 ();
 b15zdnd11an1n64x5 FILLER_103_411 ();
 b15zdnd11an1n64x5 FILLER_103_475 ();
 b15zdnd11an1n64x5 FILLER_103_539 ();
 b15zdnd11an1n64x5 FILLER_103_603 ();
 b15zdnd11an1n64x5 FILLER_103_667 ();
 b15zdnd11an1n64x5 FILLER_103_731 ();
 b15zdnd11an1n64x5 FILLER_103_795 ();
 b15zdnd11an1n32x5 FILLER_103_859 ();
 b15zdnd00an1n02x5 FILLER_103_891 ();
 b15zdnd11an1n08x5 FILLER_103_901 ();
 b15zdnd11an1n04x5 FILLER_103_909 ();
 b15zdnd00an1n02x5 FILLER_103_913 ();
 b15zdnd11an1n64x5 FILLER_103_942 ();
 b15zdnd11an1n32x5 FILLER_103_1006 ();
 b15zdnd11an1n04x5 FILLER_103_1038 ();
 b15zdnd11an1n64x5 FILLER_103_1050 ();
 b15zdnd11an1n32x5 FILLER_103_1114 ();
 b15zdnd11an1n08x5 FILLER_103_1146 ();
 b15zdnd11an1n04x5 FILLER_103_1154 ();
 b15zdnd00an1n01x5 FILLER_103_1158 ();
 b15zdnd11an1n08x5 FILLER_103_1166 ();
 b15zdnd11an1n04x5 FILLER_103_1174 ();
 b15zdnd11an1n64x5 FILLER_103_1230 ();
 b15zdnd11an1n08x5 FILLER_103_1294 ();
 b15zdnd11an1n04x5 FILLER_103_1302 ();
 b15zdnd00an1n01x5 FILLER_103_1306 ();
 b15zdnd11an1n04x5 FILLER_103_1310 ();
 b15zdnd11an1n04x5 FILLER_103_1317 ();
 b15zdnd11an1n04x5 FILLER_103_1324 ();
 b15zdnd11an1n64x5 FILLER_103_1331 ();
 b15zdnd11an1n64x5 FILLER_103_1395 ();
 b15zdnd11an1n64x5 FILLER_103_1459 ();
 b15zdnd11an1n64x5 FILLER_103_1523 ();
 b15zdnd11an1n64x5 FILLER_103_1587 ();
 b15zdnd11an1n64x5 FILLER_103_1651 ();
 b15zdnd11an1n64x5 FILLER_103_1715 ();
 b15zdnd11an1n64x5 FILLER_103_1779 ();
 b15zdnd11an1n64x5 FILLER_103_1843 ();
 b15zdnd11an1n64x5 FILLER_103_1907 ();
 b15zdnd11an1n64x5 FILLER_103_1971 ();
 b15zdnd11an1n64x5 FILLER_103_2035 ();
 b15zdnd11an1n64x5 FILLER_103_2099 ();
 b15zdnd11an1n64x5 FILLER_103_2163 ();
 b15zdnd11an1n32x5 FILLER_103_2227 ();
 b15zdnd11an1n16x5 FILLER_103_2259 ();
 b15zdnd11an1n08x5 FILLER_103_2275 ();
 b15zdnd00an1n01x5 FILLER_103_2283 ();
 b15zdnd11an1n64x5 FILLER_104_8 ();
 b15zdnd11an1n64x5 FILLER_104_72 ();
 b15zdnd11an1n64x5 FILLER_104_136 ();
 b15zdnd11an1n64x5 FILLER_104_200 ();
 b15zdnd11an1n64x5 FILLER_104_264 ();
 b15zdnd11an1n64x5 FILLER_104_328 ();
 b15zdnd11an1n64x5 FILLER_104_392 ();
 b15zdnd11an1n64x5 FILLER_104_456 ();
 b15zdnd11an1n64x5 FILLER_104_520 ();
 b15zdnd11an1n64x5 FILLER_104_584 ();
 b15zdnd11an1n64x5 FILLER_104_648 ();
 b15zdnd11an1n04x5 FILLER_104_712 ();
 b15zdnd00an1n02x5 FILLER_104_716 ();
 b15zdnd11an1n64x5 FILLER_104_726 ();
 b15zdnd11an1n64x5 FILLER_104_790 ();
 b15zdnd11an1n32x5 FILLER_104_854 ();
 b15zdnd11an1n16x5 FILLER_104_886 ();
 b15zdnd11an1n08x5 FILLER_104_902 ();
 b15zdnd11an1n04x5 FILLER_104_910 ();
 b15zdnd00an1n02x5 FILLER_104_914 ();
 b15zdnd00an1n01x5 FILLER_104_916 ();
 b15zdnd11an1n64x5 FILLER_104_920 ();
 b15zdnd11an1n64x5 FILLER_104_984 ();
 b15zdnd11an1n64x5 FILLER_104_1048 ();
 b15zdnd11an1n64x5 FILLER_104_1112 ();
 b15zdnd00an1n02x5 FILLER_104_1176 ();
 b15zdnd00an1n01x5 FILLER_104_1178 ();
 b15zdnd11an1n04x5 FILLER_104_1231 ();
 b15zdnd11an1n32x5 FILLER_104_1242 ();
 b15zdnd11an1n16x5 FILLER_104_1274 ();
 b15zdnd00an1n01x5 FILLER_104_1290 ();
 b15zdnd11an1n04x5 FILLER_104_1333 ();
 b15zdnd11an1n04x5 FILLER_104_1340 ();
 b15zdnd11an1n64x5 FILLER_104_1347 ();
 b15zdnd11an1n64x5 FILLER_104_1411 ();
 b15zdnd00an1n02x5 FILLER_104_1475 ();
 b15zdnd11an1n64x5 FILLER_104_1481 ();
 b15zdnd00an1n02x5 FILLER_104_1545 ();
 b15zdnd00an1n01x5 FILLER_104_1547 ();
 b15zdnd11an1n64x5 FILLER_104_1590 ();
 b15zdnd11an1n64x5 FILLER_104_1654 ();
 b15zdnd11an1n64x5 FILLER_104_1718 ();
 b15zdnd11an1n16x5 FILLER_104_1782 ();
 b15zdnd11an1n04x5 FILLER_104_1798 ();
 b15zdnd11an1n64x5 FILLER_104_1810 ();
 b15zdnd11an1n08x5 FILLER_104_1874 ();
 b15zdnd11an1n04x5 FILLER_104_1882 ();
 b15zdnd11an1n64x5 FILLER_104_1917 ();
 b15zdnd11an1n64x5 FILLER_104_1981 ();
 b15zdnd11an1n64x5 FILLER_104_2045 ();
 b15zdnd11an1n32x5 FILLER_104_2109 ();
 b15zdnd11an1n08x5 FILLER_104_2141 ();
 b15zdnd11an1n04x5 FILLER_104_2149 ();
 b15zdnd00an1n01x5 FILLER_104_2153 ();
 b15zdnd11an1n64x5 FILLER_104_2162 ();
 b15zdnd11an1n32x5 FILLER_104_2226 ();
 b15zdnd11an1n16x5 FILLER_104_2258 ();
 b15zdnd00an1n02x5 FILLER_104_2274 ();
 b15zdnd11an1n64x5 FILLER_105_0 ();
 b15zdnd11an1n64x5 FILLER_105_64 ();
 b15zdnd11an1n64x5 FILLER_105_128 ();
 b15zdnd11an1n64x5 FILLER_105_192 ();
 b15zdnd11an1n64x5 FILLER_105_256 ();
 b15zdnd11an1n64x5 FILLER_105_320 ();
 b15zdnd11an1n64x5 FILLER_105_384 ();
 b15zdnd11an1n64x5 FILLER_105_448 ();
 b15zdnd11an1n64x5 FILLER_105_512 ();
 b15zdnd11an1n64x5 FILLER_105_576 ();
 b15zdnd11an1n64x5 FILLER_105_640 ();
 b15zdnd11an1n64x5 FILLER_105_704 ();
 b15zdnd11an1n64x5 FILLER_105_768 ();
 b15zdnd11an1n04x5 FILLER_105_832 ();
 b15zdnd00an1n02x5 FILLER_105_836 ();
 b15zdnd00an1n01x5 FILLER_105_838 ();
 b15zdnd11an1n64x5 FILLER_105_851 ();
 b15zdnd11an1n64x5 FILLER_105_915 ();
 b15zdnd11an1n64x5 FILLER_105_979 ();
 b15zdnd11an1n32x5 FILLER_105_1043 ();
 b15zdnd11an1n16x5 FILLER_105_1075 ();
 b15zdnd11an1n08x5 FILLER_105_1091 ();
 b15zdnd00an1n01x5 FILLER_105_1099 ();
 b15zdnd11an1n64x5 FILLER_105_1112 ();
 b15zdnd11an1n16x5 FILLER_105_1176 ();
 b15zdnd11an1n04x5 FILLER_105_1192 ();
 b15zdnd00an1n02x5 FILLER_105_1196 ();
 b15zdnd11an1n04x5 FILLER_105_1201 ();
 b15zdnd11an1n16x5 FILLER_105_1208 ();
 b15zdnd00an1n01x5 FILLER_105_1224 ();
 b15zdnd11an1n32x5 FILLER_105_1232 ();
 b15zdnd11an1n16x5 FILLER_105_1264 ();
 b15zdnd11an1n08x5 FILLER_105_1280 ();
 b15zdnd00an1n02x5 FILLER_105_1288 ();
 b15zdnd11an1n64x5 FILLER_105_1342 ();
 b15zdnd11an1n64x5 FILLER_105_1406 ();
 b15zdnd11an1n64x5 FILLER_105_1470 ();
 b15zdnd11an1n64x5 FILLER_105_1534 ();
 b15zdnd11an1n64x5 FILLER_105_1598 ();
 b15zdnd11an1n64x5 FILLER_105_1662 ();
 b15zdnd11an1n64x5 FILLER_105_1726 ();
 b15zdnd11an1n64x5 FILLER_105_1790 ();
 b15zdnd11an1n16x5 FILLER_105_1854 ();
 b15zdnd11an1n08x5 FILLER_105_1870 ();
 b15zdnd11an1n04x5 FILLER_105_1878 ();
 b15zdnd00an1n02x5 FILLER_105_1882 ();
 b15zdnd11an1n64x5 FILLER_105_1898 ();
 b15zdnd11an1n64x5 FILLER_105_1962 ();
 b15zdnd11an1n64x5 FILLER_105_2026 ();
 b15zdnd11an1n64x5 FILLER_105_2090 ();
 b15zdnd11an1n08x5 FILLER_105_2154 ();
 b15zdnd11an1n04x5 FILLER_105_2162 ();
 b15zdnd00an1n02x5 FILLER_105_2166 ();
 b15zdnd11an1n64x5 FILLER_105_2195 ();
 b15zdnd11an1n16x5 FILLER_105_2259 ();
 b15zdnd11an1n08x5 FILLER_105_2275 ();
 b15zdnd00an1n01x5 FILLER_105_2283 ();
 b15zdnd11an1n64x5 FILLER_106_8 ();
 b15zdnd11an1n64x5 FILLER_106_72 ();
 b15zdnd11an1n64x5 FILLER_106_136 ();
 b15zdnd11an1n64x5 FILLER_106_200 ();
 b15zdnd11an1n64x5 FILLER_106_264 ();
 b15zdnd11an1n64x5 FILLER_106_328 ();
 b15zdnd11an1n64x5 FILLER_106_392 ();
 b15zdnd11an1n64x5 FILLER_106_456 ();
 b15zdnd11an1n64x5 FILLER_106_520 ();
 b15zdnd11an1n64x5 FILLER_106_584 ();
 b15zdnd11an1n16x5 FILLER_106_648 ();
 b15zdnd11an1n08x5 FILLER_106_664 ();
 b15zdnd11an1n04x5 FILLER_106_672 ();
 b15zdnd00an1n02x5 FILLER_106_676 ();
 b15zdnd11an1n16x5 FILLER_106_681 ();
 b15zdnd11an1n04x5 FILLER_106_697 ();
 b15zdnd00an1n02x5 FILLER_106_701 ();
 b15zdnd00an1n02x5 FILLER_106_716 ();
 b15zdnd00an1n02x5 FILLER_106_726 ();
 b15zdnd11an1n64x5 FILLER_106_731 ();
 b15zdnd11an1n64x5 FILLER_106_795 ();
 b15zdnd11an1n64x5 FILLER_106_859 ();
 b15zdnd11an1n64x5 FILLER_106_923 ();
 b15zdnd11an1n64x5 FILLER_106_987 ();
 b15zdnd11an1n64x5 FILLER_106_1051 ();
 b15zdnd11an1n32x5 FILLER_106_1115 ();
 b15zdnd11an1n16x5 FILLER_106_1147 ();
 b15zdnd11an1n08x5 FILLER_106_1163 ();
 b15zdnd00an1n02x5 FILLER_106_1171 ();
 b15zdnd11an1n16x5 FILLER_106_1180 ();
 b15zdnd00an1n02x5 FILLER_106_1196 ();
 b15zdnd00an1n01x5 FILLER_106_1198 ();
 b15zdnd11an1n04x5 FILLER_106_1202 ();
 b15zdnd11an1n32x5 FILLER_106_1209 ();
 b15zdnd11an1n16x5 FILLER_106_1241 ();
 b15zdnd00an1n01x5 FILLER_106_1257 ();
 b15zdnd11an1n16x5 FILLER_106_1265 ();
 b15zdnd11an1n08x5 FILLER_106_1281 ();
 b15zdnd11an1n04x5 FILLER_106_1296 ();
 b15zdnd00an1n01x5 FILLER_106_1300 ();
 b15zdnd11an1n08x5 FILLER_106_1353 ();
 b15zdnd11an1n04x5 FILLER_106_1361 ();
 b15zdnd00an1n02x5 FILLER_106_1365 ();
 b15zdnd00an1n01x5 FILLER_106_1367 ();
 b15zdnd11an1n32x5 FILLER_106_1376 ();
 b15zdnd11an1n08x5 FILLER_106_1422 ();
 b15zdnd00an1n02x5 FILLER_106_1430 ();
 b15zdnd11an1n64x5 FILLER_106_1444 ();
 b15zdnd11an1n64x5 FILLER_106_1508 ();
 b15zdnd11an1n64x5 FILLER_106_1572 ();
 b15zdnd11an1n64x5 FILLER_106_1636 ();
 b15zdnd11an1n64x5 FILLER_106_1700 ();
 b15zdnd11an1n64x5 FILLER_106_1764 ();
 b15zdnd11an1n64x5 FILLER_106_1828 ();
 b15zdnd00an1n02x5 FILLER_106_1892 ();
 b15zdnd00an1n01x5 FILLER_106_1894 ();
 b15zdnd11an1n64x5 FILLER_106_1898 ();
 b15zdnd11an1n64x5 FILLER_106_1962 ();
 b15zdnd11an1n32x5 FILLER_106_2026 ();
 b15zdnd11an1n04x5 FILLER_106_2058 ();
 b15zdnd00an1n02x5 FILLER_106_2062 ();
 b15zdnd00an1n01x5 FILLER_106_2064 ();
 b15zdnd11an1n64x5 FILLER_106_2074 ();
 b15zdnd11an1n16x5 FILLER_106_2138 ();
 b15zdnd11an1n64x5 FILLER_106_2162 ();
 b15zdnd11an1n32x5 FILLER_106_2226 ();
 b15zdnd11an1n16x5 FILLER_106_2258 ();
 b15zdnd00an1n02x5 FILLER_106_2274 ();
 b15zdnd11an1n64x5 FILLER_107_0 ();
 b15zdnd11an1n64x5 FILLER_107_64 ();
 b15zdnd11an1n64x5 FILLER_107_128 ();
 b15zdnd11an1n64x5 FILLER_107_192 ();
 b15zdnd11an1n64x5 FILLER_107_256 ();
 b15zdnd11an1n64x5 FILLER_107_320 ();
 b15zdnd11an1n64x5 FILLER_107_384 ();
 b15zdnd11an1n64x5 FILLER_107_448 ();
 b15zdnd11an1n32x5 FILLER_107_512 ();
 b15zdnd11an1n08x5 FILLER_107_544 ();
 b15zdnd00an1n02x5 FILLER_107_552 ();
 b15zdnd11an1n32x5 FILLER_107_571 ();
 b15zdnd11an1n08x5 FILLER_107_603 ();
 b15zdnd11an1n64x5 FILLER_107_614 ();
 b15zdnd00an1n01x5 FILLER_107_678 ();
 b15zdnd11an1n64x5 FILLER_107_692 ();
 b15zdnd11an1n64x5 FILLER_107_756 ();
 b15zdnd11an1n64x5 FILLER_107_820 ();
 b15zdnd11an1n64x5 FILLER_107_884 ();
 b15zdnd11an1n08x5 FILLER_107_948 ();
 b15zdnd11an1n04x5 FILLER_107_956 ();
 b15zdnd11an1n32x5 FILLER_107_969 ();
 b15zdnd11an1n08x5 FILLER_107_1001 ();
 b15zdnd11an1n04x5 FILLER_107_1009 ();
 b15zdnd00an1n02x5 FILLER_107_1013 ();
 b15zdnd00an1n01x5 FILLER_107_1015 ();
 b15zdnd11an1n64x5 FILLER_107_1025 ();
 b15zdnd11an1n32x5 FILLER_107_1089 ();
 b15zdnd11an1n16x5 FILLER_107_1121 ();
 b15zdnd11an1n08x5 FILLER_107_1137 ();
 b15zdnd11an1n32x5 FILLER_107_1187 ();
 b15zdnd11an1n64x5 FILLER_107_1226 ();
 b15zdnd11an1n16x5 FILLER_107_1342 ();
 b15zdnd11an1n64x5 FILLER_107_1400 ();
 b15zdnd11an1n16x5 FILLER_107_1473 ();
 b15zdnd11an1n08x5 FILLER_107_1489 ();
 b15zdnd00an1n02x5 FILLER_107_1497 ();
 b15zdnd11an1n64x5 FILLER_107_1508 ();
 b15zdnd11an1n64x5 FILLER_107_1572 ();
 b15zdnd11an1n64x5 FILLER_107_1636 ();
 b15zdnd11an1n64x5 FILLER_107_1700 ();
 b15zdnd11an1n64x5 FILLER_107_1764 ();
 b15zdnd11an1n64x5 FILLER_107_1828 ();
 b15zdnd11an1n64x5 FILLER_107_1892 ();
 b15zdnd11an1n64x5 FILLER_107_1956 ();
 b15zdnd11an1n16x5 FILLER_107_2020 ();
 b15zdnd11an1n08x5 FILLER_107_2036 ();
 b15zdnd11an1n64x5 FILLER_107_2053 ();
 b15zdnd11an1n64x5 FILLER_107_2117 ();
 b15zdnd11an1n64x5 FILLER_107_2181 ();
 b15zdnd11an1n32x5 FILLER_107_2245 ();
 b15zdnd11an1n04x5 FILLER_107_2277 ();
 b15zdnd00an1n02x5 FILLER_107_2281 ();
 b15zdnd00an1n01x5 FILLER_107_2283 ();
 b15zdnd11an1n64x5 FILLER_108_8 ();
 b15zdnd11an1n64x5 FILLER_108_72 ();
 b15zdnd11an1n64x5 FILLER_108_136 ();
 b15zdnd11an1n64x5 FILLER_108_200 ();
 b15zdnd11an1n64x5 FILLER_108_264 ();
 b15zdnd11an1n64x5 FILLER_108_328 ();
 b15zdnd11an1n64x5 FILLER_108_392 ();
 b15zdnd11an1n64x5 FILLER_108_456 ();
 b15zdnd11an1n64x5 FILLER_108_520 ();
 b15zdnd00an1n02x5 FILLER_108_584 ();
 b15zdnd00an1n01x5 FILLER_108_586 ();
 b15zdnd11an1n32x5 FILLER_108_631 ();
 b15zdnd11an1n04x5 FILLER_108_663 ();
 b15zdnd11an1n08x5 FILLER_108_709 ();
 b15zdnd00an1n01x5 FILLER_108_717 ();
 b15zdnd11an1n64x5 FILLER_108_726 ();
 b15zdnd11an1n64x5 FILLER_108_790 ();
 b15zdnd11an1n64x5 FILLER_108_854 ();
 b15zdnd11an1n64x5 FILLER_108_918 ();
 b15zdnd11an1n64x5 FILLER_108_982 ();
 b15zdnd11an1n64x5 FILLER_108_1046 ();
 b15zdnd11an1n64x5 FILLER_108_1110 ();
 b15zdnd11an1n64x5 FILLER_108_1174 ();
 b15zdnd11an1n64x5 FILLER_108_1238 ();
 b15zdnd11an1n04x5 FILLER_108_1302 ();
 b15zdnd00an1n02x5 FILLER_108_1306 ();
 b15zdnd00an1n01x5 FILLER_108_1308 ();
 b15zdnd11an1n04x5 FILLER_108_1312 ();
 b15zdnd11an1n32x5 FILLER_108_1319 ();
 b15zdnd11an1n08x5 FILLER_108_1351 ();
 b15zdnd11an1n04x5 FILLER_108_1359 ();
 b15zdnd11an1n64x5 FILLER_108_1370 ();
 b15zdnd11an1n64x5 FILLER_108_1434 ();
 b15zdnd11an1n64x5 FILLER_108_1498 ();
 b15zdnd11an1n64x5 FILLER_108_1562 ();
 b15zdnd11an1n64x5 FILLER_108_1626 ();
 b15zdnd11an1n64x5 FILLER_108_1690 ();
 b15zdnd11an1n32x5 FILLER_108_1754 ();
 b15zdnd11an1n08x5 FILLER_108_1786 ();
 b15zdnd11an1n04x5 FILLER_108_1794 ();
 b15zdnd00an1n02x5 FILLER_108_1798 ();
 b15zdnd11an1n04x5 FILLER_108_1816 ();
 b15zdnd00an1n02x5 FILLER_108_1820 ();
 b15zdnd11an1n16x5 FILLER_108_1839 ();
 b15zdnd11an1n08x5 FILLER_108_1855 ();
 b15zdnd11an1n04x5 FILLER_108_1863 ();
 b15zdnd00an1n02x5 FILLER_108_1867 ();
 b15zdnd11an1n04x5 FILLER_108_1883 ();
 b15zdnd11an1n64x5 FILLER_108_1890 ();
 b15zdnd11an1n64x5 FILLER_108_1954 ();
 b15zdnd11an1n64x5 FILLER_108_2018 ();
 b15zdnd11an1n64x5 FILLER_108_2082 ();
 b15zdnd11an1n08x5 FILLER_108_2146 ();
 b15zdnd11an1n64x5 FILLER_108_2162 ();
 b15zdnd11an1n32x5 FILLER_108_2226 ();
 b15zdnd11an1n16x5 FILLER_108_2258 ();
 b15zdnd00an1n02x5 FILLER_108_2274 ();
 b15zdnd11an1n64x5 FILLER_109_0 ();
 b15zdnd11an1n64x5 FILLER_109_64 ();
 b15zdnd11an1n32x5 FILLER_109_128 ();
 b15zdnd11an1n08x5 FILLER_109_160 ();
 b15zdnd11an1n04x5 FILLER_109_168 ();
 b15zdnd00an1n02x5 FILLER_109_172 ();
 b15zdnd00an1n01x5 FILLER_109_174 ();
 b15zdnd11an1n04x5 FILLER_109_178 ();
 b15zdnd11an1n04x5 FILLER_109_185 ();
 b15zdnd00an1n01x5 FILLER_109_189 ();
 b15zdnd11an1n64x5 FILLER_109_193 ();
 b15zdnd11an1n64x5 FILLER_109_257 ();
 b15zdnd11an1n64x5 FILLER_109_321 ();
 b15zdnd11an1n32x5 FILLER_109_385 ();
 b15zdnd00an1n02x5 FILLER_109_417 ();
 b15zdnd11an1n64x5 FILLER_109_428 ();
 b15zdnd11an1n64x5 FILLER_109_492 ();
 b15zdnd11an1n32x5 FILLER_109_556 ();
 b15zdnd11an1n08x5 FILLER_109_588 ();
 b15zdnd11an1n04x5 FILLER_109_596 ();
 b15zdnd00an1n02x5 FILLER_109_600 ();
 b15zdnd00an1n01x5 FILLER_109_602 ();
 b15zdnd11an1n04x5 FILLER_109_606 ();
 b15zdnd11an1n64x5 FILLER_109_613 ();
 b15zdnd11an1n32x5 FILLER_109_677 ();
 b15zdnd11an1n04x5 FILLER_109_709 ();
 b15zdnd00an1n01x5 FILLER_109_713 ();
 b15zdnd11an1n64x5 FILLER_109_745 ();
 b15zdnd00an1n01x5 FILLER_109_809 ();
 b15zdnd11an1n64x5 FILLER_109_822 ();
 b15zdnd11an1n64x5 FILLER_109_886 ();
 b15zdnd11an1n32x5 FILLER_109_950 ();
 b15zdnd11an1n16x5 FILLER_109_982 ();
 b15zdnd11an1n64x5 FILLER_109_1007 ();
 b15zdnd00an1n02x5 FILLER_109_1071 ();
 b15zdnd00an1n01x5 FILLER_109_1073 ();
 b15zdnd11an1n64x5 FILLER_109_1098 ();
 b15zdnd11an1n64x5 FILLER_109_1162 ();
 b15zdnd11an1n64x5 FILLER_109_1226 ();
 b15zdnd00an1n02x5 FILLER_109_1290 ();
 b15zdnd11an1n08x5 FILLER_109_1300 ();
 b15zdnd11an1n04x5 FILLER_109_1308 ();
 b15zdnd00an1n02x5 FILLER_109_1312 ();
 b15zdnd00an1n01x5 FILLER_109_1314 ();
 b15zdnd11an1n64x5 FILLER_109_1318 ();
 b15zdnd11an1n64x5 FILLER_109_1382 ();
 b15zdnd11an1n64x5 FILLER_109_1446 ();
 b15zdnd11an1n32x5 FILLER_109_1510 ();
 b15zdnd11an1n16x5 FILLER_109_1542 ();
 b15zdnd11an1n08x5 FILLER_109_1558 ();
 b15zdnd00an1n02x5 FILLER_109_1566 ();
 b15zdnd11an1n64x5 FILLER_109_1571 ();
 b15zdnd11an1n32x5 FILLER_109_1635 ();
 b15zdnd11an1n16x5 FILLER_109_1667 ();
 b15zdnd11an1n08x5 FILLER_109_1683 ();
 b15zdnd11an1n04x5 FILLER_109_1691 ();
 b15zdnd00an1n02x5 FILLER_109_1695 ();
 b15zdnd00an1n01x5 FILLER_109_1697 ();
 b15zdnd11an1n64x5 FILLER_109_1707 ();
 b15zdnd11an1n64x5 FILLER_109_1771 ();
 b15zdnd11an1n64x5 FILLER_109_1835 ();
 b15zdnd11an1n64x5 FILLER_109_1899 ();
 b15zdnd11an1n64x5 FILLER_109_1963 ();
 b15zdnd11an1n64x5 FILLER_109_2027 ();
 b15zdnd11an1n64x5 FILLER_109_2091 ();
 b15zdnd11an1n16x5 FILLER_109_2155 ();
 b15zdnd11an1n08x5 FILLER_109_2171 ();
 b15zdnd00an1n02x5 FILLER_109_2179 ();
 b15zdnd00an1n01x5 FILLER_109_2181 ();
 b15zdnd11an1n08x5 FILLER_109_2196 ();
 b15zdnd11an1n04x5 FILLER_109_2204 ();
 b15zdnd00an1n02x5 FILLER_109_2208 ();
 b15zdnd00an1n01x5 FILLER_109_2210 ();
 b15zdnd11an1n64x5 FILLER_109_2218 ();
 b15zdnd00an1n02x5 FILLER_109_2282 ();
 b15zdnd11an1n64x5 FILLER_110_8 ();
 b15zdnd11an1n64x5 FILLER_110_72 ();
 b15zdnd11an1n08x5 FILLER_110_136 ();
 b15zdnd11an1n04x5 FILLER_110_144 ();
 b15zdnd00an1n02x5 FILLER_110_148 ();
 b15zdnd11an1n64x5 FILLER_110_202 ();
 b15zdnd11an1n64x5 FILLER_110_266 ();
 b15zdnd11an1n64x5 FILLER_110_330 ();
 b15zdnd11an1n64x5 FILLER_110_394 ();
 b15zdnd11an1n16x5 FILLER_110_458 ();
 b15zdnd11an1n08x5 FILLER_110_474 ();
 b15zdnd11an1n04x5 FILLER_110_482 ();
 b15zdnd00an1n02x5 FILLER_110_486 ();
 b15zdnd11an1n64x5 FILLER_110_492 ();
 b15zdnd11an1n64x5 FILLER_110_556 ();
 b15zdnd11an1n64x5 FILLER_110_620 ();
 b15zdnd11an1n16x5 FILLER_110_684 ();
 b15zdnd00an1n02x5 FILLER_110_716 ();
 b15zdnd11an1n64x5 FILLER_110_726 ();
 b15zdnd11an1n16x5 FILLER_110_790 ();
 b15zdnd11an1n04x5 FILLER_110_806 ();
 b15zdnd00an1n02x5 FILLER_110_810 ();
 b15zdnd11an1n64x5 FILLER_110_832 ();
 b15zdnd11an1n64x5 FILLER_110_896 ();
 b15zdnd11an1n64x5 FILLER_110_960 ();
 b15zdnd11an1n64x5 FILLER_110_1024 ();
 b15zdnd11an1n64x5 FILLER_110_1088 ();
 b15zdnd11an1n64x5 FILLER_110_1152 ();
 b15zdnd11an1n64x5 FILLER_110_1216 ();
 b15zdnd11an1n04x5 FILLER_110_1280 ();
 b15zdnd00an1n02x5 FILLER_110_1284 ();
 b15zdnd00an1n01x5 FILLER_110_1286 ();
 b15zdnd11an1n64x5 FILLER_110_1295 ();
 b15zdnd11an1n64x5 FILLER_110_1359 ();
 b15zdnd11an1n64x5 FILLER_110_1423 ();
 b15zdnd11an1n32x5 FILLER_110_1487 ();
 b15zdnd11an1n08x5 FILLER_110_1519 ();
 b15zdnd00an1n01x5 FILLER_110_1527 ();
 b15zdnd11an1n04x5 FILLER_110_1570 ();
 b15zdnd11an1n04x5 FILLER_110_1577 ();
 b15zdnd11an1n64x5 FILLER_110_1584 ();
 b15zdnd11an1n64x5 FILLER_110_1648 ();
 b15zdnd11an1n16x5 FILLER_110_1712 ();
 b15zdnd11an1n04x5 FILLER_110_1728 ();
 b15zdnd00an1n02x5 FILLER_110_1732 ();
 b15zdnd11an1n16x5 FILLER_110_1743 ();
 b15zdnd00an1n01x5 FILLER_110_1759 ();
 b15zdnd11an1n04x5 FILLER_110_1776 ();
 b15zdnd11an1n64x5 FILLER_110_1789 ();
 b15zdnd11an1n64x5 FILLER_110_1853 ();
 b15zdnd11an1n64x5 FILLER_110_1917 ();
 b15zdnd11an1n64x5 FILLER_110_1981 ();
 b15zdnd11an1n64x5 FILLER_110_2045 ();
 b15zdnd11an1n32x5 FILLER_110_2109 ();
 b15zdnd11an1n08x5 FILLER_110_2141 ();
 b15zdnd11an1n04x5 FILLER_110_2149 ();
 b15zdnd00an1n01x5 FILLER_110_2153 ();
 b15zdnd11an1n16x5 FILLER_110_2162 ();
 b15zdnd11an1n08x5 FILLER_110_2178 ();
 b15zdnd00an1n01x5 FILLER_110_2186 ();
 b15zdnd11an1n64x5 FILLER_110_2201 ();
 b15zdnd11an1n08x5 FILLER_110_2265 ();
 b15zdnd00an1n02x5 FILLER_110_2273 ();
 b15zdnd00an1n01x5 FILLER_110_2275 ();
 b15zdnd11an1n64x5 FILLER_111_0 ();
 b15zdnd11an1n64x5 FILLER_111_64 ();
 b15zdnd11an1n16x5 FILLER_111_128 ();
 b15zdnd00an1n02x5 FILLER_111_144 ();
 b15zdnd11an1n04x5 FILLER_111_150 ();
 b15zdnd11an1n32x5 FILLER_111_196 ();
 b15zdnd11an1n16x5 FILLER_111_228 ();
 b15zdnd11an1n04x5 FILLER_111_244 ();
 b15zdnd00an1n02x5 FILLER_111_248 ();
 b15zdnd11an1n04x5 FILLER_111_290 ();
 b15zdnd11an1n64x5 FILLER_111_297 ();
 b15zdnd11an1n32x5 FILLER_111_361 ();
 b15zdnd11an1n08x5 FILLER_111_393 ();
 b15zdnd11an1n04x5 FILLER_111_401 ();
 b15zdnd11an1n64x5 FILLER_111_414 ();
 b15zdnd11an1n64x5 FILLER_111_478 ();
 b15zdnd11an1n64x5 FILLER_111_542 ();
 b15zdnd11an1n64x5 FILLER_111_606 ();
 b15zdnd11an1n64x5 FILLER_111_670 ();
 b15zdnd11an1n64x5 FILLER_111_734 ();
 b15zdnd11an1n64x5 FILLER_111_798 ();
 b15zdnd11an1n64x5 FILLER_111_862 ();
 b15zdnd11an1n64x5 FILLER_111_926 ();
 b15zdnd11an1n64x5 FILLER_111_990 ();
 b15zdnd11an1n64x5 FILLER_111_1054 ();
 b15zdnd11an1n64x5 FILLER_111_1118 ();
 b15zdnd11an1n64x5 FILLER_111_1182 ();
 b15zdnd11an1n32x5 FILLER_111_1246 ();
 b15zdnd11an1n04x5 FILLER_111_1278 ();
 b15zdnd00an1n01x5 FILLER_111_1282 ();
 b15zdnd11an1n64x5 FILLER_111_1307 ();
 b15zdnd11an1n32x5 FILLER_111_1371 ();
 b15zdnd11an1n16x5 FILLER_111_1403 ();
 b15zdnd11an1n04x5 FILLER_111_1419 ();
 b15zdnd00an1n02x5 FILLER_111_1423 ();
 b15zdnd11an1n64x5 FILLER_111_1436 ();
 b15zdnd11an1n32x5 FILLER_111_1500 ();
 b15zdnd11an1n16x5 FILLER_111_1532 ();
 b15zdnd11an1n32x5 FILLER_111_1600 ();
 b15zdnd11an1n16x5 FILLER_111_1632 ();
 b15zdnd00an1n02x5 FILLER_111_1648 ();
 b15zdnd11an1n08x5 FILLER_111_1653 ();
 b15zdnd11an1n04x5 FILLER_111_1661 ();
 b15zdnd00an1n02x5 FILLER_111_1665 ();
 b15zdnd00an1n01x5 FILLER_111_1667 ();
 b15zdnd11an1n32x5 FILLER_111_1710 ();
 b15zdnd11an1n16x5 FILLER_111_1742 ();
 b15zdnd11an1n08x5 FILLER_111_1758 ();
 b15zdnd11an1n04x5 FILLER_111_1766 ();
 b15zdnd00an1n02x5 FILLER_111_1770 ();
 b15zdnd00an1n01x5 FILLER_111_1772 ();
 b15zdnd11an1n64x5 FILLER_111_1804 ();
 b15zdnd11an1n64x5 FILLER_111_1868 ();
 b15zdnd11an1n64x5 FILLER_111_1932 ();
 b15zdnd11an1n64x5 FILLER_111_1996 ();
 b15zdnd11an1n64x5 FILLER_111_2060 ();
 b15zdnd11an1n64x5 FILLER_111_2124 ();
 b15zdnd11an1n64x5 FILLER_111_2188 ();
 b15zdnd11an1n32x5 FILLER_111_2252 ();
 b15zdnd11an1n64x5 FILLER_112_8 ();
 b15zdnd11an1n32x5 FILLER_112_86 ();
 b15zdnd11an1n16x5 FILLER_112_118 ();
 b15zdnd11an1n04x5 FILLER_112_134 ();
 b15zdnd00an1n02x5 FILLER_112_138 ();
 b15zdnd11an1n04x5 FILLER_112_145 ();
 b15zdnd11an1n04x5 FILLER_112_158 ();
 b15zdnd00an1n01x5 FILLER_112_162 ();
 b15zdnd11an1n64x5 FILLER_112_205 ();
 b15zdnd11an1n08x5 FILLER_112_269 ();
 b15zdnd11an1n04x5 FILLER_112_277 ();
 b15zdnd00an1n01x5 FILLER_112_281 ();
 b15zdnd11an1n64x5 FILLER_112_285 ();
 b15zdnd11an1n64x5 FILLER_112_349 ();
 b15zdnd11an1n64x5 FILLER_112_413 ();
 b15zdnd11an1n64x5 FILLER_112_477 ();
 b15zdnd11an1n64x5 FILLER_112_541 ();
 b15zdnd11an1n64x5 FILLER_112_605 ();
 b15zdnd11an1n32x5 FILLER_112_669 ();
 b15zdnd11an1n16x5 FILLER_112_701 ();
 b15zdnd00an1n01x5 FILLER_112_717 ();
 b15zdnd11an1n64x5 FILLER_112_726 ();
 b15zdnd11an1n32x5 FILLER_112_790 ();
 b15zdnd00an1n01x5 FILLER_112_822 ();
 b15zdnd11an1n64x5 FILLER_112_830 ();
 b15zdnd11an1n64x5 FILLER_112_894 ();
 b15zdnd11an1n64x5 FILLER_112_958 ();
 b15zdnd11an1n64x5 FILLER_112_1022 ();
 b15zdnd11an1n64x5 FILLER_112_1086 ();
 b15zdnd11an1n64x5 FILLER_112_1150 ();
 b15zdnd11an1n64x5 FILLER_112_1214 ();
 b15zdnd11an1n64x5 FILLER_112_1278 ();
 b15zdnd11an1n64x5 FILLER_112_1342 ();
 b15zdnd11an1n16x5 FILLER_112_1406 ();
 b15zdnd11an1n08x5 FILLER_112_1422 ();
 b15zdnd11an1n04x5 FILLER_112_1430 ();
 b15zdnd11an1n32x5 FILLER_112_1446 ();
 b15zdnd00an1n02x5 FILLER_112_1478 ();
 b15zdnd00an1n01x5 FILLER_112_1480 ();
 b15zdnd11an1n32x5 FILLER_112_1490 ();
 b15zdnd11an1n16x5 FILLER_112_1522 ();
 b15zdnd11an1n08x5 FILLER_112_1538 ();
 b15zdnd00an1n02x5 FILLER_112_1546 ();
 b15zdnd11an1n16x5 FILLER_112_1600 ();
 b15zdnd11an1n08x5 FILLER_112_1616 ();
 b15zdnd11an1n04x5 FILLER_112_1624 ();
 b15zdnd11an1n64x5 FILLER_112_1680 ();
 b15zdnd11an1n08x5 FILLER_112_1744 ();
 b15zdnd00an1n02x5 FILLER_112_1752 ();
 b15zdnd11an1n08x5 FILLER_112_1765 ();
 b15zdnd00an1n02x5 FILLER_112_1773 ();
 b15zdnd00an1n01x5 FILLER_112_1775 ();
 b15zdnd11an1n64x5 FILLER_112_1779 ();
 b15zdnd11an1n08x5 FILLER_112_1843 ();
 b15zdnd11an1n04x5 FILLER_112_1851 ();
 b15zdnd11an1n64x5 FILLER_112_1875 ();
 b15zdnd11an1n64x5 FILLER_112_1939 ();
 b15zdnd11an1n64x5 FILLER_112_2003 ();
 b15zdnd11an1n64x5 FILLER_112_2067 ();
 b15zdnd11an1n16x5 FILLER_112_2131 ();
 b15zdnd11an1n04x5 FILLER_112_2147 ();
 b15zdnd00an1n02x5 FILLER_112_2151 ();
 b15zdnd00an1n01x5 FILLER_112_2153 ();
 b15zdnd11an1n64x5 FILLER_112_2162 ();
 b15zdnd11an1n32x5 FILLER_112_2226 ();
 b15zdnd11an1n16x5 FILLER_112_2258 ();
 b15zdnd00an1n02x5 FILLER_112_2274 ();
 b15zdnd11an1n64x5 FILLER_113_0 ();
 b15zdnd11an1n64x5 FILLER_113_64 ();
 b15zdnd11an1n16x5 FILLER_113_128 ();
 b15zdnd11an1n04x5 FILLER_113_157 ();
 b15zdnd00an1n02x5 FILLER_113_161 ();
 b15zdnd11an1n64x5 FILLER_113_205 ();
 b15zdnd11an1n64x5 FILLER_113_269 ();
 b15zdnd11an1n64x5 FILLER_113_333 ();
 b15zdnd11an1n64x5 FILLER_113_397 ();
 b15zdnd11an1n64x5 FILLER_113_461 ();
 b15zdnd11an1n32x5 FILLER_113_525 ();
 b15zdnd00an1n02x5 FILLER_113_557 ();
 b15zdnd11an1n64x5 FILLER_113_562 ();
 b15zdnd11an1n64x5 FILLER_113_626 ();
 b15zdnd11an1n64x5 FILLER_113_690 ();
 b15zdnd11an1n64x5 FILLER_113_754 ();
 b15zdnd11an1n64x5 FILLER_113_818 ();
 b15zdnd11an1n64x5 FILLER_113_882 ();
 b15zdnd11an1n64x5 FILLER_113_946 ();
 b15zdnd11an1n64x5 FILLER_113_1010 ();
 b15zdnd11an1n64x5 FILLER_113_1074 ();
 b15zdnd11an1n64x5 FILLER_113_1138 ();
 b15zdnd11an1n64x5 FILLER_113_1202 ();
 b15zdnd11an1n64x5 FILLER_113_1266 ();
 b15zdnd11an1n64x5 FILLER_113_1330 ();
 b15zdnd11an1n16x5 FILLER_113_1394 ();
 b15zdnd11an1n08x5 FILLER_113_1410 ();
 b15zdnd11an1n04x5 FILLER_113_1418 ();
 b15zdnd00an1n02x5 FILLER_113_1422 ();
 b15zdnd11an1n04x5 FILLER_113_1432 ();
 b15zdnd11an1n32x5 FILLER_113_1442 ();
 b15zdnd11an1n16x5 FILLER_113_1474 ();
 b15zdnd11an1n08x5 FILLER_113_1490 ();
 b15zdnd00an1n01x5 FILLER_113_1498 ();
 b15zdnd11an1n32x5 FILLER_113_1507 ();
 b15zdnd11an1n16x5 FILLER_113_1539 ();
 b15zdnd11an1n08x5 FILLER_113_1555 ();
 b15zdnd00an1n02x5 FILLER_113_1563 ();
 b15zdnd00an1n01x5 FILLER_113_1565 ();
 b15zdnd11an1n04x5 FILLER_113_1569 ();
 b15zdnd11an1n64x5 FILLER_113_1576 ();
 b15zdnd11an1n04x5 FILLER_113_1643 ();
 b15zdnd11an1n32x5 FILLER_113_1699 ();
 b15zdnd00an1n02x5 FILLER_113_1731 ();
 b15zdnd11an1n08x5 FILLER_113_1742 ();
 b15zdnd11an1n04x5 FILLER_113_1764 ();
 b15zdnd11an1n08x5 FILLER_113_1777 ();
 b15zdnd00an1n02x5 FILLER_113_1785 ();
 b15zdnd11an1n64x5 FILLER_113_1790 ();
 b15zdnd11an1n08x5 FILLER_113_1854 ();
 b15zdnd11an1n04x5 FILLER_113_1862 ();
 b15zdnd11an1n64x5 FILLER_113_1880 ();
 b15zdnd11an1n64x5 FILLER_113_1944 ();
 b15zdnd11an1n64x5 FILLER_113_2008 ();
 b15zdnd11an1n64x5 FILLER_113_2072 ();
 b15zdnd11an1n64x5 FILLER_113_2136 ();
 b15zdnd11an1n08x5 FILLER_113_2200 ();
 b15zdnd00an1n02x5 FILLER_113_2208 ();
 b15zdnd11an1n64x5 FILLER_113_2216 ();
 b15zdnd11an1n04x5 FILLER_113_2280 ();
 b15zdnd11an1n64x5 FILLER_114_8 ();
 b15zdnd11an1n64x5 FILLER_114_72 ();
 b15zdnd11an1n08x5 FILLER_114_136 ();
 b15zdnd11an1n04x5 FILLER_114_144 ();
 b15zdnd00an1n02x5 FILLER_114_148 ();
 b15zdnd11an1n64x5 FILLER_114_192 ();
 b15zdnd11an1n64x5 FILLER_114_256 ();
 b15zdnd11an1n64x5 FILLER_114_320 ();
 b15zdnd11an1n64x5 FILLER_114_384 ();
 b15zdnd11an1n64x5 FILLER_114_448 ();
 b15zdnd11an1n08x5 FILLER_114_512 ();
 b15zdnd11an1n04x5 FILLER_114_520 ();
 b15zdnd00an1n01x5 FILLER_114_524 ();
 b15zdnd11an1n16x5 FILLER_114_532 ();
 b15zdnd00an1n01x5 FILLER_114_548 ();
 b15zdnd11an1n32x5 FILLER_114_563 ();
 b15zdnd11an1n64x5 FILLER_114_603 ();
 b15zdnd11an1n32x5 FILLER_114_667 ();
 b15zdnd11an1n16x5 FILLER_114_699 ();
 b15zdnd00an1n02x5 FILLER_114_715 ();
 b15zdnd00an1n01x5 FILLER_114_717 ();
 b15zdnd11an1n64x5 FILLER_114_726 ();
 b15zdnd11an1n64x5 FILLER_114_790 ();
 b15zdnd11an1n64x5 FILLER_114_854 ();
 b15zdnd11an1n64x5 FILLER_114_918 ();
 b15zdnd11an1n64x5 FILLER_114_982 ();
 b15zdnd11an1n64x5 FILLER_114_1046 ();
 b15zdnd11an1n64x5 FILLER_114_1110 ();
 b15zdnd11an1n16x5 FILLER_114_1174 ();
 b15zdnd11an1n04x5 FILLER_114_1190 ();
 b15zdnd00an1n02x5 FILLER_114_1194 ();
 b15zdnd11an1n64x5 FILLER_114_1205 ();
 b15zdnd11an1n64x5 FILLER_114_1269 ();
 b15zdnd11an1n64x5 FILLER_114_1333 ();
 b15zdnd11an1n64x5 FILLER_114_1397 ();
 b15zdnd11an1n64x5 FILLER_114_1461 ();
 b15zdnd11an1n32x5 FILLER_114_1525 ();
 b15zdnd11an1n16x5 FILLER_114_1557 ();
 b15zdnd11an1n64x5 FILLER_114_1576 ();
 b15zdnd11an1n08x5 FILLER_114_1640 ();
 b15zdnd00an1n01x5 FILLER_114_1648 ();
 b15zdnd11an1n16x5 FILLER_114_1652 ();
 b15zdnd00an1n01x5 FILLER_114_1668 ();
 b15zdnd11an1n04x5 FILLER_114_1672 ();
 b15zdnd11an1n16x5 FILLER_114_1679 ();
 b15zdnd11an1n08x5 FILLER_114_1695 ();
 b15zdnd11an1n04x5 FILLER_114_1703 ();
 b15zdnd00an1n02x5 FILLER_114_1707 ();
 b15zdnd11an1n32x5 FILLER_114_1751 ();
 b15zdnd11an1n04x5 FILLER_114_1783 ();
 b15zdnd11an1n16x5 FILLER_114_1795 ();
 b15zdnd11an1n32x5 FILLER_114_1827 ();
 b15zdnd11an1n16x5 FILLER_114_1859 ();
 b15zdnd00an1n02x5 FILLER_114_1875 ();
 b15zdnd00an1n01x5 FILLER_114_1877 ();
 b15zdnd11an1n04x5 FILLER_114_1881 ();
 b15zdnd11an1n64x5 FILLER_114_1888 ();
 b15zdnd11an1n64x5 FILLER_114_1952 ();
 b15zdnd11an1n16x5 FILLER_114_2016 ();
 b15zdnd11an1n08x5 FILLER_114_2032 ();
 b15zdnd11an1n04x5 FILLER_114_2040 ();
 b15zdnd00an1n02x5 FILLER_114_2044 ();
 b15zdnd00an1n01x5 FILLER_114_2046 ();
 b15zdnd11an1n64x5 FILLER_114_2050 ();
 b15zdnd11an1n32x5 FILLER_114_2114 ();
 b15zdnd11an1n08x5 FILLER_114_2146 ();
 b15zdnd11an1n64x5 FILLER_114_2162 ();
 b15zdnd11an1n32x5 FILLER_114_2226 ();
 b15zdnd11an1n16x5 FILLER_114_2258 ();
 b15zdnd00an1n02x5 FILLER_114_2274 ();
 b15zdnd11an1n64x5 FILLER_115_0 ();
 b15zdnd11an1n64x5 FILLER_115_64 ();
 b15zdnd11an1n16x5 FILLER_115_128 ();
 b15zdnd11an1n04x5 FILLER_115_144 ();
 b15zdnd00an1n02x5 FILLER_115_148 ();
 b15zdnd11an1n04x5 FILLER_115_160 ();
 b15zdnd00an1n01x5 FILLER_115_164 ();
 b15zdnd11an1n08x5 FILLER_115_170 ();
 b15zdnd00an1n01x5 FILLER_115_178 ();
 b15zdnd11an1n64x5 FILLER_115_183 ();
 b15zdnd11an1n64x5 FILLER_115_247 ();
 b15zdnd11an1n64x5 FILLER_115_311 ();
 b15zdnd11an1n64x5 FILLER_115_375 ();
 b15zdnd11an1n64x5 FILLER_115_439 ();
 b15zdnd11an1n32x5 FILLER_115_503 ();
 b15zdnd11an1n16x5 FILLER_115_535 ();
 b15zdnd11an1n64x5 FILLER_115_554 ();
 b15zdnd11an1n04x5 FILLER_115_618 ();
 b15zdnd00an1n02x5 FILLER_115_622 ();
 b15zdnd11an1n04x5 FILLER_115_652 ();
 b15zdnd11an1n64x5 FILLER_115_659 ();
 b15zdnd11an1n64x5 FILLER_115_723 ();
 b15zdnd11an1n64x5 FILLER_115_787 ();
 b15zdnd11an1n32x5 FILLER_115_851 ();
 b15zdnd11an1n16x5 FILLER_115_883 ();
 b15zdnd11an1n08x5 FILLER_115_899 ();
 b15zdnd11an1n04x5 FILLER_115_907 ();
 b15zdnd00an1n01x5 FILLER_115_911 ();
 b15zdnd11an1n04x5 FILLER_115_915 ();
 b15zdnd11an1n64x5 FILLER_115_922 ();
 b15zdnd11an1n32x5 FILLER_115_986 ();
 b15zdnd11an1n16x5 FILLER_115_1018 ();
 b15zdnd11an1n08x5 FILLER_115_1034 ();
 b15zdnd00an1n02x5 FILLER_115_1042 ();
 b15zdnd11an1n64x5 FILLER_115_1047 ();
 b15zdnd11an1n64x5 FILLER_115_1111 ();
 b15zdnd11an1n64x5 FILLER_115_1175 ();
 b15zdnd11an1n64x5 FILLER_115_1239 ();
 b15zdnd11an1n64x5 FILLER_115_1303 ();
 b15zdnd11an1n64x5 FILLER_115_1367 ();
 b15zdnd11an1n64x5 FILLER_115_1431 ();
 b15zdnd11an1n64x5 FILLER_115_1495 ();
 b15zdnd11an1n64x5 FILLER_115_1559 ();
 b15zdnd00an1n02x5 FILLER_115_1623 ();
 b15zdnd00an1n01x5 FILLER_115_1625 ();
 b15zdnd11an1n32x5 FILLER_115_1633 ();
 b15zdnd11an1n04x5 FILLER_115_1665 ();
 b15zdnd00an1n01x5 FILLER_115_1669 ();
 b15zdnd11an1n64x5 FILLER_115_1673 ();
 b15zdnd11an1n32x5 FILLER_115_1737 ();
 b15zdnd11an1n08x5 FILLER_115_1769 ();
 b15zdnd00an1n02x5 FILLER_115_1777 ();
 b15zdnd00an1n01x5 FILLER_115_1779 ();
 b15zdnd11an1n04x5 FILLER_115_1822 ();
 b15zdnd11an1n08x5 FILLER_115_1868 ();
 b15zdnd00an1n02x5 FILLER_115_1876 ();
 b15zdnd00an1n01x5 FILLER_115_1878 ();
 b15zdnd11an1n64x5 FILLER_115_1893 ();
 b15zdnd11an1n64x5 FILLER_115_1957 ();
 b15zdnd11an1n16x5 FILLER_115_2021 ();
 b15zdnd11an1n08x5 FILLER_115_2037 ();
 b15zdnd00an1n01x5 FILLER_115_2045 ();
 b15zdnd11an1n04x5 FILLER_115_2049 ();
 b15zdnd11an1n64x5 FILLER_115_2056 ();
 b15zdnd11an1n64x5 FILLER_115_2120 ();
 b15zdnd11an1n64x5 FILLER_115_2184 ();
 b15zdnd11an1n32x5 FILLER_115_2248 ();
 b15zdnd11an1n04x5 FILLER_115_2280 ();
 b15zdnd11an1n64x5 FILLER_116_8 ();
 b15zdnd11an1n64x5 FILLER_116_72 ();
 b15zdnd11an1n08x5 FILLER_116_136 ();
 b15zdnd00an1n02x5 FILLER_116_144 ();
 b15zdnd00an1n01x5 FILLER_116_146 ();
 b15zdnd11an1n64x5 FILLER_116_152 ();
 b15zdnd11an1n32x5 FILLER_116_216 ();
 b15zdnd11an1n16x5 FILLER_116_248 ();
 b15zdnd11an1n08x5 FILLER_116_264 ();
 b15zdnd11an1n04x5 FILLER_116_272 ();
 b15zdnd00an1n01x5 FILLER_116_276 ();
 b15zdnd11an1n64x5 FILLER_116_291 ();
 b15zdnd11an1n64x5 FILLER_116_355 ();
 b15zdnd00an1n02x5 FILLER_116_419 ();
 b15zdnd00an1n01x5 FILLER_116_421 ();
 b15zdnd11an1n64x5 FILLER_116_425 ();
 b15zdnd11an1n32x5 FILLER_116_489 ();
 b15zdnd11an1n16x5 FILLER_116_521 ();
 b15zdnd11an1n08x5 FILLER_116_537 ();
 b15zdnd00an1n02x5 FILLER_116_545 ();
 b15zdnd00an1n01x5 FILLER_116_547 ();
 b15zdnd11an1n64x5 FILLER_116_561 ();
 b15zdnd11an1n16x5 FILLER_116_625 ();
 b15zdnd11an1n04x5 FILLER_116_641 ();
 b15zdnd00an1n01x5 FILLER_116_645 ();
 b15zdnd11an1n64x5 FILLER_116_649 ();
 b15zdnd11an1n04x5 FILLER_116_713 ();
 b15zdnd00an1n01x5 FILLER_116_717 ();
 b15zdnd11an1n64x5 FILLER_116_726 ();
 b15zdnd11an1n32x5 FILLER_116_790 ();
 b15zdnd11an1n16x5 FILLER_116_822 ();
 b15zdnd11an1n32x5 FILLER_116_850 ();
 b15zdnd11an1n04x5 FILLER_116_882 ();
 b15zdnd00an1n02x5 FILLER_116_886 ();
 b15zdnd00an1n01x5 FILLER_116_888 ();
 b15zdnd11an1n64x5 FILLER_116_941 ();
 b15zdnd11an1n32x5 FILLER_116_1005 ();
 b15zdnd11an1n04x5 FILLER_116_1037 ();
 b15zdnd00an1n02x5 FILLER_116_1041 ();
 b15zdnd00an1n01x5 FILLER_116_1043 ();
 b15zdnd11an1n04x5 FILLER_116_1047 ();
 b15zdnd11an1n16x5 FILLER_116_1054 ();
 b15zdnd11an1n04x5 FILLER_116_1070 ();
 b15zdnd00an1n02x5 FILLER_116_1074 ();
 b15zdnd11an1n04x5 FILLER_116_1079 ();
 b15zdnd11an1n64x5 FILLER_116_1086 ();
 b15zdnd11an1n64x5 FILLER_116_1150 ();
 b15zdnd11an1n64x5 FILLER_116_1214 ();
 b15zdnd11an1n64x5 FILLER_116_1278 ();
 b15zdnd11an1n64x5 FILLER_116_1342 ();
 b15zdnd11an1n16x5 FILLER_116_1406 ();
 b15zdnd11an1n08x5 FILLER_116_1422 ();
 b15zdnd11an1n04x5 FILLER_116_1430 ();
 b15zdnd00an1n02x5 FILLER_116_1434 ();
 b15zdnd00an1n01x5 FILLER_116_1436 ();
 b15zdnd11an1n16x5 FILLER_116_1449 ();
 b15zdnd00an1n02x5 FILLER_116_1465 ();
 b15zdnd11an1n64x5 FILLER_116_1479 ();
 b15zdnd11an1n32x5 FILLER_116_1543 ();
 b15zdnd11an1n16x5 FILLER_116_1575 ();
 b15zdnd11an1n08x5 FILLER_116_1591 ();
 b15zdnd11an1n64x5 FILLER_116_1608 ();
 b15zdnd11an1n64x5 FILLER_116_1672 ();
 b15zdnd11an1n64x5 FILLER_116_1736 ();
 b15zdnd11an1n64x5 FILLER_116_1800 ();
 b15zdnd11an1n16x5 FILLER_116_1864 ();
 b15zdnd11an1n04x5 FILLER_116_1880 ();
 b15zdnd00an1n02x5 FILLER_116_1884 ();
 b15zdnd00an1n01x5 FILLER_116_1886 ();
 b15zdnd11an1n64x5 FILLER_116_1929 ();
 b15zdnd11an1n32x5 FILLER_116_1993 ();
 b15zdnd00an1n02x5 FILLER_116_2025 ();
 b15zdnd11an1n64x5 FILLER_116_2079 ();
 b15zdnd11an1n08x5 FILLER_116_2143 ();
 b15zdnd00an1n02x5 FILLER_116_2151 ();
 b15zdnd00an1n01x5 FILLER_116_2153 ();
 b15zdnd11an1n32x5 FILLER_116_2162 ();
 b15zdnd11an1n08x5 FILLER_116_2194 ();
 b15zdnd11an1n04x5 FILLER_116_2202 ();
 b15zdnd00an1n02x5 FILLER_116_2206 ();
 b15zdnd11an1n32x5 FILLER_116_2227 ();
 b15zdnd11an1n16x5 FILLER_116_2259 ();
 b15zdnd00an1n01x5 FILLER_116_2275 ();
 b15zdnd11an1n64x5 FILLER_117_0 ();
 b15zdnd11an1n64x5 FILLER_117_64 ();
 b15zdnd11an1n64x5 FILLER_117_128 ();
 b15zdnd11an1n64x5 FILLER_117_192 ();
 b15zdnd11an1n64x5 FILLER_117_256 ();
 b15zdnd11an1n64x5 FILLER_117_320 ();
 b15zdnd11an1n32x5 FILLER_117_384 ();
 b15zdnd11an1n04x5 FILLER_117_416 ();
 b15zdnd00an1n02x5 FILLER_117_420 ();
 b15zdnd11an1n04x5 FILLER_117_425 ();
 b15zdnd11an1n64x5 FILLER_117_432 ();
 b15zdnd11an1n64x5 FILLER_117_496 ();
 b15zdnd11an1n64x5 FILLER_117_560 ();
 b15zdnd11an1n64x5 FILLER_117_624 ();
 b15zdnd11an1n64x5 FILLER_117_688 ();
 b15zdnd11an1n64x5 FILLER_117_752 ();
 b15zdnd11an1n16x5 FILLER_117_816 ();
 b15zdnd11an1n04x5 FILLER_117_832 ();
 b15zdnd00an1n01x5 FILLER_117_836 ();
 b15zdnd11an1n08x5 FILLER_117_844 ();
 b15zdnd00an1n02x5 FILLER_117_852 ();
 b15zdnd11an1n04x5 FILLER_117_862 ();
 b15zdnd11an1n16x5 FILLER_117_890 ();
 b15zdnd11an1n08x5 FILLER_117_906 ();
 b15zdnd11an1n04x5 FILLER_117_914 ();
 b15zdnd00an1n01x5 FILLER_117_918 ();
 b15zdnd11an1n64x5 FILLER_117_922 ();
 b15zdnd11an1n32x5 FILLER_117_986 ();
 b15zdnd11an1n08x5 FILLER_117_1018 ();
 b15zdnd11an1n16x5 FILLER_117_1078 ();
 b15zdnd11an1n64x5 FILLER_117_1102 ();
 b15zdnd11an1n64x5 FILLER_117_1166 ();
 b15zdnd11an1n64x5 FILLER_117_1230 ();
 b15zdnd11an1n64x5 FILLER_117_1294 ();
 b15zdnd11an1n64x5 FILLER_117_1358 ();
 b15zdnd11an1n08x5 FILLER_117_1422 ();
 b15zdnd00an1n02x5 FILLER_117_1430 ();
 b15zdnd11an1n64x5 FILLER_117_1449 ();
 b15zdnd11an1n64x5 FILLER_117_1513 ();
 b15zdnd11an1n64x5 FILLER_117_1577 ();
 b15zdnd11an1n64x5 FILLER_117_1641 ();
 b15zdnd11an1n64x5 FILLER_117_1705 ();
 b15zdnd11an1n64x5 FILLER_117_1769 ();
 b15zdnd11an1n64x5 FILLER_117_1833 ();
 b15zdnd11an1n32x5 FILLER_117_1897 ();
 b15zdnd00an1n02x5 FILLER_117_1929 ();
 b15zdnd11an1n64x5 FILLER_117_1935 ();
 b15zdnd11an1n32x5 FILLER_117_1999 ();
 b15zdnd11an1n16x5 FILLER_117_2031 ();
 b15zdnd11an1n04x5 FILLER_117_2047 ();
 b15zdnd00an1n02x5 FILLER_117_2051 ();
 b15zdnd11an1n04x5 FILLER_117_2056 ();
 b15zdnd11an1n04x5 FILLER_117_2063 ();
 b15zdnd11an1n04x5 FILLER_117_2070 ();
 b15zdnd11an1n04x5 FILLER_117_2077 ();
 b15zdnd11an1n64x5 FILLER_117_2088 ();
 b15zdnd11an1n64x5 FILLER_117_2152 ();
 b15zdnd11an1n64x5 FILLER_117_2216 ();
 b15zdnd11an1n04x5 FILLER_117_2280 ();
 b15zdnd11an1n64x5 FILLER_118_8 ();
 b15zdnd11an1n64x5 FILLER_118_72 ();
 b15zdnd11an1n64x5 FILLER_118_136 ();
 b15zdnd11an1n64x5 FILLER_118_200 ();
 b15zdnd11an1n64x5 FILLER_118_264 ();
 b15zdnd11an1n64x5 FILLER_118_328 ();
 b15zdnd11an1n08x5 FILLER_118_392 ();
 b15zdnd00an1n02x5 FILLER_118_400 ();
 b15zdnd11an1n04x5 FILLER_118_454 ();
 b15zdnd11an1n64x5 FILLER_118_461 ();
 b15zdnd11an1n64x5 FILLER_118_525 ();
 b15zdnd11an1n64x5 FILLER_118_589 ();
 b15zdnd11an1n64x5 FILLER_118_653 ();
 b15zdnd00an1n01x5 FILLER_118_717 ();
 b15zdnd11an1n64x5 FILLER_118_726 ();
 b15zdnd11an1n64x5 FILLER_118_790 ();
 b15zdnd11an1n16x5 FILLER_118_854 ();
 b15zdnd00an1n02x5 FILLER_118_870 ();
 b15zdnd00an1n01x5 FILLER_118_872 ();
 b15zdnd11an1n64x5 FILLER_118_887 ();
 b15zdnd11an1n64x5 FILLER_118_951 ();
 b15zdnd11an1n32x5 FILLER_118_1015 ();
 b15zdnd11an1n04x5 FILLER_118_1047 ();
 b15zdnd00an1n02x5 FILLER_118_1051 ();
 b15zdnd00an1n01x5 FILLER_118_1053 ();
 b15zdnd11an1n64x5 FILLER_118_1106 ();
 b15zdnd11an1n16x5 FILLER_118_1170 ();
 b15zdnd00an1n02x5 FILLER_118_1186 ();
 b15zdnd00an1n01x5 FILLER_118_1188 ();
 b15zdnd11an1n64x5 FILLER_118_1197 ();
 b15zdnd11an1n08x5 FILLER_118_1261 ();
 b15zdnd00an1n02x5 FILLER_118_1269 ();
 b15zdnd00an1n01x5 FILLER_118_1271 ();
 b15zdnd11an1n64x5 FILLER_118_1288 ();
 b15zdnd11an1n64x5 FILLER_118_1352 ();
 b15zdnd11an1n16x5 FILLER_118_1416 ();
 b15zdnd11an1n64x5 FILLER_118_1450 ();
 b15zdnd11an1n64x5 FILLER_118_1514 ();
 b15zdnd11an1n64x5 FILLER_118_1578 ();
 b15zdnd11an1n64x5 FILLER_118_1642 ();
 b15zdnd11an1n64x5 FILLER_118_1706 ();
 b15zdnd11an1n64x5 FILLER_118_1770 ();
 b15zdnd11an1n16x5 FILLER_118_1834 ();
 b15zdnd11an1n08x5 FILLER_118_1850 ();
 b15zdnd11an1n08x5 FILLER_118_1870 ();
 b15zdnd11an1n04x5 FILLER_118_1878 ();
 b15zdnd00an1n01x5 FILLER_118_1882 ();
 b15zdnd11an1n04x5 FILLER_118_1886 ();
 b15zdnd00an1n02x5 FILLER_118_1890 ();
 b15zdnd00an1n01x5 FILLER_118_1892 ();
 b15zdnd11an1n64x5 FILLER_118_1896 ();
 b15zdnd11an1n64x5 FILLER_118_1960 ();
 b15zdnd11an1n08x5 FILLER_118_2024 ();
 b15zdnd00an1n02x5 FILLER_118_2032 ();
 b15zdnd11an1n04x5 FILLER_118_2086 ();
 b15zdnd11an1n32x5 FILLER_118_2093 ();
 b15zdnd11an1n16x5 FILLER_118_2125 ();
 b15zdnd11an1n08x5 FILLER_118_2141 ();
 b15zdnd11an1n04x5 FILLER_118_2149 ();
 b15zdnd00an1n01x5 FILLER_118_2153 ();
 b15zdnd11an1n32x5 FILLER_118_2162 ();
 b15zdnd11an1n16x5 FILLER_118_2194 ();
 b15zdnd00an1n02x5 FILLER_118_2210 ();
 b15zdnd00an1n01x5 FILLER_118_2212 ();
 b15zdnd11an1n04x5 FILLER_118_2218 ();
 b15zdnd11an1n04x5 FILLER_118_2225 ();
 b15zdnd00an1n02x5 FILLER_118_2274 ();
 b15zdnd11an1n64x5 FILLER_119_0 ();
 b15zdnd11an1n64x5 FILLER_119_64 ();
 b15zdnd11an1n16x5 FILLER_119_128 ();
 b15zdnd11an1n04x5 FILLER_119_144 ();
 b15zdnd11an1n64x5 FILLER_119_151 ();
 b15zdnd11an1n64x5 FILLER_119_215 ();
 b15zdnd11an1n64x5 FILLER_119_279 ();
 b15zdnd11an1n08x5 FILLER_119_343 ();
 b15zdnd11an1n04x5 FILLER_119_351 ();
 b15zdnd00an1n02x5 FILLER_119_355 ();
 b15zdnd11an1n08x5 FILLER_119_409 ();
 b15zdnd11an1n04x5 FILLER_119_417 ();
 b15zdnd11an1n04x5 FILLER_119_424 ();
 b15zdnd11an1n32x5 FILLER_119_480 ();
 b15zdnd11an1n16x5 FILLER_119_512 ();
 b15zdnd11an1n08x5 FILLER_119_528 ();
 b15zdnd11an1n04x5 FILLER_119_536 ();
 b15zdnd00an1n02x5 FILLER_119_540 ();
 b15zdnd00an1n01x5 FILLER_119_542 ();
 b15zdnd11an1n64x5 FILLER_119_560 ();
 b15zdnd11an1n32x5 FILLER_119_624 ();
 b15zdnd11an1n16x5 FILLER_119_656 ();
 b15zdnd11an1n08x5 FILLER_119_672 ();
 b15zdnd00an1n02x5 FILLER_119_680 ();
 b15zdnd11an1n16x5 FILLER_119_713 ();
 b15zdnd11an1n08x5 FILLER_119_729 ();
 b15zdnd00an1n02x5 FILLER_119_737 ();
 b15zdnd11an1n64x5 FILLER_119_742 ();
 b15zdnd11an1n16x5 FILLER_119_806 ();
 b15zdnd00an1n02x5 FILLER_119_822 ();
 b15zdnd11an1n64x5 FILLER_119_844 ();
 b15zdnd11an1n04x5 FILLER_119_908 ();
 b15zdnd11an1n04x5 FILLER_119_915 ();
 b15zdnd00an1n02x5 FILLER_119_919 ();
 b15zdnd11an1n64x5 FILLER_119_924 ();
 b15zdnd11an1n16x5 FILLER_119_988 ();
 b15zdnd11an1n08x5 FILLER_119_1004 ();
 b15zdnd11an1n04x5 FILLER_119_1012 ();
 b15zdnd00an1n02x5 FILLER_119_1016 ();
 b15zdnd00an1n01x5 FILLER_119_1018 ();
 b15zdnd11an1n04x5 FILLER_119_1071 ();
 b15zdnd00an1n02x5 FILLER_119_1075 ();
 b15zdnd11an1n64x5 FILLER_119_1080 ();
 b15zdnd11an1n08x5 FILLER_119_1144 ();
 b15zdnd00an1n02x5 FILLER_119_1152 ();
 b15zdnd00an1n01x5 FILLER_119_1154 ();
 b15zdnd11an1n16x5 FILLER_119_1158 ();
 b15zdnd00an1n01x5 FILLER_119_1174 ();
 b15zdnd11an1n64x5 FILLER_119_1202 ();
 b15zdnd11an1n64x5 FILLER_119_1266 ();
 b15zdnd11an1n32x5 FILLER_119_1330 ();
 b15zdnd11an1n16x5 FILLER_119_1362 ();
 b15zdnd11an1n04x5 FILLER_119_1378 ();
 b15zdnd00an1n02x5 FILLER_119_1382 ();
 b15zdnd11an1n32x5 FILLER_119_1404 ();
 b15zdnd11an1n08x5 FILLER_119_1436 ();
 b15zdnd11an1n04x5 FILLER_119_1444 ();
 b15zdnd00an1n01x5 FILLER_119_1448 ();
 b15zdnd11an1n64x5 FILLER_119_1456 ();
 b15zdnd11an1n64x5 FILLER_119_1520 ();
 b15zdnd11an1n64x5 FILLER_119_1584 ();
 b15zdnd11an1n64x5 FILLER_119_1648 ();
 b15zdnd11an1n32x5 FILLER_119_1712 ();
 b15zdnd11an1n16x5 FILLER_119_1744 ();
 b15zdnd11an1n04x5 FILLER_119_1760 ();
 b15zdnd00an1n02x5 FILLER_119_1764 ();
 b15zdnd00an1n01x5 FILLER_119_1766 ();
 b15zdnd11an1n16x5 FILLER_119_1781 ();
 b15zdnd11an1n08x5 FILLER_119_1797 ();
 b15zdnd00an1n01x5 FILLER_119_1805 ();
 b15zdnd11an1n32x5 FILLER_119_1827 ();
 b15zdnd11an1n04x5 FILLER_119_1859 ();
 b15zdnd11an1n32x5 FILLER_119_1907 ();
 b15zdnd11an1n16x5 FILLER_119_1939 ();
 b15zdnd11an1n08x5 FILLER_119_1955 ();
 b15zdnd11an1n04x5 FILLER_119_1963 ();
 b15zdnd11an1n64x5 FILLER_119_1971 ();
 b15zdnd11an1n04x5 FILLER_119_2035 ();
 b15zdnd00an1n01x5 FILLER_119_2039 ();
 b15zdnd11an1n64x5 FILLER_119_2092 ();
 b15zdnd11an1n32x5 FILLER_119_2156 ();
 b15zdnd11an1n08x5 FILLER_119_2188 ();
 b15zdnd00an1n02x5 FILLER_119_2196 ();
 b15zdnd00an1n01x5 FILLER_119_2198 ();
 b15zdnd11an1n16x5 FILLER_119_2251 ();
 b15zdnd00an1n02x5 FILLER_119_2267 ();
 b15zdnd00an1n01x5 FILLER_119_2269 ();
 b15zdnd11an1n08x5 FILLER_119_2274 ();
 b15zdnd00an1n02x5 FILLER_119_2282 ();
 b15zdnd11an1n64x5 FILLER_120_8 ();
 b15zdnd11an1n64x5 FILLER_120_72 ();
 b15zdnd11an1n64x5 FILLER_120_136 ();
 b15zdnd11an1n64x5 FILLER_120_200 ();
 b15zdnd11an1n32x5 FILLER_120_264 ();
 b15zdnd00an1n01x5 FILLER_120_296 ();
 b15zdnd11an1n04x5 FILLER_120_301 ();
 b15zdnd00an1n02x5 FILLER_120_305 ();
 b15zdnd00an1n01x5 FILLER_120_307 ();
 b15zdnd11an1n64x5 FILLER_120_312 ();
 b15zdnd00an1n01x5 FILLER_120_376 ();
 b15zdnd11an1n04x5 FILLER_120_380 ();
 b15zdnd11an1n64x5 FILLER_120_387 ();
 b15zdnd11an1n64x5 FILLER_120_451 ();
 b15zdnd11an1n32x5 FILLER_120_515 ();
 b15zdnd11an1n08x5 FILLER_120_547 ();
 b15zdnd11an1n04x5 FILLER_120_555 ();
 b15zdnd00an1n01x5 FILLER_120_559 ();
 b15zdnd11an1n04x5 FILLER_120_576 ();
 b15zdnd00an1n02x5 FILLER_120_580 ();
 b15zdnd11an1n64x5 FILLER_120_585 ();
 b15zdnd11an1n64x5 FILLER_120_649 ();
 b15zdnd11an1n04x5 FILLER_120_713 ();
 b15zdnd00an1n01x5 FILLER_120_717 ();
 b15zdnd00an1n02x5 FILLER_120_726 ();
 b15zdnd00an1n01x5 FILLER_120_728 ();
 b15zdnd11an1n64x5 FILLER_120_743 ();
 b15zdnd11an1n64x5 FILLER_120_807 ();
 b15zdnd11an1n16x5 FILLER_120_871 ();
 b15zdnd00an1n02x5 FILLER_120_887 ();
 b15zdnd11an1n64x5 FILLER_120_941 ();
 b15zdnd11an1n32x5 FILLER_120_1005 ();
 b15zdnd11an1n04x5 FILLER_120_1037 ();
 b15zdnd00an1n01x5 FILLER_120_1041 ();
 b15zdnd11an1n04x5 FILLER_120_1045 ();
 b15zdnd11an1n04x5 FILLER_120_1052 ();
 b15zdnd11an1n64x5 FILLER_120_1059 ();
 b15zdnd11an1n32x5 FILLER_120_1123 ();
 b15zdnd11an1n16x5 FILLER_120_1155 ();
 b15zdnd11an1n08x5 FILLER_120_1171 ();
 b15zdnd00an1n02x5 FILLER_120_1179 ();
 b15zdnd00an1n01x5 FILLER_120_1181 ();
 b15zdnd11an1n64x5 FILLER_120_1194 ();
 b15zdnd11an1n32x5 FILLER_120_1258 ();
 b15zdnd11an1n08x5 FILLER_120_1290 ();
 b15zdnd11an1n64x5 FILLER_120_1304 ();
 b15zdnd11an1n64x5 FILLER_120_1368 ();
 b15zdnd11an1n64x5 FILLER_120_1432 ();
 b15zdnd11an1n64x5 FILLER_120_1496 ();
 b15zdnd11an1n64x5 FILLER_120_1560 ();
 b15zdnd11an1n64x5 FILLER_120_1624 ();
 b15zdnd11an1n64x5 FILLER_120_1688 ();
 b15zdnd11an1n64x5 FILLER_120_1752 ();
 b15zdnd11an1n64x5 FILLER_120_1816 ();
 b15zdnd11an1n08x5 FILLER_120_1880 ();
 b15zdnd11an1n64x5 FILLER_120_1891 ();
 b15zdnd11an1n64x5 FILLER_120_1955 ();
 b15zdnd11an1n16x5 FILLER_120_2019 ();
 b15zdnd11an1n04x5 FILLER_120_2035 ();
 b15zdnd00an1n01x5 FILLER_120_2039 ();
 b15zdnd11an1n32x5 FILLER_120_2092 ();
 b15zdnd11an1n16x5 FILLER_120_2124 ();
 b15zdnd11an1n08x5 FILLER_120_2140 ();
 b15zdnd11an1n04x5 FILLER_120_2148 ();
 b15zdnd00an1n02x5 FILLER_120_2152 ();
 b15zdnd11an1n32x5 FILLER_120_2162 ();
 b15zdnd11an1n08x5 FILLER_120_2194 ();
 b15zdnd00an1n02x5 FILLER_120_2202 ();
 b15zdnd00an1n01x5 FILLER_120_2204 ();
 b15zdnd11an1n08x5 FILLER_120_2212 ();
 b15zdnd00an1n02x5 FILLER_120_2220 ();
 b15zdnd11an1n04x5 FILLER_120_2225 ();
 b15zdnd00an1n02x5 FILLER_120_2229 ();
 b15zdnd00an1n01x5 FILLER_120_2231 ();
 b15zdnd00an1n02x5 FILLER_120_2274 ();
 b15zdnd11an1n64x5 FILLER_121_0 ();
 b15zdnd11an1n64x5 FILLER_121_64 ();
 b15zdnd11an1n16x5 FILLER_121_128 ();
 b15zdnd00an1n02x5 FILLER_121_144 ();
 b15zdnd00an1n01x5 FILLER_121_146 ();
 b15zdnd11an1n64x5 FILLER_121_158 ();
 b15zdnd11an1n64x5 FILLER_121_222 ();
 b15zdnd11an1n08x5 FILLER_121_286 ();
 b15zdnd11an1n04x5 FILLER_121_294 ();
 b15zdnd00an1n02x5 FILLER_121_298 ();
 b15zdnd11an1n32x5 FILLER_121_304 ();
 b15zdnd11an1n16x5 FILLER_121_336 ();
 b15zdnd11an1n08x5 FILLER_121_352 ();
 b15zdnd11an1n04x5 FILLER_121_360 ();
 b15zdnd00an1n01x5 FILLER_121_364 ();
 b15zdnd11an1n32x5 FILLER_121_417 ();
 b15zdnd11an1n04x5 FILLER_121_449 ();
 b15zdnd11an1n64x5 FILLER_121_456 ();
 b15zdnd00an1n02x5 FILLER_121_520 ();
 b15zdnd11an1n04x5 FILLER_121_526 ();
 b15zdnd11an1n32x5 FILLER_121_534 ();
 b15zdnd11an1n16x5 FILLER_121_566 ();
 b15zdnd11an1n04x5 FILLER_121_582 ();
 b15zdnd11an1n64x5 FILLER_121_630 ();
 b15zdnd11an1n08x5 FILLER_121_694 ();
 b15zdnd00an1n02x5 FILLER_121_702 ();
 b15zdnd00an1n01x5 FILLER_121_704 ();
 b15zdnd11an1n04x5 FILLER_121_710 ();
 b15zdnd11an1n08x5 FILLER_121_717 ();
 b15zdnd00an1n02x5 FILLER_121_725 ();
 b15zdnd11an1n16x5 FILLER_121_730 ();
 b15zdnd11an1n04x5 FILLER_121_746 ();
 b15zdnd00an1n02x5 FILLER_121_750 ();
 b15zdnd00an1n01x5 FILLER_121_752 ();
 b15zdnd11an1n64x5 FILLER_121_762 ();
 b15zdnd11an1n64x5 FILLER_121_826 ();
 b15zdnd11an1n16x5 FILLER_121_890 ();
 b15zdnd11an1n08x5 FILLER_121_906 ();
 b15zdnd00an1n02x5 FILLER_121_914 ();
 b15zdnd11an1n64x5 FILLER_121_919 ();
 b15zdnd11an1n64x5 FILLER_121_983 ();
 b15zdnd11an1n64x5 FILLER_121_1047 ();
 b15zdnd11an1n32x5 FILLER_121_1111 ();
 b15zdnd00an1n01x5 FILLER_121_1143 ();
 b15zdnd11an1n32x5 FILLER_121_1155 ();
 b15zdnd11an1n16x5 FILLER_121_1187 ();
 b15zdnd00an1n02x5 FILLER_121_1203 ();
 b15zdnd11an1n32x5 FILLER_121_1217 ();
 b15zdnd11an1n16x5 FILLER_121_1249 ();
 b15zdnd11an1n04x5 FILLER_121_1265 ();
 b15zdnd00an1n02x5 FILLER_121_1269 ();
 b15zdnd00an1n01x5 FILLER_121_1271 ();
 b15zdnd11an1n64x5 FILLER_121_1317 ();
 b15zdnd11an1n64x5 FILLER_121_1381 ();
 b15zdnd11an1n64x5 FILLER_121_1445 ();
 b15zdnd11an1n64x5 FILLER_121_1509 ();
 b15zdnd11an1n32x5 FILLER_121_1573 ();
 b15zdnd11an1n16x5 FILLER_121_1605 ();
 b15zdnd11an1n04x5 FILLER_121_1621 ();
 b15zdnd00an1n02x5 FILLER_121_1625 ();
 b15zdnd11an1n64x5 FILLER_121_1636 ();
 b15zdnd11an1n64x5 FILLER_121_1700 ();
 b15zdnd11an1n64x5 FILLER_121_1764 ();
 b15zdnd11an1n08x5 FILLER_121_1828 ();
 b15zdnd11an1n04x5 FILLER_121_1836 ();
 b15zdnd11an1n64x5 FILLER_121_1860 ();
 b15zdnd11an1n64x5 FILLER_121_1924 ();
 b15zdnd11an1n64x5 FILLER_121_1988 ();
 b15zdnd11an1n04x5 FILLER_121_2052 ();
 b15zdnd00an1n02x5 FILLER_121_2056 ();
 b15zdnd11an1n04x5 FILLER_121_2061 ();
 b15zdnd11an1n04x5 FILLER_121_2068 ();
 b15zdnd11an1n64x5 FILLER_121_2075 ();
 b15zdnd11an1n64x5 FILLER_121_2139 ();
 b15zdnd11an1n16x5 FILLER_121_2203 ();
 b15zdnd11an1n08x5 FILLER_121_2219 ();
 b15zdnd00an1n02x5 FILLER_121_2227 ();
 b15zdnd11an1n16x5 FILLER_121_2232 ();
 b15zdnd11an1n32x5 FILLER_121_2252 ();
 b15zdnd11an1n64x5 FILLER_122_8 ();
 b15zdnd11an1n64x5 FILLER_122_72 ();
 b15zdnd11an1n64x5 FILLER_122_136 ();
 b15zdnd11an1n64x5 FILLER_122_200 ();
 b15zdnd11an1n64x5 FILLER_122_264 ();
 b15zdnd11an1n32x5 FILLER_122_328 ();
 b15zdnd11an1n16x5 FILLER_122_360 ();
 b15zdnd00an1n02x5 FILLER_122_376 ();
 b15zdnd11an1n04x5 FILLER_122_381 ();
 b15zdnd11an1n04x5 FILLER_122_388 ();
 b15zdnd11an1n32x5 FILLER_122_395 ();
 b15zdnd11an1n16x5 FILLER_122_427 ();
 b15zdnd00an1n02x5 FILLER_122_443 ();
 b15zdnd11an1n04x5 FILLER_122_448 ();
 b15zdnd11an1n64x5 FILLER_122_455 ();
 b15zdnd11an1n64x5 FILLER_122_519 ();
 b15zdnd11an1n16x5 FILLER_122_583 ();
 b15zdnd00an1n02x5 FILLER_122_599 ();
 b15zdnd11an1n04x5 FILLER_122_604 ();
 b15zdnd11an1n64x5 FILLER_122_611 ();
 b15zdnd11an1n16x5 FILLER_122_675 ();
 b15zdnd11an1n04x5 FILLER_122_691 ();
 b15zdnd11an1n04x5 FILLER_122_698 ();
 b15zdnd00an1n02x5 FILLER_122_716 ();
 b15zdnd00an1n02x5 FILLER_122_726 ();
 b15zdnd11an1n04x5 FILLER_122_738 ();
 b15zdnd00an1n01x5 FILLER_122_742 ();
 b15zdnd11an1n16x5 FILLER_122_763 ();
 b15zdnd00an1n02x5 FILLER_122_779 ();
 b15zdnd11an1n32x5 FILLER_122_795 ();
 b15zdnd11an1n16x5 FILLER_122_827 ();
 b15zdnd11an1n08x5 FILLER_122_843 ();
 b15zdnd00an1n01x5 FILLER_122_851 ();
 b15zdnd11an1n64x5 FILLER_122_864 ();
 b15zdnd11an1n64x5 FILLER_122_928 ();
 b15zdnd11an1n64x5 FILLER_122_992 ();
 b15zdnd11an1n64x5 FILLER_122_1056 ();
 b15zdnd11an1n64x5 FILLER_122_1120 ();
 b15zdnd11an1n64x5 FILLER_122_1184 ();
 b15zdnd11an1n04x5 FILLER_122_1248 ();
 b15zdnd00an1n02x5 FILLER_122_1252 ();
 b15zdnd00an1n01x5 FILLER_122_1254 ();
 b15zdnd11an1n64x5 FILLER_122_1262 ();
 b15zdnd11an1n64x5 FILLER_122_1326 ();
 b15zdnd11an1n32x5 FILLER_122_1390 ();
 b15zdnd11an1n16x5 FILLER_122_1422 ();
 b15zdnd11an1n64x5 FILLER_122_1445 ();
 b15zdnd11an1n64x5 FILLER_122_1509 ();
 b15zdnd11an1n64x5 FILLER_122_1573 ();
 b15zdnd11an1n64x5 FILLER_122_1637 ();
 b15zdnd11an1n64x5 FILLER_122_1701 ();
 b15zdnd11an1n64x5 FILLER_122_1765 ();
 b15zdnd11an1n32x5 FILLER_122_1829 ();
 b15zdnd11an1n04x5 FILLER_122_1861 ();
 b15zdnd00an1n02x5 FILLER_122_1865 ();
 b15zdnd00an1n01x5 FILLER_122_1867 ();
 b15zdnd11an1n64x5 FILLER_122_1885 ();
 b15zdnd11an1n64x5 FILLER_122_1949 ();
 b15zdnd11an1n32x5 FILLER_122_2013 ();
 b15zdnd11an1n16x5 FILLER_122_2045 ();
 b15zdnd11an1n04x5 FILLER_122_2061 ();
 b15zdnd11an1n64x5 FILLER_122_2068 ();
 b15zdnd11an1n16x5 FILLER_122_2132 ();
 b15zdnd11an1n04x5 FILLER_122_2148 ();
 b15zdnd00an1n02x5 FILLER_122_2152 ();
 b15zdnd11an1n16x5 FILLER_122_2162 ();
 b15zdnd00an1n02x5 FILLER_122_2178 ();
 b15zdnd00an1n01x5 FILLER_122_2180 ();
 b15zdnd11an1n64x5 FILLER_122_2188 ();
 b15zdnd11an1n16x5 FILLER_122_2252 ();
 b15zdnd11an1n08x5 FILLER_122_2268 ();
 b15zdnd11an1n16x5 FILLER_123_0 ();
 b15zdnd11an1n08x5 FILLER_123_16 ();
 b15zdnd00an1n02x5 FILLER_123_24 ();
 b15zdnd00an1n01x5 FILLER_123_26 ();
 b15zdnd11an1n64x5 FILLER_123_37 ();
 b15zdnd11an1n64x5 FILLER_123_101 ();
 b15zdnd11an1n64x5 FILLER_123_165 ();
 b15zdnd11an1n64x5 FILLER_123_229 ();
 b15zdnd11an1n64x5 FILLER_123_293 ();
 b15zdnd11an1n32x5 FILLER_123_357 ();
 b15zdnd00an1n01x5 FILLER_123_389 ();
 b15zdnd11an1n32x5 FILLER_123_393 ();
 b15zdnd00an1n01x5 FILLER_123_425 ();
 b15zdnd11an1n64x5 FILLER_123_478 ();
 b15zdnd11an1n64x5 FILLER_123_542 ();
 b15zdnd11an1n64x5 FILLER_123_606 ();
 b15zdnd11an1n16x5 FILLER_123_670 ();
 b15zdnd11an1n08x5 FILLER_123_686 ();
 b15zdnd11an1n04x5 FILLER_123_694 ();
 b15zdnd00an1n02x5 FILLER_123_698 ();
 b15zdnd11an1n08x5 FILLER_123_714 ();
 b15zdnd11an1n04x5 FILLER_123_722 ();
 b15zdnd00an1n02x5 FILLER_123_726 ();
 b15zdnd00an1n01x5 FILLER_123_728 ();
 b15zdnd11an1n64x5 FILLER_123_745 ();
 b15zdnd11an1n08x5 FILLER_123_809 ();
 b15zdnd11an1n04x5 FILLER_123_817 ();
 b15zdnd11an1n04x5 FILLER_123_828 ();
 b15zdnd00an1n02x5 FILLER_123_832 ();
 b15zdnd00an1n01x5 FILLER_123_834 ();
 b15zdnd11an1n64x5 FILLER_123_855 ();
 b15zdnd11an1n64x5 FILLER_123_919 ();
 b15zdnd11an1n64x5 FILLER_123_983 ();
 b15zdnd11an1n64x5 FILLER_123_1047 ();
 b15zdnd11an1n32x5 FILLER_123_1111 ();
 b15zdnd11an1n16x5 FILLER_123_1143 ();
 b15zdnd11an1n08x5 FILLER_123_1159 ();
 b15zdnd11an1n04x5 FILLER_123_1167 ();
 b15zdnd00an1n02x5 FILLER_123_1171 ();
 b15zdnd11an1n64x5 FILLER_123_1185 ();
 b15zdnd11an1n64x5 FILLER_123_1249 ();
 b15zdnd11an1n64x5 FILLER_123_1313 ();
 b15zdnd11an1n32x5 FILLER_123_1377 ();
 b15zdnd11an1n16x5 FILLER_123_1409 ();
 b15zdnd11an1n04x5 FILLER_123_1425 ();
 b15zdnd11an1n64x5 FILLER_123_1446 ();
 b15zdnd11an1n08x5 FILLER_123_1510 ();
 b15zdnd11an1n04x5 FILLER_123_1518 ();
 b15zdnd11an1n64x5 FILLER_123_1533 ();
 b15zdnd11an1n32x5 FILLER_123_1597 ();
 b15zdnd11an1n64x5 FILLER_123_1638 ();
 b15zdnd11an1n64x5 FILLER_123_1702 ();
 b15zdnd11an1n64x5 FILLER_123_1766 ();
 b15zdnd11an1n08x5 FILLER_123_1830 ();
 b15zdnd11an1n04x5 FILLER_123_1838 ();
 b15zdnd00an1n02x5 FILLER_123_1842 ();
 b15zdnd11an1n64x5 FILLER_123_1865 ();
 b15zdnd11an1n64x5 FILLER_123_1929 ();
 b15zdnd11an1n64x5 FILLER_123_1993 ();
 b15zdnd11an1n16x5 FILLER_123_2057 ();
 b15zdnd11an1n64x5 FILLER_123_2082 ();
 b15zdnd11an1n64x5 FILLER_123_2146 ();
 b15zdnd11an1n64x5 FILLER_123_2210 ();
 b15zdnd11an1n08x5 FILLER_123_2274 ();
 b15zdnd00an1n02x5 FILLER_123_2282 ();
 b15zdnd00an1n02x5 FILLER_124_8 ();
 b15zdnd11an1n04x5 FILLER_124_21 ();
 b15zdnd00an1n02x5 FILLER_124_25 ();
 b15zdnd00an1n01x5 FILLER_124_27 ();
 b15zdnd11an1n64x5 FILLER_124_42 ();
 b15zdnd11an1n64x5 FILLER_124_106 ();
 b15zdnd11an1n64x5 FILLER_124_170 ();
 b15zdnd11an1n16x5 FILLER_124_234 ();
 b15zdnd11an1n08x5 FILLER_124_250 ();
 b15zdnd00an1n02x5 FILLER_124_258 ();
 b15zdnd00an1n01x5 FILLER_124_260 ();
 b15zdnd11an1n16x5 FILLER_124_275 ();
 b15zdnd11an1n08x5 FILLER_124_291 ();
 b15zdnd11an1n04x5 FILLER_124_299 ();
 b15zdnd00an1n01x5 FILLER_124_303 ();
 b15zdnd11an1n64x5 FILLER_124_318 ();
 b15zdnd11an1n64x5 FILLER_124_382 ();
 b15zdnd11an1n04x5 FILLER_124_446 ();
 b15zdnd00an1n02x5 FILLER_124_450 ();
 b15zdnd11an1n64x5 FILLER_124_455 ();
 b15zdnd00an1n01x5 FILLER_124_519 ();
 b15zdnd11an1n64x5 FILLER_124_526 ();
 b15zdnd11an1n64x5 FILLER_124_590 ();
 b15zdnd11an1n32x5 FILLER_124_654 ();
 b15zdnd11an1n04x5 FILLER_124_686 ();
 b15zdnd00an1n02x5 FILLER_124_690 ();
 b15zdnd00an1n02x5 FILLER_124_716 ();
 b15zdnd11an1n64x5 FILLER_124_726 ();
 b15zdnd11an1n16x5 FILLER_124_790 ();
 b15zdnd11an1n08x5 FILLER_124_806 ();
 b15zdnd11an1n04x5 FILLER_124_814 ();
 b15zdnd11an1n32x5 FILLER_124_838 ();
 b15zdnd11an1n16x5 FILLER_124_870 ();
 b15zdnd11an1n08x5 FILLER_124_886 ();
 b15zdnd11an1n04x5 FILLER_124_894 ();
 b15zdnd00an1n02x5 FILLER_124_898 ();
 b15zdnd00an1n01x5 FILLER_124_900 ();
 b15zdnd11an1n64x5 FILLER_124_907 ();
 b15zdnd11an1n64x5 FILLER_124_971 ();
 b15zdnd11an1n64x5 FILLER_124_1035 ();
 b15zdnd11an1n64x5 FILLER_124_1099 ();
 b15zdnd11an1n08x5 FILLER_124_1163 ();
 b15zdnd11an1n04x5 FILLER_124_1171 ();
 b15zdnd00an1n02x5 FILLER_124_1175 ();
 b15zdnd00an1n01x5 FILLER_124_1177 ();
 b15zdnd11an1n64x5 FILLER_124_1190 ();
 b15zdnd11an1n64x5 FILLER_124_1254 ();
 b15zdnd11an1n32x5 FILLER_124_1318 ();
 b15zdnd11an1n16x5 FILLER_124_1350 ();
 b15zdnd11an1n08x5 FILLER_124_1366 ();
 b15zdnd00an1n02x5 FILLER_124_1374 ();
 b15zdnd00an1n01x5 FILLER_124_1376 ();
 b15zdnd11an1n64x5 FILLER_124_1394 ();
 b15zdnd11an1n32x5 FILLER_124_1458 ();
 b15zdnd11an1n16x5 FILLER_124_1490 ();
 b15zdnd11an1n08x5 FILLER_124_1506 ();
 b15zdnd00an1n01x5 FILLER_124_1514 ();
 b15zdnd11an1n64x5 FILLER_124_1524 ();
 b15zdnd11an1n64x5 FILLER_124_1588 ();
 b15zdnd11an1n64x5 FILLER_124_1652 ();
 b15zdnd11an1n64x5 FILLER_124_1716 ();
 b15zdnd00an1n02x5 FILLER_124_1780 ();
 b15zdnd11an1n64x5 FILLER_124_1802 ();
 b15zdnd11an1n64x5 FILLER_124_1866 ();
 b15zdnd11an1n64x5 FILLER_124_1930 ();
 b15zdnd11an1n64x5 FILLER_124_1994 ();
 b15zdnd11an1n64x5 FILLER_124_2058 ();
 b15zdnd11an1n32x5 FILLER_124_2122 ();
 b15zdnd11an1n64x5 FILLER_124_2162 ();
 b15zdnd11an1n32x5 FILLER_124_2226 ();
 b15zdnd11an1n16x5 FILLER_124_2258 ();
 b15zdnd00an1n02x5 FILLER_124_2274 ();
 b15zdnd11an1n16x5 FILLER_125_0 ();
 b15zdnd00an1n01x5 FILLER_125_16 ();
 b15zdnd11an1n64x5 FILLER_125_28 ();
 b15zdnd11an1n64x5 FILLER_125_92 ();
 b15zdnd11an1n04x5 FILLER_125_156 ();
 b15zdnd00an1n02x5 FILLER_125_160 ();
 b15zdnd00an1n01x5 FILLER_125_162 ();
 b15zdnd11an1n64x5 FILLER_125_168 ();
 b15zdnd11an1n64x5 FILLER_125_232 ();
 b15zdnd11an1n08x5 FILLER_125_296 ();
 b15zdnd00an1n02x5 FILLER_125_304 ();
 b15zdnd11an1n64x5 FILLER_125_310 ();
 b15zdnd11an1n64x5 FILLER_125_374 ();
 b15zdnd11an1n64x5 FILLER_125_438 ();
 b15zdnd11an1n64x5 FILLER_125_502 ();
 b15zdnd11an1n64x5 FILLER_125_566 ();
 b15zdnd11an1n64x5 FILLER_125_630 ();
 b15zdnd11an1n04x5 FILLER_125_694 ();
 b15zdnd00an1n01x5 FILLER_125_698 ();
 b15zdnd11an1n64x5 FILLER_125_715 ();
 b15zdnd11an1n64x5 FILLER_125_779 ();
 b15zdnd11an1n64x5 FILLER_125_843 ();
 b15zdnd11an1n64x5 FILLER_125_907 ();
 b15zdnd11an1n64x5 FILLER_125_971 ();
 b15zdnd11an1n64x5 FILLER_125_1035 ();
 b15zdnd11an1n64x5 FILLER_125_1099 ();
 b15zdnd11an1n08x5 FILLER_125_1163 ();
 b15zdnd00an1n02x5 FILLER_125_1171 ();
 b15zdnd11an1n64x5 FILLER_125_1184 ();
 b15zdnd11an1n08x5 FILLER_125_1248 ();
 b15zdnd00an1n02x5 FILLER_125_1256 ();
 b15zdnd11an1n32x5 FILLER_125_1265 ();
 b15zdnd11an1n16x5 FILLER_125_1297 ();
 b15zdnd11an1n04x5 FILLER_125_1313 ();
 b15zdnd00an1n02x5 FILLER_125_1317 ();
 b15zdnd00an1n01x5 FILLER_125_1319 ();
 b15zdnd11an1n64x5 FILLER_125_1337 ();
 b15zdnd11an1n32x5 FILLER_125_1401 ();
 b15zdnd00an1n02x5 FILLER_125_1433 ();
 b15zdnd00an1n01x5 FILLER_125_1435 ();
 b15zdnd11an1n64x5 FILLER_125_1441 ();
 b15zdnd11an1n04x5 FILLER_125_1505 ();
 b15zdnd00an1n02x5 FILLER_125_1509 ();
 b15zdnd11an1n64x5 FILLER_125_1520 ();
 b15zdnd11an1n64x5 FILLER_125_1584 ();
 b15zdnd11an1n64x5 FILLER_125_1648 ();
 b15zdnd11an1n64x5 FILLER_125_1712 ();
 b15zdnd11an1n64x5 FILLER_125_1776 ();
 b15zdnd11an1n64x5 FILLER_125_1840 ();
 b15zdnd11an1n64x5 FILLER_125_1904 ();
 b15zdnd11an1n64x5 FILLER_125_1968 ();
 b15zdnd11an1n64x5 FILLER_125_2032 ();
 b15zdnd11an1n64x5 FILLER_125_2096 ();
 b15zdnd11an1n64x5 FILLER_125_2160 ();
 b15zdnd11an1n32x5 FILLER_125_2224 ();
 b15zdnd11an1n16x5 FILLER_125_2256 ();
 b15zdnd11an1n08x5 FILLER_125_2272 ();
 b15zdnd11an1n04x5 FILLER_125_2280 ();
 b15zdnd11an1n64x5 FILLER_126_8 ();
 b15zdnd11an1n64x5 FILLER_126_72 ();
 b15zdnd11an1n64x5 FILLER_126_136 ();
 b15zdnd11an1n64x5 FILLER_126_200 ();
 b15zdnd11an1n64x5 FILLER_126_264 ();
 b15zdnd11an1n64x5 FILLER_126_328 ();
 b15zdnd11an1n64x5 FILLER_126_392 ();
 b15zdnd11an1n16x5 FILLER_126_456 ();
 b15zdnd11an1n04x5 FILLER_126_472 ();
 b15zdnd00an1n01x5 FILLER_126_476 ();
 b15zdnd11an1n32x5 FILLER_126_485 ();
 b15zdnd11an1n04x5 FILLER_126_525 ();
 b15zdnd11an1n64x5 FILLER_126_533 ();
 b15zdnd11an1n64x5 FILLER_126_597 ();
 b15zdnd11an1n32x5 FILLER_126_661 ();
 b15zdnd11an1n16x5 FILLER_126_693 ();
 b15zdnd11an1n08x5 FILLER_126_709 ();
 b15zdnd00an1n01x5 FILLER_126_717 ();
 b15zdnd11an1n16x5 FILLER_126_726 ();
 b15zdnd00an1n01x5 FILLER_126_742 ();
 b15zdnd11an1n04x5 FILLER_126_763 ();
 b15zdnd11an1n64x5 FILLER_126_776 ();
 b15zdnd11an1n64x5 FILLER_126_840 ();
 b15zdnd11an1n64x5 FILLER_126_904 ();
 b15zdnd11an1n64x5 FILLER_126_968 ();
 b15zdnd11an1n64x5 FILLER_126_1032 ();
 b15zdnd11an1n64x5 FILLER_126_1096 ();
 b15zdnd11an1n08x5 FILLER_126_1160 ();
 b15zdnd11an1n04x5 FILLER_126_1168 ();
 b15zdnd00an1n02x5 FILLER_126_1172 ();
 b15zdnd11an1n64x5 FILLER_126_1185 ();
 b15zdnd11an1n04x5 FILLER_126_1249 ();
 b15zdnd00an1n02x5 FILLER_126_1253 ();
 b15zdnd11an1n08x5 FILLER_126_1265 ();
 b15zdnd11an1n04x5 FILLER_126_1273 ();
 b15zdnd00an1n02x5 FILLER_126_1277 ();
 b15zdnd11an1n16x5 FILLER_126_1289 ();
 b15zdnd11an1n08x5 FILLER_126_1305 ();
 b15zdnd11an1n64x5 FILLER_126_1325 ();
 b15zdnd11an1n64x5 FILLER_126_1389 ();
 b15zdnd11an1n64x5 FILLER_126_1453 ();
 b15zdnd11an1n64x5 FILLER_126_1517 ();
 b15zdnd11an1n32x5 FILLER_126_1581 ();
 b15zdnd11an1n08x5 FILLER_126_1613 ();
 b15zdnd11an1n04x5 FILLER_126_1621 ();
 b15zdnd00an1n02x5 FILLER_126_1625 ();
 b15zdnd11an1n64x5 FILLER_126_1636 ();
 b15zdnd11an1n16x5 FILLER_126_1700 ();
 b15zdnd11an1n04x5 FILLER_126_1716 ();
 b15zdnd00an1n01x5 FILLER_126_1720 ();
 b15zdnd11an1n64x5 FILLER_126_1742 ();
 b15zdnd11an1n64x5 FILLER_126_1806 ();
 b15zdnd11an1n16x5 FILLER_126_1870 ();
 b15zdnd00an1n02x5 FILLER_126_1886 ();
 b15zdnd11an1n64x5 FILLER_126_1930 ();
 b15zdnd11an1n64x5 FILLER_126_1994 ();
 b15zdnd11an1n64x5 FILLER_126_2058 ();
 b15zdnd11an1n32x5 FILLER_126_2122 ();
 b15zdnd11an1n64x5 FILLER_126_2162 ();
 b15zdnd11an1n32x5 FILLER_126_2226 ();
 b15zdnd11an1n16x5 FILLER_126_2258 ();
 b15zdnd00an1n02x5 FILLER_126_2274 ();
 b15zdnd11an1n64x5 FILLER_127_0 ();
 b15zdnd11an1n64x5 FILLER_127_64 ();
 b15zdnd11an1n64x5 FILLER_127_128 ();
 b15zdnd11an1n64x5 FILLER_127_192 ();
 b15zdnd11an1n64x5 FILLER_127_256 ();
 b15zdnd11an1n64x5 FILLER_127_320 ();
 b15zdnd11an1n64x5 FILLER_127_384 ();
 b15zdnd11an1n64x5 FILLER_127_448 ();
 b15zdnd11an1n64x5 FILLER_127_512 ();
 b15zdnd11an1n16x5 FILLER_127_576 ();
 b15zdnd11an1n08x5 FILLER_127_592 ();
 b15zdnd00an1n02x5 FILLER_127_600 ();
 b15zdnd00an1n01x5 FILLER_127_602 ();
 b15zdnd11an1n64x5 FILLER_127_615 ();
 b15zdnd11an1n64x5 FILLER_127_679 ();
 b15zdnd11an1n64x5 FILLER_127_743 ();
 b15zdnd11an1n64x5 FILLER_127_807 ();
 b15zdnd11an1n08x5 FILLER_127_871 ();
 b15zdnd00an1n01x5 FILLER_127_879 ();
 b15zdnd11an1n08x5 FILLER_127_892 ();
 b15zdnd00an1n02x5 FILLER_127_900 ();
 b15zdnd11an1n64x5 FILLER_127_916 ();
 b15zdnd11an1n64x5 FILLER_127_980 ();
 b15zdnd11an1n64x5 FILLER_127_1044 ();
 b15zdnd11an1n64x5 FILLER_127_1108 ();
 b15zdnd11an1n64x5 FILLER_127_1172 ();
 b15zdnd11an1n08x5 FILLER_127_1236 ();
 b15zdnd11an1n04x5 FILLER_127_1244 ();
 b15zdnd00an1n02x5 FILLER_127_1248 ();
 b15zdnd11an1n64x5 FILLER_127_1256 ();
 b15zdnd11an1n64x5 FILLER_127_1320 ();
 b15zdnd11an1n64x5 FILLER_127_1384 ();
 b15zdnd11an1n64x5 FILLER_127_1448 ();
 b15zdnd11an1n64x5 FILLER_127_1512 ();
 b15zdnd11an1n64x5 FILLER_127_1576 ();
 b15zdnd11an1n64x5 FILLER_127_1640 ();
 b15zdnd11an1n64x5 FILLER_127_1704 ();
 b15zdnd11an1n64x5 FILLER_127_1768 ();
 b15zdnd11an1n64x5 FILLER_127_1832 ();
 b15zdnd11an1n64x5 FILLER_127_1896 ();
 b15zdnd11an1n64x5 FILLER_127_1960 ();
 b15zdnd11an1n64x5 FILLER_127_2024 ();
 b15zdnd11an1n64x5 FILLER_127_2088 ();
 b15zdnd11an1n64x5 FILLER_127_2152 ();
 b15zdnd11an1n64x5 FILLER_127_2216 ();
 b15zdnd11an1n04x5 FILLER_127_2280 ();
 b15zdnd11an1n64x5 FILLER_128_8 ();
 b15zdnd11an1n64x5 FILLER_128_72 ();
 b15zdnd11an1n64x5 FILLER_128_136 ();
 b15zdnd11an1n64x5 FILLER_128_200 ();
 b15zdnd11an1n64x5 FILLER_128_264 ();
 b15zdnd11an1n64x5 FILLER_128_328 ();
 b15zdnd11an1n64x5 FILLER_128_392 ();
 b15zdnd11an1n64x5 FILLER_128_456 ();
 b15zdnd11an1n64x5 FILLER_128_520 ();
 b15zdnd11an1n64x5 FILLER_128_584 ();
 b15zdnd11an1n32x5 FILLER_128_648 ();
 b15zdnd11an1n16x5 FILLER_128_680 ();
 b15zdnd00an1n02x5 FILLER_128_696 ();
 b15zdnd00an1n01x5 FILLER_128_698 ();
 b15zdnd11an1n04x5 FILLER_128_711 ();
 b15zdnd00an1n02x5 FILLER_128_715 ();
 b15zdnd00an1n01x5 FILLER_128_717 ();
 b15zdnd11an1n64x5 FILLER_128_726 ();
 b15zdnd11an1n32x5 FILLER_128_790 ();
 b15zdnd11an1n16x5 FILLER_128_822 ();
 b15zdnd11an1n04x5 FILLER_128_838 ();
 b15zdnd11an1n04x5 FILLER_128_849 ();
 b15zdnd00an1n02x5 FILLER_128_853 ();
 b15zdnd11an1n64x5 FILLER_128_875 ();
 b15zdnd11an1n64x5 FILLER_128_939 ();
 b15zdnd11an1n64x5 FILLER_128_1003 ();
 b15zdnd11an1n64x5 FILLER_128_1067 ();
 b15zdnd11an1n04x5 FILLER_128_1131 ();
 b15zdnd00an1n01x5 FILLER_128_1135 ();
 b15zdnd11an1n64x5 FILLER_128_1145 ();
 b15zdnd11an1n64x5 FILLER_128_1209 ();
 b15zdnd11an1n04x5 FILLER_128_1273 ();
 b15zdnd00an1n01x5 FILLER_128_1277 ();
 b15zdnd11an1n16x5 FILLER_128_1294 ();
 b15zdnd11an1n04x5 FILLER_128_1310 ();
 b15zdnd11an1n64x5 FILLER_128_1326 ();
 b15zdnd11an1n64x5 FILLER_128_1390 ();
 b15zdnd11an1n64x5 FILLER_128_1454 ();
 b15zdnd11an1n64x5 FILLER_128_1518 ();
 b15zdnd11an1n64x5 FILLER_128_1582 ();
 b15zdnd11an1n64x5 FILLER_128_1646 ();
 b15zdnd11an1n64x5 FILLER_128_1710 ();
 b15zdnd11an1n64x5 FILLER_128_1774 ();
 b15zdnd11an1n64x5 FILLER_128_1838 ();
 b15zdnd11an1n64x5 FILLER_128_1902 ();
 b15zdnd11an1n64x5 FILLER_128_1966 ();
 b15zdnd11an1n16x5 FILLER_128_2030 ();
 b15zdnd11an1n08x5 FILLER_128_2046 ();
 b15zdnd11an1n04x5 FILLER_128_2054 ();
 b15zdnd00an1n01x5 FILLER_128_2058 ();
 b15zdnd11an1n64x5 FILLER_128_2067 ();
 b15zdnd11an1n16x5 FILLER_128_2131 ();
 b15zdnd11an1n04x5 FILLER_128_2147 ();
 b15zdnd00an1n02x5 FILLER_128_2151 ();
 b15zdnd00an1n01x5 FILLER_128_2153 ();
 b15zdnd11an1n08x5 FILLER_128_2162 ();
 b15zdnd00an1n01x5 FILLER_128_2170 ();
 b15zdnd11an1n64x5 FILLER_128_2178 ();
 b15zdnd11an1n32x5 FILLER_128_2242 ();
 b15zdnd00an1n02x5 FILLER_128_2274 ();
 b15zdnd11an1n64x5 FILLER_129_0 ();
 b15zdnd00an1n02x5 FILLER_129_64 ();
 b15zdnd00an1n01x5 FILLER_129_66 ();
 b15zdnd11an1n64x5 FILLER_129_76 ();
 b15zdnd11an1n16x5 FILLER_129_140 ();
 b15zdnd11an1n08x5 FILLER_129_156 ();
 b15zdnd11an1n04x5 FILLER_129_164 ();
 b15zdnd11an1n64x5 FILLER_129_210 ();
 b15zdnd11an1n64x5 FILLER_129_274 ();
 b15zdnd11an1n64x5 FILLER_129_338 ();
 b15zdnd11an1n64x5 FILLER_129_402 ();
 b15zdnd11an1n64x5 FILLER_129_466 ();
 b15zdnd11an1n64x5 FILLER_129_530 ();
 b15zdnd11an1n64x5 FILLER_129_594 ();
 b15zdnd11an1n32x5 FILLER_129_658 ();
 b15zdnd11an1n08x5 FILLER_129_690 ();
 b15zdnd00an1n02x5 FILLER_129_698 ();
 b15zdnd11an1n64x5 FILLER_129_714 ();
 b15zdnd11an1n32x5 FILLER_129_778 ();
 b15zdnd11an1n08x5 FILLER_129_810 ();
 b15zdnd11an1n04x5 FILLER_129_818 ();
 b15zdnd00an1n02x5 FILLER_129_822 ();
 b15zdnd11an1n04x5 FILLER_129_848 ();
 b15zdnd11an1n64x5 FILLER_129_859 ();
 b15zdnd11an1n64x5 FILLER_129_923 ();
 b15zdnd11an1n16x5 FILLER_129_987 ();
 b15zdnd11an1n08x5 FILLER_129_1003 ();
 b15zdnd00an1n02x5 FILLER_129_1011 ();
 b15zdnd00an1n01x5 FILLER_129_1013 ();
 b15zdnd11an1n64x5 FILLER_129_1038 ();
 b15zdnd11an1n32x5 FILLER_129_1102 ();
 b15zdnd11an1n16x5 FILLER_129_1134 ();
 b15zdnd11an1n08x5 FILLER_129_1150 ();
 b15zdnd11an1n04x5 FILLER_129_1158 ();
 b15zdnd00an1n01x5 FILLER_129_1162 ();
 b15zdnd11an1n32x5 FILLER_129_1175 ();
 b15zdnd11an1n16x5 FILLER_129_1207 ();
 b15zdnd11an1n08x5 FILLER_129_1223 ();
 b15zdnd00an1n02x5 FILLER_129_1231 ();
 b15zdnd11an1n64x5 FILLER_129_1239 ();
 b15zdnd11an1n64x5 FILLER_129_1303 ();
 b15zdnd11an1n64x5 FILLER_129_1367 ();
 b15zdnd11an1n16x5 FILLER_129_1431 ();
 b15zdnd11an1n08x5 FILLER_129_1447 ();
 b15zdnd11an1n04x5 FILLER_129_1455 ();
 b15zdnd11an1n32x5 FILLER_129_1479 ();
 b15zdnd11an1n16x5 FILLER_129_1511 ();
 b15zdnd11an1n04x5 FILLER_129_1527 ();
 b15zdnd11an1n64x5 FILLER_129_1542 ();
 b15zdnd11an1n64x5 FILLER_129_1606 ();
 b15zdnd11an1n64x5 FILLER_129_1670 ();
 b15zdnd11an1n64x5 FILLER_129_1734 ();
 b15zdnd11an1n64x5 FILLER_129_1798 ();
 b15zdnd11an1n64x5 FILLER_129_1862 ();
 b15zdnd00an1n02x5 FILLER_129_1926 ();
 b15zdnd11an1n64x5 FILLER_129_1931 ();
 b15zdnd11an1n64x5 FILLER_129_1995 ();
 b15zdnd11an1n64x5 FILLER_129_2059 ();
 b15zdnd11an1n64x5 FILLER_129_2123 ();
 b15zdnd11an1n64x5 FILLER_129_2187 ();
 b15zdnd11an1n32x5 FILLER_129_2251 ();
 b15zdnd00an1n01x5 FILLER_129_2283 ();
 b15zdnd11an1n64x5 FILLER_130_8 ();
 b15zdnd11an1n04x5 FILLER_130_72 ();
 b15zdnd11an1n64x5 FILLER_130_121 ();
 b15zdnd00an1n02x5 FILLER_130_185 ();
 b15zdnd00an1n01x5 FILLER_130_187 ();
 b15zdnd11an1n16x5 FILLER_130_192 ();
 b15zdnd11an1n04x5 FILLER_130_208 ();
 b15zdnd00an1n01x5 FILLER_130_212 ();
 b15zdnd11an1n64x5 FILLER_130_265 ();
 b15zdnd11an1n64x5 FILLER_130_329 ();
 b15zdnd11an1n64x5 FILLER_130_393 ();
 b15zdnd11an1n64x5 FILLER_130_457 ();
 b15zdnd11an1n64x5 FILLER_130_521 ();
 b15zdnd11an1n64x5 FILLER_130_585 ();
 b15zdnd11an1n32x5 FILLER_130_649 ();
 b15zdnd11an1n16x5 FILLER_130_681 ();
 b15zdnd00an1n02x5 FILLER_130_697 ();
 b15zdnd00an1n01x5 FILLER_130_699 ();
 b15zdnd00an1n02x5 FILLER_130_716 ();
 b15zdnd11an1n64x5 FILLER_130_726 ();
 b15zdnd11an1n64x5 FILLER_130_790 ();
 b15zdnd11an1n64x5 FILLER_130_854 ();
 b15zdnd11an1n64x5 FILLER_130_918 ();
 b15zdnd11an1n64x5 FILLER_130_982 ();
 b15zdnd11an1n64x5 FILLER_130_1046 ();
 b15zdnd11an1n64x5 FILLER_130_1110 ();
 b15zdnd11an1n64x5 FILLER_130_1174 ();
 b15zdnd11an1n64x5 FILLER_130_1238 ();
 b15zdnd11an1n16x5 FILLER_130_1302 ();
 b15zdnd00an1n01x5 FILLER_130_1318 ();
 b15zdnd11an1n64x5 FILLER_130_1333 ();
 b15zdnd11an1n64x5 FILLER_130_1397 ();
 b15zdnd11an1n64x5 FILLER_130_1461 ();
 b15zdnd11an1n08x5 FILLER_130_1525 ();
 b15zdnd00an1n01x5 FILLER_130_1533 ();
 b15zdnd11an1n64x5 FILLER_130_1543 ();
 b15zdnd11an1n64x5 FILLER_130_1607 ();
 b15zdnd11an1n64x5 FILLER_130_1671 ();
 b15zdnd11an1n16x5 FILLER_130_1735 ();
 b15zdnd11an1n08x5 FILLER_130_1751 ();
 b15zdnd00an1n01x5 FILLER_130_1759 ();
 b15zdnd11an1n64x5 FILLER_130_1768 ();
 b15zdnd11an1n64x5 FILLER_130_1832 ();
 b15zdnd11an1n08x5 FILLER_130_1896 ();
 b15zdnd00an1n01x5 FILLER_130_1904 ();
 b15zdnd11an1n64x5 FILLER_130_1933 ();
 b15zdnd11an1n64x5 FILLER_130_1997 ();
 b15zdnd11an1n64x5 FILLER_130_2061 ();
 b15zdnd11an1n16x5 FILLER_130_2125 ();
 b15zdnd11an1n08x5 FILLER_130_2141 ();
 b15zdnd11an1n04x5 FILLER_130_2149 ();
 b15zdnd00an1n01x5 FILLER_130_2153 ();
 b15zdnd11an1n64x5 FILLER_130_2162 ();
 b15zdnd11an1n32x5 FILLER_130_2226 ();
 b15zdnd11an1n04x5 FILLER_130_2258 ();
 b15zdnd00an1n01x5 FILLER_130_2262 ();
 b15zdnd11an1n08x5 FILLER_130_2267 ();
 b15zdnd00an1n01x5 FILLER_130_2275 ();
 b15zdnd11an1n64x5 FILLER_131_0 ();
 b15zdnd11an1n64x5 FILLER_131_64 ();
 b15zdnd11an1n64x5 FILLER_131_128 ();
 b15zdnd11an1n32x5 FILLER_131_192 ();
 b15zdnd11an1n08x5 FILLER_131_224 ();
 b15zdnd00an1n01x5 FILLER_131_232 ();
 b15zdnd11an1n04x5 FILLER_131_236 ();
 b15zdnd11an1n64x5 FILLER_131_243 ();
 b15zdnd11an1n64x5 FILLER_131_307 ();
 b15zdnd11an1n64x5 FILLER_131_371 ();
 b15zdnd11an1n64x5 FILLER_131_435 ();
 b15zdnd11an1n64x5 FILLER_131_499 ();
 b15zdnd11an1n64x5 FILLER_131_563 ();
 b15zdnd11an1n64x5 FILLER_131_627 ();
 b15zdnd11an1n64x5 FILLER_131_691 ();
 b15zdnd11an1n64x5 FILLER_131_755 ();
 b15zdnd11an1n64x5 FILLER_131_819 ();
 b15zdnd11an1n64x5 FILLER_131_883 ();
 b15zdnd11an1n64x5 FILLER_131_947 ();
 b15zdnd11an1n64x5 FILLER_131_1011 ();
 b15zdnd11an1n64x5 FILLER_131_1075 ();
 b15zdnd11an1n64x5 FILLER_131_1139 ();
 b15zdnd11an1n64x5 FILLER_131_1203 ();
 b15zdnd11an1n64x5 FILLER_131_1267 ();
 b15zdnd11an1n64x5 FILLER_131_1331 ();
 b15zdnd11an1n64x5 FILLER_131_1395 ();
 b15zdnd11an1n64x5 FILLER_131_1459 ();
 b15zdnd11an1n32x5 FILLER_131_1523 ();
 b15zdnd11an1n16x5 FILLER_131_1555 ();
 b15zdnd00an1n01x5 FILLER_131_1571 ();
 b15zdnd11an1n64x5 FILLER_131_1575 ();
 b15zdnd11an1n64x5 FILLER_131_1639 ();
 b15zdnd11an1n64x5 FILLER_131_1703 ();
 b15zdnd11an1n64x5 FILLER_131_1767 ();
 b15zdnd11an1n64x5 FILLER_131_1831 ();
 b15zdnd11an1n16x5 FILLER_131_1895 ();
 b15zdnd11an1n08x5 FILLER_131_1911 ();
 b15zdnd11an1n04x5 FILLER_131_1919 ();
 b15zdnd00an1n01x5 FILLER_131_1923 ();
 b15zdnd11an1n64x5 FILLER_131_1927 ();
 b15zdnd11an1n64x5 FILLER_131_1991 ();
 b15zdnd11an1n64x5 FILLER_131_2055 ();
 b15zdnd11an1n64x5 FILLER_131_2119 ();
 b15zdnd11an1n64x5 FILLER_131_2183 ();
 b15zdnd11an1n32x5 FILLER_131_2247 ();
 b15zdnd11an1n04x5 FILLER_131_2279 ();
 b15zdnd00an1n01x5 FILLER_131_2283 ();
 b15zdnd11an1n16x5 FILLER_132_8 ();
 b15zdnd11an1n08x5 FILLER_132_24 ();
 b15zdnd11an1n04x5 FILLER_132_32 ();
 b15zdnd11an1n08x5 FILLER_132_40 ();
 b15zdnd11an1n04x5 FILLER_132_48 ();
 b15zdnd00an1n01x5 FILLER_132_52 ();
 b15zdnd11an1n04x5 FILLER_132_56 ();
 b15zdnd11an1n64x5 FILLER_132_63 ();
 b15zdnd11an1n32x5 FILLER_132_127 ();
 b15zdnd11an1n08x5 FILLER_132_159 ();
 b15zdnd11an1n16x5 FILLER_132_170 ();
 b15zdnd11an1n04x5 FILLER_132_186 ();
 b15zdnd11an1n08x5 FILLER_132_232 ();
 b15zdnd00an1n01x5 FILLER_132_240 ();
 b15zdnd11an1n64x5 FILLER_132_248 ();
 b15zdnd11an1n64x5 FILLER_132_312 ();
 b15zdnd11an1n64x5 FILLER_132_376 ();
 b15zdnd11an1n64x5 FILLER_132_440 ();
 b15zdnd11an1n64x5 FILLER_132_504 ();
 b15zdnd11an1n64x5 FILLER_132_568 ();
 b15zdnd11an1n64x5 FILLER_132_632 ();
 b15zdnd11an1n16x5 FILLER_132_696 ();
 b15zdnd11an1n04x5 FILLER_132_712 ();
 b15zdnd00an1n02x5 FILLER_132_716 ();
 b15zdnd00an1n02x5 FILLER_132_726 ();
 b15zdnd11an1n64x5 FILLER_132_742 ();
 b15zdnd11an1n64x5 FILLER_132_806 ();
 b15zdnd11an1n64x5 FILLER_132_870 ();
 b15zdnd11an1n64x5 FILLER_132_934 ();
 b15zdnd11an1n64x5 FILLER_132_998 ();
 b15zdnd11an1n64x5 FILLER_132_1062 ();
 b15zdnd11an1n64x5 FILLER_132_1126 ();
 b15zdnd11an1n64x5 FILLER_132_1190 ();
 b15zdnd11an1n64x5 FILLER_132_1254 ();
 b15zdnd11an1n64x5 FILLER_132_1318 ();
 b15zdnd11an1n64x5 FILLER_132_1382 ();
 b15zdnd11an1n64x5 FILLER_132_1446 ();
 b15zdnd11an1n32x5 FILLER_132_1510 ();
 b15zdnd11an1n16x5 FILLER_132_1542 ();
 b15zdnd11an1n08x5 FILLER_132_1558 ();
 b15zdnd11an1n04x5 FILLER_132_1566 ();
 b15zdnd00an1n02x5 FILLER_132_1570 ();
 b15zdnd11an1n32x5 FILLER_132_1599 ();
 b15zdnd11an1n16x5 FILLER_132_1631 ();
 b15zdnd11an1n08x5 FILLER_132_1647 ();
 b15zdnd11an1n04x5 FILLER_132_1655 ();
 b15zdnd00an1n01x5 FILLER_132_1659 ();
 b15zdnd11an1n04x5 FILLER_132_1663 ();
 b15zdnd11an1n64x5 FILLER_132_1670 ();
 b15zdnd11an1n64x5 FILLER_132_1734 ();
 b15zdnd11an1n64x5 FILLER_132_1798 ();
 b15zdnd11an1n64x5 FILLER_132_1862 ();
 b15zdnd11an1n64x5 FILLER_132_1926 ();
 b15zdnd11an1n64x5 FILLER_132_1990 ();
 b15zdnd11an1n64x5 FILLER_132_2054 ();
 b15zdnd11an1n32x5 FILLER_132_2118 ();
 b15zdnd11an1n04x5 FILLER_132_2150 ();
 b15zdnd11an1n08x5 FILLER_132_2162 ();
 b15zdnd11an1n04x5 FILLER_132_2170 ();
 b15zdnd00an1n01x5 FILLER_132_2174 ();
 b15zdnd11an1n32x5 FILLER_132_2193 ();
 b15zdnd11an1n16x5 FILLER_132_2225 ();
 b15zdnd00an1n01x5 FILLER_132_2241 ();
 b15zdnd11an1n04x5 FILLER_132_2253 ();
 b15zdnd11an1n08x5 FILLER_132_2268 ();
 b15zdnd11an1n16x5 FILLER_133_0 ();
 b15zdnd00an1n01x5 FILLER_133_16 ();
 b15zdnd11an1n04x5 FILLER_133_21 ();
 b15zdnd00an1n02x5 FILLER_133_25 ();
 b15zdnd11an1n64x5 FILLER_133_69 ();
 b15zdnd11an1n04x5 FILLER_133_133 ();
 b15zdnd00an1n02x5 FILLER_133_137 ();
 b15zdnd00an1n01x5 FILLER_133_139 ();
 b15zdnd11an1n32x5 FILLER_133_192 ();
 b15zdnd11an1n08x5 FILLER_133_224 ();
 b15zdnd00an1n02x5 FILLER_133_232 ();
 b15zdnd11an1n64x5 FILLER_133_237 ();
 b15zdnd11an1n64x5 FILLER_133_301 ();
 b15zdnd11an1n64x5 FILLER_133_365 ();
 b15zdnd11an1n64x5 FILLER_133_429 ();
 b15zdnd11an1n32x5 FILLER_133_493 ();
 b15zdnd11an1n04x5 FILLER_133_525 ();
 b15zdnd11an1n64x5 FILLER_133_537 ();
 b15zdnd11an1n64x5 FILLER_133_601 ();
 b15zdnd11an1n64x5 FILLER_133_665 ();
 b15zdnd11an1n32x5 FILLER_133_729 ();
 b15zdnd11an1n16x5 FILLER_133_761 ();
 b15zdnd11an1n04x5 FILLER_133_777 ();
 b15zdnd00an1n02x5 FILLER_133_781 ();
 b15zdnd11an1n64x5 FILLER_133_814 ();
 b15zdnd11an1n64x5 FILLER_133_878 ();
 b15zdnd11an1n64x5 FILLER_133_942 ();
 b15zdnd11an1n64x5 FILLER_133_1006 ();
 b15zdnd11an1n64x5 FILLER_133_1070 ();
 b15zdnd11an1n64x5 FILLER_133_1134 ();
 b15zdnd11an1n64x5 FILLER_133_1198 ();
 b15zdnd11an1n32x5 FILLER_133_1262 ();
 b15zdnd11an1n16x5 FILLER_133_1294 ();
 b15zdnd11an1n08x5 FILLER_133_1310 ();
 b15zdnd00an1n02x5 FILLER_133_1318 ();
 b15zdnd00an1n01x5 FILLER_133_1320 ();
 b15zdnd11an1n32x5 FILLER_133_1333 ();
 b15zdnd11an1n04x5 FILLER_133_1365 ();
 b15zdnd00an1n01x5 FILLER_133_1369 ();
 b15zdnd11an1n64x5 FILLER_133_1392 ();
 b15zdnd11an1n64x5 FILLER_133_1456 ();
 b15zdnd11an1n32x5 FILLER_133_1520 ();
 b15zdnd00an1n02x5 FILLER_133_1552 ();
 b15zdnd00an1n01x5 FILLER_133_1554 ();
 b15zdnd11an1n32x5 FILLER_133_1607 ();
 b15zdnd00an1n02x5 FILLER_133_1639 ();
 b15zdnd00an1n01x5 FILLER_133_1641 ();
 b15zdnd11an1n64x5 FILLER_133_1694 ();
 b15zdnd11an1n64x5 FILLER_133_1758 ();
 b15zdnd11an1n64x5 FILLER_133_1822 ();
 b15zdnd11an1n64x5 FILLER_133_1886 ();
 b15zdnd11an1n64x5 FILLER_133_1950 ();
 b15zdnd11an1n64x5 FILLER_133_2014 ();
 b15zdnd11an1n64x5 FILLER_133_2078 ();
 b15zdnd11an1n64x5 FILLER_133_2142 ();
 b15zdnd11an1n64x5 FILLER_133_2206 ();
 b15zdnd11an1n08x5 FILLER_133_2270 ();
 b15zdnd11an1n04x5 FILLER_133_2278 ();
 b15zdnd00an1n02x5 FILLER_133_2282 ();
 b15zdnd11an1n16x5 FILLER_134_8 ();
 b15zdnd11an1n08x5 FILLER_134_24 ();
 b15zdnd00an1n01x5 FILLER_134_32 ();
 b15zdnd11an1n04x5 FILLER_134_85 ();
 b15zdnd11an1n04x5 FILLER_134_115 ();
 b15zdnd11an1n32x5 FILLER_134_124 ();
 b15zdnd00an1n02x5 FILLER_134_156 ();
 b15zdnd00an1n01x5 FILLER_134_158 ();
 b15zdnd11an1n04x5 FILLER_134_162 ();
 b15zdnd11an1n64x5 FILLER_134_169 ();
 b15zdnd11an1n08x5 FILLER_134_233 ();
 b15zdnd11an1n64x5 FILLER_134_246 ();
 b15zdnd11an1n64x5 FILLER_134_310 ();
 b15zdnd11an1n64x5 FILLER_134_374 ();
 b15zdnd11an1n64x5 FILLER_134_438 ();
 b15zdnd11an1n64x5 FILLER_134_502 ();
 b15zdnd11an1n64x5 FILLER_134_566 ();
 b15zdnd11an1n64x5 FILLER_134_630 ();
 b15zdnd11an1n16x5 FILLER_134_694 ();
 b15zdnd11an1n08x5 FILLER_134_710 ();
 b15zdnd11an1n64x5 FILLER_134_726 ();
 b15zdnd11an1n64x5 FILLER_134_790 ();
 b15zdnd11an1n64x5 FILLER_134_854 ();
 b15zdnd11an1n64x5 FILLER_134_918 ();
 b15zdnd11an1n64x5 FILLER_134_982 ();
 b15zdnd11an1n64x5 FILLER_134_1046 ();
 b15zdnd11an1n16x5 FILLER_134_1110 ();
 b15zdnd11an1n08x5 FILLER_134_1126 ();
 b15zdnd11an1n04x5 FILLER_134_1134 ();
 b15zdnd00an1n02x5 FILLER_134_1138 ();
 b15zdnd11an1n64x5 FILLER_134_1148 ();
 b15zdnd11an1n64x5 FILLER_134_1212 ();
 b15zdnd11an1n64x5 FILLER_134_1276 ();
 b15zdnd11an1n64x5 FILLER_134_1340 ();
 b15zdnd11an1n64x5 FILLER_134_1404 ();
 b15zdnd11an1n64x5 FILLER_134_1468 ();
 b15zdnd11an1n16x5 FILLER_134_1532 ();
 b15zdnd11an1n04x5 FILLER_134_1548 ();
 b15zdnd00an1n02x5 FILLER_134_1552 ();
 b15zdnd11an1n32x5 FILLER_134_1606 ();
 b15zdnd11an1n04x5 FILLER_134_1638 ();
 b15zdnd11an1n16x5 FILLER_134_1694 ();
 b15zdnd00an1n01x5 FILLER_134_1710 ();
 b15zdnd11an1n64x5 FILLER_134_1720 ();
 b15zdnd11an1n64x5 FILLER_134_1784 ();
 b15zdnd11an1n64x5 FILLER_134_1848 ();
 b15zdnd11an1n64x5 FILLER_134_1912 ();
 b15zdnd11an1n64x5 FILLER_134_1976 ();
 b15zdnd11an1n64x5 FILLER_134_2040 ();
 b15zdnd11an1n32x5 FILLER_134_2104 ();
 b15zdnd11an1n16x5 FILLER_134_2136 ();
 b15zdnd00an1n02x5 FILLER_134_2152 ();
 b15zdnd11an1n32x5 FILLER_134_2162 ();
 b15zdnd11an1n08x5 FILLER_134_2194 ();
 b15zdnd11an1n04x5 FILLER_134_2202 ();
 b15zdnd11an1n32x5 FILLER_134_2228 ();
 b15zdnd11an1n16x5 FILLER_134_2260 ();
 b15zdnd11an1n32x5 FILLER_135_0 ();
 b15zdnd11an1n16x5 FILLER_135_32 ();
 b15zdnd11an1n04x5 FILLER_135_48 ();
 b15zdnd00an1n02x5 FILLER_135_52 ();
 b15zdnd00an1n01x5 FILLER_135_54 ();
 b15zdnd11an1n16x5 FILLER_135_58 ();
 b15zdnd11an1n08x5 FILLER_135_74 ();
 b15zdnd11an1n04x5 FILLER_135_82 ();
 b15zdnd00an1n01x5 FILLER_135_86 ();
 b15zdnd11an1n64x5 FILLER_135_107 ();
 b15zdnd11an1n64x5 FILLER_135_171 ();
 b15zdnd11an1n64x5 FILLER_135_235 ();
 b15zdnd11an1n64x5 FILLER_135_299 ();
 b15zdnd11an1n64x5 FILLER_135_363 ();
 b15zdnd11an1n64x5 FILLER_135_427 ();
 b15zdnd11an1n64x5 FILLER_135_491 ();
 b15zdnd11an1n64x5 FILLER_135_555 ();
 b15zdnd11an1n64x5 FILLER_135_619 ();
 b15zdnd11an1n64x5 FILLER_135_683 ();
 b15zdnd11an1n64x5 FILLER_135_747 ();
 b15zdnd11an1n64x5 FILLER_135_811 ();
 b15zdnd11an1n64x5 FILLER_135_875 ();
 b15zdnd11an1n64x5 FILLER_135_939 ();
 b15zdnd11an1n64x5 FILLER_135_1003 ();
 b15zdnd11an1n64x5 FILLER_135_1067 ();
 b15zdnd11an1n32x5 FILLER_135_1131 ();
 b15zdnd11an1n16x5 FILLER_135_1163 ();
 b15zdnd11an1n08x5 FILLER_135_1179 ();
 b15zdnd11an1n04x5 FILLER_135_1187 ();
 b15zdnd00an1n02x5 FILLER_135_1191 ();
 b15zdnd11an1n16x5 FILLER_135_1206 ();
 b15zdnd11an1n04x5 FILLER_135_1222 ();
 b15zdnd11an1n64x5 FILLER_135_1238 ();
 b15zdnd11an1n64x5 FILLER_135_1302 ();
 b15zdnd11an1n64x5 FILLER_135_1366 ();
 b15zdnd11an1n64x5 FILLER_135_1430 ();
 b15zdnd11an1n64x5 FILLER_135_1494 ();
 b15zdnd11an1n08x5 FILLER_135_1558 ();
 b15zdnd11an1n04x5 FILLER_135_1566 ();
 b15zdnd00an1n02x5 FILLER_135_1570 ();
 b15zdnd00an1n01x5 FILLER_135_1572 ();
 b15zdnd11an1n04x5 FILLER_135_1576 ();
 b15zdnd11an1n04x5 FILLER_135_1583 ();
 b15zdnd11an1n64x5 FILLER_135_1590 ();
 b15zdnd11an1n04x5 FILLER_135_1654 ();
 b15zdnd00an1n02x5 FILLER_135_1658 ();
 b15zdnd11an1n04x5 FILLER_135_1663 ();
 b15zdnd11an1n04x5 FILLER_135_1670 ();
 b15zdnd11an1n32x5 FILLER_135_1677 ();
 b15zdnd00an1n01x5 FILLER_135_1709 ();
 b15zdnd11an1n64x5 FILLER_135_1719 ();
 b15zdnd11an1n64x5 FILLER_135_1783 ();
 b15zdnd11an1n64x5 FILLER_135_1847 ();
 b15zdnd11an1n64x5 FILLER_135_1911 ();
 b15zdnd11an1n64x5 FILLER_135_1975 ();
 b15zdnd11an1n16x5 FILLER_135_2039 ();
 b15zdnd00an1n01x5 FILLER_135_2055 ();
 b15zdnd11an1n64x5 FILLER_135_2060 ();
 b15zdnd11an1n64x5 FILLER_135_2124 ();
 b15zdnd11an1n64x5 FILLER_135_2188 ();
 b15zdnd11an1n32x5 FILLER_135_2252 ();
 b15zdnd11an1n64x5 FILLER_136_8 ();
 b15zdnd11an1n64x5 FILLER_136_72 ();
 b15zdnd11an1n64x5 FILLER_136_136 ();
 b15zdnd11an1n64x5 FILLER_136_200 ();
 b15zdnd11an1n64x5 FILLER_136_264 ();
 b15zdnd11an1n64x5 FILLER_136_328 ();
 b15zdnd11an1n64x5 FILLER_136_392 ();
 b15zdnd11an1n64x5 FILLER_136_456 ();
 b15zdnd11an1n32x5 FILLER_136_520 ();
 b15zdnd11an1n08x5 FILLER_136_552 ();
 b15zdnd11an1n04x5 FILLER_136_560 ();
 b15zdnd00an1n01x5 FILLER_136_564 ();
 b15zdnd11an1n64x5 FILLER_136_585 ();
 b15zdnd11an1n32x5 FILLER_136_649 ();
 b15zdnd00an1n02x5 FILLER_136_681 ();
 b15zdnd11an1n16x5 FILLER_136_689 ();
 b15zdnd11an1n08x5 FILLER_136_705 ();
 b15zdnd11an1n04x5 FILLER_136_713 ();
 b15zdnd00an1n01x5 FILLER_136_717 ();
 b15zdnd11an1n64x5 FILLER_136_726 ();
 b15zdnd11an1n64x5 FILLER_136_790 ();
 b15zdnd11an1n64x5 FILLER_136_854 ();
 b15zdnd11an1n32x5 FILLER_136_918 ();
 b15zdnd11an1n16x5 FILLER_136_950 ();
 b15zdnd00an1n01x5 FILLER_136_966 ();
 b15zdnd11an1n64x5 FILLER_136_981 ();
 b15zdnd11an1n64x5 FILLER_136_1045 ();
 b15zdnd11an1n64x5 FILLER_136_1109 ();
 b15zdnd11an1n16x5 FILLER_136_1173 ();
 b15zdnd11an1n04x5 FILLER_136_1189 ();
 b15zdnd00an1n02x5 FILLER_136_1193 ();
 b15zdnd11an1n16x5 FILLER_136_1211 ();
 b15zdnd11an1n04x5 FILLER_136_1227 ();
 b15zdnd11an1n64x5 FILLER_136_1241 ();
 b15zdnd11an1n16x5 FILLER_136_1305 ();
 b15zdnd11an1n08x5 FILLER_136_1321 ();
 b15zdnd11an1n64x5 FILLER_136_1349 ();
 b15zdnd11an1n04x5 FILLER_136_1413 ();
 b15zdnd11an1n32x5 FILLER_136_1431 ();
 b15zdnd11an1n08x5 FILLER_136_1463 ();
 b15zdnd11an1n04x5 FILLER_136_1471 ();
 b15zdnd00an1n01x5 FILLER_136_1475 ();
 b15zdnd11an1n64x5 FILLER_136_1485 ();
 b15zdnd11an1n16x5 FILLER_136_1549 ();
 b15zdnd11an1n08x5 FILLER_136_1565 ();
 b15zdnd00an1n01x5 FILLER_136_1573 ();
 b15zdnd11an1n04x5 FILLER_136_1577 ();
 b15zdnd11an1n04x5 FILLER_136_1584 ();
 b15zdnd11an1n64x5 FILLER_136_1591 ();
 b15zdnd11an1n08x5 FILLER_136_1655 ();
 b15zdnd11an1n04x5 FILLER_136_1663 ();
 b15zdnd11an1n32x5 FILLER_136_1670 ();
 b15zdnd00an1n02x5 FILLER_136_1702 ();
 b15zdnd00an1n01x5 FILLER_136_1704 ();
 b15zdnd11an1n64x5 FILLER_136_1714 ();
 b15zdnd11an1n32x5 FILLER_136_1778 ();
 b15zdnd11an1n16x5 FILLER_136_1810 ();
 b15zdnd11an1n08x5 FILLER_136_1826 ();
 b15zdnd11an1n04x5 FILLER_136_1834 ();
 b15zdnd11an1n04x5 FILLER_136_1850 ();
 b15zdnd11an1n64x5 FILLER_136_1868 ();
 b15zdnd11an1n64x5 FILLER_136_1932 ();
 b15zdnd11an1n32x5 FILLER_136_1996 ();
 b15zdnd11an1n16x5 FILLER_136_2028 ();
 b15zdnd11an1n04x5 FILLER_136_2044 ();
 b15zdnd00an1n02x5 FILLER_136_2048 ();
 b15zdnd00an1n01x5 FILLER_136_2050 ();
 b15zdnd11an1n04x5 FILLER_136_2055 ();
 b15zdnd11an1n04x5 FILLER_136_2065 ();
 b15zdnd11an1n64x5 FILLER_136_2073 ();
 b15zdnd11an1n16x5 FILLER_136_2137 ();
 b15zdnd00an1n01x5 FILLER_136_2153 ();
 b15zdnd11an1n16x5 FILLER_136_2162 ();
 b15zdnd11an1n04x5 FILLER_136_2178 ();
 b15zdnd00an1n01x5 FILLER_136_2182 ();
 b15zdnd11an1n16x5 FILLER_136_2186 ();
 b15zdnd11an1n08x5 FILLER_136_2202 ();
 b15zdnd11an1n04x5 FILLER_136_2210 ();
 b15zdnd11an1n04x5 FILLER_136_2228 ();
 b15zdnd11an1n32x5 FILLER_136_2244 ();
 b15zdnd11an1n64x5 FILLER_137_0 ();
 b15zdnd11an1n64x5 FILLER_137_64 ();
 b15zdnd11an1n64x5 FILLER_137_128 ();
 b15zdnd11an1n08x5 FILLER_137_192 ();
 b15zdnd11an1n32x5 FILLER_137_208 ();
 b15zdnd00an1n02x5 FILLER_137_240 ();
 b15zdnd11an1n16x5 FILLER_137_249 ();
 b15zdnd00an1n02x5 FILLER_137_265 ();
 b15zdnd00an1n01x5 FILLER_137_267 ();
 b15zdnd11an1n32x5 FILLER_137_282 ();
 b15zdnd11an1n08x5 FILLER_137_314 ();
 b15zdnd00an1n02x5 FILLER_137_322 ();
 b15zdnd00an1n01x5 FILLER_137_324 ();
 b15zdnd11an1n64x5 FILLER_137_346 ();
 b15zdnd11an1n64x5 FILLER_137_410 ();
 b15zdnd11an1n64x5 FILLER_137_474 ();
 b15zdnd11an1n64x5 FILLER_137_538 ();
 b15zdnd11an1n64x5 FILLER_137_602 ();
 b15zdnd11an1n64x5 FILLER_137_666 ();
 b15zdnd11an1n64x5 FILLER_137_730 ();
 b15zdnd11an1n64x5 FILLER_137_794 ();
 b15zdnd11an1n64x5 FILLER_137_858 ();
 b15zdnd11an1n16x5 FILLER_137_922 ();
 b15zdnd11an1n08x5 FILLER_137_938 ();
 b15zdnd11an1n04x5 FILLER_137_946 ();
 b15zdnd11an1n04x5 FILLER_137_967 ();
 b15zdnd11an1n04x5 FILLER_137_978 ();
 b15zdnd11an1n64x5 FILLER_137_997 ();
 b15zdnd11an1n64x5 FILLER_137_1061 ();
 b15zdnd11an1n08x5 FILLER_137_1125 ();
 b15zdnd11an1n04x5 FILLER_137_1133 ();
 b15zdnd11an1n32x5 FILLER_137_1146 ();
 b15zdnd11an1n08x5 FILLER_137_1178 ();
 b15zdnd11an1n04x5 FILLER_137_1186 ();
 b15zdnd00an1n02x5 FILLER_137_1190 ();
 b15zdnd00an1n01x5 FILLER_137_1192 ();
 b15zdnd11an1n64x5 FILLER_137_1207 ();
 b15zdnd11an1n64x5 FILLER_137_1271 ();
 b15zdnd11an1n64x5 FILLER_137_1335 ();
 b15zdnd11an1n08x5 FILLER_137_1399 ();
 b15zdnd11an1n04x5 FILLER_137_1407 ();
 b15zdnd11an1n64x5 FILLER_137_1443 ();
 b15zdnd11an1n64x5 FILLER_137_1507 ();
 b15zdnd11an1n64x5 FILLER_137_1571 ();
 b15zdnd11an1n64x5 FILLER_137_1635 ();
 b15zdnd11an1n32x5 FILLER_137_1699 ();
 b15zdnd11an1n64x5 FILLER_137_1740 ();
 b15zdnd11an1n04x5 FILLER_137_1804 ();
 b15zdnd11an1n04x5 FILLER_137_1824 ();
 b15zdnd00an1n02x5 FILLER_137_1828 ();
 b15zdnd11an1n08x5 FILLER_137_1846 ();
 b15zdnd11an1n04x5 FILLER_137_1854 ();
 b15zdnd00an1n02x5 FILLER_137_1858 ();
 b15zdnd00an1n01x5 FILLER_137_1860 ();
 b15zdnd11an1n04x5 FILLER_137_1864 ();
 b15zdnd11an1n16x5 FILLER_137_1882 ();
 b15zdnd11an1n08x5 FILLER_137_1898 ();
 b15zdnd11an1n04x5 FILLER_137_1906 ();
 b15zdnd00an1n01x5 FILLER_137_1910 ();
 b15zdnd11an1n64x5 FILLER_137_1914 ();
 b15zdnd11an1n64x5 FILLER_137_1978 ();
 b15zdnd00an1n02x5 FILLER_137_2042 ();
 b15zdnd11an1n64x5 FILLER_137_2048 ();
 b15zdnd11an1n32x5 FILLER_137_2112 ();
 b15zdnd11an1n08x5 FILLER_137_2144 ();
 b15zdnd11an1n04x5 FILLER_137_2152 ();
 b15zdnd00an1n01x5 FILLER_137_2156 ();
 b15zdnd11an1n04x5 FILLER_137_2209 ();
 b15zdnd00an1n01x5 FILLER_137_2213 ();
 b15zdnd11an1n32x5 FILLER_137_2225 ();
 b15zdnd11an1n16x5 FILLER_137_2257 ();
 b15zdnd11an1n08x5 FILLER_137_2273 ();
 b15zdnd00an1n02x5 FILLER_137_2281 ();
 b15zdnd00an1n01x5 FILLER_137_2283 ();
 b15zdnd11an1n64x5 FILLER_138_8 ();
 b15zdnd00an1n02x5 FILLER_138_72 ();
 b15zdnd00an1n01x5 FILLER_138_74 ();
 b15zdnd11an1n64x5 FILLER_138_95 ();
 b15zdnd11an1n64x5 FILLER_138_159 ();
 b15zdnd11an1n64x5 FILLER_138_223 ();
 b15zdnd11an1n08x5 FILLER_138_287 ();
 b15zdnd00an1n02x5 FILLER_138_295 ();
 b15zdnd11an1n64x5 FILLER_138_304 ();
 b15zdnd11an1n64x5 FILLER_138_368 ();
 b15zdnd11an1n64x5 FILLER_138_432 ();
 b15zdnd11an1n64x5 FILLER_138_496 ();
 b15zdnd11an1n64x5 FILLER_138_560 ();
 b15zdnd11an1n64x5 FILLER_138_624 ();
 b15zdnd11an1n16x5 FILLER_138_688 ();
 b15zdnd11an1n08x5 FILLER_138_704 ();
 b15zdnd11an1n04x5 FILLER_138_712 ();
 b15zdnd00an1n02x5 FILLER_138_716 ();
 b15zdnd11an1n64x5 FILLER_138_726 ();
 b15zdnd11an1n64x5 FILLER_138_790 ();
 b15zdnd11an1n64x5 FILLER_138_854 ();
 b15zdnd11an1n16x5 FILLER_138_918 ();
 b15zdnd11an1n04x5 FILLER_138_934 ();
 b15zdnd11an1n32x5 FILLER_138_969 ();
 b15zdnd11an1n16x5 FILLER_138_1001 ();
 b15zdnd00an1n01x5 FILLER_138_1017 ();
 b15zdnd11an1n64x5 FILLER_138_1049 ();
 b15zdnd11an1n08x5 FILLER_138_1113 ();
 b15zdnd11an1n04x5 FILLER_138_1121 ();
 b15zdnd00an1n02x5 FILLER_138_1125 ();
 b15zdnd00an1n01x5 FILLER_138_1127 ();
 b15zdnd11an1n04x5 FILLER_138_1152 ();
 b15zdnd11an1n64x5 FILLER_138_1165 ();
 b15zdnd11an1n64x5 FILLER_138_1229 ();
 b15zdnd11an1n64x5 FILLER_138_1293 ();
 b15zdnd11an1n64x5 FILLER_138_1357 ();
 b15zdnd11an1n64x5 FILLER_138_1421 ();
 b15zdnd11an1n64x5 FILLER_138_1485 ();
 b15zdnd11an1n64x5 FILLER_138_1549 ();
 b15zdnd11an1n64x5 FILLER_138_1613 ();
 b15zdnd11an1n64x5 FILLER_138_1677 ();
 b15zdnd11an1n08x5 FILLER_138_1741 ();
 b15zdnd11an1n04x5 FILLER_138_1749 ();
 b15zdnd00an1n02x5 FILLER_138_1753 ();
 b15zdnd00an1n01x5 FILLER_138_1755 ();
 b15zdnd11an1n32x5 FILLER_138_1798 ();
 b15zdnd11an1n64x5 FILLER_138_1833 ();
 b15zdnd11an1n32x5 FILLER_138_1897 ();
 b15zdnd11an1n08x5 FILLER_138_1929 ();
 b15zdnd11an1n04x5 FILLER_138_1937 ();
 b15zdnd00an1n02x5 FILLER_138_1941 ();
 b15zdnd00an1n01x5 FILLER_138_1943 ();
 b15zdnd11an1n16x5 FILLER_138_1958 ();
 b15zdnd11an1n04x5 FILLER_138_2016 ();
 b15zdnd11an1n64x5 FILLER_138_2034 ();
 b15zdnd11an1n32x5 FILLER_138_2098 ();
 b15zdnd11an1n16x5 FILLER_138_2130 ();
 b15zdnd11an1n08x5 FILLER_138_2146 ();
 b15zdnd11an1n16x5 FILLER_138_2162 ();
 b15zdnd11an1n04x5 FILLER_138_2178 ();
 b15zdnd11an1n64x5 FILLER_138_2185 ();
 b15zdnd11an1n16x5 FILLER_138_2249 ();
 b15zdnd11an1n08x5 FILLER_138_2265 ();
 b15zdnd00an1n02x5 FILLER_138_2273 ();
 b15zdnd00an1n01x5 FILLER_138_2275 ();
 b15zdnd11an1n64x5 FILLER_139_0 ();
 b15zdnd11an1n64x5 FILLER_139_64 ();
 b15zdnd11an1n16x5 FILLER_139_128 ();
 b15zdnd11an1n04x5 FILLER_139_144 ();
 b15zdnd00an1n02x5 FILLER_139_148 ();
 b15zdnd00an1n01x5 FILLER_139_150 ();
 b15zdnd11an1n64x5 FILLER_139_193 ();
 b15zdnd11an1n16x5 FILLER_139_257 ();
 b15zdnd11an1n04x5 FILLER_139_273 ();
 b15zdnd00an1n02x5 FILLER_139_277 ();
 b15zdnd00an1n01x5 FILLER_139_279 ();
 b15zdnd11an1n16x5 FILLER_139_285 ();
 b15zdnd11an1n08x5 FILLER_139_301 ();
 b15zdnd00an1n01x5 FILLER_139_309 ();
 b15zdnd11an1n64x5 FILLER_139_320 ();
 b15zdnd11an1n64x5 FILLER_139_384 ();
 b15zdnd11an1n64x5 FILLER_139_448 ();
 b15zdnd11an1n32x5 FILLER_139_512 ();
 b15zdnd11an1n16x5 FILLER_139_544 ();
 b15zdnd11an1n08x5 FILLER_139_560 ();
 b15zdnd00an1n01x5 FILLER_139_568 ();
 b15zdnd11an1n04x5 FILLER_139_585 ();
 b15zdnd11an1n64x5 FILLER_139_603 ();
 b15zdnd11an1n64x5 FILLER_139_667 ();
 b15zdnd11an1n16x5 FILLER_139_731 ();
 b15zdnd11an1n04x5 FILLER_139_747 ();
 b15zdnd00an1n02x5 FILLER_139_751 ();
 b15zdnd11an1n64x5 FILLER_139_760 ();
 b15zdnd11an1n64x5 FILLER_139_824 ();
 b15zdnd11an1n64x5 FILLER_139_888 ();
 b15zdnd11an1n32x5 FILLER_139_952 ();
 b15zdnd00an1n02x5 FILLER_139_984 ();
 b15zdnd11an1n64x5 FILLER_139_995 ();
 b15zdnd11an1n16x5 FILLER_139_1059 ();
 b15zdnd11an1n08x5 FILLER_139_1075 ();
 b15zdnd00an1n02x5 FILLER_139_1083 ();
 b15zdnd00an1n01x5 FILLER_139_1085 ();
 b15zdnd11an1n08x5 FILLER_139_1100 ();
 b15zdnd11an1n04x5 FILLER_139_1108 ();
 b15zdnd00an1n01x5 FILLER_139_1112 ();
 b15zdnd11an1n64x5 FILLER_139_1122 ();
 b15zdnd11an1n64x5 FILLER_139_1186 ();
 b15zdnd11an1n64x5 FILLER_139_1250 ();
 b15zdnd11an1n64x5 FILLER_139_1314 ();
 b15zdnd11an1n32x5 FILLER_139_1378 ();
 b15zdnd11an1n08x5 FILLER_139_1410 ();
 b15zdnd00an1n02x5 FILLER_139_1418 ();
 b15zdnd11an1n64x5 FILLER_139_1431 ();
 b15zdnd11an1n64x5 FILLER_139_1495 ();
 b15zdnd11an1n64x5 FILLER_139_1559 ();
 b15zdnd11an1n64x5 FILLER_139_1623 ();
 b15zdnd11an1n64x5 FILLER_139_1687 ();
 b15zdnd11an1n32x5 FILLER_139_1751 ();
 b15zdnd11an1n08x5 FILLER_139_1783 ();
 b15zdnd00an1n01x5 FILLER_139_1791 ();
 b15zdnd11an1n04x5 FILLER_139_1808 ();
 b15zdnd00an1n02x5 FILLER_139_1812 ();
 b15zdnd11an1n04x5 FILLER_139_1827 ();
 b15zdnd11an1n04x5 FILLER_139_1844 ();
 b15zdnd11an1n64x5 FILLER_139_1851 ();
 b15zdnd11an1n16x5 FILLER_139_1915 ();
 b15zdnd11an1n04x5 FILLER_139_1931 ();
 b15zdnd00an1n02x5 FILLER_139_1935 ();
 b15zdnd00an1n01x5 FILLER_139_1937 ();
 b15zdnd11an1n16x5 FILLER_139_1980 ();
 b15zdnd11an1n04x5 FILLER_139_1996 ();
 b15zdnd00an1n01x5 FILLER_139_2000 ();
 b15zdnd11an1n08x5 FILLER_139_2045 ();
 b15zdnd11an1n04x5 FILLER_139_2053 ();
 b15zdnd00an1n01x5 FILLER_139_2057 ();
 b15zdnd11an1n64x5 FILLER_139_2062 ();
 b15zdnd11an1n32x5 FILLER_139_2126 ();
 b15zdnd11an1n16x5 FILLER_139_2158 ();
 b15zdnd11an1n04x5 FILLER_139_2174 ();
 b15zdnd00an1n02x5 FILLER_139_2178 ();
 b15zdnd00an1n01x5 FILLER_139_2180 ();
 b15zdnd11an1n16x5 FILLER_139_2184 ();
 b15zdnd11an1n04x5 FILLER_139_2200 ();
 b15zdnd00an1n02x5 FILLER_139_2204 ();
 b15zdnd11an1n04x5 FILLER_139_2248 ();
 b15zdnd00an1n02x5 FILLER_139_2252 ();
 b15zdnd11an1n16x5 FILLER_139_2265 ();
 b15zdnd00an1n02x5 FILLER_139_2281 ();
 b15zdnd00an1n01x5 FILLER_139_2283 ();
 b15zdnd11an1n32x5 FILLER_140_8 ();
 b15zdnd11an1n16x5 FILLER_140_40 ();
 b15zdnd11an1n08x5 FILLER_140_56 ();
 b15zdnd00an1n02x5 FILLER_140_64 ();
 b15zdnd00an1n01x5 FILLER_140_66 ();
 b15zdnd11an1n32x5 FILLER_140_81 ();
 b15zdnd11an1n08x5 FILLER_140_113 ();
 b15zdnd00an1n02x5 FILLER_140_121 ();
 b15zdnd00an1n01x5 FILLER_140_123 ();
 b15zdnd11an1n32x5 FILLER_140_139 ();
 b15zdnd11an1n16x5 FILLER_140_171 ();
 b15zdnd11an1n04x5 FILLER_140_187 ();
 b15zdnd00an1n01x5 FILLER_140_191 ();
 b15zdnd11an1n64x5 FILLER_140_202 ();
 b15zdnd11an1n32x5 FILLER_140_266 ();
 b15zdnd11an1n16x5 FILLER_140_298 ();
 b15zdnd11an1n08x5 FILLER_140_314 ();
 b15zdnd00an1n02x5 FILLER_140_322 ();
 b15zdnd11an1n64x5 FILLER_140_333 ();
 b15zdnd11an1n64x5 FILLER_140_397 ();
 b15zdnd11an1n64x5 FILLER_140_461 ();
 b15zdnd11an1n16x5 FILLER_140_525 ();
 b15zdnd11an1n08x5 FILLER_140_541 ();
 b15zdnd00an1n02x5 FILLER_140_549 ();
 b15zdnd11an1n04x5 FILLER_140_564 ();
 b15zdnd11an1n04x5 FILLER_140_580 ();
 b15zdnd00an1n02x5 FILLER_140_584 ();
 b15zdnd11an1n64x5 FILLER_140_618 ();
 b15zdnd11an1n32x5 FILLER_140_682 ();
 b15zdnd11an1n04x5 FILLER_140_714 ();
 b15zdnd11an1n08x5 FILLER_140_726 ();
 b15zdnd00an1n02x5 FILLER_140_734 ();
 b15zdnd11an1n64x5 FILLER_140_767 ();
 b15zdnd00an1n02x5 FILLER_140_831 ();
 b15zdnd00an1n01x5 FILLER_140_833 ();
 b15zdnd11an1n08x5 FILLER_140_879 ();
 b15zdnd11an1n04x5 FILLER_140_887 ();
 b15zdnd00an1n02x5 FILLER_140_891 ();
 b15zdnd11an1n64x5 FILLER_140_913 ();
 b15zdnd11an1n64x5 FILLER_140_977 ();
 b15zdnd11an1n16x5 FILLER_140_1041 ();
 b15zdnd00an1n02x5 FILLER_140_1057 ();
 b15zdnd00an1n01x5 FILLER_140_1059 ();
 b15zdnd11an1n04x5 FILLER_140_1077 ();
 b15zdnd11an1n64x5 FILLER_140_1091 ();
 b15zdnd11an1n04x5 FILLER_140_1155 ();
 b15zdnd00an1n01x5 FILLER_140_1159 ();
 b15zdnd11an1n32x5 FILLER_140_1171 ();
 b15zdnd11an1n16x5 FILLER_140_1203 ();
 b15zdnd11an1n04x5 FILLER_140_1219 ();
 b15zdnd11an1n64x5 FILLER_140_1239 ();
 b15zdnd11an1n16x5 FILLER_140_1303 ();
 b15zdnd11an1n08x5 FILLER_140_1319 ();
 b15zdnd00an1n02x5 FILLER_140_1327 ();
 b15zdnd11an1n64x5 FILLER_140_1346 ();
 b15zdnd11an1n16x5 FILLER_140_1410 ();
 b15zdnd11an1n04x5 FILLER_140_1426 ();
 b15zdnd11an1n64x5 FILLER_140_1433 ();
 b15zdnd11an1n64x5 FILLER_140_1497 ();
 b15zdnd11an1n64x5 FILLER_140_1561 ();
 b15zdnd11an1n64x5 FILLER_140_1625 ();
 b15zdnd11an1n64x5 FILLER_140_1689 ();
 b15zdnd11an1n64x5 FILLER_140_1753 ();
 b15zdnd11an1n64x5 FILLER_140_1817 ();
 b15zdnd11an1n32x5 FILLER_140_1881 ();
 b15zdnd11an1n16x5 FILLER_140_1913 ();
 b15zdnd00an1n02x5 FILLER_140_1929 ();
 b15zdnd11an1n16x5 FILLER_140_1945 ();
 b15zdnd11an1n04x5 FILLER_140_1961 ();
 b15zdnd11an1n04x5 FILLER_140_1968 ();
 b15zdnd11an1n16x5 FILLER_140_1975 ();
 b15zdnd11an1n08x5 FILLER_140_1991 ();
 b15zdnd11an1n08x5 FILLER_140_2007 ();
 b15zdnd11an1n04x5 FILLER_140_2018 ();
 b15zdnd11an1n04x5 FILLER_140_2025 ();
 b15zdnd11an1n64x5 FILLER_140_2032 ();
 b15zdnd11an1n16x5 FILLER_140_2096 ();
 b15zdnd11an1n04x5 FILLER_140_2112 ();
 b15zdnd00an1n01x5 FILLER_140_2116 ();
 b15zdnd11an1n16x5 FILLER_140_2127 ();
 b15zdnd11an1n08x5 FILLER_140_2143 ();
 b15zdnd00an1n02x5 FILLER_140_2151 ();
 b15zdnd00an1n01x5 FILLER_140_2153 ();
 b15zdnd11an1n32x5 FILLER_140_2162 ();
 b15zdnd11an1n04x5 FILLER_140_2194 ();
 b15zdnd00an1n02x5 FILLER_140_2198 ();
 b15zdnd11an1n16x5 FILLER_140_2214 ();
 b15zdnd11an1n08x5 FILLER_140_2230 ();
 b15zdnd11an1n04x5 FILLER_140_2238 ();
 b15zdnd11an1n16x5 FILLER_140_2253 ();
 b15zdnd11an1n04x5 FILLER_140_2269 ();
 b15zdnd00an1n02x5 FILLER_140_2273 ();
 b15zdnd00an1n01x5 FILLER_140_2275 ();
 b15zdnd11an1n64x5 FILLER_141_0 ();
 b15zdnd11an1n08x5 FILLER_141_64 ();
 b15zdnd11an1n04x5 FILLER_141_72 ();
 b15zdnd11an1n64x5 FILLER_141_96 ();
 b15zdnd11an1n32x5 FILLER_141_160 ();
 b15zdnd11an1n08x5 FILLER_141_192 ();
 b15zdnd00an1n01x5 FILLER_141_200 ();
 b15zdnd11an1n64x5 FILLER_141_243 ();
 b15zdnd11an1n64x5 FILLER_141_307 ();
 b15zdnd11an1n64x5 FILLER_141_371 ();
 b15zdnd11an1n64x5 FILLER_141_435 ();
 b15zdnd11an1n04x5 FILLER_141_499 ();
 b15zdnd00an1n02x5 FILLER_141_503 ();
 b15zdnd11an1n04x5 FILLER_141_519 ();
 b15zdnd11an1n08x5 FILLER_141_531 ();
 b15zdnd11an1n04x5 FILLER_141_539 ();
 b15zdnd11an1n04x5 FILLER_141_546 ();
 b15zdnd11an1n16x5 FILLER_141_560 ();
 b15zdnd11an1n64x5 FILLER_141_596 ();
 b15zdnd11an1n64x5 FILLER_141_660 ();
 b15zdnd11an1n64x5 FILLER_141_724 ();
 b15zdnd11an1n64x5 FILLER_141_788 ();
 b15zdnd11an1n64x5 FILLER_141_852 ();
 b15zdnd11an1n04x5 FILLER_141_916 ();
 b15zdnd00an1n02x5 FILLER_141_920 ();
 b15zdnd11an1n16x5 FILLER_141_938 ();
 b15zdnd11an1n08x5 FILLER_141_954 ();
 b15zdnd11an1n04x5 FILLER_141_962 ();
 b15zdnd11an1n32x5 FILLER_141_975 ();
 b15zdnd11an1n16x5 FILLER_141_1007 ();
 b15zdnd11an1n08x5 FILLER_141_1023 ();
 b15zdnd00an1n02x5 FILLER_141_1031 ();
 b15zdnd11an1n04x5 FILLER_141_1040 ();
 b15zdnd00an1n01x5 FILLER_141_1044 ();
 b15zdnd11an1n08x5 FILLER_141_1057 ();
 b15zdnd00an1n01x5 FILLER_141_1065 ();
 b15zdnd11an1n16x5 FILLER_141_1097 ();
 b15zdnd11an1n08x5 FILLER_141_1113 ();
 b15zdnd00an1n01x5 FILLER_141_1121 ();
 b15zdnd11an1n16x5 FILLER_141_1131 ();
 b15zdnd11an1n08x5 FILLER_141_1147 ();
 b15zdnd00an1n02x5 FILLER_141_1155 ();
 b15zdnd11an1n64x5 FILLER_141_1166 ();
 b15zdnd11an1n16x5 FILLER_141_1230 ();
 b15zdnd11an1n16x5 FILLER_141_1260 ();
 b15zdnd11an1n08x5 FILLER_141_1276 ();
 b15zdnd00an1n02x5 FILLER_141_1284 ();
 b15zdnd00an1n01x5 FILLER_141_1286 ();
 b15zdnd11an1n04x5 FILLER_141_1304 ();
 b15zdnd11an1n64x5 FILLER_141_1328 ();
 b15zdnd11an1n32x5 FILLER_141_1392 ();
 b15zdnd11an1n04x5 FILLER_141_1424 ();
 b15zdnd00an1n01x5 FILLER_141_1428 ();
 b15zdnd11an1n04x5 FILLER_141_1432 ();
 b15zdnd11an1n64x5 FILLER_141_1439 ();
 b15zdnd11an1n08x5 FILLER_141_1503 ();
 b15zdnd00an1n01x5 FILLER_141_1511 ();
 b15zdnd11an1n64x5 FILLER_141_1518 ();
 b15zdnd11an1n64x5 FILLER_141_1582 ();
 b15zdnd11an1n64x5 FILLER_141_1646 ();
 b15zdnd11an1n64x5 FILLER_141_1710 ();
 b15zdnd11an1n64x5 FILLER_141_1774 ();
 b15zdnd11an1n64x5 FILLER_141_1838 ();
 b15zdnd11an1n64x5 FILLER_141_1902 ();
 b15zdnd11an1n64x5 FILLER_141_1966 ();
 b15zdnd11an1n64x5 FILLER_141_2030 ();
 b15zdnd11an1n64x5 FILLER_141_2094 ();
 b15zdnd11an1n64x5 FILLER_141_2158 ();
 b15zdnd11an1n32x5 FILLER_141_2222 ();
 b15zdnd11an1n16x5 FILLER_141_2254 ();
 b15zdnd11an1n08x5 FILLER_141_2270 ();
 b15zdnd11an1n04x5 FILLER_141_2278 ();
 b15zdnd00an1n02x5 FILLER_141_2282 ();
 b15zdnd11an1n64x5 FILLER_142_8 ();
 b15zdnd11an1n64x5 FILLER_142_72 ();
 b15zdnd11an1n64x5 FILLER_142_136 ();
 b15zdnd11an1n32x5 FILLER_142_200 ();
 b15zdnd11an1n04x5 FILLER_142_232 ();
 b15zdnd11an1n64x5 FILLER_142_252 ();
 b15zdnd11an1n64x5 FILLER_142_316 ();
 b15zdnd11an1n64x5 FILLER_142_380 ();
 b15zdnd11an1n64x5 FILLER_142_444 ();
 b15zdnd11an1n16x5 FILLER_142_508 ();
 b15zdnd00an1n02x5 FILLER_142_524 ();
 b15zdnd11an1n04x5 FILLER_142_532 ();
 b15zdnd00an1n02x5 FILLER_142_536 ();
 b15zdnd00an1n01x5 FILLER_142_538 ();
 b15zdnd11an1n04x5 FILLER_142_545 ();
 b15zdnd00an1n02x5 FILLER_142_549 ();
 b15zdnd00an1n01x5 FILLER_142_551 ();
 b15zdnd11an1n16x5 FILLER_142_555 ();
 b15zdnd11an1n08x5 FILLER_142_571 ();
 b15zdnd00an1n02x5 FILLER_142_579 ();
 b15zdnd00an1n01x5 FILLER_142_581 ();
 b15zdnd11an1n64x5 FILLER_142_596 ();
 b15zdnd11an1n04x5 FILLER_142_660 ();
 b15zdnd00an1n02x5 FILLER_142_664 ();
 b15zdnd00an1n01x5 FILLER_142_666 ();
 b15zdnd11an1n16x5 FILLER_142_678 ();
 b15zdnd11an1n04x5 FILLER_142_694 ();
 b15zdnd11an1n08x5 FILLER_142_710 ();
 b15zdnd11an1n64x5 FILLER_142_726 ();
 b15zdnd11an1n04x5 FILLER_142_790 ();
 b15zdnd00an1n02x5 FILLER_142_794 ();
 b15zdnd11an1n08x5 FILLER_142_820 ();
 b15zdnd00an1n02x5 FILLER_142_828 ();
 b15zdnd11an1n32x5 FILLER_142_838 ();
 b15zdnd11an1n16x5 FILLER_142_870 ();
 b15zdnd11an1n04x5 FILLER_142_886 ();
 b15zdnd00an1n02x5 FILLER_142_890 ();
 b15zdnd00an1n01x5 FILLER_142_892 ();
 b15zdnd11an1n16x5 FILLER_142_902 ();
 b15zdnd00an1n01x5 FILLER_142_918 ();
 b15zdnd11an1n64x5 FILLER_142_930 ();
 b15zdnd11an1n32x5 FILLER_142_994 ();
 b15zdnd11an1n16x5 FILLER_142_1026 ();
 b15zdnd11an1n08x5 FILLER_142_1042 ();
 b15zdnd00an1n02x5 FILLER_142_1050 ();
 b15zdnd11an1n04x5 FILLER_142_1083 ();
 b15zdnd11an1n64x5 FILLER_142_1101 ();
 b15zdnd11an1n64x5 FILLER_142_1165 ();
 b15zdnd11an1n04x5 FILLER_142_1229 ();
 b15zdnd00an1n02x5 FILLER_142_1233 ();
 b15zdnd11an1n32x5 FILLER_142_1247 ();
 b15zdnd11an1n08x5 FILLER_142_1279 ();
 b15zdnd11an1n04x5 FILLER_142_1287 ();
 b15zdnd00an1n02x5 FILLER_142_1291 ();
 b15zdnd11an1n64x5 FILLER_142_1313 ();
 b15zdnd11an1n32x5 FILLER_142_1377 ();
 b15zdnd00an1n01x5 FILLER_142_1409 ();
 b15zdnd11an1n32x5 FILLER_142_1462 ();
 b15zdnd11an1n16x5 FILLER_142_1494 ();
 b15zdnd11an1n04x5 FILLER_142_1510 ();
 b15zdnd00an1n02x5 FILLER_142_1514 ();
 b15zdnd11an1n64x5 FILLER_142_1522 ();
 b15zdnd11an1n64x5 FILLER_142_1586 ();
 b15zdnd11an1n64x5 FILLER_142_1650 ();
 b15zdnd11an1n64x5 FILLER_142_1714 ();
 b15zdnd11an1n64x5 FILLER_142_1778 ();
 b15zdnd11an1n16x5 FILLER_142_1842 ();
 b15zdnd11an1n04x5 FILLER_142_1858 ();
 b15zdnd11an1n64x5 FILLER_142_1869 ();
 b15zdnd11an1n64x5 FILLER_142_1933 ();
 b15zdnd11an1n64x5 FILLER_142_1997 ();
 b15zdnd11an1n64x5 FILLER_142_2061 ();
 b15zdnd11an1n16x5 FILLER_142_2125 ();
 b15zdnd11an1n08x5 FILLER_142_2141 ();
 b15zdnd11an1n04x5 FILLER_142_2149 ();
 b15zdnd00an1n01x5 FILLER_142_2153 ();
 b15zdnd11an1n32x5 FILLER_142_2162 ();
 b15zdnd11an1n08x5 FILLER_142_2194 ();
 b15zdnd00an1n02x5 FILLER_142_2202 ();
 b15zdnd00an1n01x5 FILLER_142_2204 ();
 b15zdnd11an1n32x5 FILLER_142_2223 ();
 b15zdnd11an1n16x5 FILLER_142_2255 ();
 b15zdnd11an1n04x5 FILLER_142_2271 ();
 b15zdnd00an1n01x5 FILLER_142_2275 ();
 b15zdnd11an1n64x5 FILLER_143_0 ();
 b15zdnd11an1n32x5 FILLER_143_64 ();
 b15zdnd11an1n16x5 FILLER_143_96 ();
 b15zdnd11an1n04x5 FILLER_143_112 ();
 b15zdnd00an1n02x5 FILLER_143_116 ();
 b15zdnd00an1n01x5 FILLER_143_118 ();
 b15zdnd11an1n64x5 FILLER_143_161 ();
 b15zdnd11an1n64x5 FILLER_143_225 ();
 b15zdnd11an1n64x5 FILLER_143_289 ();
 b15zdnd11an1n16x5 FILLER_143_353 ();
 b15zdnd00an1n02x5 FILLER_143_369 ();
 b15zdnd11an1n64x5 FILLER_143_382 ();
 b15zdnd11an1n64x5 FILLER_143_446 ();
 b15zdnd11an1n08x5 FILLER_143_510 ();
 b15zdnd00an1n01x5 FILLER_143_518 ();
 b15zdnd11an1n04x5 FILLER_143_526 ();
 b15zdnd11an1n08x5 FILLER_143_537 ();
 b15zdnd00an1n01x5 FILLER_143_545 ();
 b15zdnd11an1n64x5 FILLER_143_552 ();
 b15zdnd00an1n02x5 FILLER_143_616 ();
 b15zdnd11an1n32x5 FILLER_143_624 ();
 b15zdnd11an1n08x5 FILLER_143_656 ();
 b15zdnd00an1n02x5 FILLER_143_664 ();
 b15zdnd00an1n01x5 FILLER_143_666 ();
 b15zdnd11an1n64x5 FILLER_143_670 ();
 b15zdnd11an1n32x5 FILLER_143_734 ();
 b15zdnd11an1n16x5 FILLER_143_766 ();
 b15zdnd11an1n04x5 FILLER_143_782 ();
 b15zdnd00an1n01x5 FILLER_143_786 ();
 b15zdnd11an1n04x5 FILLER_143_790 ();
 b15zdnd11an1n08x5 FILLER_143_807 ();
 b15zdnd00an1n02x5 FILLER_143_815 ();
 b15zdnd11an1n04x5 FILLER_143_820 ();
 b15zdnd00an1n02x5 FILLER_143_824 ();
 b15zdnd00an1n01x5 FILLER_143_826 ();
 b15zdnd11an1n64x5 FILLER_143_835 ();
 b15zdnd00an1n02x5 FILLER_143_899 ();
 b15zdnd11an1n04x5 FILLER_143_910 ();
 b15zdnd11an1n64x5 FILLER_143_925 ();
 b15zdnd11an1n64x5 FILLER_143_989 ();
 b15zdnd11an1n32x5 FILLER_143_1053 ();
 b15zdnd11an1n16x5 FILLER_143_1085 ();
 b15zdnd11an1n08x5 FILLER_143_1101 ();
 b15zdnd00an1n02x5 FILLER_143_1109 ();
 b15zdnd00an1n01x5 FILLER_143_1111 ();
 b15zdnd11an1n64x5 FILLER_143_1128 ();
 b15zdnd11an1n64x5 FILLER_143_1192 ();
 b15zdnd11an1n32x5 FILLER_143_1256 ();
 b15zdnd11an1n08x5 FILLER_143_1288 ();
 b15zdnd00an1n02x5 FILLER_143_1296 ();
 b15zdnd00an1n01x5 FILLER_143_1298 ();
 b15zdnd11an1n08x5 FILLER_143_1316 ();
 b15zdnd11an1n04x5 FILLER_143_1324 ();
 b15zdnd00an1n02x5 FILLER_143_1328 ();
 b15zdnd00an1n01x5 FILLER_143_1330 ();
 b15zdnd11an1n64x5 FILLER_143_1338 ();
 b15zdnd11an1n64x5 FILLER_143_1402 ();
 b15zdnd11an1n32x5 FILLER_143_1466 ();
 b15zdnd11an1n04x5 FILLER_143_1498 ();
 b15zdnd00an1n02x5 FILLER_143_1502 ();
 b15zdnd11an1n04x5 FILLER_143_1525 ();
 b15zdnd11an1n64x5 FILLER_143_1546 ();
 b15zdnd11an1n64x5 FILLER_143_1610 ();
 b15zdnd11an1n64x5 FILLER_143_1674 ();
 b15zdnd11an1n64x5 FILLER_143_1738 ();
 b15zdnd11an1n64x5 FILLER_143_1802 ();
 b15zdnd11an1n64x5 FILLER_143_1866 ();
 b15zdnd11an1n64x5 FILLER_143_1930 ();
 b15zdnd11an1n64x5 FILLER_143_1994 ();
 b15zdnd11an1n64x5 FILLER_143_2058 ();
 b15zdnd11an1n64x5 FILLER_143_2122 ();
 b15zdnd11an1n64x5 FILLER_143_2186 ();
 b15zdnd11an1n32x5 FILLER_143_2250 ();
 b15zdnd00an1n02x5 FILLER_143_2282 ();
 b15zdnd11an1n64x5 FILLER_144_8 ();
 b15zdnd11an1n64x5 FILLER_144_72 ();
 b15zdnd11an1n32x5 FILLER_144_136 ();
 b15zdnd11an1n16x5 FILLER_144_168 ();
 b15zdnd11an1n08x5 FILLER_144_184 ();
 b15zdnd11an1n04x5 FILLER_144_192 ();
 b15zdnd00an1n02x5 FILLER_144_196 ();
 b15zdnd00an1n01x5 FILLER_144_198 ();
 b15zdnd11an1n64x5 FILLER_144_251 ();
 b15zdnd11an1n64x5 FILLER_144_315 ();
 b15zdnd11an1n08x5 FILLER_144_379 ();
 b15zdnd00an1n02x5 FILLER_144_387 ();
 b15zdnd00an1n01x5 FILLER_144_389 ();
 b15zdnd11an1n64x5 FILLER_144_442 ();
 b15zdnd11an1n04x5 FILLER_144_506 ();
 b15zdnd00an1n02x5 FILLER_144_510 ();
 b15zdnd11an1n04x5 FILLER_144_517 ();
 b15zdnd00an1n02x5 FILLER_144_521 ();
 b15zdnd11an1n32x5 FILLER_144_555 ();
 b15zdnd11an1n16x5 FILLER_144_587 ();
 b15zdnd11an1n08x5 FILLER_144_603 ();
 b15zdnd11an1n04x5 FILLER_144_611 ();
 b15zdnd00an1n02x5 FILLER_144_615 ();
 b15zdnd00an1n01x5 FILLER_144_617 ();
 b15zdnd11an1n16x5 FILLER_144_627 ();
 b15zdnd11an1n16x5 FILLER_144_687 ();
 b15zdnd00an1n02x5 FILLER_144_703 ();
 b15zdnd00an1n01x5 FILLER_144_705 ();
 b15zdnd11an1n04x5 FILLER_144_713 ();
 b15zdnd00an1n01x5 FILLER_144_717 ();
 b15zdnd11an1n32x5 FILLER_144_726 ();
 b15zdnd11an1n16x5 FILLER_144_758 ();
 b15zdnd00an1n02x5 FILLER_144_774 ();
 b15zdnd00an1n01x5 FILLER_144_776 ();
 b15zdnd11an1n04x5 FILLER_144_790 ();
 b15zdnd11an1n08x5 FILLER_144_810 ();
 b15zdnd00an1n02x5 FILLER_144_818 ();
 b15zdnd11an1n16x5 FILLER_144_840 ();
 b15zdnd11an1n08x5 FILLER_144_856 ();
 b15zdnd00an1n02x5 FILLER_144_864 ();
 b15zdnd11an1n64x5 FILLER_144_880 ();
 b15zdnd11an1n64x5 FILLER_144_944 ();
 b15zdnd11an1n64x5 FILLER_144_1008 ();
 b15zdnd11an1n32x5 FILLER_144_1072 ();
 b15zdnd11an1n04x5 FILLER_144_1104 ();
 b15zdnd00an1n01x5 FILLER_144_1108 ();
 b15zdnd11an1n64x5 FILLER_144_1123 ();
 b15zdnd11an1n64x5 FILLER_144_1187 ();
 b15zdnd11an1n16x5 FILLER_144_1251 ();
 b15zdnd11an1n08x5 FILLER_144_1267 ();
 b15zdnd11an1n08x5 FILLER_144_1299 ();
 b15zdnd11an1n64x5 FILLER_144_1321 ();
 b15zdnd11an1n32x5 FILLER_144_1385 ();
 b15zdnd11an1n08x5 FILLER_144_1417 ();
 b15zdnd00an1n01x5 FILLER_144_1425 ();
 b15zdnd11an1n04x5 FILLER_144_1431 ();
 b15zdnd11an1n32x5 FILLER_144_1455 ();
 b15zdnd11an1n04x5 FILLER_144_1487 ();
 b15zdnd00an1n01x5 FILLER_144_1491 ();
 b15zdnd11an1n64x5 FILLER_144_1512 ();
 b15zdnd11an1n64x5 FILLER_144_1576 ();
 b15zdnd11an1n64x5 FILLER_144_1640 ();
 b15zdnd11an1n08x5 FILLER_144_1704 ();
 b15zdnd11an1n04x5 FILLER_144_1712 ();
 b15zdnd00an1n01x5 FILLER_144_1716 ();
 b15zdnd11an1n64x5 FILLER_144_1733 ();
 b15zdnd11an1n32x5 FILLER_144_1797 ();
 b15zdnd11an1n04x5 FILLER_144_1829 ();
 b15zdnd11an1n64x5 FILLER_144_1841 ();
 b15zdnd11an1n64x5 FILLER_144_1905 ();
 b15zdnd11an1n64x5 FILLER_144_1969 ();
 b15zdnd11an1n64x5 FILLER_144_2033 ();
 b15zdnd11an1n32x5 FILLER_144_2097 ();
 b15zdnd11an1n16x5 FILLER_144_2138 ();
 b15zdnd11an1n32x5 FILLER_144_2162 ();
 b15zdnd11an1n04x5 FILLER_144_2194 ();
 b15zdnd11an1n04x5 FILLER_144_2203 ();
 b15zdnd11an1n32x5 FILLER_144_2210 ();
 b15zdnd11an1n16x5 FILLER_144_2242 ();
 b15zdnd11an1n04x5 FILLER_144_2258 ();
 b15zdnd00an1n01x5 FILLER_144_2262 ();
 b15zdnd11an1n08x5 FILLER_144_2267 ();
 b15zdnd00an1n01x5 FILLER_144_2275 ();
 b15zdnd11an1n64x5 FILLER_145_0 ();
 b15zdnd11an1n64x5 FILLER_145_64 ();
 b15zdnd11an1n64x5 FILLER_145_128 ();
 b15zdnd11an1n16x5 FILLER_145_192 ();
 b15zdnd11an1n08x5 FILLER_145_208 ();
 b15zdnd00an1n02x5 FILLER_145_216 ();
 b15zdnd00an1n01x5 FILLER_145_218 ();
 b15zdnd11an1n04x5 FILLER_145_222 ();
 b15zdnd11an1n04x5 FILLER_145_229 ();
 b15zdnd11an1n64x5 FILLER_145_236 ();
 b15zdnd11an1n64x5 FILLER_145_300 ();
 b15zdnd11an1n32x5 FILLER_145_364 ();
 b15zdnd11an1n08x5 FILLER_145_396 ();
 b15zdnd11an1n04x5 FILLER_145_404 ();
 b15zdnd00an1n02x5 FILLER_145_408 ();
 b15zdnd11an1n04x5 FILLER_145_413 ();
 b15zdnd11an1n64x5 FILLER_145_420 ();
 b15zdnd11an1n08x5 FILLER_145_484 ();
 b15zdnd11an1n04x5 FILLER_145_492 ();
 b15zdnd00an1n02x5 FILLER_145_496 ();
 b15zdnd11an1n16x5 FILLER_145_510 ();
 b15zdnd11an1n08x5 FILLER_145_526 ();
 b15zdnd11an1n04x5 FILLER_145_534 ();
 b15zdnd11an1n32x5 FILLER_145_570 ();
 b15zdnd11an1n16x5 FILLER_145_602 ();
 b15zdnd11an1n08x5 FILLER_145_618 ();
 b15zdnd11an1n16x5 FILLER_145_640 ();
 b15zdnd00an1n01x5 FILLER_145_656 ();
 b15zdnd11an1n04x5 FILLER_145_660 ();
 b15zdnd11an1n32x5 FILLER_145_667 ();
 b15zdnd11an1n32x5 FILLER_145_710 ();
 b15zdnd11an1n04x5 FILLER_145_742 ();
 b15zdnd11an1n04x5 FILLER_145_754 ();
 b15zdnd11an1n04x5 FILLER_145_789 ();
 b15zdnd00an1n02x5 FILLER_145_793 ();
 b15zdnd11an1n16x5 FILLER_145_837 ();
 b15zdnd00an1n02x5 FILLER_145_853 ();
 b15zdnd11an1n16x5 FILLER_145_858 ();
 b15zdnd11an1n64x5 FILLER_145_894 ();
 b15zdnd11an1n64x5 FILLER_145_958 ();
 b15zdnd11an1n64x5 FILLER_145_1022 ();
 b15zdnd11an1n64x5 FILLER_145_1086 ();
 b15zdnd11an1n04x5 FILLER_145_1150 ();
 b15zdnd00an1n02x5 FILLER_145_1154 ();
 b15zdnd11an1n64x5 FILLER_145_1164 ();
 b15zdnd11an1n32x5 FILLER_145_1228 ();
 b15zdnd11an1n16x5 FILLER_145_1260 ();
 b15zdnd11an1n08x5 FILLER_145_1276 ();
 b15zdnd11an1n64x5 FILLER_145_1304 ();
 b15zdnd11an1n64x5 FILLER_145_1368 ();
 b15zdnd11an1n08x5 FILLER_145_1432 ();
 b15zdnd00an1n01x5 FILLER_145_1440 ();
 b15zdnd11an1n64x5 FILLER_145_1448 ();
 b15zdnd11an1n64x5 FILLER_145_1512 ();
 b15zdnd11an1n64x5 FILLER_145_1576 ();
 b15zdnd11an1n64x5 FILLER_145_1640 ();
 b15zdnd11an1n64x5 FILLER_145_1704 ();
 b15zdnd11an1n32x5 FILLER_145_1768 ();
 b15zdnd11an1n16x5 FILLER_145_1800 ();
 b15zdnd11an1n04x5 FILLER_145_1816 ();
 b15zdnd00an1n01x5 FILLER_145_1820 ();
 b15zdnd11an1n64x5 FILLER_145_1836 ();
 b15zdnd11an1n08x5 FILLER_145_1900 ();
 b15zdnd00an1n01x5 FILLER_145_1908 ();
 b15zdnd11an1n64x5 FILLER_145_1921 ();
 b15zdnd11an1n64x5 FILLER_145_1985 ();
 b15zdnd11an1n64x5 FILLER_145_2049 ();
 b15zdnd11an1n64x5 FILLER_145_2113 ();
 b15zdnd11an1n16x5 FILLER_145_2177 ();
 b15zdnd11an1n08x5 FILLER_145_2193 ();
 b15zdnd11an1n04x5 FILLER_145_2201 ();
 b15zdnd11an1n64x5 FILLER_145_2212 ();
 b15zdnd11an1n08x5 FILLER_145_2276 ();
 b15zdnd11an1n64x5 FILLER_146_8 ();
 b15zdnd11an1n64x5 FILLER_146_72 ();
 b15zdnd11an1n64x5 FILLER_146_136 ();
 b15zdnd11an1n64x5 FILLER_146_200 ();
 b15zdnd11an1n64x5 FILLER_146_264 ();
 b15zdnd11an1n04x5 FILLER_146_328 ();
 b15zdnd00an1n01x5 FILLER_146_332 ();
 b15zdnd11an1n32x5 FILLER_146_358 ();
 b15zdnd11an1n16x5 FILLER_146_390 ();
 b15zdnd11an1n08x5 FILLER_146_406 ();
 b15zdnd11an1n04x5 FILLER_146_414 ();
 b15zdnd11an1n64x5 FILLER_146_421 ();
 b15zdnd11an1n64x5 FILLER_146_485 ();
 b15zdnd11an1n64x5 FILLER_146_549 ();
 b15zdnd11an1n32x5 FILLER_146_613 ();
 b15zdnd11an1n16x5 FILLER_146_645 ();
 b15zdnd11an1n04x5 FILLER_146_661 ();
 b15zdnd00an1n02x5 FILLER_146_665 ();
 b15zdnd00an1n01x5 FILLER_146_667 ();
 b15zdnd11an1n32x5 FILLER_146_676 ();
 b15zdnd11an1n08x5 FILLER_146_708 ();
 b15zdnd00an1n02x5 FILLER_146_716 ();
 b15zdnd11an1n64x5 FILLER_146_726 ();
 b15zdnd00an1n02x5 FILLER_146_790 ();
 b15zdnd00an1n01x5 FILLER_146_792 ();
 b15zdnd11an1n08x5 FILLER_146_837 ();
 b15zdnd11an1n04x5 FILLER_146_845 ();
 b15zdnd11an1n08x5 FILLER_146_862 ();
 b15zdnd11an1n64x5 FILLER_146_886 ();
 b15zdnd11an1n64x5 FILLER_146_950 ();
 b15zdnd11an1n64x5 FILLER_146_1014 ();
 b15zdnd11an1n64x5 FILLER_146_1078 ();
 b15zdnd11an1n64x5 FILLER_146_1142 ();
 b15zdnd11an1n64x5 FILLER_146_1206 ();
 b15zdnd11an1n04x5 FILLER_146_1270 ();
 b15zdnd00an1n02x5 FILLER_146_1274 ();
 b15zdnd11an1n64x5 FILLER_146_1290 ();
 b15zdnd11an1n64x5 FILLER_146_1354 ();
 b15zdnd11an1n64x5 FILLER_146_1418 ();
 b15zdnd11an1n32x5 FILLER_146_1482 ();
 b15zdnd11an1n08x5 FILLER_146_1514 ();
 b15zdnd00an1n02x5 FILLER_146_1522 ();
 b15zdnd00an1n01x5 FILLER_146_1524 ();
 b15zdnd11an1n08x5 FILLER_146_1530 ();
 b15zdnd00an1n01x5 FILLER_146_1538 ();
 b15zdnd11an1n04x5 FILLER_146_1553 ();
 b15zdnd00an1n02x5 FILLER_146_1557 ();
 b15zdnd11an1n64x5 FILLER_146_1573 ();
 b15zdnd11an1n64x5 FILLER_146_1637 ();
 b15zdnd11an1n64x5 FILLER_146_1701 ();
 b15zdnd11an1n64x5 FILLER_146_1765 ();
 b15zdnd11an1n64x5 FILLER_146_1829 ();
 b15zdnd11an1n64x5 FILLER_146_1893 ();
 b15zdnd11an1n64x5 FILLER_146_1957 ();
 b15zdnd11an1n64x5 FILLER_146_2021 ();
 b15zdnd11an1n64x5 FILLER_146_2085 ();
 b15zdnd11an1n04x5 FILLER_146_2149 ();
 b15zdnd00an1n01x5 FILLER_146_2153 ();
 b15zdnd11an1n64x5 FILLER_146_2162 ();
 b15zdnd11an1n32x5 FILLER_146_2226 ();
 b15zdnd11an1n16x5 FILLER_146_2258 ();
 b15zdnd00an1n02x5 FILLER_146_2274 ();
 b15zdnd11an1n32x5 FILLER_147_0 ();
 b15zdnd11an1n04x5 FILLER_147_32 ();
 b15zdnd00an1n01x5 FILLER_147_36 ();
 b15zdnd11an1n64x5 FILLER_147_41 ();
 b15zdnd11an1n64x5 FILLER_147_105 ();
 b15zdnd11an1n64x5 FILLER_147_169 ();
 b15zdnd11an1n64x5 FILLER_147_233 ();
 b15zdnd11an1n32x5 FILLER_147_297 ();
 b15zdnd11an1n08x5 FILLER_147_329 ();
 b15zdnd11an1n04x5 FILLER_147_337 ();
 b15zdnd11an1n16x5 FILLER_147_383 ();
 b15zdnd11an1n04x5 FILLER_147_399 ();
 b15zdnd00an1n02x5 FILLER_147_403 ();
 b15zdnd00an1n01x5 FILLER_147_405 ();
 b15zdnd11an1n32x5 FILLER_147_412 ();
 b15zdnd11an1n16x5 FILLER_147_444 ();
 b15zdnd11an1n04x5 FILLER_147_460 ();
 b15zdnd00an1n02x5 FILLER_147_464 ();
 b15zdnd11an1n64x5 FILLER_147_477 ();
 b15zdnd11an1n64x5 FILLER_147_541 ();
 b15zdnd11an1n08x5 FILLER_147_605 ();
 b15zdnd11an1n04x5 FILLER_147_613 ();
 b15zdnd00an1n02x5 FILLER_147_617 ();
 b15zdnd00an1n01x5 FILLER_147_619 ();
 b15zdnd11an1n32x5 FILLER_147_626 ();
 b15zdnd11an1n16x5 FILLER_147_658 ();
 b15zdnd00an1n02x5 FILLER_147_674 ();
 b15zdnd00an1n01x5 FILLER_147_676 ();
 b15zdnd11an1n64x5 FILLER_147_683 ();
 b15zdnd11an1n32x5 FILLER_147_747 ();
 b15zdnd11an1n16x5 FILLER_147_779 ();
 b15zdnd11an1n08x5 FILLER_147_795 ();
 b15zdnd00an1n01x5 FILLER_147_803 ();
 b15zdnd11an1n08x5 FILLER_147_807 ();
 b15zdnd00an1n01x5 FILLER_147_815 ();
 b15zdnd11an1n16x5 FILLER_147_819 ();
 b15zdnd11an1n04x5 FILLER_147_835 ();
 b15zdnd00an1n02x5 FILLER_147_839 ();
 b15zdnd00an1n01x5 FILLER_147_841 ();
 b15zdnd11an1n64x5 FILLER_147_884 ();
 b15zdnd11an1n04x5 FILLER_147_948 ();
 b15zdnd11an1n64x5 FILLER_147_966 ();
 b15zdnd11an1n64x5 FILLER_147_1030 ();
 b15zdnd11an1n64x5 FILLER_147_1094 ();
 b15zdnd11an1n64x5 FILLER_147_1158 ();
 b15zdnd11an1n64x5 FILLER_147_1222 ();
 b15zdnd11an1n08x5 FILLER_147_1286 ();
 b15zdnd11an1n04x5 FILLER_147_1294 ();
 b15zdnd00an1n02x5 FILLER_147_1298 ();
 b15zdnd11an1n64x5 FILLER_147_1320 ();
 b15zdnd11an1n16x5 FILLER_147_1384 ();
 b15zdnd11an1n08x5 FILLER_147_1400 ();
 b15zdnd11an1n04x5 FILLER_147_1408 ();
 b15zdnd00an1n02x5 FILLER_147_1412 ();
 b15zdnd11an1n32x5 FILLER_147_1431 ();
 b15zdnd11an1n08x5 FILLER_147_1463 ();
 b15zdnd00an1n02x5 FILLER_147_1471 ();
 b15zdnd11an1n64x5 FILLER_147_1481 ();
 b15zdnd11an1n64x5 FILLER_147_1545 ();
 b15zdnd11an1n64x5 FILLER_147_1609 ();
 b15zdnd11an1n64x5 FILLER_147_1673 ();
 b15zdnd11an1n64x5 FILLER_147_1737 ();
 b15zdnd11an1n32x5 FILLER_147_1801 ();
 b15zdnd11an1n08x5 FILLER_147_1833 ();
 b15zdnd11an1n04x5 FILLER_147_1841 ();
 b15zdnd00an1n02x5 FILLER_147_1845 ();
 b15zdnd11an1n08x5 FILLER_147_1865 ();
 b15zdnd00an1n02x5 FILLER_147_1873 ();
 b15zdnd11an1n64x5 FILLER_147_1917 ();
 b15zdnd11an1n64x5 FILLER_147_1981 ();
 b15zdnd11an1n64x5 FILLER_147_2045 ();
 b15zdnd11an1n64x5 FILLER_147_2109 ();
 b15zdnd11an1n64x5 FILLER_147_2173 ();
 b15zdnd11an1n32x5 FILLER_147_2237 ();
 b15zdnd11an1n08x5 FILLER_147_2269 ();
 b15zdnd11an1n04x5 FILLER_147_2277 ();
 b15zdnd00an1n02x5 FILLER_147_2281 ();
 b15zdnd00an1n01x5 FILLER_147_2283 ();
 b15zdnd11an1n64x5 FILLER_148_8 ();
 b15zdnd11an1n64x5 FILLER_148_72 ();
 b15zdnd11an1n64x5 FILLER_148_136 ();
 b15zdnd11an1n64x5 FILLER_148_200 ();
 b15zdnd11an1n64x5 FILLER_148_264 ();
 b15zdnd11an1n08x5 FILLER_148_328 ();
 b15zdnd00an1n01x5 FILLER_148_336 ();
 b15zdnd11an1n04x5 FILLER_148_342 ();
 b15zdnd11an1n16x5 FILLER_148_398 ();
 b15zdnd11an1n04x5 FILLER_148_414 ();
 b15zdnd00an1n01x5 FILLER_148_418 ();
 b15zdnd11an1n64x5 FILLER_148_426 ();
 b15zdnd11an1n64x5 FILLER_148_490 ();
 b15zdnd11an1n16x5 FILLER_148_554 ();
 b15zdnd11an1n04x5 FILLER_148_570 ();
 b15zdnd00an1n01x5 FILLER_148_574 ();
 b15zdnd11an1n16x5 FILLER_148_579 ();
 b15zdnd11an1n08x5 FILLER_148_595 ();
 b15zdnd11an1n04x5 FILLER_148_603 ();
 b15zdnd11an1n64x5 FILLER_148_611 ();
 b15zdnd11an1n32x5 FILLER_148_675 ();
 b15zdnd11an1n08x5 FILLER_148_707 ();
 b15zdnd00an1n02x5 FILLER_148_715 ();
 b15zdnd00an1n01x5 FILLER_148_717 ();
 b15zdnd11an1n64x5 FILLER_148_726 ();
 b15zdnd11an1n16x5 FILLER_148_790 ();
 b15zdnd11an1n08x5 FILLER_148_806 ();
 b15zdnd00an1n02x5 FILLER_148_814 ();
 b15zdnd00an1n01x5 FILLER_148_816 ();
 b15zdnd11an1n16x5 FILLER_148_820 ();
 b15zdnd11an1n08x5 FILLER_148_836 ();
 b15zdnd00an1n02x5 FILLER_148_844 ();
 b15zdnd00an1n01x5 FILLER_148_846 ();
 b15zdnd11an1n04x5 FILLER_148_857 ();
 b15zdnd11an1n64x5 FILLER_148_864 ();
 b15zdnd11an1n64x5 FILLER_148_928 ();
 b15zdnd11an1n64x5 FILLER_148_992 ();
 b15zdnd11an1n64x5 FILLER_148_1056 ();
 b15zdnd11an1n64x5 FILLER_148_1120 ();
 b15zdnd11an1n64x5 FILLER_148_1184 ();
 b15zdnd11an1n32x5 FILLER_148_1248 ();
 b15zdnd11an1n08x5 FILLER_148_1280 ();
 b15zdnd11an1n04x5 FILLER_148_1288 ();
 b15zdnd11an1n64x5 FILLER_148_1304 ();
 b15zdnd11an1n64x5 FILLER_148_1368 ();
 b15zdnd11an1n64x5 FILLER_148_1432 ();
 b15zdnd11an1n64x5 FILLER_148_1496 ();
 b15zdnd11an1n64x5 FILLER_148_1560 ();
 b15zdnd11an1n64x5 FILLER_148_1624 ();
 b15zdnd11an1n64x5 FILLER_148_1688 ();
 b15zdnd11an1n64x5 FILLER_148_1752 ();
 b15zdnd11an1n64x5 FILLER_148_1816 ();
 b15zdnd11an1n64x5 FILLER_148_1880 ();
 b15zdnd11an1n64x5 FILLER_148_1944 ();
 b15zdnd11an1n64x5 FILLER_148_2008 ();
 b15zdnd11an1n64x5 FILLER_148_2072 ();
 b15zdnd11an1n16x5 FILLER_148_2136 ();
 b15zdnd00an1n02x5 FILLER_148_2152 ();
 b15zdnd11an1n32x5 FILLER_148_2162 ();
 b15zdnd11an1n16x5 FILLER_148_2194 ();
 b15zdnd11an1n04x5 FILLER_148_2210 ();
 b15zdnd00an1n02x5 FILLER_148_2214 ();
 b15zdnd11an1n32x5 FILLER_148_2238 ();
 b15zdnd11an1n04x5 FILLER_148_2270 ();
 b15zdnd00an1n02x5 FILLER_148_2274 ();
 b15zdnd11an1n64x5 FILLER_149_0 ();
 b15zdnd11an1n64x5 FILLER_149_64 ();
 b15zdnd11an1n64x5 FILLER_149_128 ();
 b15zdnd11an1n64x5 FILLER_149_192 ();
 b15zdnd11an1n64x5 FILLER_149_256 ();
 b15zdnd11an1n32x5 FILLER_149_320 ();
 b15zdnd11an1n08x5 FILLER_149_352 ();
 b15zdnd11an1n04x5 FILLER_149_360 ();
 b15zdnd00an1n02x5 FILLER_149_364 ();
 b15zdnd11an1n04x5 FILLER_149_369 ();
 b15zdnd11an1n16x5 FILLER_149_376 ();
 b15zdnd11an1n08x5 FILLER_149_392 ();
 b15zdnd11an1n04x5 FILLER_149_400 ();
 b15zdnd11an1n64x5 FILLER_149_413 ();
 b15zdnd11an1n64x5 FILLER_149_477 ();
 b15zdnd11an1n16x5 FILLER_149_541 ();
 b15zdnd11an1n08x5 FILLER_149_557 ();
 b15zdnd11an1n04x5 FILLER_149_565 ();
 b15zdnd00an1n02x5 FILLER_149_569 ();
 b15zdnd11an1n04x5 FILLER_149_580 ();
 b15zdnd00an1n02x5 FILLER_149_584 ();
 b15zdnd00an1n01x5 FILLER_149_586 ();
 b15zdnd11an1n16x5 FILLER_149_593 ();
 b15zdnd11an1n04x5 FILLER_149_609 ();
 b15zdnd00an1n02x5 FILLER_149_613 ();
 b15zdnd00an1n01x5 FILLER_149_615 ();
 b15zdnd11an1n64x5 FILLER_149_648 ();
 b15zdnd11an1n64x5 FILLER_149_712 ();
 b15zdnd11an1n64x5 FILLER_149_776 ();
 b15zdnd11an1n64x5 FILLER_149_840 ();
 b15zdnd11an1n64x5 FILLER_149_904 ();
 b15zdnd11an1n64x5 FILLER_149_968 ();
 b15zdnd11an1n64x5 FILLER_149_1032 ();
 b15zdnd11an1n64x5 FILLER_149_1096 ();
 b15zdnd11an1n64x5 FILLER_149_1160 ();
 b15zdnd11an1n64x5 FILLER_149_1224 ();
 b15zdnd11an1n64x5 FILLER_149_1288 ();
 b15zdnd11an1n64x5 FILLER_149_1352 ();
 b15zdnd11an1n64x5 FILLER_149_1416 ();
 b15zdnd11an1n64x5 FILLER_149_1480 ();
 b15zdnd11an1n64x5 FILLER_149_1544 ();
 b15zdnd11an1n64x5 FILLER_149_1608 ();
 b15zdnd11an1n64x5 FILLER_149_1672 ();
 b15zdnd11an1n32x5 FILLER_149_1736 ();
 b15zdnd00an1n01x5 FILLER_149_1768 ();
 b15zdnd11an1n64x5 FILLER_149_1775 ();
 b15zdnd11an1n64x5 FILLER_149_1839 ();
 b15zdnd11an1n64x5 FILLER_149_1903 ();
 b15zdnd11an1n64x5 FILLER_149_1967 ();
 b15zdnd11an1n64x5 FILLER_149_2031 ();
 b15zdnd11an1n32x5 FILLER_149_2095 ();
 b15zdnd00an1n02x5 FILLER_149_2127 ();
 b15zdnd00an1n01x5 FILLER_149_2129 ();
 b15zdnd11an1n04x5 FILLER_149_2133 ();
 b15zdnd11an1n32x5 FILLER_149_2140 ();
 b15zdnd11an1n16x5 FILLER_149_2172 ();
 b15zdnd00an1n02x5 FILLER_149_2188 ();
 b15zdnd00an1n01x5 FILLER_149_2190 ();
 b15zdnd11an1n64x5 FILLER_149_2200 ();
 b15zdnd11an1n16x5 FILLER_149_2264 ();
 b15zdnd11an1n04x5 FILLER_149_2280 ();
 b15zdnd11an1n64x5 FILLER_150_8 ();
 b15zdnd11an1n64x5 FILLER_150_72 ();
 b15zdnd11an1n64x5 FILLER_150_136 ();
 b15zdnd11an1n32x5 FILLER_150_200 ();
 b15zdnd11an1n16x5 FILLER_150_232 ();
 b15zdnd11an1n04x5 FILLER_150_248 ();
 b15zdnd00an1n01x5 FILLER_150_252 ();
 b15zdnd11an1n64x5 FILLER_150_295 ();
 b15zdnd11an1n08x5 FILLER_150_359 ();
 b15zdnd11an1n04x5 FILLER_150_367 ();
 b15zdnd11an1n64x5 FILLER_150_374 ();
 b15zdnd11an1n64x5 FILLER_150_438 ();
 b15zdnd11an1n16x5 FILLER_150_502 ();
 b15zdnd00an1n01x5 FILLER_150_518 ();
 b15zdnd11an1n32x5 FILLER_150_529 ();
 b15zdnd11an1n08x5 FILLER_150_561 ();
 b15zdnd11an1n64x5 FILLER_150_593 ();
 b15zdnd11an1n32x5 FILLER_150_657 ();
 b15zdnd11an1n16x5 FILLER_150_689 ();
 b15zdnd11an1n08x5 FILLER_150_705 ();
 b15zdnd11an1n04x5 FILLER_150_713 ();
 b15zdnd00an1n01x5 FILLER_150_717 ();
 b15zdnd11an1n64x5 FILLER_150_726 ();
 b15zdnd11an1n16x5 FILLER_150_790 ();
 b15zdnd11an1n04x5 FILLER_150_806 ();
 b15zdnd00an1n02x5 FILLER_150_810 ();
 b15zdnd11an1n64x5 FILLER_150_824 ();
 b15zdnd11an1n32x5 FILLER_150_888 ();
 b15zdnd11an1n08x5 FILLER_150_920 ();
 b15zdnd00an1n02x5 FILLER_150_928 ();
 b15zdnd00an1n01x5 FILLER_150_930 ();
 b15zdnd11an1n64x5 FILLER_150_973 ();
 b15zdnd11an1n64x5 FILLER_150_1037 ();
 b15zdnd11an1n64x5 FILLER_150_1101 ();
 b15zdnd11an1n64x5 FILLER_150_1165 ();
 b15zdnd11an1n32x5 FILLER_150_1229 ();
 b15zdnd11an1n08x5 FILLER_150_1261 ();
 b15zdnd11an1n04x5 FILLER_150_1269 ();
 b15zdnd00an1n02x5 FILLER_150_1273 ();
 b15zdnd00an1n01x5 FILLER_150_1275 ();
 b15zdnd11an1n32x5 FILLER_150_1288 ();
 b15zdnd11an1n04x5 FILLER_150_1323 ();
 b15zdnd11an1n64x5 FILLER_150_1330 ();
 b15zdnd11an1n64x5 FILLER_150_1394 ();
 b15zdnd11an1n64x5 FILLER_150_1458 ();
 b15zdnd11an1n32x5 FILLER_150_1522 ();
 b15zdnd11an1n08x5 FILLER_150_1554 ();
 b15zdnd11an1n04x5 FILLER_150_1562 ();
 b15zdnd11an1n64x5 FILLER_150_1574 ();
 b15zdnd11an1n64x5 FILLER_150_1638 ();
 b15zdnd11an1n64x5 FILLER_150_1702 ();
 b15zdnd11an1n64x5 FILLER_150_1766 ();
 b15zdnd11an1n32x5 FILLER_150_1830 ();
 b15zdnd11an1n08x5 FILLER_150_1862 ();
 b15zdnd11an1n64x5 FILLER_150_1915 ();
 b15zdnd11an1n64x5 FILLER_150_1979 ();
 b15zdnd11an1n64x5 FILLER_150_2043 ();
 b15zdnd11an1n04x5 FILLER_150_2107 ();
 b15zdnd11an1n08x5 FILLER_150_2143 ();
 b15zdnd00an1n02x5 FILLER_150_2151 ();
 b15zdnd00an1n01x5 FILLER_150_2153 ();
 b15zdnd11an1n64x5 FILLER_150_2162 ();
 b15zdnd11an1n32x5 FILLER_150_2226 ();
 b15zdnd11an1n16x5 FILLER_150_2258 ();
 b15zdnd00an1n02x5 FILLER_150_2274 ();
 b15zdnd11an1n64x5 FILLER_151_0 ();
 b15zdnd11an1n64x5 FILLER_151_64 ();
 b15zdnd11an1n64x5 FILLER_151_128 ();
 b15zdnd11an1n64x5 FILLER_151_192 ();
 b15zdnd11an1n64x5 FILLER_151_256 ();
 b15zdnd11an1n64x5 FILLER_151_320 ();
 b15zdnd11an1n64x5 FILLER_151_384 ();
 b15zdnd11an1n64x5 FILLER_151_448 ();
 b15zdnd11an1n08x5 FILLER_151_512 ();
 b15zdnd11an1n04x5 FILLER_151_520 ();
 b15zdnd00an1n02x5 FILLER_151_524 ();
 b15zdnd00an1n01x5 FILLER_151_526 ();
 b15zdnd11an1n04x5 FILLER_151_542 ();
 b15zdnd11an1n64x5 FILLER_151_557 ();
 b15zdnd11an1n64x5 FILLER_151_621 ();
 b15zdnd11an1n64x5 FILLER_151_685 ();
 b15zdnd11an1n64x5 FILLER_151_749 ();
 b15zdnd11an1n64x5 FILLER_151_813 ();
 b15zdnd11an1n64x5 FILLER_151_877 ();
 b15zdnd11an1n64x5 FILLER_151_983 ();
 b15zdnd11an1n64x5 FILLER_151_1047 ();
 b15zdnd11an1n64x5 FILLER_151_1111 ();
 b15zdnd11an1n64x5 FILLER_151_1175 ();
 b15zdnd11an1n32x5 FILLER_151_1239 ();
 b15zdnd11an1n08x5 FILLER_151_1271 ();
 b15zdnd11an1n04x5 FILLER_151_1279 ();
 b15zdnd00an1n02x5 FILLER_151_1283 ();
 b15zdnd00an1n01x5 FILLER_151_1285 ();
 b15zdnd11an1n04x5 FILLER_151_1298 ();
 b15zdnd11an1n64x5 FILLER_151_1354 ();
 b15zdnd11an1n64x5 FILLER_151_1418 ();
 b15zdnd11an1n64x5 FILLER_151_1482 ();
 b15zdnd11an1n64x5 FILLER_151_1546 ();
 b15zdnd11an1n64x5 FILLER_151_1610 ();
 b15zdnd11an1n64x5 FILLER_151_1674 ();
 b15zdnd11an1n64x5 FILLER_151_1738 ();
 b15zdnd11an1n64x5 FILLER_151_1802 ();
 b15zdnd11an1n64x5 FILLER_151_1866 ();
 b15zdnd11an1n64x5 FILLER_151_1930 ();
 b15zdnd11an1n64x5 FILLER_151_1994 ();
 b15zdnd11an1n64x5 FILLER_151_2058 ();
 b15zdnd11an1n16x5 FILLER_151_2122 ();
 b15zdnd00an1n02x5 FILLER_151_2138 ();
 b15zdnd00an1n01x5 FILLER_151_2140 ();
 b15zdnd11an1n64x5 FILLER_151_2144 ();
 b15zdnd11an1n64x5 FILLER_151_2208 ();
 b15zdnd11an1n08x5 FILLER_151_2272 ();
 b15zdnd11an1n04x5 FILLER_151_2280 ();
 b15zdnd11an1n64x5 FILLER_152_8 ();
 b15zdnd11an1n64x5 FILLER_152_72 ();
 b15zdnd11an1n64x5 FILLER_152_136 ();
 b15zdnd11an1n64x5 FILLER_152_200 ();
 b15zdnd11an1n64x5 FILLER_152_264 ();
 b15zdnd11an1n64x5 FILLER_152_328 ();
 b15zdnd11an1n64x5 FILLER_152_392 ();
 b15zdnd11an1n64x5 FILLER_152_456 ();
 b15zdnd11an1n32x5 FILLER_152_520 ();
 b15zdnd00an1n01x5 FILLER_152_552 ();
 b15zdnd11an1n64x5 FILLER_152_564 ();
 b15zdnd11an1n64x5 FILLER_152_628 ();
 b15zdnd11an1n16x5 FILLER_152_692 ();
 b15zdnd11an1n08x5 FILLER_152_708 ();
 b15zdnd00an1n02x5 FILLER_152_716 ();
 b15zdnd11an1n64x5 FILLER_152_726 ();
 b15zdnd11an1n64x5 FILLER_152_790 ();
 b15zdnd11an1n64x5 FILLER_152_854 ();
 b15zdnd11an1n64x5 FILLER_152_918 ();
 b15zdnd11an1n64x5 FILLER_152_982 ();
 b15zdnd11an1n64x5 FILLER_152_1046 ();
 b15zdnd11an1n64x5 FILLER_152_1110 ();
 b15zdnd11an1n64x5 FILLER_152_1174 ();
 b15zdnd11an1n64x5 FILLER_152_1238 ();
 b15zdnd11an1n08x5 FILLER_152_1302 ();
 b15zdnd00an1n01x5 FILLER_152_1310 ();
 b15zdnd11an1n08x5 FILLER_152_1318 ();
 b15zdnd00an1n01x5 FILLER_152_1326 ();
 b15zdnd11an1n08x5 FILLER_152_1330 ();
 b15zdnd11an1n04x5 FILLER_152_1338 ();
 b15zdnd11an1n32x5 FILLER_152_1384 ();
 b15zdnd11an1n64x5 FILLER_152_1420 ();
 b15zdnd11an1n32x5 FILLER_152_1484 ();
 b15zdnd11an1n16x5 FILLER_152_1516 ();
 b15zdnd11an1n04x5 FILLER_152_1532 ();
 b15zdnd11an1n64x5 FILLER_152_1540 ();
 b15zdnd11an1n64x5 FILLER_152_1604 ();
 b15zdnd11an1n64x5 FILLER_152_1668 ();
 b15zdnd11an1n64x5 FILLER_152_1732 ();
 b15zdnd11an1n64x5 FILLER_152_1796 ();
 b15zdnd11an1n64x5 FILLER_152_1860 ();
 b15zdnd11an1n64x5 FILLER_152_1924 ();
 b15zdnd11an1n64x5 FILLER_152_1988 ();
 b15zdnd11an1n32x5 FILLER_152_2052 ();
 b15zdnd11an1n08x5 FILLER_152_2084 ();
 b15zdnd11an1n16x5 FILLER_152_2123 ();
 b15zdnd11an1n08x5 FILLER_152_2139 ();
 b15zdnd11an1n04x5 FILLER_152_2147 ();
 b15zdnd00an1n02x5 FILLER_152_2151 ();
 b15zdnd00an1n01x5 FILLER_152_2153 ();
 b15zdnd11an1n64x5 FILLER_152_2162 ();
 b15zdnd11an1n32x5 FILLER_152_2226 ();
 b15zdnd11an1n16x5 FILLER_152_2258 ();
 b15zdnd00an1n02x5 FILLER_152_2274 ();
 b15zdnd11an1n64x5 FILLER_153_0 ();
 b15zdnd11an1n64x5 FILLER_153_64 ();
 b15zdnd11an1n16x5 FILLER_153_128 ();
 b15zdnd11an1n08x5 FILLER_153_144 ();
 b15zdnd11an1n04x5 FILLER_153_152 ();
 b15zdnd00an1n02x5 FILLER_153_156 ();
 b15zdnd11an1n64x5 FILLER_153_164 ();
 b15zdnd11an1n04x5 FILLER_153_228 ();
 b15zdnd00an1n02x5 FILLER_153_232 ();
 b15zdnd11an1n64x5 FILLER_153_237 ();
 b15zdnd11an1n64x5 FILLER_153_301 ();
 b15zdnd11an1n64x5 FILLER_153_365 ();
 b15zdnd11an1n64x5 FILLER_153_429 ();
 b15zdnd11an1n16x5 FILLER_153_493 ();
 b15zdnd11an1n04x5 FILLER_153_509 ();
 b15zdnd00an1n02x5 FILLER_153_513 ();
 b15zdnd00an1n01x5 FILLER_153_515 ();
 b15zdnd11an1n16x5 FILLER_153_520 ();
 b15zdnd00an1n02x5 FILLER_153_536 ();
 b15zdnd11an1n64x5 FILLER_153_549 ();
 b15zdnd11an1n64x5 FILLER_153_613 ();
 b15zdnd11an1n64x5 FILLER_153_677 ();
 b15zdnd11an1n64x5 FILLER_153_741 ();
 b15zdnd11an1n64x5 FILLER_153_805 ();
 b15zdnd11an1n64x5 FILLER_153_869 ();
 b15zdnd11an1n64x5 FILLER_153_933 ();
 b15zdnd11an1n64x5 FILLER_153_997 ();
 b15zdnd11an1n64x5 FILLER_153_1061 ();
 b15zdnd11an1n64x5 FILLER_153_1125 ();
 b15zdnd11an1n64x5 FILLER_153_1189 ();
 b15zdnd11an1n64x5 FILLER_153_1253 ();
 b15zdnd11an1n64x5 FILLER_153_1317 ();
 b15zdnd11an1n64x5 FILLER_153_1381 ();
 b15zdnd11an1n64x5 FILLER_153_1445 ();
 b15zdnd11an1n32x5 FILLER_153_1509 ();
 b15zdnd11an1n16x5 FILLER_153_1541 ();
 b15zdnd11an1n08x5 FILLER_153_1557 ();
 b15zdnd11an1n08x5 FILLER_153_1582 ();
 b15zdnd11an1n04x5 FILLER_153_1590 ();
 b15zdnd00an1n01x5 FILLER_153_1594 ();
 b15zdnd11an1n64x5 FILLER_153_1600 ();
 b15zdnd11an1n32x5 FILLER_153_1664 ();
 b15zdnd11an1n16x5 FILLER_153_1696 ();
 b15zdnd11an1n08x5 FILLER_153_1712 ();
 b15zdnd11an1n04x5 FILLER_153_1720 ();
 b15zdnd11an1n04x5 FILLER_153_1730 ();
 b15zdnd11an1n32x5 FILLER_153_1741 ();
 b15zdnd11an1n04x5 FILLER_153_1773 ();
 b15zdnd11an1n64x5 FILLER_153_1783 ();
 b15zdnd11an1n64x5 FILLER_153_1847 ();
 b15zdnd11an1n16x5 FILLER_153_1911 ();
 b15zdnd00an1n02x5 FILLER_153_1927 ();
 b15zdnd11an1n64x5 FILLER_153_1973 ();
 b15zdnd11an1n64x5 FILLER_153_2037 ();
 b15zdnd00an1n02x5 FILLER_153_2101 ();
 b15zdnd11an1n64x5 FILLER_153_2145 ();
 b15zdnd11an1n64x5 FILLER_153_2209 ();
 b15zdnd11an1n08x5 FILLER_153_2273 ();
 b15zdnd00an1n02x5 FILLER_153_2281 ();
 b15zdnd00an1n01x5 FILLER_153_2283 ();
 b15zdnd11an1n08x5 FILLER_154_8 ();
 b15zdnd11an1n04x5 FILLER_154_16 ();
 b15zdnd00an1n01x5 FILLER_154_20 ();
 b15zdnd11an1n64x5 FILLER_154_25 ();
 b15zdnd11an1n64x5 FILLER_154_89 ();
 b15zdnd11an1n32x5 FILLER_154_153 ();
 b15zdnd11an1n08x5 FILLER_154_185 ();
 b15zdnd11an1n04x5 FILLER_154_193 ();
 b15zdnd00an1n01x5 FILLER_154_197 ();
 b15zdnd11an1n64x5 FILLER_154_238 ();
 b15zdnd11an1n64x5 FILLER_154_302 ();
 b15zdnd11an1n64x5 FILLER_154_366 ();
 b15zdnd11an1n64x5 FILLER_154_430 ();
 b15zdnd11an1n64x5 FILLER_154_494 ();
 b15zdnd11an1n64x5 FILLER_154_558 ();
 b15zdnd11an1n64x5 FILLER_154_622 ();
 b15zdnd11an1n32x5 FILLER_154_686 ();
 b15zdnd11an1n64x5 FILLER_154_726 ();
 b15zdnd11an1n64x5 FILLER_154_790 ();
 b15zdnd11an1n64x5 FILLER_154_854 ();
 b15zdnd11an1n64x5 FILLER_154_918 ();
 b15zdnd11an1n64x5 FILLER_154_982 ();
 b15zdnd11an1n64x5 FILLER_154_1046 ();
 b15zdnd11an1n64x5 FILLER_154_1110 ();
 b15zdnd11an1n64x5 FILLER_154_1174 ();
 b15zdnd11an1n64x5 FILLER_154_1238 ();
 b15zdnd11an1n64x5 FILLER_154_1302 ();
 b15zdnd11an1n64x5 FILLER_154_1366 ();
 b15zdnd11an1n64x5 FILLER_154_1430 ();
 b15zdnd11an1n64x5 FILLER_154_1494 ();
 b15zdnd11an1n08x5 FILLER_154_1558 ();
 b15zdnd11an1n04x5 FILLER_154_1566 ();
 b15zdnd00an1n02x5 FILLER_154_1570 ();
 b15zdnd11an1n64x5 FILLER_154_1593 ();
 b15zdnd11an1n64x5 FILLER_154_1657 ();
 b15zdnd11an1n32x5 FILLER_154_1721 ();
 b15zdnd11an1n16x5 FILLER_154_1753 ();
 b15zdnd11an1n08x5 FILLER_154_1769 ();
 b15zdnd00an1n02x5 FILLER_154_1777 ();
 b15zdnd11an1n08x5 FILLER_154_1786 ();
 b15zdnd11an1n04x5 FILLER_154_1794 ();
 b15zdnd00an1n02x5 FILLER_154_1798 ();
 b15zdnd11an1n64x5 FILLER_154_1806 ();
 b15zdnd11an1n64x5 FILLER_154_1870 ();
 b15zdnd11an1n08x5 FILLER_154_1934 ();
 b15zdnd00an1n02x5 FILLER_154_1942 ();
 b15zdnd11an1n04x5 FILLER_154_1947 ();
 b15zdnd11an1n04x5 FILLER_154_1954 ();
 b15zdnd11an1n64x5 FILLER_154_1961 ();
 b15zdnd11an1n32x5 FILLER_154_2025 ();
 b15zdnd11an1n16x5 FILLER_154_2057 ();
 b15zdnd00an1n02x5 FILLER_154_2073 ();
 b15zdnd00an1n01x5 FILLER_154_2075 ();
 b15zdnd11an1n32x5 FILLER_154_2121 ();
 b15zdnd00an1n01x5 FILLER_154_2153 ();
 b15zdnd11an1n64x5 FILLER_154_2162 ();
 b15zdnd11an1n32x5 FILLER_154_2226 ();
 b15zdnd11an1n16x5 FILLER_154_2258 ();
 b15zdnd00an1n02x5 FILLER_154_2274 ();
 b15zdnd11an1n64x5 FILLER_155_0 ();
 b15zdnd11an1n64x5 FILLER_155_64 ();
 b15zdnd11an1n16x5 FILLER_155_128 ();
 b15zdnd11an1n08x5 FILLER_155_144 ();
 b15zdnd00an1n02x5 FILLER_155_152 ();
 b15zdnd00an1n01x5 FILLER_155_154 ();
 b15zdnd11an1n64x5 FILLER_155_165 ();
 b15zdnd11an1n04x5 FILLER_155_229 ();
 b15zdnd00an1n01x5 FILLER_155_233 ();
 b15zdnd11an1n32x5 FILLER_155_237 ();
 b15zdnd11an1n08x5 FILLER_155_269 ();
 b15zdnd11an1n04x5 FILLER_155_277 ();
 b15zdnd00an1n02x5 FILLER_155_281 ();
 b15zdnd00an1n01x5 FILLER_155_283 ();
 b15zdnd11an1n64x5 FILLER_155_336 ();
 b15zdnd11an1n64x5 FILLER_155_400 ();
 b15zdnd11an1n64x5 FILLER_155_464 ();
 b15zdnd11an1n64x5 FILLER_155_528 ();
 b15zdnd11an1n64x5 FILLER_155_592 ();
 b15zdnd11an1n64x5 FILLER_155_656 ();
 b15zdnd11an1n64x5 FILLER_155_720 ();
 b15zdnd11an1n64x5 FILLER_155_784 ();
 b15zdnd11an1n64x5 FILLER_155_848 ();
 b15zdnd11an1n64x5 FILLER_155_912 ();
 b15zdnd11an1n64x5 FILLER_155_976 ();
 b15zdnd11an1n64x5 FILLER_155_1040 ();
 b15zdnd11an1n64x5 FILLER_155_1104 ();
 b15zdnd11an1n64x5 FILLER_155_1168 ();
 b15zdnd11an1n64x5 FILLER_155_1232 ();
 b15zdnd11an1n64x5 FILLER_155_1296 ();
 b15zdnd11an1n64x5 FILLER_155_1360 ();
 b15zdnd11an1n32x5 FILLER_155_1424 ();
 b15zdnd11an1n04x5 FILLER_155_1456 ();
 b15zdnd00an1n02x5 FILLER_155_1460 ();
 b15zdnd11an1n64x5 FILLER_155_1504 ();
 b15zdnd11an1n64x5 FILLER_155_1568 ();
 b15zdnd11an1n64x5 FILLER_155_1632 ();
 b15zdnd11an1n16x5 FILLER_155_1696 ();
 b15zdnd11an1n08x5 FILLER_155_1712 ();
 b15zdnd11an1n04x5 FILLER_155_1720 ();
 b15zdnd00an1n01x5 FILLER_155_1724 ();
 b15zdnd11an1n32x5 FILLER_155_1739 ();
 b15zdnd11an1n16x5 FILLER_155_1771 ();
 b15zdnd11an1n08x5 FILLER_155_1787 ();
 b15zdnd00an1n02x5 FILLER_155_1795 ();
 b15zdnd00an1n01x5 FILLER_155_1797 ();
 b15zdnd11an1n64x5 FILLER_155_1801 ();
 b15zdnd11an1n64x5 FILLER_155_1865 ();
 b15zdnd11an1n64x5 FILLER_155_1929 ();
 b15zdnd11an1n64x5 FILLER_155_1993 ();
 b15zdnd11an1n64x5 FILLER_155_2057 ();
 b15zdnd11an1n64x5 FILLER_155_2121 ();
 b15zdnd11an1n64x5 FILLER_155_2185 ();
 b15zdnd11an1n32x5 FILLER_155_2249 ();
 b15zdnd00an1n02x5 FILLER_155_2281 ();
 b15zdnd00an1n01x5 FILLER_155_2283 ();
 b15zdnd11an1n64x5 FILLER_156_8 ();
 b15zdnd11an1n64x5 FILLER_156_72 ();
 b15zdnd11an1n64x5 FILLER_156_136 ();
 b15zdnd11an1n64x5 FILLER_156_200 ();
 b15zdnd11an1n32x5 FILLER_156_264 ();
 b15zdnd11an1n04x5 FILLER_156_296 ();
 b15zdnd11an1n04x5 FILLER_156_303 ();
 b15zdnd11an1n04x5 FILLER_156_310 ();
 b15zdnd11an1n04x5 FILLER_156_317 ();
 b15zdnd11an1n64x5 FILLER_156_324 ();
 b15zdnd11an1n32x5 FILLER_156_388 ();
 b15zdnd11an1n04x5 FILLER_156_420 ();
 b15zdnd00an1n02x5 FILLER_156_424 ();
 b15zdnd11an1n64x5 FILLER_156_434 ();
 b15zdnd11an1n32x5 FILLER_156_498 ();
 b15zdnd11an1n16x5 FILLER_156_530 ();
 b15zdnd11an1n08x5 FILLER_156_546 ();
 b15zdnd11an1n04x5 FILLER_156_554 ();
 b15zdnd00an1n01x5 FILLER_156_558 ();
 b15zdnd11an1n64x5 FILLER_156_573 ();
 b15zdnd11an1n64x5 FILLER_156_637 ();
 b15zdnd11an1n16x5 FILLER_156_701 ();
 b15zdnd00an1n01x5 FILLER_156_717 ();
 b15zdnd11an1n64x5 FILLER_156_726 ();
 b15zdnd11an1n32x5 FILLER_156_790 ();
 b15zdnd11an1n16x5 FILLER_156_822 ();
 b15zdnd11an1n08x5 FILLER_156_838 ();
 b15zdnd00an1n02x5 FILLER_156_846 ();
 b15zdnd11an1n64x5 FILLER_156_868 ();
 b15zdnd11an1n16x5 FILLER_156_932 ();
 b15zdnd11an1n08x5 FILLER_156_948 ();
 b15zdnd00an1n02x5 FILLER_156_956 ();
 b15zdnd00an1n01x5 FILLER_156_958 ();
 b15zdnd11an1n64x5 FILLER_156_972 ();
 b15zdnd11an1n64x5 FILLER_156_1036 ();
 b15zdnd11an1n64x5 FILLER_156_1100 ();
 b15zdnd11an1n64x5 FILLER_156_1164 ();
 b15zdnd11an1n64x5 FILLER_156_1228 ();
 b15zdnd11an1n64x5 FILLER_156_1292 ();
 b15zdnd11an1n64x5 FILLER_156_1356 ();
 b15zdnd11an1n64x5 FILLER_156_1420 ();
 b15zdnd11an1n64x5 FILLER_156_1484 ();
 b15zdnd11an1n64x5 FILLER_156_1548 ();
 b15zdnd11an1n64x5 FILLER_156_1612 ();
 b15zdnd11an1n32x5 FILLER_156_1676 ();
 b15zdnd00an1n02x5 FILLER_156_1708 ();
 b15zdnd00an1n01x5 FILLER_156_1710 ();
 b15zdnd11an1n04x5 FILLER_156_1714 ();
 b15zdnd11an1n32x5 FILLER_156_1732 ();
 b15zdnd11an1n16x5 FILLER_156_1764 ();
 b15zdnd00an1n02x5 FILLER_156_1780 ();
 b15zdnd00an1n01x5 FILLER_156_1782 ();
 b15zdnd11an1n32x5 FILLER_156_1825 ();
 b15zdnd11an1n16x5 FILLER_156_1857 ();
 b15zdnd11an1n08x5 FILLER_156_1873 ();
 b15zdnd11an1n64x5 FILLER_156_1884 ();
 b15zdnd11an1n64x5 FILLER_156_1948 ();
 b15zdnd11an1n64x5 FILLER_156_2012 ();
 b15zdnd11an1n64x5 FILLER_156_2076 ();
 b15zdnd11an1n08x5 FILLER_156_2140 ();
 b15zdnd11an1n04x5 FILLER_156_2148 ();
 b15zdnd00an1n02x5 FILLER_156_2152 ();
 b15zdnd11an1n64x5 FILLER_156_2162 ();
 b15zdnd11an1n32x5 FILLER_156_2226 ();
 b15zdnd11an1n16x5 FILLER_156_2258 ();
 b15zdnd00an1n02x5 FILLER_156_2274 ();
 b15zdnd11an1n64x5 FILLER_157_0 ();
 b15zdnd11an1n64x5 FILLER_157_64 ();
 b15zdnd11an1n64x5 FILLER_157_128 ();
 b15zdnd11an1n64x5 FILLER_157_192 ();
 b15zdnd11an1n32x5 FILLER_157_256 ();
 b15zdnd11an1n16x5 FILLER_157_288 ();
 b15zdnd11an1n04x5 FILLER_157_304 ();
 b15zdnd00an1n02x5 FILLER_157_308 ();
 b15zdnd11an1n64x5 FILLER_157_313 ();
 b15zdnd11an1n16x5 FILLER_157_377 ();
 b15zdnd11an1n08x5 FILLER_157_393 ();
 b15zdnd11an1n04x5 FILLER_157_401 ();
 b15zdnd00an1n02x5 FILLER_157_405 ();
 b15zdnd11an1n64x5 FILLER_157_446 ();
 b15zdnd11an1n64x5 FILLER_157_510 ();
 b15zdnd11an1n64x5 FILLER_157_574 ();
 b15zdnd11an1n16x5 FILLER_157_638 ();
 b15zdnd11an1n64x5 FILLER_157_662 ();
 b15zdnd11an1n64x5 FILLER_157_726 ();
 b15zdnd11an1n64x5 FILLER_157_790 ();
 b15zdnd11an1n64x5 FILLER_157_854 ();
 b15zdnd11an1n64x5 FILLER_157_918 ();
 b15zdnd11an1n64x5 FILLER_157_982 ();
 b15zdnd11an1n64x5 FILLER_157_1046 ();
 b15zdnd11an1n32x5 FILLER_157_1110 ();
 b15zdnd00an1n01x5 FILLER_157_1142 ();
 b15zdnd11an1n64x5 FILLER_157_1146 ();
 b15zdnd11an1n64x5 FILLER_157_1210 ();
 b15zdnd11an1n64x5 FILLER_157_1274 ();
 b15zdnd11an1n64x5 FILLER_157_1338 ();
 b15zdnd11an1n64x5 FILLER_157_1402 ();
 b15zdnd11an1n64x5 FILLER_157_1466 ();
 b15zdnd11an1n64x5 FILLER_157_1530 ();
 b15zdnd11an1n64x5 FILLER_157_1594 ();
 b15zdnd11an1n32x5 FILLER_157_1658 ();
 b15zdnd11an1n04x5 FILLER_157_1690 ();
 b15zdnd11an1n64x5 FILLER_157_1720 ();
 b15zdnd00an1n02x5 FILLER_157_1784 ();
 b15zdnd00an1n01x5 FILLER_157_1786 ();
 b15zdnd11an1n32x5 FILLER_157_1801 ();
 b15zdnd11an1n04x5 FILLER_157_1833 ();
 b15zdnd00an1n01x5 FILLER_157_1837 ();
 b15zdnd11an1n04x5 FILLER_157_1882 ();
 b15zdnd11an1n04x5 FILLER_157_1889 ();
 b15zdnd11an1n64x5 FILLER_157_1896 ();
 b15zdnd11an1n64x5 FILLER_157_1960 ();
 b15zdnd11an1n32x5 FILLER_157_2024 ();
 b15zdnd11an1n08x5 FILLER_157_2056 ();
 b15zdnd00an1n02x5 FILLER_157_2064 ();
 b15zdnd00an1n01x5 FILLER_157_2066 ();
 b15zdnd11an1n04x5 FILLER_157_2099 ();
 b15zdnd11an1n64x5 FILLER_157_2106 ();
 b15zdnd11an1n16x5 FILLER_157_2170 ();
 b15zdnd11an1n08x5 FILLER_157_2186 ();
 b15zdnd11an1n04x5 FILLER_157_2194 ();
 b15zdnd00an1n02x5 FILLER_157_2198 ();
 b15zdnd00an1n01x5 FILLER_157_2200 ();
 b15zdnd11an1n64x5 FILLER_157_2206 ();
 b15zdnd11an1n08x5 FILLER_157_2270 ();
 b15zdnd11an1n04x5 FILLER_157_2278 ();
 b15zdnd00an1n02x5 FILLER_157_2282 ();
 b15zdnd11an1n64x5 FILLER_158_8 ();
 b15zdnd11an1n64x5 FILLER_158_72 ();
 b15zdnd11an1n64x5 FILLER_158_136 ();
 b15zdnd11an1n64x5 FILLER_158_200 ();
 b15zdnd11an1n64x5 FILLER_158_264 ();
 b15zdnd11an1n64x5 FILLER_158_328 ();
 b15zdnd11an1n32x5 FILLER_158_392 ();
 b15zdnd11an1n16x5 FILLER_158_424 ();
 b15zdnd00an1n02x5 FILLER_158_440 ();
 b15zdnd00an1n01x5 FILLER_158_442 ();
 b15zdnd11an1n32x5 FILLER_158_451 ();
 b15zdnd11an1n16x5 FILLER_158_483 ();
 b15zdnd11an1n08x5 FILLER_158_499 ();
 b15zdnd11an1n04x5 FILLER_158_507 ();
 b15zdnd11an1n64x5 FILLER_158_538 ();
 b15zdnd11an1n64x5 FILLER_158_602 ();
 b15zdnd11an1n32x5 FILLER_158_666 ();
 b15zdnd11an1n16x5 FILLER_158_698 ();
 b15zdnd11an1n04x5 FILLER_158_714 ();
 b15zdnd11an1n64x5 FILLER_158_726 ();
 b15zdnd11an1n64x5 FILLER_158_790 ();
 b15zdnd11an1n64x5 FILLER_158_854 ();
 b15zdnd11an1n64x5 FILLER_158_918 ();
 b15zdnd00an1n01x5 FILLER_158_982 ();
 b15zdnd11an1n04x5 FILLER_158_986 ();
 b15zdnd11an1n64x5 FILLER_158_993 ();
 b15zdnd11an1n32x5 FILLER_158_1057 ();
 b15zdnd11an1n16x5 FILLER_158_1089 ();
 b15zdnd11an1n08x5 FILLER_158_1105 ();
 b15zdnd11an1n04x5 FILLER_158_1113 ();
 b15zdnd00an1n01x5 FILLER_158_1117 ();
 b15zdnd11an1n64x5 FILLER_158_1170 ();
 b15zdnd11an1n64x5 FILLER_158_1234 ();
 b15zdnd11an1n64x5 FILLER_158_1298 ();
 b15zdnd11an1n64x5 FILLER_158_1362 ();
 b15zdnd11an1n64x5 FILLER_158_1426 ();
 b15zdnd11an1n64x5 FILLER_158_1490 ();
 b15zdnd11an1n32x5 FILLER_158_1554 ();
 b15zdnd11an1n16x5 FILLER_158_1586 ();
 b15zdnd11an1n08x5 FILLER_158_1602 ();
 b15zdnd00an1n01x5 FILLER_158_1610 ();
 b15zdnd11an1n16x5 FILLER_158_1619 ();
 b15zdnd11an1n08x5 FILLER_158_1635 ();
 b15zdnd11an1n04x5 FILLER_158_1643 ();
 b15zdnd00an1n02x5 FILLER_158_1647 ();
 b15zdnd00an1n01x5 FILLER_158_1649 ();
 b15zdnd11an1n32x5 FILLER_158_1660 ();
 b15zdnd11an1n16x5 FILLER_158_1692 ();
 b15zdnd11an1n08x5 FILLER_158_1708 ();
 b15zdnd00an1n02x5 FILLER_158_1716 ();
 b15zdnd11an1n32x5 FILLER_158_1739 ();
 b15zdnd11an1n08x5 FILLER_158_1771 ();
 b15zdnd11an1n04x5 FILLER_158_1779 ();
 b15zdnd00an1n02x5 FILLER_158_1783 ();
 b15zdnd00an1n01x5 FILLER_158_1785 ();
 b15zdnd11an1n64x5 FILLER_158_1789 ();
 b15zdnd11an1n64x5 FILLER_158_1853 ();
 b15zdnd11an1n64x5 FILLER_158_1917 ();
 b15zdnd11an1n64x5 FILLER_158_1981 ();
 b15zdnd11an1n32x5 FILLER_158_2045 ();
 b15zdnd11an1n16x5 FILLER_158_2077 ();
 b15zdnd00an1n02x5 FILLER_158_2093 ();
 b15zdnd11an1n16x5 FILLER_158_2098 ();
 b15zdnd11an1n04x5 FILLER_158_2114 ();
 b15zdnd00an1n02x5 FILLER_158_2118 ();
 b15zdnd11an1n16x5 FILLER_158_2134 ();
 b15zdnd11an1n04x5 FILLER_158_2150 ();
 b15zdnd11an1n32x5 FILLER_158_2162 ();
 b15zdnd00an1n01x5 FILLER_158_2194 ();
 b15zdnd11an1n64x5 FILLER_158_2206 ();
 b15zdnd11an1n04x5 FILLER_158_2270 ();
 b15zdnd00an1n02x5 FILLER_158_2274 ();
 b15zdnd11an1n64x5 FILLER_159_0 ();
 b15zdnd11an1n64x5 FILLER_159_64 ();
 b15zdnd11an1n64x5 FILLER_159_128 ();
 b15zdnd11an1n64x5 FILLER_159_192 ();
 b15zdnd11an1n64x5 FILLER_159_256 ();
 b15zdnd11an1n64x5 FILLER_159_320 ();
 b15zdnd11an1n64x5 FILLER_159_384 ();
 b15zdnd11an1n32x5 FILLER_159_448 ();
 b15zdnd11an1n16x5 FILLER_159_480 ();
 b15zdnd11an1n08x5 FILLER_159_496 ();
 b15zdnd11an1n04x5 FILLER_159_504 ();
 b15zdnd00an1n02x5 FILLER_159_508 ();
 b15zdnd11an1n64x5 FILLER_159_513 ();
 b15zdnd11an1n64x5 FILLER_159_577 ();
 b15zdnd11an1n64x5 FILLER_159_641 ();
 b15zdnd11an1n64x5 FILLER_159_705 ();
 b15zdnd11an1n64x5 FILLER_159_769 ();
 b15zdnd11an1n64x5 FILLER_159_833 ();
 b15zdnd11an1n32x5 FILLER_159_897 ();
 b15zdnd11an1n16x5 FILLER_159_929 ();
 b15zdnd11an1n08x5 FILLER_159_945 ();
 b15zdnd11an1n04x5 FILLER_159_953 ();
 b15zdnd00an1n02x5 FILLER_159_957 ();
 b15zdnd00an1n01x5 FILLER_159_959 ();
 b15zdnd11an1n32x5 FILLER_159_1012 ();
 b15zdnd11an1n16x5 FILLER_159_1053 ();
 b15zdnd00an1n02x5 FILLER_159_1069 ();
 b15zdnd11an1n32x5 FILLER_159_1080 ();
 b15zdnd11an1n64x5 FILLER_159_1164 ();
 b15zdnd11an1n64x5 FILLER_159_1228 ();
 b15zdnd11an1n64x5 FILLER_159_1292 ();
 b15zdnd11an1n64x5 FILLER_159_1356 ();
 b15zdnd11an1n64x5 FILLER_159_1420 ();
 b15zdnd11an1n64x5 FILLER_159_1484 ();
 b15zdnd11an1n64x5 FILLER_159_1548 ();
 b15zdnd11an1n32x5 FILLER_159_1612 ();
 b15zdnd11an1n16x5 FILLER_159_1644 ();
 b15zdnd11an1n04x5 FILLER_159_1660 ();
 b15zdnd00an1n01x5 FILLER_159_1664 ();
 b15zdnd11an1n32x5 FILLER_159_1668 ();
 b15zdnd11an1n16x5 FILLER_159_1700 ();
 b15zdnd11an1n08x5 FILLER_159_1716 ();
 b15zdnd11an1n04x5 FILLER_159_1724 ();
 b15zdnd00an1n02x5 FILLER_159_1728 ();
 b15zdnd11an1n32x5 FILLER_159_1746 ();
 b15zdnd11an1n08x5 FILLER_159_1778 ();
 b15zdnd00an1n01x5 FILLER_159_1786 ();
 b15zdnd11an1n64x5 FILLER_159_1800 ();
 b15zdnd11an1n64x5 FILLER_159_1864 ();
 b15zdnd11an1n64x5 FILLER_159_1928 ();
 b15zdnd11an1n32x5 FILLER_159_1992 ();
 b15zdnd11an1n16x5 FILLER_159_2024 ();
 b15zdnd11an1n08x5 FILLER_159_2040 ();
 b15zdnd00an1n01x5 FILLER_159_2048 ();
 b15zdnd11an1n04x5 FILLER_159_2089 ();
 b15zdnd11an1n64x5 FILLER_159_2096 ();
 b15zdnd11an1n32x5 FILLER_159_2160 ();
 b15zdnd11an1n08x5 FILLER_159_2192 ();
 b15zdnd11an1n04x5 FILLER_159_2200 ();
 b15zdnd00an1n02x5 FILLER_159_2204 ();
 b15zdnd00an1n01x5 FILLER_159_2206 ();
 b15zdnd11an1n08x5 FILLER_159_2210 ();
 b15zdnd00an1n02x5 FILLER_159_2218 ();
 b15zdnd00an1n01x5 FILLER_159_2220 ();
 b15zdnd11an1n32x5 FILLER_159_2224 ();
 b15zdnd11an1n16x5 FILLER_159_2256 ();
 b15zdnd11an1n08x5 FILLER_159_2272 ();
 b15zdnd11an1n04x5 FILLER_159_2280 ();
 b15zdnd11an1n64x5 FILLER_160_8 ();
 b15zdnd11an1n64x5 FILLER_160_72 ();
 b15zdnd11an1n16x5 FILLER_160_136 ();
 b15zdnd11an1n04x5 FILLER_160_152 ();
 b15zdnd00an1n02x5 FILLER_160_156 ();
 b15zdnd11an1n64x5 FILLER_160_162 ();
 b15zdnd11an1n64x5 FILLER_160_226 ();
 b15zdnd11an1n64x5 FILLER_160_290 ();
 b15zdnd11an1n64x5 FILLER_160_354 ();
 b15zdnd11an1n64x5 FILLER_160_418 ();
 b15zdnd11an1n64x5 FILLER_160_482 ();
 b15zdnd11an1n64x5 FILLER_160_546 ();
 b15zdnd11an1n64x5 FILLER_160_610 ();
 b15zdnd11an1n32x5 FILLER_160_674 ();
 b15zdnd11an1n08x5 FILLER_160_706 ();
 b15zdnd11an1n04x5 FILLER_160_714 ();
 b15zdnd11an1n64x5 FILLER_160_726 ();
 b15zdnd11an1n64x5 FILLER_160_790 ();
 b15zdnd11an1n64x5 FILLER_160_854 ();
 b15zdnd11an1n32x5 FILLER_160_918 ();
 b15zdnd11an1n08x5 FILLER_160_950 ();
 b15zdnd11an1n04x5 FILLER_160_958 ();
 b15zdnd00an1n02x5 FILLER_160_962 ();
 b15zdnd11an1n64x5 FILLER_160_1016 ();
 b15zdnd11an1n32x5 FILLER_160_1080 ();
 b15zdnd11an1n16x5 FILLER_160_1112 ();
 b15zdnd00an1n02x5 FILLER_160_1128 ();
 b15zdnd00an1n01x5 FILLER_160_1130 ();
 b15zdnd11an1n04x5 FILLER_160_1134 ();
 b15zdnd11an1n04x5 FILLER_160_1141 ();
 b15zdnd11an1n64x5 FILLER_160_1148 ();
 b15zdnd11an1n64x5 FILLER_160_1212 ();
 b15zdnd11an1n08x5 FILLER_160_1276 ();
 b15zdnd11an1n04x5 FILLER_160_1284 ();
 b15zdnd00an1n01x5 FILLER_160_1288 ();
 b15zdnd11an1n64x5 FILLER_160_1310 ();
 b15zdnd11an1n64x5 FILLER_160_1374 ();
 b15zdnd11an1n64x5 FILLER_160_1438 ();
 b15zdnd11an1n64x5 FILLER_160_1502 ();
 b15zdnd11an1n64x5 FILLER_160_1566 ();
 b15zdnd11an1n64x5 FILLER_160_1630 ();
 b15zdnd11an1n16x5 FILLER_160_1694 ();
 b15zdnd11an1n08x5 FILLER_160_1727 ();
 b15zdnd11an1n64x5 FILLER_160_1743 ();
 b15zdnd11an1n32x5 FILLER_160_1807 ();
 b15zdnd11an1n16x5 FILLER_160_1839 ();
 b15zdnd11an1n04x5 FILLER_160_1855 ();
 b15zdnd00an1n02x5 FILLER_160_1859 ();
 b15zdnd11an1n64x5 FILLER_160_1881 ();
 b15zdnd11an1n32x5 FILLER_160_1945 ();
 b15zdnd11an1n08x5 FILLER_160_1977 ();
 b15zdnd11an1n04x5 FILLER_160_1985 ();
 b15zdnd00an1n01x5 FILLER_160_1989 ();
 b15zdnd11an1n64x5 FILLER_160_2016 ();
 b15zdnd11an1n04x5 FILLER_160_2080 ();
 b15zdnd00an1n01x5 FILLER_160_2084 ();
 b15zdnd11an1n32x5 FILLER_160_2088 ();
 b15zdnd11an1n08x5 FILLER_160_2120 ();
 b15zdnd00an1n02x5 FILLER_160_2128 ();
 b15zdnd00an1n02x5 FILLER_160_2152 ();
 b15zdnd11an1n32x5 FILLER_160_2162 ();
 b15zdnd11an1n08x5 FILLER_160_2194 ();
 b15zdnd00an1n02x5 FILLER_160_2202 ();
 b15zdnd11an1n08x5 FILLER_160_2217 ();
 b15zdnd11an1n32x5 FILLER_160_2237 ();
 b15zdnd11an1n04x5 FILLER_160_2269 ();
 b15zdnd00an1n02x5 FILLER_160_2273 ();
 b15zdnd00an1n01x5 FILLER_160_2275 ();
 b15zdnd11an1n64x5 FILLER_161_0 ();
 b15zdnd11an1n64x5 FILLER_161_64 ();
 b15zdnd11an1n16x5 FILLER_161_128 ();
 b15zdnd11an1n08x5 FILLER_161_158 ();
 b15zdnd00an1n02x5 FILLER_161_166 ();
 b15zdnd00an1n01x5 FILLER_161_168 ();
 b15zdnd11an1n64x5 FILLER_161_172 ();
 b15zdnd11an1n64x5 FILLER_161_236 ();
 b15zdnd11an1n64x5 FILLER_161_300 ();
 b15zdnd11an1n64x5 FILLER_161_364 ();
 b15zdnd11an1n64x5 FILLER_161_428 ();
 b15zdnd11an1n64x5 FILLER_161_492 ();
 b15zdnd11an1n08x5 FILLER_161_556 ();
 b15zdnd11an1n04x5 FILLER_161_564 ();
 b15zdnd00an1n01x5 FILLER_161_568 ();
 b15zdnd11an1n64x5 FILLER_161_573 ();
 b15zdnd11an1n64x5 FILLER_161_637 ();
 b15zdnd11an1n64x5 FILLER_161_701 ();
 b15zdnd11an1n64x5 FILLER_161_765 ();
 b15zdnd11an1n64x5 FILLER_161_829 ();
 b15zdnd11an1n64x5 FILLER_161_893 ();
 b15zdnd11an1n16x5 FILLER_161_957 ();
 b15zdnd11an1n04x5 FILLER_161_973 ();
 b15zdnd11an1n04x5 FILLER_161_980 ();
 b15zdnd11an1n04x5 FILLER_161_987 ();
 b15zdnd11an1n64x5 FILLER_161_994 ();
 b15zdnd11an1n64x5 FILLER_161_1058 ();
 b15zdnd11an1n16x5 FILLER_161_1122 ();
 b15zdnd11an1n04x5 FILLER_161_1141 ();
 b15zdnd11an1n64x5 FILLER_161_1148 ();
 b15zdnd11an1n32x5 FILLER_161_1212 ();
 b15zdnd11an1n08x5 FILLER_161_1244 ();
 b15zdnd00an1n02x5 FILLER_161_1252 ();
 b15zdnd11an1n64x5 FILLER_161_1280 ();
 b15zdnd11an1n64x5 FILLER_161_1344 ();
 b15zdnd11an1n64x5 FILLER_161_1408 ();
 b15zdnd11an1n64x5 FILLER_161_1472 ();
 b15zdnd11an1n32x5 FILLER_161_1536 ();
 b15zdnd11an1n16x5 FILLER_161_1568 ();
 b15zdnd11an1n04x5 FILLER_161_1584 ();
 b15zdnd11an1n64x5 FILLER_161_1592 ();
 b15zdnd11an1n64x5 FILLER_161_1656 ();
 b15zdnd11an1n64x5 FILLER_161_1720 ();
 b15zdnd11an1n32x5 FILLER_161_1784 ();
 b15zdnd11an1n16x5 FILLER_161_1816 ();
 b15zdnd11an1n04x5 FILLER_161_1832 ();
 b15zdnd00an1n02x5 FILLER_161_1836 ();
 b15zdnd11an1n64x5 FILLER_161_1844 ();
 b15zdnd11an1n32x5 FILLER_161_1908 ();
 b15zdnd11an1n16x5 FILLER_161_1940 ();
 b15zdnd11an1n08x5 FILLER_161_1956 ();
 b15zdnd11an1n64x5 FILLER_161_1967 ();
 b15zdnd11an1n64x5 FILLER_161_2031 ();
 b15zdnd11an1n64x5 FILLER_161_2095 ();
 b15zdnd11an1n32x5 FILLER_161_2159 ();
 b15zdnd11an1n08x5 FILLER_161_2191 ();
 b15zdnd11an1n04x5 FILLER_161_2241 ();
 b15zdnd11an1n16x5 FILLER_161_2259 ();
 b15zdnd11an1n08x5 FILLER_161_2275 ();
 b15zdnd00an1n01x5 FILLER_161_2283 ();
 b15zdnd11an1n64x5 FILLER_162_8 ();
 b15zdnd11an1n64x5 FILLER_162_72 ();
 b15zdnd11an1n08x5 FILLER_162_136 ();
 b15zdnd00an1n01x5 FILLER_162_144 ();
 b15zdnd11an1n64x5 FILLER_162_152 ();
 b15zdnd11an1n64x5 FILLER_162_216 ();
 b15zdnd11an1n16x5 FILLER_162_280 ();
 b15zdnd00an1n02x5 FILLER_162_296 ();
 b15zdnd00an1n01x5 FILLER_162_298 ();
 b15zdnd11an1n64x5 FILLER_162_304 ();
 b15zdnd11an1n64x5 FILLER_162_368 ();
 b15zdnd11an1n64x5 FILLER_162_432 ();
 b15zdnd11an1n32x5 FILLER_162_496 ();
 b15zdnd11an1n16x5 FILLER_162_528 ();
 b15zdnd11an1n08x5 FILLER_162_544 ();
 b15zdnd11an1n04x5 FILLER_162_552 ();
 b15zdnd00an1n02x5 FILLER_162_556 ();
 b15zdnd00an1n01x5 FILLER_162_558 ();
 b15zdnd11an1n64x5 FILLER_162_563 ();
 b15zdnd11an1n64x5 FILLER_162_627 ();
 b15zdnd11an1n16x5 FILLER_162_691 ();
 b15zdnd11an1n08x5 FILLER_162_707 ();
 b15zdnd00an1n02x5 FILLER_162_715 ();
 b15zdnd00an1n01x5 FILLER_162_717 ();
 b15zdnd11an1n64x5 FILLER_162_726 ();
 b15zdnd11an1n16x5 FILLER_162_790 ();
 b15zdnd11an1n08x5 FILLER_162_806 ();
 b15zdnd11an1n04x5 FILLER_162_814 ();
 b15zdnd00an1n02x5 FILLER_162_818 ();
 b15zdnd11an1n64x5 FILLER_162_827 ();
 b15zdnd11an1n64x5 FILLER_162_891 ();
 b15zdnd11an1n32x5 FILLER_162_955 ();
 b15zdnd00an1n02x5 FILLER_162_987 ();
 b15zdnd11an1n64x5 FILLER_162_992 ();
 b15zdnd11an1n32x5 FILLER_162_1056 ();
 b15zdnd11an1n16x5 FILLER_162_1088 ();
 b15zdnd11an1n08x5 FILLER_162_1104 ();
 b15zdnd11an1n04x5 FILLER_162_1139 ();
 b15zdnd11an1n08x5 FILLER_162_1146 ();
 b15zdnd00an1n02x5 FILLER_162_1154 ();
 b15zdnd00an1n01x5 FILLER_162_1156 ();
 b15zdnd11an1n64x5 FILLER_162_1183 ();
 b15zdnd11an1n64x5 FILLER_162_1247 ();
 b15zdnd11an1n64x5 FILLER_162_1311 ();
 b15zdnd11an1n32x5 FILLER_162_1375 ();
 b15zdnd11an1n16x5 FILLER_162_1407 ();
 b15zdnd00an1n02x5 FILLER_162_1423 ();
 b15zdnd11an1n32x5 FILLER_162_1428 ();
 b15zdnd11an1n16x5 FILLER_162_1460 ();
 b15zdnd00an1n02x5 FILLER_162_1476 ();
 b15zdnd00an1n01x5 FILLER_162_1478 ();
 b15zdnd11an1n64x5 FILLER_162_1484 ();
 b15zdnd11an1n64x5 FILLER_162_1548 ();
 b15zdnd11an1n64x5 FILLER_162_1612 ();
 b15zdnd11an1n16x5 FILLER_162_1676 ();
 b15zdnd11an1n04x5 FILLER_162_1692 ();
 b15zdnd00an1n02x5 FILLER_162_1696 ();
 b15zdnd11an1n64x5 FILLER_162_1706 ();
 b15zdnd11an1n64x5 FILLER_162_1770 ();
 b15zdnd11an1n64x5 FILLER_162_1834 ();
 b15zdnd11an1n32x5 FILLER_162_1898 ();
 b15zdnd11an1n08x5 FILLER_162_1930 ();
 b15zdnd11an1n32x5 FILLER_162_1990 ();
 b15zdnd11an1n16x5 FILLER_162_2022 ();
 b15zdnd00an1n01x5 FILLER_162_2038 ();
 b15zdnd11an1n64x5 FILLER_162_2060 ();
 b15zdnd11an1n16x5 FILLER_162_2124 ();
 b15zdnd11an1n08x5 FILLER_162_2140 ();
 b15zdnd11an1n04x5 FILLER_162_2148 ();
 b15zdnd00an1n02x5 FILLER_162_2152 ();
 b15zdnd11an1n16x5 FILLER_162_2162 ();
 b15zdnd11an1n08x5 FILLER_162_2178 ();
 b15zdnd00an1n01x5 FILLER_162_2186 ();
 b15zdnd11an1n32x5 FILLER_162_2239 ();
 b15zdnd11an1n04x5 FILLER_162_2271 ();
 b15zdnd00an1n01x5 FILLER_162_2275 ();
 b15zdnd11an1n64x5 FILLER_163_0 ();
 b15zdnd11an1n64x5 FILLER_163_64 ();
 b15zdnd11an1n64x5 FILLER_163_128 ();
 b15zdnd11an1n64x5 FILLER_163_192 ();
 b15zdnd11an1n64x5 FILLER_163_256 ();
 b15zdnd11an1n64x5 FILLER_163_320 ();
 b15zdnd11an1n64x5 FILLER_163_384 ();
 b15zdnd11an1n64x5 FILLER_163_448 ();
 b15zdnd11an1n64x5 FILLER_163_512 ();
 b15zdnd11an1n64x5 FILLER_163_576 ();
 b15zdnd11an1n64x5 FILLER_163_640 ();
 b15zdnd11an1n32x5 FILLER_163_704 ();
 b15zdnd11an1n04x5 FILLER_163_736 ();
 b15zdnd00an1n02x5 FILLER_163_740 ();
 b15zdnd11an1n64x5 FILLER_163_746 ();
 b15zdnd11an1n64x5 FILLER_163_810 ();
 b15zdnd11an1n64x5 FILLER_163_874 ();
 b15zdnd11an1n64x5 FILLER_163_938 ();
 b15zdnd11an1n64x5 FILLER_163_1002 ();
 b15zdnd11an1n04x5 FILLER_163_1066 ();
 b15zdnd00an1n02x5 FILLER_163_1070 ();
 b15zdnd11an1n16x5 FILLER_163_1081 ();
 b15zdnd11an1n08x5 FILLER_163_1097 ();
 b15zdnd11an1n04x5 FILLER_163_1105 ();
 b15zdnd00an1n02x5 FILLER_163_1109 ();
 b15zdnd00an1n01x5 FILLER_163_1111 ();
 b15zdnd11an1n04x5 FILLER_163_1115 ();
 b15zdnd11an1n64x5 FILLER_163_1171 ();
 b15zdnd11an1n64x5 FILLER_163_1235 ();
 b15zdnd11an1n64x5 FILLER_163_1299 ();
 b15zdnd11an1n16x5 FILLER_163_1363 ();
 b15zdnd11an1n08x5 FILLER_163_1379 ();
 b15zdnd00an1n02x5 FILLER_163_1387 ();
 b15zdnd00an1n01x5 FILLER_163_1389 ();
 b15zdnd11an1n04x5 FILLER_163_1395 ();
 b15zdnd11an1n16x5 FILLER_163_1451 ();
 b15zdnd11an1n08x5 FILLER_163_1467 ();
 b15zdnd00an1n02x5 FILLER_163_1475 ();
 b15zdnd00an1n01x5 FILLER_163_1477 ();
 b15zdnd11an1n32x5 FILLER_163_1520 ();
 b15zdnd00an1n01x5 FILLER_163_1552 ();
 b15zdnd11an1n32x5 FILLER_163_1561 ();
 b15zdnd11an1n16x5 FILLER_163_1593 ();
 b15zdnd11an1n64x5 FILLER_163_1661 ();
 b15zdnd11an1n64x5 FILLER_163_1725 ();
 b15zdnd11an1n64x5 FILLER_163_1789 ();
 b15zdnd11an1n64x5 FILLER_163_1853 ();
 b15zdnd11an1n32x5 FILLER_163_1917 ();
 b15zdnd11an1n08x5 FILLER_163_1949 ();
 b15zdnd11an1n04x5 FILLER_163_1960 ();
 b15zdnd11an1n64x5 FILLER_163_1967 ();
 b15zdnd11an1n64x5 FILLER_163_2031 ();
 b15zdnd11an1n64x5 FILLER_163_2095 ();
 b15zdnd11an1n32x5 FILLER_163_2159 ();
 b15zdnd11an1n04x5 FILLER_163_2191 ();
 b15zdnd00an1n01x5 FILLER_163_2195 ();
 b15zdnd11an1n04x5 FILLER_163_2209 ();
 b15zdnd11an1n64x5 FILLER_163_2216 ();
 b15zdnd11an1n04x5 FILLER_163_2280 ();
 b15zdnd11an1n64x5 FILLER_164_8 ();
 b15zdnd11an1n64x5 FILLER_164_72 ();
 b15zdnd11an1n64x5 FILLER_164_136 ();
 b15zdnd11an1n64x5 FILLER_164_200 ();
 b15zdnd11an1n16x5 FILLER_164_264 ();
 b15zdnd11an1n08x5 FILLER_164_280 ();
 b15zdnd11an1n04x5 FILLER_164_288 ();
 b15zdnd11an1n64x5 FILLER_164_307 ();
 b15zdnd11an1n64x5 FILLER_164_371 ();
 b15zdnd11an1n32x5 FILLER_164_435 ();
 b15zdnd11an1n16x5 FILLER_164_467 ();
 b15zdnd11an1n08x5 FILLER_164_483 ();
 b15zdnd00an1n02x5 FILLER_164_491 ();
 b15zdnd00an1n01x5 FILLER_164_493 ();
 b15zdnd11an1n64x5 FILLER_164_497 ();
 b15zdnd11an1n64x5 FILLER_164_561 ();
 b15zdnd11an1n64x5 FILLER_164_625 ();
 b15zdnd11an1n16x5 FILLER_164_689 ();
 b15zdnd11an1n08x5 FILLER_164_705 ();
 b15zdnd11an1n04x5 FILLER_164_713 ();
 b15zdnd00an1n01x5 FILLER_164_717 ();
 b15zdnd11an1n64x5 FILLER_164_726 ();
 b15zdnd11an1n64x5 FILLER_164_790 ();
 b15zdnd11an1n64x5 FILLER_164_854 ();
 b15zdnd11an1n64x5 FILLER_164_918 ();
 b15zdnd11an1n04x5 FILLER_164_982 ();
 b15zdnd00an1n02x5 FILLER_164_986 ();
 b15zdnd11an1n64x5 FILLER_164_991 ();
 b15zdnd11an1n64x5 FILLER_164_1055 ();
 b15zdnd11an1n16x5 FILLER_164_1119 ();
 b15zdnd11an1n08x5 FILLER_164_1135 ();
 b15zdnd00an1n01x5 FILLER_164_1143 ();
 b15zdnd11an1n16x5 FILLER_164_1147 ();
 b15zdnd11an1n08x5 FILLER_164_1163 ();
 b15zdnd00an1n02x5 FILLER_164_1171 ();
 b15zdnd11an1n64x5 FILLER_164_1193 ();
 b15zdnd11an1n32x5 FILLER_164_1257 ();
 b15zdnd00an1n02x5 FILLER_164_1289 ();
 b15zdnd11an1n64x5 FILLER_164_1297 ();
 b15zdnd11an1n32x5 FILLER_164_1361 ();
 b15zdnd11an1n16x5 FILLER_164_1393 ();
 b15zdnd11an1n08x5 FILLER_164_1409 ();
 b15zdnd11an1n04x5 FILLER_164_1417 ();
 b15zdnd00an1n02x5 FILLER_164_1421 ();
 b15zdnd00an1n01x5 FILLER_164_1423 ();
 b15zdnd11an1n04x5 FILLER_164_1427 ();
 b15zdnd11an1n32x5 FILLER_164_1434 ();
 b15zdnd11an1n08x5 FILLER_164_1466 ();
 b15zdnd00an1n02x5 FILLER_164_1474 ();
 b15zdnd00an1n01x5 FILLER_164_1476 ();
 b15zdnd11an1n64x5 FILLER_164_1487 ();
 b15zdnd11an1n64x5 FILLER_164_1551 ();
 b15zdnd11an1n08x5 FILLER_164_1615 ();
 b15zdnd11an1n04x5 FILLER_164_1623 ();
 b15zdnd11an1n04x5 FILLER_164_1630 ();
 b15zdnd11an1n04x5 FILLER_164_1637 ();
 b15zdnd11an1n64x5 FILLER_164_1644 ();
 b15zdnd11an1n64x5 FILLER_164_1708 ();
 b15zdnd11an1n16x5 FILLER_164_1772 ();
 b15zdnd11an1n04x5 FILLER_164_1788 ();
 b15zdnd00an1n02x5 FILLER_164_1792 ();
 b15zdnd00an1n01x5 FILLER_164_1794 ();
 b15zdnd11an1n04x5 FILLER_164_1816 ();
 b15zdnd11an1n64x5 FILLER_164_1832 ();
 b15zdnd11an1n64x5 FILLER_164_1908 ();
 b15zdnd11an1n64x5 FILLER_164_1972 ();
 b15zdnd11an1n64x5 FILLER_164_2036 ();
 b15zdnd11an1n32x5 FILLER_164_2100 ();
 b15zdnd11an1n16x5 FILLER_164_2132 ();
 b15zdnd11an1n04x5 FILLER_164_2148 ();
 b15zdnd00an1n02x5 FILLER_164_2152 ();
 b15zdnd11an1n32x5 FILLER_164_2162 ();
 b15zdnd00an1n02x5 FILLER_164_2194 ();
 b15zdnd11an1n08x5 FILLER_164_2206 ();
 b15zdnd11an1n04x5 FILLER_164_2214 ();
 b15zdnd11an1n04x5 FILLER_164_2225 ();
 b15zdnd11an1n32x5 FILLER_164_2233 ();
 b15zdnd11an1n08x5 FILLER_164_2265 ();
 b15zdnd00an1n02x5 FILLER_164_2273 ();
 b15zdnd00an1n01x5 FILLER_164_2275 ();
 b15zdnd11an1n64x5 FILLER_165_0 ();
 b15zdnd11an1n64x5 FILLER_165_64 ();
 b15zdnd11an1n08x5 FILLER_165_128 ();
 b15zdnd11an1n04x5 FILLER_165_136 ();
 b15zdnd00an1n02x5 FILLER_165_140 ();
 b15zdnd11an1n04x5 FILLER_165_155 ();
 b15zdnd11an1n64x5 FILLER_165_167 ();
 b15zdnd11an1n64x5 FILLER_165_231 ();
 b15zdnd11an1n32x5 FILLER_165_295 ();
 b15zdnd11an1n08x5 FILLER_165_327 ();
 b15zdnd00an1n01x5 FILLER_165_335 ();
 b15zdnd11an1n64x5 FILLER_165_350 ();
 b15zdnd11an1n32x5 FILLER_165_414 ();
 b15zdnd11an1n16x5 FILLER_165_446 ();
 b15zdnd11an1n04x5 FILLER_165_462 ();
 b15zdnd00an1n01x5 FILLER_165_466 ();
 b15zdnd11an1n64x5 FILLER_165_519 ();
 b15zdnd11an1n64x5 FILLER_165_583 ();
 b15zdnd11an1n16x5 FILLER_165_647 ();
 b15zdnd11an1n08x5 FILLER_165_663 ();
 b15zdnd00an1n02x5 FILLER_165_671 ();
 b15zdnd11an1n08x5 FILLER_165_676 ();
 b15zdnd11an1n04x5 FILLER_165_684 ();
 b15zdnd00an1n02x5 FILLER_165_688 ();
 b15zdnd11an1n64x5 FILLER_165_693 ();
 b15zdnd11an1n64x5 FILLER_165_757 ();
 b15zdnd11an1n64x5 FILLER_165_821 ();
 b15zdnd11an1n64x5 FILLER_165_885 ();
 b15zdnd11an1n08x5 FILLER_165_949 ();
 b15zdnd11an1n04x5 FILLER_165_957 ();
 b15zdnd11an1n64x5 FILLER_165_1013 ();
 b15zdnd11an1n32x5 FILLER_165_1077 ();
 b15zdnd11an1n16x5 FILLER_165_1109 ();
 b15zdnd11an1n08x5 FILLER_165_1125 ();
 b15zdnd11an1n04x5 FILLER_165_1133 ();
 b15zdnd00an1n02x5 FILLER_165_1137 ();
 b15zdnd00an1n01x5 FILLER_165_1139 ();
 b15zdnd11an1n64x5 FILLER_165_1143 ();
 b15zdnd11an1n64x5 FILLER_165_1207 ();
 b15zdnd11an1n64x5 FILLER_165_1271 ();
 b15zdnd11an1n64x5 FILLER_165_1335 ();
 b15zdnd11an1n64x5 FILLER_165_1399 ();
 b15zdnd11an1n16x5 FILLER_165_1463 ();
 b15zdnd11an1n08x5 FILLER_165_1479 ();
 b15zdnd11an1n04x5 FILLER_165_1487 ();
 b15zdnd00an1n02x5 FILLER_165_1491 ();
 b15zdnd00an1n01x5 FILLER_165_1493 ();
 b15zdnd11an1n64x5 FILLER_165_1514 ();
 b15zdnd11an1n64x5 FILLER_165_1578 ();
 b15zdnd11an1n64x5 FILLER_165_1642 ();
 b15zdnd11an1n64x5 FILLER_165_1706 ();
 b15zdnd11an1n32x5 FILLER_165_1770 ();
 b15zdnd11an1n04x5 FILLER_165_1802 ();
 b15zdnd00an1n01x5 FILLER_165_1806 ();
 b15zdnd11an1n08x5 FILLER_165_1814 ();
 b15zdnd00an1n02x5 FILLER_165_1822 ();
 b15zdnd00an1n01x5 FILLER_165_1824 ();
 b15zdnd11an1n64x5 FILLER_165_1831 ();
 b15zdnd11an1n64x5 FILLER_165_1895 ();
 b15zdnd11an1n64x5 FILLER_165_1959 ();
 b15zdnd11an1n64x5 FILLER_165_2023 ();
 b15zdnd11an1n64x5 FILLER_165_2087 ();
 b15zdnd11an1n64x5 FILLER_165_2151 ();
 b15zdnd11an1n64x5 FILLER_165_2215 ();
 b15zdnd11an1n04x5 FILLER_165_2279 ();
 b15zdnd00an1n01x5 FILLER_165_2283 ();
 b15zdnd11an1n64x5 FILLER_166_8 ();
 b15zdnd11an1n64x5 FILLER_166_72 ();
 b15zdnd11an1n08x5 FILLER_166_136 ();
 b15zdnd11an1n04x5 FILLER_166_150 ();
 b15zdnd11an1n04x5 FILLER_166_163 ();
 b15zdnd11an1n64x5 FILLER_166_173 ();
 b15zdnd11an1n32x5 FILLER_166_237 ();
 b15zdnd11an1n16x5 FILLER_166_269 ();
 b15zdnd11an1n08x5 FILLER_166_285 ();
 b15zdnd11an1n04x5 FILLER_166_293 ();
 b15zdnd00an1n02x5 FILLER_166_297 ();
 b15zdnd00an1n01x5 FILLER_166_299 ();
 b15zdnd11an1n08x5 FILLER_166_342 ();
 b15zdnd11an1n04x5 FILLER_166_350 ();
 b15zdnd11an1n32x5 FILLER_166_396 ();
 b15zdnd11an1n08x5 FILLER_166_428 ();
 b15zdnd00an1n02x5 FILLER_166_436 ();
 b15zdnd11an1n32x5 FILLER_166_441 ();
 b15zdnd11an1n08x5 FILLER_166_473 ();
 b15zdnd11an1n04x5 FILLER_166_481 ();
 b15zdnd00an1n01x5 FILLER_166_485 ();
 b15zdnd11an1n04x5 FILLER_166_489 ();
 b15zdnd11an1n64x5 FILLER_166_496 ();
 b15zdnd11an1n32x5 FILLER_166_560 ();
 b15zdnd11an1n08x5 FILLER_166_592 ();
 b15zdnd00an1n02x5 FILLER_166_600 ();
 b15zdnd00an1n01x5 FILLER_166_602 ();
 b15zdnd11an1n16x5 FILLER_166_606 ();
 b15zdnd11an1n04x5 FILLER_166_622 ();
 b15zdnd00an1n02x5 FILLER_166_626 ();
 b15zdnd11an1n08x5 FILLER_166_648 ();
 b15zdnd11an1n04x5 FILLER_166_656 ();
 b15zdnd00an1n02x5 FILLER_166_660 ();
 b15zdnd00an1n01x5 FILLER_166_662 ();
 b15zdnd00an1n02x5 FILLER_166_715 ();
 b15zdnd00an1n01x5 FILLER_166_717 ();
 b15zdnd11an1n08x5 FILLER_166_726 ();
 b15zdnd00an1n01x5 FILLER_166_734 ();
 b15zdnd11an1n64x5 FILLER_166_743 ();
 b15zdnd11an1n04x5 FILLER_166_807 ();
 b15zdnd00an1n02x5 FILLER_166_811 ();
 b15zdnd11an1n04x5 FILLER_166_836 ();
 b15zdnd11an1n32x5 FILLER_166_854 ();
 b15zdnd11an1n04x5 FILLER_166_886 ();
 b15zdnd00an1n02x5 FILLER_166_890 ();
 b15zdnd00an1n01x5 FILLER_166_892 ();
 b15zdnd11an1n32x5 FILLER_166_902 ();
 b15zdnd11an1n16x5 FILLER_166_934 ();
 b15zdnd11an1n08x5 FILLER_166_950 ();
 b15zdnd11an1n04x5 FILLER_166_958 ();
 b15zdnd11an1n64x5 FILLER_166_1014 ();
 b15zdnd11an1n64x5 FILLER_166_1078 ();
 b15zdnd11an1n64x5 FILLER_166_1142 ();
 b15zdnd11an1n64x5 FILLER_166_1206 ();
 b15zdnd11an1n64x5 FILLER_166_1270 ();
 b15zdnd11an1n32x5 FILLER_166_1334 ();
 b15zdnd11an1n16x5 FILLER_166_1366 ();
 b15zdnd00an1n02x5 FILLER_166_1382 ();
 b15zdnd11an1n04x5 FILLER_166_1387 ();
 b15zdnd11an1n64x5 FILLER_166_1394 ();
 b15zdnd11an1n32x5 FILLER_166_1458 ();
 b15zdnd11an1n16x5 FILLER_166_1490 ();
 b15zdnd11an1n08x5 FILLER_166_1506 ();
 b15zdnd00an1n02x5 FILLER_166_1514 ();
 b15zdnd00an1n01x5 FILLER_166_1516 ();
 b15zdnd11an1n64x5 FILLER_166_1525 ();
 b15zdnd11an1n64x5 FILLER_166_1589 ();
 b15zdnd11an1n64x5 FILLER_166_1653 ();
 b15zdnd11an1n64x5 FILLER_166_1717 ();
 b15zdnd11an1n64x5 FILLER_166_1781 ();
 b15zdnd11an1n64x5 FILLER_166_1845 ();
 b15zdnd11an1n64x5 FILLER_166_1909 ();
 b15zdnd11an1n64x5 FILLER_166_1973 ();
 b15zdnd11an1n64x5 FILLER_166_2037 ();
 b15zdnd11an1n32x5 FILLER_166_2101 ();
 b15zdnd11an1n16x5 FILLER_166_2133 ();
 b15zdnd11an1n04x5 FILLER_166_2149 ();
 b15zdnd00an1n01x5 FILLER_166_2153 ();
 b15zdnd11an1n64x5 FILLER_166_2162 ();
 b15zdnd11an1n32x5 FILLER_166_2226 ();
 b15zdnd11an1n16x5 FILLER_166_2258 ();
 b15zdnd00an1n02x5 FILLER_166_2274 ();
 b15zdnd11an1n64x5 FILLER_167_0 ();
 b15zdnd11an1n64x5 FILLER_167_64 ();
 b15zdnd11an1n16x5 FILLER_167_128 ();
 b15zdnd11an1n08x5 FILLER_167_144 ();
 b15zdnd11an1n04x5 FILLER_167_152 ();
 b15zdnd11an1n08x5 FILLER_167_198 ();
 b15zdnd11an1n04x5 FILLER_167_206 ();
 b15zdnd11an1n16x5 FILLER_167_252 ();
 b15zdnd00an1n02x5 FILLER_167_268 ();
 b15zdnd11an1n04x5 FILLER_167_273 ();
 b15zdnd11an1n64x5 FILLER_167_280 ();
 b15zdnd11an1n64x5 FILLER_167_344 ();
 b15zdnd00an1n02x5 FILLER_167_408 ();
 b15zdnd00an1n01x5 FILLER_167_410 ();
 b15zdnd11an1n64x5 FILLER_167_463 ();
 b15zdnd11an1n32x5 FILLER_167_527 ();
 b15zdnd11an1n16x5 FILLER_167_559 ();
 b15zdnd11an1n08x5 FILLER_167_575 ();
 b15zdnd11an1n32x5 FILLER_167_635 ();
 b15zdnd11an1n04x5 FILLER_167_670 ();
 b15zdnd11an1n04x5 FILLER_167_677 ();
 b15zdnd11an1n32x5 FILLER_167_733 ();
 b15zdnd00an1n01x5 FILLER_167_765 ();
 b15zdnd11an1n64x5 FILLER_167_770 ();
 b15zdnd11an1n16x5 FILLER_167_834 ();
 b15zdnd00an1n02x5 FILLER_167_850 ();
 b15zdnd11an1n16x5 FILLER_167_876 ();
 b15zdnd00an1n01x5 FILLER_167_892 ();
 b15zdnd11an1n04x5 FILLER_167_902 ();
 b15zdnd11an1n64x5 FILLER_167_915 ();
 b15zdnd00an1n02x5 FILLER_167_979 ();
 b15zdnd00an1n01x5 FILLER_167_981 ();
 b15zdnd11an1n04x5 FILLER_167_985 ();
 b15zdnd11an1n04x5 FILLER_167_992 ();
 b15zdnd11an1n64x5 FILLER_167_999 ();
 b15zdnd11an1n64x5 FILLER_167_1063 ();
 b15zdnd11an1n08x5 FILLER_167_1127 ();
 b15zdnd00an1n02x5 FILLER_167_1135 ();
 b15zdnd00an1n01x5 FILLER_167_1137 ();
 b15zdnd11an1n64x5 FILLER_167_1141 ();
 b15zdnd11an1n64x5 FILLER_167_1205 ();
 b15zdnd11an1n04x5 FILLER_167_1269 ();
 b15zdnd00an1n01x5 FILLER_167_1273 ();
 b15zdnd11an1n32x5 FILLER_167_1279 ();
 b15zdnd11an1n16x5 FILLER_167_1311 ();
 b15zdnd11an1n08x5 FILLER_167_1327 ();
 b15zdnd11an1n16x5 FILLER_167_1339 ();
 b15zdnd11an1n08x5 FILLER_167_1355 ();
 b15zdnd00an1n02x5 FILLER_167_1363 ();
 b15zdnd00an1n01x5 FILLER_167_1365 ();
 b15zdnd11an1n64x5 FILLER_167_1418 ();
 b15zdnd11an1n32x5 FILLER_167_1482 ();
 b15zdnd11an1n16x5 FILLER_167_1514 ();
 b15zdnd11an1n04x5 FILLER_167_1530 ();
 b15zdnd11an1n04x5 FILLER_167_1537 ();
 b15zdnd11an1n04x5 FILLER_167_1544 ();
 b15zdnd11an1n64x5 FILLER_167_1551 ();
 b15zdnd11an1n64x5 FILLER_167_1615 ();
 b15zdnd11an1n32x5 FILLER_167_1679 ();
 b15zdnd11an1n16x5 FILLER_167_1711 ();
 b15zdnd11an1n08x5 FILLER_167_1727 ();
 b15zdnd11an1n04x5 FILLER_167_1735 ();
 b15zdnd00an1n02x5 FILLER_167_1739 ();
 b15zdnd00an1n01x5 FILLER_167_1741 ();
 b15zdnd11an1n64x5 FILLER_167_1759 ();
 b15zdnd11an1n32x5 FILLER_167_1823 ();
 b15zdnd11an1n16x5 FILLER_167_1855 ();
 b15zdnd11an1n04x5 FILLER_167_1871 ();
 b15zdnd00an1n01x5 FILLER_167_1875 ();
 b15zdnd11an1n64x5 FILLER_167_1890 ();
 b15zdnd11an1n64x5 FILLER_167_1954 ();
 b15zdnd11an1n64x5 FILLER_167_2018 ();
 b15zdnd11an1n64x5 FILLER_167_2082 ();
 b15zdnd11an1n16x5 FILLER_167_2146 ();
 b15zdnd11an1n08x5 FILLER_167_2162 ();
 b15zdnd11an1n04x5 FILLER_167_2170 ();
 b15zdnd00an1n02x5 FILLER_167_2174 ();
 b15zdnd11an1n64x5 FILLER_167_2190 ();
 b15zdnd11an1n16x5 FILLER_167_2254 ();
 b15zdnd11an1n08x5 FILLER_167_2270 ();
 b15zdnd11an1n04x5 FILLER_167_2278 ();
 b15zdnd00an1n02x5 FILLER_167_2282 ();
 b15zdnd11an1n64x5 FILLER_168_8 ();
 b15zdnd11an1n64x5 FILLER_168_72 ();
 b15zdnd11an1n64x5 FILLER_168_136 ();
 b15zdnd11an1n32x5 FILLER_168_200 ();
 b15zdnd11an1n16x5 FILLER_168_232 ();
 b15zdnd00an1n02x5 FILLER_168_248 ();
 b15zdnd11an1n64x5 FILLER_168_302 ();
 b15zdnd11an1n64x5 FILLER_168_366 ();
 b15zdnd11an1n04x5 FILLER_168_433 ();
 b15zdnd11an1n64x5 FILLER_168_440 ();
 b15zdnd11an1n32x5 FILLER_168_504 ();
 b15zdnd11an1n08x5 FILLER_168_536 ();
 b15zdnd11an1n04x5 FILLER_168_544 ();
 b15zdnd00an1n02x5 FILLER_168_548 ();
 b15zdnd11an1n32x5 FILLER_168_555 ();
 b15zdnd11an1n08x5 FILLER_168_587 ();
 b15zdnd11an1n04x5 FILLER_168_595 ();
 b15zdnd11an1n04x5 FILLER_168_602 ();
 b15zdnd11an1n32x5 FILLER_168_609 ();
 b15zdnd11an1n04x5 FILLER_168_641 ();
 b15zdnd00an1n02x5 FILLER_168_645 ();
 b15zdnd00an1n01x5 FILLER_168_647 ();
 b15zdnd11an1n04x5 FILLER_168_700 ();
 b15zdnd11an1n04x5 FILLER_168_707 ();
 b15zdnd11an1n04x5 FILLER_168_714 ();
 b15zdnd11an1n64x5 FILLER_168_726 ();
 b15zdnd11an1n64x5 FILLER_168_790 ();
 b15zdnd11an1n64x5 FILLER_168_854 ();
 b15zdnd11an1n64x5 FILLER_168_918 ();
 b15zdnd11an1n04x5 FILLER_168_982 ();
 b15zdnd00an1n01x5 FILLER_168_986 ();
 b15zdnd11an1n04x5 FILLER_168_990 ();
 b15zdnd11an1n64x5 FILLER_168_997 ();
 b15zdnd11an1n32x5 FILLER_168_1061 ();
 b15zdnd11an1n16x5 FILLER_168_1093 ();
 b15zdnd00an1n02x5 FILLER_168_1109 ();
 b15zdnd11an1n64x5 FILLER_168_1163 ();
 b15zdnd11an1n16x5 FILLER_168_1227 ();
 b15zdnd00an1n01x5 FILLER_168_1243 ();
 b15zdnd11an1n16x5 FILLER_168_1255 ();
 b15zdnd11an1n08x5 FILLER_168_1271 ();
 b15zdnd00an1n02x5 FILLER_168_1279 ();
 b15zdnd00an1n01x5 FILLER_168_1281 ();
 b15zdnd11an1n32x5 FILLER_168_1294 ();
 b15zdnd00an1n02x5 FILLER_168_1326 ();
 b15zdnd11an1n08x5 FILLER_168_1332 ();
 b15zdnd11an1n16x5 FILLER_168_1344 ();
 b15zdnd11an1n64x5 FILLER_168_1412 ();
 b15zdnd11an1n32x5 FILLER_168_1476 ();
 b15zdnd11an1n08x5 FILLER_168_1508 ();
 b15zdnd11an1n64x5 FILLER_168_1568 ();
 b15zdnd11an1n64x5 FILLER_168_1632 ();
 b15zdnd11an1n64x5 FILLER_168_1696 ();
 b15zdnd11an1n64x5 FILLER_168_1760 ();
 b15zdnd11an1n64x5 FILLER_168_1824 ();
 b15zdnd11an1n64x5 FILLER_168_1888 ();
 b15zdnd11an1n64x5 FILLER_168_1952 ();
 b15zdnd11an1n64x5 FILLER_168_2016 ();
 b15zdnd11an1n64x5 FILLER_168_2080 ();
 b15zdnd11an1n08x5 FILLER_168_2144 ();
 b15zdnd00an1n02x5 FILLER_168_2152 ();
 b15zdnd11an1n64x5 FILLER_168_2162 ();
 b15zdnd11an1n32x5 FILLER_168_2226 ();
 b15zdnd11an1n16x5 FILLER_168_2258 ();
 b15zdnd00an1n02x5 FILLER_168_2274 ();
 b15zdnd11an1n64x5 FILLER_169_0 ();
 b15zdnd11an1n64x5 FILLER_169_64 ();
 b15zdnd11an1n32x5 FILLER_169_128 ();
 b15zdnd11an1n04x5 FILLER_169_160 ();
 b15zdnd11an1n64x5 FILLER_169_206 ();
 b15zdnd00an1n01x5 FILLER_169_270 ();
 b15zdnd11an1n16x5 FILLER_169_274 ();
 b15zdnd11an1n04x5 FILLER_169_290 ();
 b15zdnd11an1n64x5 FILLER_169_302 ();
 b15zdnd11an1n64x5 FILLER_169_366 ();
 b15zdnd11an1n64x5 FILLER_169_430 ();
 b15zdnd11an1n64x5 FILLER_169_494 ();
 b15zdnd11an1n64x5 FILLER_169_558 ();
 b15zdnd11an1n08x5 FILLER_169_622 ();
 b15zdnd00an1n02x5 FILLER_169_630 ();
 b15zdnd11an1n16x5 FILLER_169_658 ();
 b15zdnd11an1n08x5 FILLER_169_677 ();
 b15zdnd11an1n04x5 FILLER_169_685 ();
 b15zdnd11an1n08x5 FILLER_169_692 ();
 b15zdnd11an1n04x5 FILLER_169_700 ();
 b15zdnd00an1n02x5 FILLER_169_704 ();
 b15zdnd00an1n01x5 FILLER_169_706 ();
 b15zdnd11an1n64x5 FILLER_169_710 ();
 b15zdnd11an1n32x5 FILLER_169_774 ();
 b15zdnd11an1n16x5 FILLER_169_806 ();
 b15zdnd11an1n08x5 FILLER_169_822 ();
 b15zdnd11an1n04x5 FILLER_169_830 ();
 b15zdnd11an1n64x5 FILLER_169_856 ();
 b15zdnd11an1n64x5 FILLER_169_920 ();
 b15zdnd11an1n64x5 FILLER_169_984 ();
 b15zdnd11an1n64x5 FILLER_169_1048 ();
 b15zdnd11an1n16x5 FILLER_169_1112 ();
 b15zdnd00an1n02x5 FILLER_169_1128 ();
 b15zdnd11an1n04x5 FILLER_169_1133 ();
 b15zdnd11an1n64x5 FILLER_169_1140 ();
 b15zdnd11an1n32x5 FILLER_169_1204 ();
 b15zdnd11an1n08x5 FILLER_169_1236 ();
 b15zdnd00an1n02x5 FILLER_169_1244 ();
 b15zdnd00an1n01x5 FILLER_169_1246 ();
 b15zdnd11an1n04x5 FILLER_169_1261 ();
 b15zdnd11an1n64x5 FILLER_169_1276 ();
 b15zdnd11an1n32x5 FILLER_169_1340 ();
 b15zdnd11an1n04x5 FILLER_169_1372 ();
 b15zdnd00an1n02x5 FILLER_169_1376 ();
 b15zdnd11an1n04x5 FILLER_169_1381 ();
 b15zdnd11an1n04x5 FILLER_169_1388 ();
 b15zdnd11an1n04x5 FILLER_169_1395 ();
 b15zdnd11an1n64x5 FILLER_169_1402 ();
 b15zdnd11an1n32x5 FILLER_169_1466 ();
 b15zdnd11an1n16x5 FILLER_169_1498 ();
 b15zdnd00an1n01x5 FILLER_169_1514 ();
 b15zdnd11an1n32x5 FILLER_169_1567 ();
 b15zdnd11an1n04x5 FILLER_169_1599 ();
 b15zdnd00an1n02x5 FILLER_169_1603 ();
 b15zdnd00an1n01x5 FILLER_169_1605 ();
 b15zdnd11an1n64x5 FILLER_169_1610 ();
 b15zdnd11an1n64x5 FILLER_169_1674 ();
 b15zdnd11an1n32x5 FILLER_169_1738 ();
 b15zdnd11an1n16x5 FILLER_169_1770 ();
 b15zdnd11an1n04x5 FILLER_169_1786 ();
 b15zdnd00an1n02x5 FILLER_169_1790 ();
 b15zdnd11an1n64x5 FILLER_169_1809 ();
 b15zdnd11an1n64x5 FILLER_169_1873 ();
 b15zdnd11an1n64x5 FILLER_169_1937 ();
 b15zdnd11an1n64x5 FILLER_169_2001 ();
 b15zdnd11an1n64x5 FILLER_169_2065 ();
 b15zdnd11an1n64x5 FILLER_169_2129 ();
 b15zdnd11an1n64x5 FILLER_169_2193 ();
 b15zdnd11an1n16x5 FILLER_169_2257 ();
 b15zdnd11an1n08x5 FILLER_169_2273 ();
 b15zdnd00an1n02x5 FILLER_169_2281 ();
 b15zdnd00an1n01x5 FILLER_169_2283 ();
 b15zdnd11an1n64x5 FILLER_170_8 ();
 b15zdnd11an1n64x5 FILLER_170_72 ();
 b15zdnd11an1n16x5 FILLER_170_136 ();
 b15zdnd11an1n08x5 FILLER_170_152 ();
 b15zdnd11an1n04x5 FILLER_170_160 ();
 b15zdnd00an1n02x5 FILLER_170_164 ();
 b15zdnd11an1n64x5 FILLER_170_208 ();
 b15zdnd11an1n04x5 FILLER_170_272 ();
 b15zdnd00an1n02x5 FILLER_170_276 ();
 b15zdnd11an1n64x5 FILLER_170_317 ();
 b15zdnd11an1n64x5 FILLER_170_381 ();
 b15zdnd11an1n64x5 FILLER_170_445 ();
 b15zdnd11an1n64x5 FILLER_170_509 ();
 b15zdnd11an1n64x5 FILLER_170_573 ();
 b15zdnd11an1n32x5 FILLER_170_664 ();
 b15zdnd11an1n16x5 FILLER_170_696 ();
 b15zdnd11an1n04x5 FILLER_170_712 ();
 b15zdnd00an1n02x5 FILLER_170_716 ();
 b15zdnd11an1n64x5 FILLER_170_726 ();
 b15zdnd11an1n16x5 FILLER_170_790 ();
 b15zdnd11an1n08x5 FILLER_170_806 ();
 b15zdnd11an1n04x5 FILLER_170_814 ();
 b15zdnd11an1n08x5 FILLER_170_830 ();
 b15zdnd11an1n04x5 FILLER_170_838 ();
 b15zdnd11an1n64x5 FILLER_170_873 ();
 b15zdnd11an1n64x5 FILLER_170_937 ();
 b15zdnd11an1n64x5 FILLER_170_1001 ();
 b15zdnd11an1n64x5 FILLER_170_1065 ();
 b15zdnd11an1n64x5 FILLER_170_1129 ();
 b15zdnd11an1n64x5 FILLER_170_1193 ();
 b15zdnd11an1n64x5 FILLER_170_1257 ();
 b15zdnd11an1n64x5 FILLER_170_1321 ();
 b15zdnd00an1n01x5 FILLER_170_1385 ();
 b15zdnd11an1n04x5 FILLER_170_1389 ();
 b15zdnd11an1n64x5 FILLER_170_1420 ();
 b15zdnd11an1n32x5 FILLER_170_1484 ();
 b15zdnd11an1n16x5 FILLER_170_1516 ();
 b15zdnd00an1n01x5 FILLER_170_1532 ();
 b15zdnd11an1n04x5 FILLER_170_1536 ();
 b15zdnd00an1n01x5 FILLER_170_1540 ();
 b15zdnd11an1n64x5 FILLER_170_1544 ();
 b15zdnd11an1n64x5 FILLER_170_1608 ();
 b15zdnd11an1n08x5 FILLER_170_1672 ();
 b15zdnd11an1n04x5 FILLER_170_1680 ();
 b15zdnd00an1n01x5 FILLER_170_1684 ();
 b15zdnd11an1n64x5 FILLER_170_1690 ();
 b15zdnd11an1n64x5 FILLER_170_1754 ();
 b15zdnd11an1n64x5 FILLER_170_1818 ();
 b15zdnd11an1n64x5 FILLER_170_1882 ();
 b15zdnd11an1n64x5 FILLER_170_1946 ();
 b15zdnd11an1n32x5 FILLER_170_2010 ();
 b15zdnd11an1n08x5 FILLER_170_2042 ();
 b15zdnd11an1n04x5 FILLER_170_2050 ();
 b15zdnd11an1n32x5 FILLER_170_2096 ();
 b15zdnd11an1n16x5 FILLER_170_2128 ();
 b15zdnd11an1n08x5 FILLER_170_2144 ();
 b15zdnd00an1n02x5 FILLER_170_2152 ();
 b15zdnd11an1n64x5 FILLER_170_2162 ();
 b15zdnd11an1n32x5 FILLER_170_2226 ();
 b15zdnd11an1n16x5 FILLER_170_2258 ();
 b15zdnd00an1n02x5 FILLER_170_2274 ();
 b15zdnd11an1n64x5 FILLER_171_0 ();
 b15zdnd11an1n64x5 FILLER_171_64 ();
 b15zdnd11an1n64x5 FILLER_171_128 ();
 b15zdnd11an1n64x5 FILLER_171_192 ();
 b15zdnd11an1n16x5 FILLER_171_256 ();
 b15zdnd11an1n08x5 FILLER_171_272 ();
 b15zdnd00an1n01x5 FILLER_171_280 ();
 b15zdnd11an1n64x5 FILLER_171_285 ();
 b15zdnd11an1n64x5 FILLER_171_349 ();
 b15zdnd11an1n64x5 FILLER_171_413 ();
 b15zdnd11an1n64x5 FILLER_171_477 ();
 b15zdnd11an1n64x5 FILLER_171_541 ();
 b15zdnd11an1n32x5 FILLER_171_605 ();
 b15zdnd00an1n02x5 FILLER_171_637 ();
 b15zdnd11an1n64x5 FILLER_171_642 ();
 b15zdnd11an1n64x5 FILLER_171_706 ();
 b15zdnd11an1n64x5 FILLER_171_770 ();
 b15zdnd11an1n64x5 FILLER_171_834 ();
 b15zdnd11an1n64x5 FILLER_171_898 ();
 b15zdnd11an1n64x5 FILLER_171_962 ();
 b15zdnd11an1n64x5 FILLER_171_1026 ();
 b15zdnd11an1n64x5 FILLER_171_1090 ();
 b15zdnd11an1n64x5 FILLER_171_1154 ();
 b15zdnd11an1n64x5 FILLER_171_1218 ();
 b15zdnd11an1n64x5 FILLER_171_1282 ();
 b15zdnd11an1n64x5 FILLER_171_1346 ();
 b15zdnd11an1n64x5 FILLER_171_1410 ();
 b15zdnd11an1n64x5 FILLER_171_1474 ();
 b15zdnd00an1n01x5 FILLER_171_1538 ();
 b15zdnd11an1n64x5 FILLER_171_1542 ();
 b15zdnd11an1n64x5 FILLER_171_1606 ();
 b15zdnd11an1n64x5 FILLER_171_1670 ();
 b15zdnd11an1n64x5 FILLER_171_1734 ();
 b15zdnd11an1n64x5 FILLER_171_1798 ();
 b15zdnd11an1n64x5 FILLER_171_1862 ();
 b15zdnd11an1n64x5 FILLER_171_1926 ();
 b15zdnd11an1n64x5 FILLER_171_1990 ();
 b15zdnd11an1n64x5 FILLER_171_2054 ();
 b15zdnd11an1n64x5 FILLER_171_2118 ();
 b15zdnd11an1n04x5 FILLER_171_2182 ();
 b15zdnd00an1n02x5 FILLER_171_2186 ();
 b15zdnd00an1n01x5 FILLER_171_2188 ();
 b15zdnd11an1n64x5 FILLER_171_2201 ();
 b15zdnd11an1n16x5 FILLER_171_2265 ();
 b15zdnd00an1n02x5 FILLER_171_2281 ();
 b15zdnd00an1n01x5 FILLER_171_2283 ();
 b15zdnd11an1n64x5 FILLER_172_8 ();
 b15zdnd11an1n64x5 FILLER_172_72 ();
 b15zdnd11an1n64x5 FILLER_172_136 ();
 b15zdnd11an1n64x5 FILLER_172_200 ();
 b15zdnd11an1n16x5 FILLER_172_264 ();
 b15zdnd11an1n04x5 FILLER_172_280 ();
 b15zdnd11an1n64x5 FILLER_172_326 ();
 b15zdnd11an1n64x5 FILLER_172_390 ();
 b15zdnd11an1n64x5 FILLER_172_454 ();
 b15zdnd11an1n64x5 FILLER_172_518 ();
 b15zdnd11an1n64x5 FILLER_172_582 ();
 b15zdnd11an1n64x5 FILLER_172_646 ();
 b15zdnd11an1n08x5 FILLER_172_710 ();
 b15zdnd11an1n32x5 FILLER_172_726 ();
 b15zdnd11an1n16x5 FILLER_172_758 ();
 b15zdnd11an1n08x5 FILLER_172_774 ();
 b15zdnd00an1n02x5 FILLER_172_782 ();
 b15zdnd11an1n16x5 FILLER_172_792 ();
 b15zdnd11an1n04x5 FILLER_172_808 ();
 b15zdnd00an1n01x5 FILLER_172_812 ();
 b15zdnd11an1n32x5 FILLER_172_824 ();
 b15zdnd11an1n08x5 FILLER_172_856 ();
 b15zdnd11an1n64x5 FILLER_172_875 ();
 b15zdnd11an1n64x5 FILLER_172_939 ();
 b15zdnd11an1n64x5 FILLER_172_1003 ();
 b15zdnd11an1n64x5 FILLER_172_1067 ();
 b15zdnd11an1n64x5 FILLER_172_1131 ();
 b15zdnd11an1n64x5 FILLER_172_1195 ();
 b15zdnd11an1n64x5 FILLER_172_1259 ();
 b15zdnd11an1n64x5 FILLER_172_1323 ();
 b15zdnd11an1n64x5 FILLER_172_1387 ();
 b15zdnd11an1n64x5 FILLER_172_1451 ();
 b15zdnd11an1n64x5 FILLER_172_1515 ();
 b15zdnd11an1n64x5 FILLER_172_1579 ();
 b15zdnd11an1n64x5 FILLER_172_1643 ();
 b15zdnd11an1n64x5 FILLER_172_1707 ();
 b15zdnd11an1n32x5 FILLER_172_1771 ();
 b15zdnd11an1n08x5 FILLER_172_1803 ();
 b15zdnd11an1n64x5 FILLER_172_1819 ();
 b15zdnd11an1n64x5 FILLER_172_1883 ();
 b15zdnd11an1n64x5 FILLER_172_1947 ();
 b15zdnd11an1n64x5 FILLER_172_2011 ();
 b15zdnd11an1n64x5 FILLER_172_2075 ();
 b15zdnd11an1n08x5 FILLER_172_2139 ();
 b15zdnd11an1n04x5 FILLER_172_2147 ();
 b15zdnd00an1n02x5 FILLER_172_2151 ();
 b15zdnd00an1n01x5 FILLER_172_2153 ();
 b15zdnd11an1n64x5 FILLER_172_2162 ();
 b15zdnd11an1n32x5 FILLER_172_2226 ();
 b15zdnd11an1n16x5 FILLER_172_2258 ();
 b15zdnd00an1n02x5 FILLER_172_2274 ();
 b15zdnd11an1n64x5 FILLER_173_0 ();
 b15zdnd11an1n64x5 FILLER_173_64 ();
 b15zdnd11an1n08x5 FILLER_173_128 ();
 b15zdnd11an1n64x5 FILLER_173_188 ();
 b15zdnd11an1n32x5 FILLER_173_252 ();
 b15zdnd11an1n16x5 FILLER_173_284 ();
 b15zdnd11an1n04x5 FILLER_173_300 ();
 b15zdnd00an1n02x5 FILLER_173_304 ();
 b15zdnd11an1n08x5 FILLER_173_309 ();
 b15zdnd00an1n01x5 FILLER_173_317 ();
 b15zdnd11an1n64x5 FILLER_173_360 ();
 b15zdnd11an1n04x5 FILLER_173_424 ();
 b15zdnd00an1n01x5 FILLER_173_428 ();
 b15zdnd11an1n64x5 FILLER_173_444 ();
 b15zdnd11an1n08x5 FILLER_173_528 ();
 b15zdnd11an1n04x5 FILLER_173_536 ();
 b15zdnd00an1n02x5 FILLER_173_540 ();
 b15zdnd00an1n01x5 FILLER_173_542 ();
 b15zdnd11an1n64x5 FILLER_173_563 ();
 b15zdnd11an1n16x5 FILLER_173_627 ();
 b15zdnd11an1n08x5 FILLER_173_643 ();
 b15zdnd11an1n04x5 FILLER_173_651 ();
 b15zdnd11an1n64x5 FILLER_173_664 ();
 b15zdnd11an1n64x5 FILLER_173_728 ();
 b15zdnd11an1n08x5 FILLER_173_792 ();
 b15zdnd00an1n01x5 FILLER_173_800 ();
 b15zdnd11an1n64x5 FILLER_173_817 ();
 b15zdnd11an1n64x5 FILLER_173_881 ();
 b15zdnd11an1n64x5 FILLER_173_945 ();
 b15zdnd11an1n64x5 FILLER_173_1009 ();
 b15zdnd11an1n64x5 FILLER_173_1073 ();
 b15zdnd11an1n64x5 FILLER_173_1137 ();
 b15zdnd11an1n04x5 FILLER_173_1201 ();
 b15zdnd00an1n02x5 FILLER_173_1205 ();
 b15zdnd11an1n64x5 FILLER_173_1216 ();
 b15zdnd11an1n64x5 FILLER_173_1280 ();
 b15zdnd11an1n64x5 FILLER_173_1344 ();
 b15zdnd11an1n64x5 FILLER_173_1408 ();
 b15zdnd11an1n64x5 FILLER_173_1472 ();
 b15zdnd11an1n16x5 FILLER_173_1536 ();
 b15zdnd11an1n04x5 FILLER_173_1552 ();
 b15zdnd00an1n01x5 FILLER_173_1556 ();
 b15zdnd11an1n64x5 FILLER_173_1565 ();
 b15zdnd11an1n08x5 FILLER_173_1629 ();
 b15zdnd11an1n64x5 FILLER_173_1651 ();
 b15zdnd11an1n64x5 FILLER_173_1715 ();
 b15zdnd11an1n08x5 FILLER_173_1779 ();
 b15zdnd00an1n02x5 FILLER_173_1787 ();
 b15zdnd00an1n01x5 FILLER_173_1789 ();
 b15zdnd11an1n64x5 FILLER_173_1810 ();
 b15zdnd11an1n64x5 FILLER_173_1874 ();
 b15zdnd11an1n64x5 FILLER_173_1938 ();
 b15zdnd11an1n64x5 FILLER_173_2002 ();
 b15zdnd11an1n64x5 FILLER_173_2066 ();
 b15zdnd11an1n64x5 FILLER_173_2130 ();
 b15zdnd11an1n16x5 FILLER_173_2194 ();
 b15zdnd11an1n04x5 FILLER_173_2210 ();
 b15zdnd11an1n32x5 FILLER_173_2236 ();
 b15zdnd11an1n16x5 FILLER_173_2268 ();
 b15zdnd11an1n64x5 FILLER_174_8 ();
 b15zdnd11an1n64x5 FILLER_174_72 ();
 b15zdnd11an1n16x5 FILLER_174_136 ();
 b15zdnd11an1n04x5 FILLER_174_152 ();
 b15zdnd00an1n02x5 FILLER_174_156 ();
 b15zdnd00an1n01x5 FILLER_174_158 ();
 b15zdnd11an1n04x5 FILLER_174_162 ();
 b15zdnd11an1n64x5 FILLER_174_169 ();
 b15zdnd11an1n32x5 FILLER_174_233 ();
 b15zdnd11an1n04x5 FILLER_174_265 ();
 b15zdnd00an1n01x5 FILLER_174_269 ();
 b15zdnd11an1n64x5 FILLER_174_310 ();
 b15zdnd11an1n64x5 FILLER_174_374 ();
 b15zdnd11an1n64x5 FILLER_174_438 ();
 b15zdnd11an1n16x5 FILLER_174_502 ();
 b15zdnd00an1n01x5 FILLER_174_518 ();
 b15zdnd11an1n64x5 FILLER_174_535 ();
 b15zdnd11an1n64x5 FILLER_174_599 ();
 b15zdnd11an1n32x5 FILLER_174_663 ();
 b15zdnd11an1n16x5 FILLER_174_695 ();
 b15zdnd11an1n04x5 FILLER_174_711 ();
 b15zdnd00an1n02x5 FILLER_174_715 ();
 b15zdnd00an1n01x5 FILLER_174_717 ();
 b15zdnd11an1n64x5 FILLER_174_726 ();
 b15zdnd11an1n08x5 FILLER_174_790 ();
 b15zdnd00an1n02x5 FILLER_174_798 ();
 b15zdnd00an1n01x5 FILLER_174_800 ();
 b15zdnd11an1n04x5 FILLER_174_808 ();
 b15zdnd11an1n64x5 FILLER_174_818 ();
 b15zdnd11an1n16x5 FILLER_174_882 ();
 b15zdnd11an1n08x5 FILLER_174_898 ();
 b15zdnd11an1n04x5 FILLER_174_906 ();
 b15zdnd00an1n02x5 FILLER_174_910 ();
 b15zdnd11an1n64x5 FILLER_174_918 ();
 b15zdnd11an1n64x5 FILLER_174_982 ();
 b15zdnd11an1n64x5 FILLER_174_1046 ();
 b15zdnd11an1n64x5 FILLER_174_1110 ();
 b15zdnd11an1n64x5 FILLER_174_1174 ();
 b15zdnd11an1n16x5 FILLER_174_1238 ();
 b15zdnd11an1n04x5 FILLER_174_1254 ();
 b15zdnd00an1n02x5 FILLER_174_1258 ();
 b15zdnd00an1n01x5 FILLER_174_1260 ();
 b15zdnd11an1n32x5 FILLER_174_1264 ();
 b15zdnd11an1n08x5 FILLER_174_1296 ();
 b15zdnd11an1n04x5 FILLER_174_1304 ();
 b15zdnd11an1n64x5 FILLER_174_1328 ();
 b15zdnd11an1n64x5 FILLER_174_1392 ();
 b15zdnd11an1n64x5 FILLER_174_1456 ();
 b15zdnd11an1n16x5 FILLER_174_1520 ();
 b15zdnd11an1n08x5 FILLER_174_1536 ();
 b15zdnd00an1n02x5 FILLER_174_1544 ();
 b15zdnd00an1n01x5 FILLER_174_1546 ();
 b15zdnd11an1n32x5 FILLER_174_1571 ();
 b15zdnd11an1n08x5 FILLER_174_1607 ();
 b15zdnd00an1n02x5 FILLER_174_1615 ();
 b15zdnd00an1n01x5 FILLER_174_1617 ();
 b15zdnd11an1n64x5 FILLER_174_1635 ();
 b15zdnd11an1n64x5 FILLER_174_1699 ();
 b15zdnd11an1n08x5 FILLER_174_1763 ();
 b15zdnd11an1n04x5 FILLER_174_1771 ();
 b15zdnd00an1n02x5 FILLER_174_1775 ();
 b15zdnd11an1n04x5 FILLER_174_1799 ();
 b15zdnd11an1n64x5 FILLER_174_1811 ();
 b15zdnd11an1n16x5 FILLER_174_1875 ();
 b15zdnd11an1n04x5 FILLER_174_1891 ();
 b15zdnd11an1n16x5 FILLER_174_1912 ();
 b15zdnd11an1n04x5 FILLER_174_1928 ();
 b15zdnd00an1n02x5 FILLER_174_1932 ();
 b15zdnd00an1n01x5 FILLER_174_1934 ();
 b15zdnd11an1n64x5 FILLER_174_1938 ();
 b15zdnd11an1n64x5 FILLER_174_2002 ();
 b15zdnd11an1n08x5 FILLER_174_2066 ();
 b15zdnd11an1n04x5 FILLER_174_2074 ();
 b15zdnd11an1n16x5 FILLER_174_2084 ();
 b15zdnd11an1n08x5 FILLER_174_2100 ();
 b15zdnd00an1n01x5 FILLER_174_2108 ();
 b15zdnd11an1n32x5 FILLER_174_2117 ();
 b15zdnd11an1n04x5 FILLER_174_2149 ();
 b15zdnd00an1n01x5 FILLER_174_2153 ();
 b15zdnd11an1n64x5 FILLER_174_2162 ();
 b15zdnd11an1n32x5 FILLER_174_2226 ();
 b15zdnd11an1n16x5 FILLER_174_2258 ();
 b15zdnd00an1n02x5 FILLER_174_2274 ();
 b15zdnd11an1n64x5 FILLER_175_0 ();
 b15zdnd11an1n64x5 FILLER_175_64 ();
 b15zdnd11an1n16x5 FILLER_175_128 ();
 b15zdnd11an1n08x5 FILLER_175_144 ();
 b15zdnd11an1n04x5 FILLER_175_152 ();
 b15zdnd00an1n02x5 FILLER_175_156 ();
 b15zdnd00an1n01x5 FILLER_175_158 ();
 b15zdnd11an1n64x5 FILLER_175_162 ();
 b15zdnd11an1n64x5 FILLER_175_226 ();
 b15zdnd11an1n16x5 FILLER_175_290 ();
 b15zdnd00an1n02x5 FILLER_175_306 ();
 b15zdnd11an1n64x5 FILLER_175_311 ();
 b15zdnd11an1n08x5 FILLER_175_375 ();
 b15zdnd00an1n02x5 FILLER_175_383 ();
 b15zdnd11an1n32x5 FILLER_175_388 ();
 b15zdnd00an1n02x5 FILLER_175_420 ();
 b15zdnd11an1n64x5 FILLER_175_438 ();
 b15zdnd11an1n64x5 FILLER_175_502 ();
 b15zdnd11an1n64x5 FILLER_175_566 ();
 b15zdnd11an1n64x5 FILLER_175_630 ();
 b15zdnd11an1n64x5 FILLER_175_694 ();
 b15zdnd11an1n64x5 FILLER_175_758 ();
 b15zdnd11an1n04x5 FILLER_175_822 ();
 b15zdnd00an1n02x5 FILLER_175_826 ();
 b15zdnd00an1n01x5 FILLER_175_828 ();
 b15zdnd11an1n64x5 FILLER_175_836 ();
 b15zdnd11an1n64x5 FILLER_175_900 ();
 b15zdnd11an1n64x5 FILLER_175_964 ();
 b15zdnd11an1n64x5 FILLER_175_1028 ();
 b15zdnd11an1n64x5 FILLER_175_1092 ();
 b15zdnd11an1n64x5 FILLER_175_1156 ();
 b15zdnd11an1n08x5 FILLER_175_1220 ();
 b15zdnd11an1n04x5 FILLER_175_1228 ();
 b15zdnd00an1n02x5 FILLER_175_1232 ();
 b15zdnd00an1n01x5 FILLER_175_1234 ();
 b15zdnd11an1n64x5 FILLER_175_1287 ();
 b15zdnd11an1n64x5 FILLER_175_1351 ();
 b15zdnd11an1n64x5 FILLER_175_1415 ();
 b15zdnd11an1n64x5 FILLER_175_1479 ();
 b15zdnd11an1n32x5 FILLER_175_1543 ();
 b15zdnd11an1n16x5 FILLER_175_1575 ();
 b15zdnd11an1n04x5 FILLER_175_1591 ();
 b15zdnd00an1n01x5 FILLER_175_1595 ();
 b15zdnd11an1n32x5 FILLER_175_1604 ();
 b15zdnd11an1n08x5 FILLER_175_1636 ();
 b15zdnd00an1n02x5 FILLER_175_1644 ();
 b15zdnd11an1n64x5 FILLER_175_1656 ();
 b15zdnd11an1n08x5 FILLER_175_1720 ();
 b15zdnd11an1n04x5 FILLER_175_1728 ();
 b15zdnd00an1n01x5 FILLER_175_1732 ();
 b15zdnd11an1n64x5 FILLER_175_1747 ();
 b15zdnd11an1n64x5 FILLER_175_1811 ();
 b15zdnd11an1n32x5 FILLER_175_1875 ();
 b15zdnd11an1n16x5 FILLER_175_1907 ();
 b15zdnd11an1n04x5 FILLER_175_1923 ();
 b15zdnd00an1n01x5 FILLER_175_1927 ();
 b15zdnd11an1n64x5 FILLER_175_1948 ();
 b15zdnd11an1n64x5 FILLER_175_2012 ();
 b15zdnd11an1n64x5 FILLER_175_2076 ();
 b15zdnd11an1n64x5 FILLER_175_2140 ();
 b15zdnd11an1n64x5 FILLER_175_2204 ();
 b15zdnd11an1n16x5 FILLER_175_2268 ();
 b15zdnd11an1n16x5 FILLER_176_8 ();
 b15zdnd11an1n04x5 FILLER_176_24 ();
 b15zdnd11an1n64x5 FILLER_176_42 ();
 b15zdnd11an1n64x5 FILLER_176_106 ();
 b15zdnd11an1n64x5 FILLER_176_170 ();
 b15zdnd11an1n64x5 FILLER_176_234 ();
 b15zdnd11an1n64x5 FILLER_176_298 ();
 b15zdnd11an1n16x5 FILLER_176_362 ();
 b15zdnd11an1n04x5 FILLER_176_378 ();
 b15zdnd11an1n04x5 FILLER_176_385 ();
 b15zdnd00an1n02x5 FILLER_176_389 ();
 b15zdnd00an1n01x5 FILLER_176_391 ();
 b15zdnd11an1n64x5 FILLER_176_395 ();
 b15zdnd11an1n64x5 FILLER_176_459 ();
 b15zdnd11an1n64x5 FILLER_176_523 ();
 b15zdnd11an1n64x5 FILLER_176_587 ();
 b15zdnd11an1n64x5 FILLER_176_651 ();
 b15zdnd00an1n02x5 FILLER_176_715 ();
 b15zdnd00an1n01x5 FILLER_176_717 ();
 b15zdnd11an1n32x5 FILLER_176_726 ();
 b15zdnd11an1n16x5 FILLER_176_758 ();
 b15zdnd11an1n64x5 FILLER_176_780 ();
 b15zdnd11an1n32x5 FILLER_176_844 ();
 b15zdnd11an1n04x5 FILLER_176_876 ();
 b15zdnd00an1n01x5 FILLER_176_880 ();
 b15zdnd11an1n64x5 FILLER_176_886 ();
 b15zdnd11an1n64x5 FILLER_176_950 ();
 b15zdnd11an1n64x5 FILLER_176_1014 ();
 b15zdnd11an1n64x5 FILLER_176_1078 ();
 b15zdnd11an1n64x5 FILLER_176_1142 ();
 b15zdnd11an1n32x5 FILLER_176_1206 ();
 b15zdnd11an1n08x5 FILLER_176_1238 ();
 b15zdnd11an1n04x5 FILLER_176_1246 ();
 b15zdnd00an1n02x5 FILLER_176_1250 ();
 b15zdnd00an1n01x5 FILLER_176_1252 ();
 b15zdnd11an1n04x5 FILLER_176_1256 ();
 b15zdnd11an1n64x5 FILLER_176_1263 ();
 b15zdnd11an1n64x5 FILLER_176_1327 ();
 b15zdnd11an1n64x5 FILLER_176_1391 ();
 b15zdnd11an1n64x5 FILLER_176_1455 ();
 b15zdnd11an1n64x5 FILLER_176_1519 ();
 b15zdnd11an1n64x5 FILLER_176_1583 ();
 b15zdnd11an1n64x5 FILLER_176_1647 ();
 b15zdnd11an1n64x5 FILLER_176_1711 ();
 b15zdnd11an1n04x5 FILLER_176_1775 ();
 b15zdnd00an1n01x5 FILLER_176_1779 ();
 b15zdnd11an1n64x5 FILLER_176_1800 ();
 b15zdnd11an1n64x5 FILLER_176_1864 ();
 b15zdnd11an1n16x5 FILLER_176_1928 ();
 b15zdnd11an1n64x5 FILLER_176_1947 ();
 b15zdnd11an1n64x5 FILLER_176_2011 ();
 b15zdnd00an1n02x5 FILLER_176_2075 ();
 b15zdnd11an1n64x5 FILLER_176_2085 ();
 b15zdnd11an1n04x5 FILLER_176_2149 ();
 b15zdnd00an1n01x5 FILLER_176_2153 ();
 b15zdnd11an1n64x5 FILLER_176_2162 ();
 b15zdnd11an1n32x5 FILLER_176_2226 ();
 b15zdnd11an1n16x5 FILLER_176_2258 ();
 b15zdnd00an1n02x5 FILLER_176_2274 ();
 b15zdnd11an1n16x5 FILLER_177_0 ();
 b15zdnd11an1n08x5 FILLER_177_16 ();
 b15zdnd11an1n04x5 FILLER_177_24 ();
 b15zdnd00an1n01x5 FILLER_177_28 ();
 b15zdnd11an1n64x5 FILLER_177_40 ();
 b15zdnd11an1n64x5 FILLER_177_104 ();
 b15zdnd11an1n64x5 FILLER_177_168 ();
 b15zdnd11an1n64x5 FILLER_177_232 ();
 b15zdnd11an1n08x5 FILLER_177_296 ();
 b15zdnd00an1n02x5 FILLER_177_304 ();
 b15zdnd11an1n32x5 FILLER_177_318 ();
 b15zdnd00an1n02x5 FILLER_177_350 ();
 b15zdnd00an1n01x5 FILLER_177_352 ();
 b15zdnd11an1n64x5 FILLER_177_405 ();
 b15zdnd11an1n64x5 FILLER_177_469 ();
 b15zdnd11an1n64x5 FILLER_177_533 ();
 b15zdnd11an1n64x5 FILLER_177_597 ();
 b15zdnd11an1n64x5 FILLER_177_661 ();
 b15zdnd11an1n64x5 FILLER_177_725 ();
 b15zdnd11an1n64x5 FILLER_177_789 ();
 b15zdnd11an1n64x5 FILLER_177_853 ();
 b15zdnd11an1n64x5 FILLER_177_917 ();
 b15zdnd11an1n64x5 FILLER_177_981 ();
 b15zdnd11an1n64x5 FILLER_177_1045 ();
 b15zdnd11an1n64x5 FILLER_177_1109 ();
 b15zdnd11an1n64x5 FILLER_177_1173 ();
 b15zdnd11an1n64x5 FILLER_177_1237 ();
 b15zdnd11an1n64x5 FILLER_177_1301 ();
 b15zdnd11an1n64x5 FILLER_177_1365 ();
 b15zdnd11an1n64x5 FILLER_177_1429 ();
 b15zdnd11an1n64x5 FILLER_177_1493 ();
 b15zdnd11an1n64x5 FILLER_177_1557 ();
 b15zdnd11an1n64x5 FILLER_177_1621 ();
 b15zdnd11an1n64x5 FILLER_177_1685 ();
 b15zdnd11an1n64x5 FILLER_177_1749 ();
 b15zdnd11an1n64x5 FILLER_177_1813 ();
 b15zdnd11an1n32x5 FILLER_177_1877 ();
 b15zdnd00an1n02x5 FILLER_177_1909 ();
 b15zdnd11an1n04x5 FILLER_177_1963 ();
 b15zdnd11an1n64x5 FILLER_177_1970 ();
 b15zdnd11an1n32x5 FILLER_177_2034 ();
 b15zdnd11an1n08x5 FILLER_177_2066 ();
 b15zdnd00an1n02x5 FILLER_177_2074 ();
 b15zdnd11an1n64x5 FILLER_177_2086 ();
 b15zdnd11an1n32x5 FILLER_177_2150 ();
 b15zdnd00an1n02x5 FILLER_177_2182 ();
 b15zdnd11an1n04x5 FILLER_177_2195 ();
 b15zdnd11an1n64x5 FILLER_177_2206 ();
 b15zdnd11an1n08x5 FILLER_177_2270 ();
 b15zdnd11an1n04x5 FILLER_177_2278 ();
 b15zdnd00an1n02x5 FILLER_177_2282 ();
 b15zdnd11an1n64x5 FILLER_178_8 ();
 b15zdnd11an1n64x5 FILLER_178_72 ();
 b15zdnd11an1n64x5 FILLER_178_136 ();
 b15zdnd11an1n64x5 FILLER_178_200 ();
 b15zdnd11an1n64x5 FILLER_178_264 ();
 b15zdnd11an1n64x5 FILLER_178_328 ();
 b15zdnd11an1n64x5 FILLER_178_392 ();
 b15zdnd11an1n64x5 FILLER_178_456 ();
 b15zdnd11an1n64x5 FILLER_178_520 ();
 b15zdnd11an1n64x5 FILLER_178_584 ();
 b15zdnd11an1n16x5 FILLER_178_648 ();
 b15zdnd11an1n32x5 FILLER_178_673 ();
 b15zdnd11an1n08x5 FILLER_178_705 ();
 b15zdnd11an1n04x5 FILLER_178_713 ();
 b15zdnd00an1n01x5 FILLER_178_717 ();
 b15zdnd11an1n64x5 FILLER_178_726 ();
 b15zdnd11an1n64x5 FILLER_178_790 ();
 b15zdnd11an1n64x5 FILLER_178_854 ();
 b15zdnd11an1n64x5 FILLER_178_918 ();
 b15zdnd11an1n64x5 FILLER_178_982 ();
 b15zdnd11an1n64x5 FILLER_178_1046 ();
 b15zdnd11an1n64x5 FILLER_178_1110 ();
 b15zdnd11an1n64x5 FILLER_178_1174 ();
 b15zdnd11an1n64x5 FILLER_178_1238 ();
 b15zdnd11an1n64x5 FILLER_178_1302 ();
 b15zdnd11an1n64x5 FILLER_178_1366 ();
 b15zdnd00an1n02x5 FILLER_178_1430 ();
 b15zdnd11an1n32x5 FILLER_178_1441 ();
 b15zdnd11an1n08x5 FILLER_178_1473 ();
 b15zdnd11an1n04x5 FILLER_178_1481 ();
 b15zdnd00an1n02x5 FILLER_178_1485 ();
 b15zdnd00an1n01x5 FILLER_178_1487 ();
 b15zdnd11an1n64x5 FILLER_178_1497 ();
 b15zdnd11an1n64x5 FILLER_178_1561 ();
 b15zdnd11an1n64x5 FILLER_178_1625 ();
 b15zdnd11an1n04x5 FILLER_178_1689 ();
 b15zdnd00an1n01x5 FILLER_178_1693 ();
 b15zdnd11an1n64x5 FILLER_178_1697 ();
 b15zdnd11an1n64x5 FILLER_178_1761 ();
 b15zdnd11an1n64x5 FILLER_178_1825 ();
 b15zdnd11an1n64x5 FILLER_178_1889 ();
 b15zdnd11an1n64x5 FILLER_178_1953 ();
 b15zdnd11an1n32x5 FILLER_178_2017 ();
 b15zdnd11an1n16x5 FILLER_178_2049 ();
 b15zdnd11an1n04x5 FILLER_178_2065 ();
 b15zdnd11an1n64x5 FILLER_178_2089 ();
 b15zdnd00an1n01x5 FILLER_178_2153 ();
 b15zdnd11an1n64x5 FILLER_178_2162 ();
 b15zdnd11an1n32x5 FILLER_178_2226 ();
 b15zdnd11an1n16x5 FILLER_178_2258 ();
 b15zdnd00an1n02x5 FILLER_178_2274 ();
 b15zdnd11an1n64x5 FILLER_179_0 ();
 b15zdnd11an1n64x5 FILLER_179_64 ();
 b15zdnd11an1n64x5 FILLER_179_128 ();
 b15zdnd11an1n64x5 FILLER_179_192 ();
 b15zdnd11an1n64x5 FILLER_179_256 ();
 b15zdnd11an1n64x5 FILLER_179_320 ();
 b15zdnd11an1n64x5 FILLER_179_384 ();
 b15zdnd11an1n32x5 FILLER_179_448 ();
 b15zdnd11an1n16x5 FILLER_179_480 ();
 b15zdnd11an1n04x5 FILLER_179_496 ();
 b15zdnd00an1n02x5 FILLER_179_500 ();
 b15zdnd00an1n01x5 FILLER_179_502 ();
 b15zdnd11an1n64x5 FILLER_179_510 ();
 b15zdnd11an1n64x5 FILLER_179_574 ();
 b15zdnd11an1n64x5 FILLER_179_638 ();
 b15zdnd11an1n64x5 FILLER_179_702 ();
 b15zdnd11an1n64x5 FILLER_179_766 ();
 b15zdnd11an1n64x5 FILLER_179_830 ();
 b15zdnd11an1n64x5 FILLER_179_894 ();
 b15zdnd11an1n64x5 FILLER_179_958 ();
 b15zdnd11an1n64x5 FILLER_179_1022 ();
 b15zdnd11an1n32x5 FILLER_179_1086 ();
 b15zdnd00an1n02x5 FILLER_179_1118 ();
 b15zdnd00an1n01x5 FILLER_179_1120 ();
 b15zdnd11an1n64x5 FILLER_179_1130 ();
 b15zdnd11an1n64x5 FILLER_179_1194 ();
 b15zdnd11an1n64x5 FILLER_179_1258 ();
 b15zdnd11an1n64x5 FILLER_179_1322 ();
 b15zdnd11an1n64x5 FILLER_179_1386 ();
 b15zdnd11an1n64x5 FILLER_179_1450 ();
 b15zdnd11an1n64x5 FILLER_179_1514 ();
 b15zdnd11an1n64x5 FILLER_179_1578 ();
 b15zdnd11an1n08x5 FILLER_179_1642 ();
 b15zdnd00an1n02x5 FILLER_179_1650 ();
 b15zdnd00an1n01x5 FILLER_179_1652 ();
 b15zdnd11an1n04x5 FILLER_179_1664 ();
 b15zdnd11an1n64x5 FILLER_179_1720 ();
 b15zdnd11an1n16x5 FILLER_179_1784 ();
 b15zdnd11an1n08x5 FILLER_179_1800 ();
 b15zdnd11an1n04x5 FILLER_179_1808 ();
 b15zdnd00an1n02x5 FILLER_179_1812 ();
 b15zdnd00an1n01x5 FILLER_179_1814 ();
 b15zdnd11an1n16x5 FILLER_179_1818 ();
 b15zdnd11an1n04x5 FILLER_179_1837 ();
 b15zdnd11an1n64x5 FILLER_179_1844 ();
 b15zdnd11an1n64x5 FILLER_179_1908 ();
 b15zdnd11an1n64x5 FILLER_179_1972 ();
 b15zdnd11an1n32x5 FILLER_179_2036 ();
 b15zdnd11an1n08x5 FILLER_179_2068 ();
 b15zdnd11an1n04x5 FILLER_179_2076 ();
 b15zdnd00an1n02x5 FILLER_179_2080 ();
 b15zdnd00an1n01x5 FILLER_179_2082 ();
 b15zdnd11an1n04x5 FILLER_179_2123 ();
 b15zdnd11an1n32x5 FILLER_179_2130 ();
 b15zdnd11an1n16x5 FILLER_179_2162 ();
 b15zdnd11an1n08x5 FILLER_179_2178 ();
 b15zdnd11an1n04x5 FILLER_179_2191 ();
 b15zdnd11an1n64x5 FILLER_179_2202 ();
 b15zdnd11an1n16x5 FILLER_179_2266 ();
 b15zdnd00an1n02x5 FILLER_179_2282 ();
 b15zdnd11an1n64x5 FILLER_180_8 ();
 b15zdnd11an1n64x5 FILLER_180_72 ();
 b15zdnd11an1n64x5 FILLER_180_136 ();
 b15zdnd11an1n64x5 FILLER_180_200 ();
 b15zdnd11an1n64x5 FILLER_180_264 ();
 b15zdnd11an1n64x5 FILLER_180_328 ();
 b15zdnd11an1n64x5 FILLER_180_392 ();
 b15zdnd11an1n64x5 FILLER_180_456 ();
 b15zdnd11an1n64x5 FILLER_180_520 ();
 b15zdnd11an1n64x5 FILLER_180_584 ();
 b15zdnd11an1n64x5 FILLER_180_648 ();
 b15zdnd11an1n04x5 FILLER_180_712 ();
 b15zdnd00an1n02x5 FILLER_180_716 ();
 b15zdnd11an1n64x5 FILLER_180_726 ();
 b15zdnd11an1n64x5 FILLER_180_790 ();
 b15zdnd11an1n32x5 FILLER_180_854 ();
 b15zdnd11an1n16x5 FILLER_180_886 ();
 b15zdnd11an1n04x5 FILLER_180_902 ();
 b15zdnd00an1n02x5 FILLER_180_906 ();
 b15zdnd00an1n01x5 FILLER_180_908 ();
 b15zdnd11an1n64x5 FILLER_180_921 ();
 b15zdnd11an1n64x5 FILLER_180_985 ();
 b15zdnd11an1n64x5 FILLER_180_1049 ();
 b15zdnd11an1n64x5 FILLER_180_1113 ();
 b15zdnd11an1n64x5 FILLER_180_1177 ();
 b15zdnd11an1n64x5 FILLER_180_1241 ();
 b15zdnd11an1n64x5 FILLER_180_1305 ();
 b15zdnd11an1n64x5 FILLER_180_1369 ();
 b15zdnd11an1n32x5 FILLER_180_1433 ();
 b15zdnd11an1n04x5 FILLER_180_1465 ();
 b15zdnd00an1n01x5 FILLER_180_1469 ();
 b15zdnd11an1n64x5 FILLER_180_1479 ();
 b15zdnd11an1n64x5 FILLER_180_1543 ();
 b15zdnd11an1n64x5 FILLER_180_1607 ();
 b15zdnd11an1n08x5 FILLER_180_1671 ();
 b15zdnd11an1n04x5 FILLER_180_1679 ();
 b15zdnd00an1n02x5 FILLER_180_1683 ();
 b15zdnd00an1n01x5 FILLER_180_1685 ();
 b15zdnd11an1n04x5 FILLER_180_1689 ();
 b15zdnd11an1n64x5 FILLER_180_1696 ();
 b15zdnd11an1n16x5 FILLER_180_1760 ();
 b15zdnd11an1n08x5 FILLER_180_1776 ();
 b15zdnd11an1n04x5 FILLER_180_1784 ();
 b15zdnd00an1n02x5 FILLER_180_1788 ();
 b15zdnd00an1n01x5 FILLER_180_1790 ();
 b15zdnd11an1n64x5 FILLER_180_1843 ();
 b15zdnd11an1n64x5 FILLER_180_1907 ();
 b15zdnd11an1n64x5 FILLER_180_1971 ();
 b15zdnd11an1n64x5 FILLER_180_2035 ();
 b15zdnd11an1n16x5 FILLER_180_2099 ();
 b15zdnd11an1n04x5 FILLER_180_2115 ();
 b15zdnd11an1n32x5 FILLER_180_2122 ();
 b15zdnd11an1n64x5 FILLER_180_2162 ();
 b15zdnd11an1n32x5 FILLER_180_2226 ();
 b15zdnd11an1n16x5 FILLER_180_2258 ();
 b15zdnd00an1n02x5 FILLER_180_2274 ();
 b15zdnd11an1n04x5 FILLER_181_0 ();
 b15zdnd00an1n01x5 FILLER_181_4 ();
 b15zdnd11an1n16x5 FILLER_181_16 ();
 b15zdnd00an1n02x5 FILLER_181_32 ();
 b15zdnd00an1n01x5 FILLER_181_34 ();
 b15zdnd11an1n64x5 FILLER_181_49 ();
 b15zdnd11an1n64x5 FILLER_181_113 ();
 b15zdnd11an1n64x5 FILLER_181_177 ();
 b15zdnd11an1n64x5 FILLER_181_241 ();
 b15zdnd11an1n64x5 FILLER_181_305 ();
 b15zdnd11an1n64x5 FILLER_181_369 ();
 b15zdnd11an1n16x5 FILLER_181_433 ();
 b15zdnd11an1n64x5 FILLER_181_460 ();
 b15zdnd11an1n64x5 FILLER_181_524 ();
 b15zdnd11an1n64x5 FILLER_181_588 ();
 b15zdnd11an1n64x5 FILLER_181_652 ();
 b15zdnd11an1n64x5 FILLER_181_716 ();
 b15zdnd11an1n64x5 FILLER_181_780 ();
 b15zdnd11an1n64x5 FILLER_181_844 ();
 b15zdnd11an1n64x5 FILLER_181_908 ();
 b15zdnd11an1n64x5 FILLER_181_972 ();
 b15zdnd11an1n64x5 FILLER_181_1036 ();
 b15zdnd11an1n64x5 FILLER_181_1100 ();
 b15zdnd11an1n64x5 FILLER_181_1164 ();
 b15zdnd11an1n64x5 FILLER_181_1228 ();
 b15zdnd11an1n64x5 FILLER_181_1292 ();
 b15zdnd11an1n64x5 FILLER_181_1356 ();
 b15zdnd11an1n64x5 FILLER_181_1420 ();
 b15zdnd11an1n64x5 FILLER_181_1484 ();
 b15zdnd11an1n64x5 FILLER_181_1548 ();
 b15zdnd11an1n64x5 FILLER_181_1612 ();
 b15zdnd11an1n16x5 FILLER_181_1676 ();
 b15zdnd11an1n08x5 FILLER_181_1692 ();
 b15zdnd11an1n04x5 FILLER_181_1700 ();
 b15zdnd00an1n02x5 FILLER_181_1704 ();
 b15zdnd00an1n01x5 FILLER_181_1706 ();
 b15zdnd11an1n16x5 FILLER_181_1721 ();
 b15zdnd00an1n02x5 FILLER_181_1737 ();
 b15zdnd00an1n01x5 FILLER_181_1739 ();
 b15zdnd11an1n04x5 FILLER_181_1746 ();
 b15zdnd00an1n01x5 FILLER_181_1750 ();
 b15zdnd11an1n64x5 FILLER_181_1793 ();
 b15zdnd11an1n64x5 FILLER_181_1857 ();
 b15zdnd11an1n64x5 FILLER_181_1921 ();
 b15zdnd11an1n32x5 FILLER_181_1985 ();
 b15zdnd11an1n16x5 FILLER_181_2017 ();
 b15zdnd00an1n02x5 FILLER_181_2033 ();
 b15zdnd00an1n01x5 FILLER_181_2035 ();
 b15zdnd11an1n04x5 FILLER_181_2039 ();
 b15zdnd11an1n16x5 FILLER_181_2046 ();
 b15zdnd11an1n08x5 FILLER_181_2062 ();
 b15zdnd11an1n04x5 FILLER_181_2070 ();
 b15zdnd00an1n02x5 FILLER_181_2074 ();
 b15zdnd00an1n01x5 FILLER_181_2076 ();
 b15zdnd11an1n64x5 FILLER_181_2085 ();
 b15zdnd11an1n32x5 FILLER_181_2149 ();
 b15zdnd11an1n16x5 FILLER_181_2181 ();
 b15zdnd11an1n04x5 FILLER_181_2197 ();
 b15zdnd00an1n01x5 FILLER_181_2201 ();
 b15zdnd11an1n32x5 FILLER_181_2207 ();
 b15zdnd11an1n08x5 FILLER_181_2239 ();
 b15zdnd00an1n02x5 FILLER_181_2247 ();
 b15zdnd00an1n01x5 FILLER_181_2249 ();
 b15zdnd11an1n16x5 FILLER_181_2264 ();
 b15zdnd11an1n04x5 FILLER_181_2280 ();
 b15zdnd11an1n64x5 FILLER_182_8 ();
 b15zdnd11an1n32x5 FILLER_182_72 ();
 b15zdnd11an1n16x5 FILLER_182_104 ();
 b15zdnd11an1n08x5 FILLER_182_120 ();
 b15zdnd11an1n04x5 FILLER_182_128 ();
 b15zdnd00an1n02x5 FILLER_182_132 ();
 b15zdnd00an1n01x5 FILLER_182_134 ();
 b15zdnd11an1n64x5 FILLER_182_157 ();
 b15zdnd11an1n32x5 FILLER_182_221 ();
 b15zdnd11an1n08x5 FILLER_182_253 ();
 b15zdnd11an1n64x5 FILLER_182_269 ();
 b15zdnd11an1n64x5 FILLER_182_333 ();
 b15zdnd11an1n64x5 FILLER_182_397 ();
 b15zdnd11an1n64x5 FILLER_182_461 ();
 b15zdnd11an1n64x5 FILLER_182_525 ();
 b15zdnd11an1n64x5 FILLER_182_589 ();
 b15zdnd11an1n64x5 FILLER_182_653 ();
 b15zdnd00an1n01x5 FILLER_182_717 ();
 b15zdnd11an1n32x5 FILLER_182_726 ();
 b15zdnd00an1n01x5 FILLER_182_758 ();
 b15zdnd11an1n64x5 FILLER_182_773 ();
 b15zdnd11an1n64x5 FILLER_182_837 ();
 b15zdnd11an1n64x5 FILLER_182_901 ();
 b15zdnd11an1n32x5 FILLER_182_965 ();
 b15zdnd11an1n16x5 FILLER_182_997 ();
 b15zdnd11an1n08x5 FILLER_182_1013 ();
 b15zdnd11an1n64x5 FILLER_182_1041 ();
 b15zdnd11an1n64x5 FILLER_182_1105 ();
 b15zdnd11an1n64x5 FILLER_182_1169 ();
 b15zdnd11an1n64x5 FILLER_182_1233 ();
 b15zdnd11an1n64x5 FILLER_182_1297 ();
 b15zdnd11an1n64x5 FILLER_182_1361 ();
 b15zdnd11an1n64x5 FILLER_182_1425 ();
 b15zdnd11an1n64x5 FILLER_182_1489 ();
 b15zdnd11an1n64x5 FILLER_182_1553 ();
 b15zdnd11an1n64x5 FILLER_182_1617 ();
 b15zdnd11an1n64x5 FILLER_182_1681 ();
 b15zdnd11an1n64x5 FILLER_182_1745 ();
 b15zdnd11an1n64x5 FILLER_182_1809 ();
 b15zdnd11an1n32x5 FILLER_182_1873 ();
 b15zdnd11an1n08x5 FILLER_182_1905 ();
 b15zdnd00an1n02x5 FILLER_182_1913 ();
 b15zdnd00an1n01x5 FILLER_182_1915 ();
 b15zdnd11an1n64x5 FILLER_182_1937 ();
 b15zdnd11an1n08x5 FILLER_182_2001 ();
 b15zdnd11an1n04x5 FILLER_182_2009 ();
 b15zdnd00an1n01x5 FILLER_182_2013 ();
 b15zdnd11an1n16x5 FILLER_182_2046 ();
 b15zdnd00an1n02x5 FILLER_182_2062 ();
 b15zdnd00an1n01x5 FILLER_182_2064 ();
 b15zdnd11an1n04x5 FILLER_182_2069 ();
 b15zdnd00an1n02x5 FILLER_182_2073 ();
 b15zdnd11an1n08x5 FILLER_182_2078 ();
 b15zdnd00an1n02x5 FILLER_182_2086 ();
 b15zdnd00an1n01x5 FILLER_182_2088 ();
 b15zdnd11an1n32x5 FILLER_182_2094 ();
 b15zdnd11an1n16x5 FILLER_182_2126 ();
 b15zdnd11an1n08x5 FILLER_182_2142 ();
 b15zdnd11an1n04x5 FILLER_182_2150 ();
 b15zdnd11an1n64x5 FILLER_182_2162 ();
 b15zdnd11an1n16x5 FILLER_182_2226 ();
 b15zdnd11an1n08x5 FILLER_182_2242 ();
 b15zdnd11an1n04x5 FILLER_182_2250 ();
 b15zdnd00an1n01x5 FILLER_182_2254 ();
 b15zdnd11an1n08x5 FILLER_182_2266 ();
 b15zdnd00an1n02x5 FILLER_182_2274 ();
 b15zdnd11an1n64x5 FILLER_183_0 ();
 b15zdnd11an1n64x5 FILLER_183_64 ();
 b15zdnd11an1n16x5 FILLER_183_128 ();
 b15zdnd11an1n04x5 FILLER_183_144 ();
 b15zdnd11an1n64x5 FILLER_183_162 ();
 b15zdnd11an1n64x5 FILLER_183_226 ();
 b15zdnd11an1n08x5 FILLER_183_290 ();
 b15zdnd11an1n04x5 FILLER_183_298 ();
 b15zdnd11an1n64x5 FILLER_183_313 ();
 b15zdnd11an1n64x5 FILLER_183_377 ();
 b15zdnd11an1n32x5 FILLER_183_441 ();
 b15zdnd11an1n16x5 FILLER_183_493 ();
 b15zdnd11an1n08x5 FILLER_183_509 ();
 b15zdnd00an1n01x5 FILLER_183_517 ();
 b15zdnd11an1n64x5 FILLER_183_534 ();
 b15zdnd11an1n32x5 FILLER_183_598 ();
 b15zdnd11an1n16x5 FILLER_183_630 ();
 b15zdnd11an1n08x5 FILLER_183_646 ();
 b15zdnd00an1n01x5 FILLER_183_654 ();
 b15zdnd11an1n64x5 FILLER_183_664 ();
 b15zdnd11an1n64x5 FILLER_183_728 ();
 b15zdnd11an1n16x5 FILLER_183_792 ();
 b15zdnd00an1n02x5 FILLER_183_808 ();
 b15zdnd11an1n64x5 FILLER_183_827 ();
 b15zdnd11an1n64x5 FILLER_183_891 ();
 b15zdnd11an1n32x5 FILLER_183_955 ();
 b15zdnd11an1n16x5 FILLER_183_987 ();
 b15zdnd00an1n01x5 FILLER_183_1003 ();
 b15zdnd11an1n64x5 FILLER_183_1020 ();
 b15zdnd11an1n64x5 FILLER_183_1084 ();
 b15zdnd11an1n64x5 FILLER_183_1148 ();
 b15zdnd11an1n04x5 FILLER_183_1212 ();
 b15zdnd00an1n02x5 FILLER_183_1216 ();
 b15zdnd11an1n64x5 FILLER_183_1232 ();
 b15zdnd11an1n16x5 FILLER_183_1296 ();
 b15zdnd11an1n08x5 FILLER_183_1312 ();
 b15zdnd11an1n04x5 FILLER_183_1320 ();
 b15zdnd00an1n02x5 FILLER_183_1324 ();
 b15zdnd11an1n64x5 FILLER_183_1343 ();
 b15zdnd11an1n64x5 FILLER_183_1407 ();
 b15zdnd11an1n64x5 FILLER_183_1471 ();
 b15zdnd11an1n64x5 FILLER_183_1535 ();
 b15zdnd11an1n08x5 FILLER_183_1599 ();
 b15zdnd11an1n04x5 FILLER_183_1607 ();
 b15zdnd11an1n64x5 FILLER_183_1615 ();
 b15zdnd11an1n64x5 FILLER_183_1679 ();
 b15zdnd11an1n64x5 FILLER_183_1743 ();
 b15zdnd11an1n32x5 FILLER_183_1807 ();
 b15zdnd11an1n04x5 FILLER_183_1839 ();
 b15zdnd11an1n64x5 FILLER_183_1851 ();
 b15zdnd11an1n64x5 FILLER_183_1915 ();
 b15zdnd11an1n64x5 FILLER_183_1979 ();
 b15zdnd11an1n16x5 FILLER_183_2043 ();
 b15zdnd11an1n08x5 FILLER_183_2059 ();
 b15zdnd11an1n04x5 FILLER_183_2067 ();
 b15zdnd00an1n01x5 FILLER_183_2071 ();
 b15zdnd11an1n04x5 FILLER_183_2084 ();
 b15zdnd11an1n64x5 FILLER_183_2100 ();
 b15zdnd11an1n64x5 FILLER_183_2164 ();
 b15zdnd11an1n32x5 FILLER_183_2228 ();
 b15zdnd00an1n02x5 FILLER_183_2260 ();
 b15zdnd11an1n16x5 FILLER_183_2266 ();
 b15zdnd00an1n02x5 FILLER_183_2282 ();
 b15zdnd11an1n64x5 FILLER_184_8 ();
 b15zdnd11an1n64x5 FILLER_184_72 ();
 b15zdnd11an1n64x5 FILLER_184_136 ();
 b15zdnd11an1n64x5 FILLER_184_200 ();
 b15zdnd11an1n64x5 FILLER_184_264 ();
 b15zdnd11an1n64x5 FILLER_184_328 ();
 b15zdnd11an1n64x5 FILLER_184_392 ();
 b15zdnd11an1n64x5 FILLER_184_456 ();
 b15zdnd11an1n32x5 FILLER_184_520 ();
 b15zdnd11an1n04x5 FILLER_184_566 ();
 b15zdnd11an1n04x5 FILLER_184_593 ();
 b15zdnd11an1n64x5 FILLER_184_617 ();
 b15zdnd11an1n32x5 FILLER_184_681 ();
 b15zdnd11an1n04x5 FILLER_184_713 ();
 b15zdnd00an1n01x5 FILLER_184_717 ();
 b15zdnd11an1n64x5 FILLER_184_726 ();
 b15zdnd11an1n64x5 FILLER_184_790 ();
 b15zdnd11an1n64x5 FILLER_184_854 ();
 b15zdnd11an1n64x5 FILLER_184_918 ();
 b15zdnd11an1n64x5 FILLER_184_982 ();
 b15zdnd11an1n16x5 FILLER_184_1046 ();
 b15zdnd11an1n04x5 FILLER_184_1062 ();
 b15zdnd00an1n02x5 FILLER_184_1066 ();
 b15zdnd11an1n64x5 FILLER_184_1082 ();
 b15zdnd11an1n16x5 FILLER_184_1146 ();
 b15zdnd11an1n08x5 FILLER_184_1162 ();
 b15zdnd00an1n02x5 FILLER_184_1170 ();
 b15zdnd00an1n01x5 FILLER_184_1172 ();
 b15zdnd11an1n32x5 FILLER_184_1189 ();
 b15zdnd11an1n04x5 FILLER_184_1221 ();
 b15zdnd00an1n01x5 FILLER_184_1225 ();
 b15zdnd11an1n32x5 FILLER_184_1235 ();
 b15zdnd11an1n16x5 FILLER_184_1267 ();
 b15zdnd11an1n04x5 FILLER_184_1283 ();
 b15zdnd00an1n01x5 FILLER_184_1287 ();
 b15zdnd11an1n32x5 FILLER_184_1308 ();
 b15zdnd00an1n02x5 FILLER_184_1340 ();
 b15zdnd11an1n64x5 FILLER_184_1356 ();
 b15zdnd11an1n64x5 FILLER_184_1420 ();
 b15zdnd11an1n64x5 FILLER_184_1484 ();
 b15zdnd11an1n32x5 FILLER_184_1548 ();
 b15zdnd11an1n16x5 FILLER_184_1580 ();
 b15zdnd11an1n08x5 FILLER_184_1596 ();
 b15zdnd11an1n04x5 FILLER_184_1604 ();
 b15zdnd00an1n01x5 FILLER_184_1608 ();
 b15zdnd11an1n04x5 FILLER_184_1613 ();
 b15zdnd11an1n04x5 FILLER_184_1621 ();
 b15zdnd11an1n64x5 FILLER_184_1629 ();
 b15zdnd11an1n64x5 FILLER_184_1693 ();
 b15zdnd11an1n64x5 FILLER_184_1757 ();
 b15zdnd11an1n64x5 FILLER_184_1821 ();
 b15zdnd11an1n16x5 FILLER_184_1885 ();
 b15zdnd11an1n08x5 FILLER_184_1901 ();
 b15zdnd11an1n04x5 FILLER_184_1909 ();
 b15zdnd11an1n64x5 FILLER_184_1919 ();
 b15zdnd11an1n64x5 FILLER_184_1983 ();
 b15zdnd11an1n64x5 FILLER_184_2047 ();
 b15zdnd11an1n32x5 FILLER_184_2111 ();
 b15zdnd11an1n08x5 FILLER_184_2143 ();
 b15zdnd00an1n02x5 FILLER_184_2151 ();
 b15zdnd00an1n01x5 FILLER_184_2153 ();
 b15zdnd11an1n32x5 FILLER_184_2162 ();
 b15zdnd11an1n04x5 FILLER_184_2197 ();
 b15zdnd11an1n64x5 FILLER_184_2204 ();
 b15zdnd11an1n08x5 FILLER_184_2268 ();
 b15zdnd11an1n64x5 FILLER_185_0 ();
 b15zdnd11an1n64x5 FILLER_185_64 ();
 b15zdnd11an1n64x5 FILLER_185_128 ();
 b15zdnd11an1n64x5 FILLER_185_192 ();
 b15zdnd11an1n64x5 FILLER_185_256 ();
 b15zdnd11an1n64x5 FILLER_185_320 ();
 b15zdnd11an1n64x5 FILLER_185_384 ();
 b15zdnd11an1n04x5 FILLER_185_448 ();
 b15zdnd11an1n32x5 FILLER_185_459 ();
 b15zdnd11an1n16x5 FILLER_185_491 ();
 b15zdnd11an1n04x5 FILLER_185_507 ();
 b15zdnd00an1n02x5 FILLER_185_511 ();
 b15zdnd00an1n01x5 FILLER_185_513 ();
 b15zdnd11an1n04x5 FILLER_185_537 ();
 b15zdnd11an1n64x5 FILLER_185_547 ();
 b15zdnd11an1n64x5 FILLER_185_611 ();
 b15zdnd11an1n64x5 FILLER_185_675 ();
 b15zdnd11an1n64x5 FILLER_185_739 ();
 b15zdnd11an1n64x5 FILLER_185_803 ();
 b15zdnd11an1n64x5 FILLER_185_867 ();
 b15zdnd11an1n16x5 FILLER_185_931 ();
 b15zdnd11an1n04x5 FILLER_185_947 ();
 b15zdnd00an1n02x5 FILLER_185_951 ();
 b15zdnd11an1n04x5 FILLER_185_970 ();
 b15zdnd11an1n04x5 FILLER_185_994 ();
 b15zdnd11an1n04x5 FILLER_185_1010 ();
 b15zdnd00an1n01x5 FILLER_185_1014 ();
 b15zdnd11an1n04x5 FILLER_185_1046 ();
 b15zdnd11an1n04x5 FILLER_185_1062 ();
 b15zdnd00an1n02x5 FILLER_185_1066 ();
 b15zdnd11an1n08x5 FILLER_185_1080 ();
 b15zdnd11an1n04x5 FILLER_185_1088 ();
 b15zdnd00an1n01x5 FILLER_185_1092 ();
 b15zdnd11an1n16x5 FILLER_185_1107 ();
 b15zdnd11an1n04x5 FILLER_185_1143 ();
 b15zdnd00an1n02x5 FILLER_185_1147 ();
 b15zdnd11an1n16x5 FILLER_185_1155 ();
 b15zdnd11an1n04x5 FILLER_185_1171 ();
 b15zdnd11an1n04x5 FILLER_185_1187 ();
 b15zdnd11an1n64x5 FILLER_185_1196 ();
 b15zdnd11an1n64x5 FILLER_185_1260 ();
 b15zdnd11an1n64x5 FILLER_185_1350 ();
 b15zdnd11an1n64x5 FILLER_185_1414 ();
 b15zdnd11an1n64x5 FILLER_185_1478 ();
 b15zdnd11an1n64x5 FILLER_185_1542 ();
 b15zdnd11an1n04x5 FILLER_185_1606 ();
 b15zdnd11an1n08x5 FILLER_185_1614 ();
 b15zdnd11an1n04x5 FILLER_185_1622 ();
 b15zdnd11an1n64x5 FILLER_185_1630 ();
 b15zdnd00an1n02x5 FILLER_185_1694 ();
 b15zdnd11an1n04x5 FILLER_185_1708 ();
 b15zdnd11an1n64x5 FILLER_185_1732 ();
 b15zdnd11an1n64x5 FILLER_185_1796 ();
 b15zdnd11an1n64x5 FILLER_185_1860 ();
 b15zdnd11an1n64x5 FILLER_185_1924 ();
 b15zdnd11an1n64x5 FILLER_185_1988 ();
 b15zdnd11an1n64x5 FILLER_185_2052 ();
 b15zdnd11an1n32x5 FILLER_185_2116 ();
 b15zdnd11an1n16x5 FILLER_185_2148 ();
 b15zdnd11an1n08x5 FILLER_185_2164 ();
 b15zdnd11an1n04x5 FILLER_185_2172 ();
 b15zdnd11an1n16x5 FILLER_185_2228 ();
 b15zdnd00an1n02x5 FILLER_185_2244 ();
 b15zdnd11an1n32x5 FILLER_185_2250 ();
 b15zdnd00an1n02x5 FILLER_185_2282 ();
 b15zdnd11an1n64x5 FILLER_186_8 ();
 b15zdnd11an1n64x5 FILLER_186_72 ();
 b15zdnd11an1n64x5 FILLER_186_136 ();
 b15zdnd11an1n64x5 FILLER_186_200 ();
 b15zdnd11an1n32x5 FILLER_186_264 ();
 b15zdnd11an1n04x5 FILLER_186_296 ();
 b15zdnd00an1n02x5 FILLER_186_300 ();
 b15zdnd00an1n01x5 FILLER_186_302 ();
 b15zdnd11an1n64x5 FILLER_186_307 ();
 b15zdnd11an1n64x5 FILLER_186_371 ();
 b15zdnd11an1n64x5 FILLER_186_435 ();
 b15zdnd11an1n08x5 FILLER_186_499 ();
 b15zdnd00an1n02x5 FILLER_186_507 ();
 b15zdnd00an1n01x5 FILLER_186_509 ();
 b15zdnd11an1n04x5 FILLER_186_526 ();
 b15zdnd00an1n02x5 FILLER_186_530 ();
 b15zdnd11an1n64x5 FILLER_186_548 ();
 b15zdnd11an1n64x5 FILLER_186_612 ();
 b15zdnd11an1n32x5 FILLER_186_676 ();
 b15zdnd11an1n08x5 FILLER_186_708 ();
 b15zdnd00an1n02x5 FILLER_186_716 ();
 b15zdnd11an1n64x5 FILLER_186_726 ();
 b15zdnd11an1n64x5 FILLER_186_790 ();
 b15zdnd11an1n64x5 FILLER_186_854 ();
 b15zdnd11an1n32x5 FILLER_186_918 ();
 b15zdnd11an1n16x5 FILLER_186_950 ();
 b15zdnd11an1n08x5 FILLER_186_966 ();
 b15zdnd00an1n01x5 FILLER_186_974 ();
 b15zdnd11an1n16x5 FILLER_186_988 ();
 b15zdnd11an1n04x5 FILLER_186_1004 ();
 b15zdnd11an1n16x5 FILLER_186_1022 ();
 b15zdnd11an1n08x5 FILLER_186_1052 ();
 b15zdnd00an1n02x5 FILLER_186_1060 ();
 b15zdnd11an1n16x5 FILLER_186_1073 ();
 b15zdnd11an1n16x5 FILLER_186_1103 ();
 b15zdnd11an1n08x5 FILLER_186_1133 ();
 b15zdnd00an1n02x5 FILLER_186_1141 ();
 b15zdnd00an1n01x5 FILLER_186_1143 ();
 b15zdnd11an1n64x5 FILLER_186_1156 ();
 b15zdnd11an1n64x5 FILLER_186_1220 ();
 b15zdnd11an1n64x5 FILLER_186_1284 ();
 b15zdnd11an1n64x5 FILLER_186_1348 ();
 b15zdnd11an1n64x5 FILLER_186_1412 ();
 b15zdnd11an1n64x5 FILLER_186_1476 ();
 b15zdnd11an1n64x5 FILLER_186_1540 ();
 b15zdnd11an1n16x5 FILLER_186_1604 ();
 b15zdnd11an1n08x5 FILLER_186_1620 ();
 b15zdnd11an1n04x5 FILLER_186_1628 ();
 b15zdnd00an1n01x5 FILLER_186_1632 ();
 b15zdnd11an1n32x5 FILLER_186_1640 ();
 b15zdnd11an1n16x5 FILLER_186_1672 ();
 b15zdnd11an1n04x5 FILLER_186_1688 ();
 b15zdnd00an1n02x5 FILLER_186_1692 ();
 b15zdnd11an1n64x5 FILLER_186_1699 ();
 b15zdnd11an1n64x5 FILLER_186_1763 ();
 b15zdnd11an1n64x5 FILLER_186_1827 ();
 b15zdnd11an1n64x5 FILLER_186_1891 ();
 b15zdnd11an1n64x5 FILLER_186_1955 ();
 b15zdnd11an1n64x5 FILLER_186_2019 ();
 b15zdnd11an1n64x5 FILLER_186_2083 ();
 b15zdnd11an1n04x5 FILLER_186_2147 ();
 b15zdnd00an1n02x5 FILLER_186_2151 ();
 b15zdnd00an1n01x5 FILLER_186_2153 ();
 b15zdnd11an1n16x5 FILLER_186_2162 ();
 b15zdnd11an1n08x5 FILLER_186_2178 ();
 b15zdnd11an1n04x5 FILLER_186_2186 ();
 b15zdnd11an1n04x5 FILLER_186_2197 ();
 b15zdnd11an1n08x5 FILLER_186_2204 ();
 b15zdnd00an1n02x5 FILLER_186_2212 ();
 b15zdnd00an1n01x5 FILLER_186_2214 ();
 b15zdnd11an1n08x5 FILLER_186_2236 ();
 b15zdnd00an1n02x5 FILLER_186_2244 ();
 b15zdnd11an1n16x5 FILLER_186_2250 ();
 b15zdnd11an1n08x5 FILLER_186_2266 ();
 b15zdnd00an1n02x5 FILLER_186_2274 ();
 b15zdnd11an1n64x5 FILLER_187_0 ();
 b15zdnd11an1n64x5 FILLER_187_64 ();
 b15zdnd11an1n64x5 FILLER_187_128 ();
 b15zdnd11an1n32x5 FILLER_187_192 ();
 b15zdnd11an1n16x5 FILLER_187_224 ();
 b15zdnd11an1n08x5 FILLER_187_240 ();
 b15zdnd00an1n01x5 FILLER_187_248 ();
 b15zdnd11an1n64x5 FILLER_187_254 ();
 b15zdnd11an1n64x5 FILLER_187_318 ();
 b15zdnd11an1n64x5 FILLER_187_382 ();
 b15zdnd11an1n64x5 FILLER_187_446 ();
 b15zdnd11an1n32x5 FILLER_187_510 ();
 b15zdnd11an1n16x5 FILLER_187_542 ();
 b15zdnd11an1n08x5 FILLER_187_558 ();
 b15zdnd00an1n01x5 FILLER_187_566 ();
 b15zdnd11an1n64x5 FILLER_187_573 ();
 b15zdnd11an1n64x5 FILLER_187_637 ();
 b15zdnd11an1n64x5 FILLER_187_701 ();
 b15zdnd11an1n16x5 FILLER_187_765 ();
 b15zdnd11an1n08x5 FILLER_187_781 ();
 b15zdnd11an1n04x5 FILLER_187_789 ();
 b15zdnd00an1n01x5 FILLER_187_793 ();
 b15zdnd11an1n64x5 FILLER_187_803 ();
 b15zdnd11an1n16x5 FILLER_187_867 ();
 b15zdnd00an1n01x5 FILLER_187_883 ();
 b15zdnd11an1n64x5 FILLER_187_898 ();
 b15zdnd11an1n64x5 FILLER_187_962 ();
 b15zdnd11an1n64x5 FILLER_187_1026 ();
 b15zdnd11an1n64x5 FILLER_187_1090 ();
 b15zdnd11an1n64x5 FILLER_187_1154 ();
 b15zdnd11an1n64x5 FILLER_187_1218 ();
 b15zdnd11an1n64x5 FILLER_187_1282 ();
 b15zdnd11an1n32x5 FILLER_187_1346 ();
 b15zdnd11an1n16x5 FILLER_187_1378 ();
 b15zdnd11an1n08x5 FILLER_187_1394 ();
 b15zdnd11an1n04x5 FILLER_187_1402 ();
 b15zdnd00an1n02x5 FILLER_187_1406 ();
 b15zdnd00an1n01x5 FILLER_187_1408 ();
 b15zdnd11an1n08x5 FILLER_187_1461 ();
 b15zdnd11an1n04x5 FILLER_187_1469 ();
 b15zdnd11an1n32x5 FILLER_187_1481 ();
 b15zdnd11an1n16x5 FILLER_187_1513 ();
 b15zdnd11an1n04x5 FILLER_187_1529 ();
 b15zdnd00an1n01x5 FILLER_187_1533 ();
 b15zdnd11an1n64x5 FILLER_187_1537 ();
 b15zdnd11an1n16x5 FILLER_187_1601 ();
 b15zdnd11an1n08x5 FILLER_187_1617 ();
 b15zdnd00an1n02x5 FILLER_187_1625 ();
 b15zdnd11an1n08x5 FILLER_187_1636 ();
 b15zdnd11an1n04x5 FILLER_187_1644 ();
 b15zdnd00an1n01x5 FILLER_187_1648 ();
 b15zdnd11an1n64x5 FILLER_187_1669 ();
 b15zdnd11an1n16x5 FILLER_187_1733 ();
 b15zdnd00an1n02x5 FILLER_187_1749 ();
 b15zdnd00an1n01x5 FILLER_187_1751 ();
 b15zdnd11an1n04x5 FILLER_187_1761 ();
 b15zdnd11an1n08x5 FILLER_187_1771 ();
 b15zdnd00an1n02x5 FILLER_187_1779 ();
 b15zdnd00an1n01x5 FILLER_187_1781 ();
 b15zdnd11an1n64x5 FILLER_187_1799 ();
 b15zdnd11an1n64x5 FILLER_187_1863 ();
 b15zdnd11an1n64x5 FILLER_187_1927 ();
 b15zdnd11an1n64x5 FILLER_187_1991 ();
 b15zdnd11an1n64x5 FILLER_187_2055 ();
 b15zdnd11an1n64x5 FILLER_187_2119 ();
 b15zdnd11an1n32x5 FILLER_187_2183 ();
 b15zdnd11an1n16x5 FILLER_187_2236 ();
 b15zdnd11an1n08x5 FILLER_187_2252 ();
 b15zdnd11an1n04x5 FILLER_187_2260 ();
 b15zdnd00an1n02x5 FILLER_187_2264 ();
 b15zdnd00an1n01x5 FILLER_187_2266 ();
 b15zdnd11an1n04x5 FILLER_187_2278 ();
 b15zdnd00an1n02x5 FILLER_187_2282 ();
 b15zdnd11an1n64x5 FILLER_188_8 ();
 b15zdnd11an1n64x5 FILLER_188_72 ();
 b15zdnd11an1n64x5 FILLER_188_136 ();
 b15zdnd11an1n32x5 FILLER_188_200 ();
 b15zdnd00an1n02x5 FILLER_188_232 ();
 b15zdnd11an1n04x5 FILLER_188_240 ();
 b15zdnd11an1n04x5 FILLER_188_248 ();
 b15zdnd11an1n04x5 FILLER_188_258 ();
 b15zdnd11an1n16x5 FILLER_188_272 ();
 b15zdnd11an1n04x5 FILLER_188_288 ();
 b15zdnd00an1n02x5 FILLER_188_292 ();
 b15zdnd11an1n64x5 FILLER_188_298 ();
 b15zdnd11an1n64x5 FILLER_188_362 ();
 b15zdnd11an1n64x5 FILLER_188_426 ();
 b15zdnd11an1n64x5 FILLER_188_490 ();
 b15zdnd11an1n32x5 FILLER_188_554 ();
 b15zdnd11an1n08x5 FILLER_188_638 ();
 b15zdnd11an1n32x5 FILLER_188_649 ();
 b15zdnd00an1n01x5 FILLER_188_681 ();
 b15zdnd11an1n16x5 FILLER_188_692 ();
 b15zdnd11an1n08x5 FILLER_188_708 ();
 b15zdnd00an1n02x5 FILLER_188_716 ();
 b15zdnd11an1n64x5 FILLER_188_726 ();
 b15zdnd11an1n64x5 FILLER_188_790 ();
 b15zdnd11an1n64x5 FILLER_188_854 ();
 b15zdnd11an1n64x5 FILLER_188_918 ();
 b15zdnd11an1n64x5 FILLER_188_982 ();
 b15zdnd11an1n64x5 FILLER_188_1046 ();
 b15zdnd11an1n64x5 FILLER_188_1110 ();
 b15zdnd00an1n02x5 FILLER_188_1174 ();
 b15zdnd00an1n01x5 FILLER_188_1176 ();
 b15zdnd11an1n32x5 FILLER_188_1201 ();
 b15zdnd11an1n16x5 FILLER_188_1233 ();
 b15zdnd11an1n08x5 FILLER_188_1249 ();
 b15zdnd00an1n01x5 FILLER_188_1257 ();
 b15zdnd11an1n64x5 FILLER_188_1272 ();
 b15zdnd11an1n64x5 FILLER_188_1336 ();
 b15zdnd11an1n08x5 FILLER_188_1400 ();
 b15zdnd00an1n02x5 FILLER_188_1408 ();
 b15zdnd00an1n01x5 FILLER_188_1410 ();
 b15zdnd11an1n04x5 FILLER_188_1419 ();
 b15zdnd00an1n02x5 FILLER_188_1423 ();
 b15zdnd00an1n01x5 FILLER_188_1425 ();
 b15zdnd11an1n04x5 FILLER_188_1429 ();
 b15zdnd11an1n64x5 FILLER_188_1436 ();
 b15zdnd11an1n32x5 FILLER_188_1500 ();
 b15zdnd00an1n01x5 FILLER_188_1532 ();
 b15zdnd11an1n64x5 FILLER_188_1536 ();
 b15zdnd11an1n16x5 FILLER_188_1600 ();
 b15zdnd00an1n02x5 FILLER_188_1616 ();
 b15zdnd11an1n64x5 FILLER_188_1626 ();
 b15zdnd11an1n64x5 FILLER_188_1690 ();
 b15zdnd11an1n08x5 FILLER_188_1754 ();
 b15zdnd00an1n01x5 FILLER_188_1762 ();
 b15zdnd11an1n64x5 FILLER_188_1769 ();
 b15zdnd11an1n32x5 FILLER_188_1833 ();
 b15zdnd11an1n16x5 FILLER_188_1865 ();
 b15zdnd11an1n08x5 FILLER_188_1881 ();
 b15zdnd00an1n02x5 FILLER_188_1889 ();
 b15zdnd11an1n64x5 FILLER_188_1933 ();
 b15zdnd11an1n64x5 FILLER_188_1997 ();
 b15zdnd11an1n64x5 FILLER_188_2061 ();
 b15zdnd11an1n16x5 FILLER_188_2125 ();
 b15zdnd11an1n08x5 FILLER_188_2141 ();
 b15zdnd11an1n04x5 FILLER_188_2149 ();
 b15zdnd00an1n01x5 FILLER_188_2153 ();
 b15zdnd11an1n64x5 FILLER_188_2162 ();
 b15zdnd11an1n16x5 FILLER_188_2226 ();
 b15zdnd11an1n08x5 FILLER_188_2242 ();
 b15zdnd11an1n04x5 FILLER_188_2250 ();
 b15zdnd00an1n01x5 FILLER_188_2254 ();
 b15zdnd11an1n04x5 FILLER_188_2269 ();
 b15zdnd00an1n02x5 FILLER_188_2273 ();
 b15zdnd00an1n01x5 FILLER_188_2275 ();
 b15zdnd11an1n64x5 FILLER_189_0 ();
 b15zdnd11an1n08x5 FILLER_189_64 ();
 b15zdnd11an1n04x5 FILLER_189_72 ();
 b15zdnd11an1n64x5 FILLER_189_83 ();
 b15zdnd11an1n64x5 FILLER_189_147 ();
 b15zdnd11an1n04x5 FILLER_189_211 ();
 b15zdnd11an1n08x5 FILLER_189_218 ();
 b15zdnd00an1n02x5 FILLER_189_226 ();
 b15zdnd11an1n04x5 FILLER_189_233 ();
 b15zdnd00an1n02x5 FILLER_189_237 ();
 b15zdnd11an1n04x5 FILLER_189_257 ();
 b15zdnd11an1n08x5 FILLER_189_265 ();
 b15zdnd00an1n02x5 FILLER_189_273 ();
 b15zdnd11an1n32x5 FILLER_189_317 ();
 b15zdnd11an1n08x5 FILLER_189_349 ();
 b15zdnd00an1n01x5 FILLER_189_357 ();
 b15zdnd11an1n64x5 FILLER_189_372 ();
 b15zdnd11an1n08x5 FILLER_189_436 ();
 b15zdnd00an1n02x5 FILLER_189_444 ();
 b15zdnd11an1n64x5 FILLER_189_462 ();
 b15zdnd11an1n32x5 FILLER_189_526 ();
 b15zdnd11an1n32x5 FILLER_189_566 ();
 b15zdnd11an1n08x5 FILLER_189_598 ();
 b15zdnd11an1n04x5 FILLER_189_609 ();
 b15zdnd11an1n04x5 FILLER_189_616 ();
 b15zdnd00an1n01x5 FILLER_189_620 ();
 b15zdnd11an1n08x5 FILLER_189_673 ();
 b15zdnd11an1n16x5 FILLER_189_733 ();
 b15zdnd11an1n08x5 FILLER_189_749 ();
 b15zdnd11an1n04x5 FILLER_189_757 ();
 b15zdnd00an1n01x5 FILLER_189_761 ();
 b15zdnd11an1n16x5 FILLER_189_766 ();
 b15zdnd11an1n64x5 FILLER_189_786 ();
 b15zdnd11an1n08x5 FILLER_189_850 ();
 b15zdnd00an1n02x5 FILLER_189_858 ();
 b15zdnd00an1n01x5 FILLER_189_860 ();
 b15zdnd11an1n16x5 FILLER_189_881 ();
 b15zdnd11an1n04x5 FILLER_189_897 ();
 b15zdnd11an1n32x5 FILLER_189_904 ();
 b15zdnd11an1n16x5 FILLER_189_936 ();
 b15zdnd11an1n04x5 FILLER_189_952 ();
 b15zdnd00an1n02x5 FILLER_189_956 ();
 b15zdnd00an1n01x5 FILLER_189_958 ();
 b15zdnd11an1n04x5 FILLER_189_990 ();
 b15zdnd11an1n16x5 FILLER_189_997 ();
 b15zdnd11an1n08x5 FILLER_189_1013 ();
 b15zdnd11an1n04x5 FILLER_189_1021 ();
 b15zdnd00an1n01x5 FILLER_189_1025 ();
 b15zdnd11an1n64x5 FILLER_189_1037 ();
 b15zdnd11an1n08x5 FILLER_189_1101 ();
 b15zdnd11an1n04x5 FILLER_189_1109 ();
 b15zdnd11an1n64x5 FILLER_189_1116 ();
 b15zdnd11an1n64x5 FILLER_189_1180 ();
 b15zdnd11an1n08x5 FILLER_189_1244 ();
 b15zdnd11an1n32x5 FILLER_189_1272 ();
 b15zdnd11an1n16x5 FILLER_189_1304 ();
 b15zdnd11an1n04x5 FILLER_189_1320 ();
 b15zdnd00an1n02x5 FILLER_189_1324 ();
 b15zdnd11an1n32x5 FILLER_189_1331 ();
 b15zdnd11an1n16x5 FILLER_189_1363 ();
 b15zdnd11an1n04x5 FILLER_189_1379 ();
 b15zdnd00an1n02x5 FILLER_189_1383 ();
 b15zdnd11an1n04x5 FILLER_189_1388 ();
 b15zdnd11an1n32x5 FILLER_189_1395 ();
 b15zdnd11an1n08x5 FILLER_189_1427 ();
 b15zdnd11an1n64x5 FILLER_189_1438 ();
 b15zdnd11an1n04x5 FILLER_189_1502 ();
 b15zdnd00an1n02x5 FILLER_189_1506 ();
 b15zdnd11an1n16x5 FILLER_189_1560 ();
 b15zdnd11an1n08x5 FILLER_189_1576 ();
 b15zdnd11an1n04x5 FILLER_189_1584 ();
 b15zdnd11an1n64x5 FILLER_189_1592 ();
 b15zdnd11an1n64x5 FILLER_189_1656 ();
 b15zdnd11an1n16x5 FILLER_189_1720 ();
 b15zdnd11an1n08x5 FILLER_189_1736 ();
 b15zdnd00an1n02x5 FILLER_189_1744 ();
 b15zdnd11an1n16x5 FILLER_189_1764 ();
 b15zdnd11an1n08x5 FILLER_189_1780 ();
 b15zdnd00an1n01x5 FILLER_189_1788 ();
 b15zdnd11an1n64x5 FILLER_189_1800 ();
 b15zdnd11an1n32x5 FILLER_189_1864 ();
 b15zdnd11an1n08x5 FILLER_189_1896 ();
 b15zdnd00an1n01x5 FILLER_189_1904 ();
 b15zdnd11an1n64x5 FILLER_189_1908 ();
 b15zdnd11an1n64x5 FILLER_189_1972 ();
 b15zdnd11an1n64x5 FILLER_189_2036 ();
 b15zdnd11an1n64x5 FILLER_189_2100 ();
 b15zdnd11an1n32x5 FILLER_189_2164 ();
 b15zdnd11an1n08x5 FILLER_189_2196 ();
 b15zdnd11an1n04x5 FILLER_189_2204 ();
 b15zdnd00an1n02x5 FILLER_189_2208 ();
 b15zdnd11an1n04x5 FILLER_189_2218 ();
 b15zdnd11an1n32x5 FILLER_189_2226 ();
 b15zdnd11an1n16x5 FILLER_189_2258 ();
 b15zdnd11an1n08x5 FILLER_189_2274 ();
 b15zdnd00an1n02x5 FILLER_189_2282 ();
 b15zdnd11an1n64x5 FILLER_190_8 ();
 b15zdnd11an1n64x5 FILLER_190_72 ();
 b15zdnd11an1n64x5 FILLER_190_136 ();
 b15zdnd11an1n64x5 FILLER_190_200 ();
 b15zdnd11an1n32x5 FILLER_190_264 ();
 b15zdnd11an1n08x5 FILLER_190_296 ();
 b15zdnd11an1n64x5 FILLER_190_326 ();
 b15zdnd11an1n64x5 FILLER_190_390 ();
 b15zdnd11an1n08x5 FILLER_190_454 ();
 b15zdnd11an1n64x5 FILLER_190_476 ();
 b15zdnd11an1n16x5 FILLER_190_540 ();
 b15zdnd11an1n08x5 FILLER_190_556 ();
 b15zdnd00an1n02x5 FILLER_190_564 ();
 b15zdnd11an1n32x5 FILLER_190_576 ();
 b15zdnd00an1n02x5 FILLER_190_608 ();
 b15zdnd00an1n01x5 FILLER_190_610 ();
 b15zdnd11an1n16x5 FILLER_190_614 ();
 b15zdnd11an1n04x5 FILLER_190_630 ();
 b15zdnd00an1n02x5 FILLER_190_634 ();
 b15zdnd00an1n01x5 FILLER_190_636 ();
 b15zdnd11an1n08x5 FILLER_190_689 ();
 b15zdnd11an1n04x5 FILLER_190_697 ();
 b15zdnd11an1n04x5 FILLER_190_704 ();
 b15zdnd11an1n04x5 FILLER_190_711 ();
 b15zdnd00an1n02x5 FILLER_190_715 ();
 b15zdnd00an1n01x5 FILLER_190_717 ();
 b15zdnd11an1n64x5 FILLER_190_726 ();
 b15zdnd11an1n16x5 FILLER_190_790 ();
 b15zdnd00an1n02x5 FILLER_190_806 ();
 b15zdnd00an1n01x5 FILLER_190_808 ();
 b15zdnd11an1n32x5 FILLER_190_823 ();
 b15zdnd11an1n16x5 FILLER_190_855 ();
 b15zdnd11an1n04x5 FILLER_190_871 ();
 b15zdnd00an1n02x5 FILLER_190_875 ();
 b15zdnd00an1n01x5 FILLER_190_877 ();
 b15zdnd11an1n04x5 FILLER_190_930 ();
 b15zdnd11an1n64x5 FILLER_190_945 ();
 b15zdnd11an1n32x5 FILLER_190_1009 ();
 b15zdnd11an1n08x5 FILLER_190_1041 ();
 b15zdnd00an1n01x5 FILLER_190_1049 ();
 b15zdnd11an1n32x5 FILLER_190_1057 ();
 b15zdnd11an1n16x5 FILLER_190_1089 ();
 b15zdnd00an1n01x5 FILLER_190_1105 ();
 b15zdnd11an1n64x5 FILLER_190_1109 ();
 b15zdnd11an1n64x5 FILLER_190_1173 ();
 b15zdnd11an1n64x5 FILLER_190_1237 ();
 b15zdnd11an1n64x5 FILLER_190_1301 ();
 b15zdnd00an1n02x5 FILLER_190_1365 ();
 b15zdnd11an1n64x5 FILLER_190_1419 ();
 b15zdnd11an1n16x5 FILLER_190_1483 ();
 b15zdnd11an1n04x5 FILLER_190_1499 ();
 b15zdnd00an1n02x5 FILLER_190_1503 ();
 b15zdnd00an1n01x5 FILLER_190_1505 ();
 b15zdnd11an1n64x5 FILLER_190_1558 ();
 b15zdnd11an1n64x5 FILLER_190_1622 ();
 b15zdnd11an1n64x5 FILLER_190_1686 ();
 b15zdnd11an1n64x5 FILLER_190_1750 ();
 b15zdnd11an1n64x5 FILLER_190_1814 ();
 b15zdnd00an1n02x5 FILLER_190_1878 ();
 b15zdnd11an1n04x5 FILLER_190_1908 ();
 b15zdnd11an1n64x5 FILLER_190_1915 ();
 b15zdnd11an1n64x5 FILLER_190_1979 ();
 b15zdnd11an1n64x5 FILLER_190_2043 ();
 b15zdnd11an1n32x5 FILLER_190_2107 ();
 b15zdnd11an1n08x5 FILLER_190_2139 ();
 b15zdnd11an1n04x5 FILLER_190_2147 ();
 b15zdnd00an1n02x5 FILLER_190_2151 ();
 b15zdnd00an1n01x5 FILLER_190_2153 ();
 b15zdnd11an1n32x5 FILLER_190_2162 ();
 b15zdnd11an1n16x5 FILLER_190_2194 ();
 b15zdnd00an1n02x5 FILLER_190_2210 ();
 b15zdnd11an1n32x5 FILLER_190_2226 ();
 b15zdnd11an1n16x5 FILLER_190_2258 ();
 b15zdnd00an1n02x5 FILLER_190_2274 ();
 b15zdnd11an1n64x5 FILLER_191_0 ();
 b15zdnd11an1n64x5 FILLER_191_64 ();
 b15zdnd11an1n64x5 FILLER_191_128 ();
 b15zdnd11an1n64x5 FILLER_191_192 ();
 b15zdnd11an1n16x5 FILLER_191_256 ();
 b15zdnd11an1n04x5 FILLER_191_272 ();
 b15zdnd00an1n01x5 FILLER_191_276 ();
 b15zdnd11an1n08x5 FILLER_191_319 ();
 b15zdnd11an1n16x5 FILLER_191_330 ();
 b15zdnd11an1n08x5 FILLER_191_346 ();
 b15zdnd11an1n64x5 FILLER_191_365 ();
 b15zdnd11an1n16x5 FILLER_191_429 ();
 b15zdnd00an1n02x5 FILLER_191_445 ();
 b15zdnd00an1n01x5 FILLER_191_447 ();
 b15zdnd11an1n64x5 FILLER_191_460 ();
 b15zdnd11an1n64x5 FILLER_191_524 ();
 b15zdnd11an1n32x5 FILLER_191_588 ();
 b15zdnd11an1n16x5 FILLER_191_620 ();
 b15zdnd11an1n04x5 FILLER_191_636 ();
 b15zdnd00an1n01x5 FILLER_191_640 ();
 b15zdnd11an1n04x5 FILLER_191_644 ();
 b15zdnd11an1n04x5 FILLER_191_651 ();
 b15zdnd00an1n02x5 FILLER_191_655 ();
 b15zdnd11an1n04x5 FILLER_191_660 ();
 b15zdnd11an1n32x5 FILLER_191_667 ();
 b15zdnd11an1n08x5 FILLER_191_699 ();
 b15zdnd11an1n64x5 FILLER_191_710 ();
 b15zdnd11an1n32x5 FILLER_191_774 ();
 b15zdnd11an1n08x5 FILLER_191_806 ();
 b15zdnd11an1n04x5 FILLER_191_814 ();
 b15zdnd00an1n02x5 FILLER_191_818 ();
 b15zdnd00an1n01x5 FILLER_191_820 ();
 b15zdnd11an1n08x5 FILLER_191_841 ();
 b15zdnd00an1n02x5 FILLER_191_849 ();
 b15zdnd00an1n01x5 FILLER_191_851 ();
 b15zdnd11an1n16x5 FILLER_191_872 ();
 b15zdnd11an1n08x5 FILLER_191_888 ();
 b15zdnd00an1n02x5 FILLER_191_896 ();
 b15zdnd11an1n04x5 FILLER_191_901 ();
 b15zdnd11an1n64x5 FILLER_191_908 ();
 b15zdnd11an1n32x5 FILLER_191_972 ();
 b15zdnd11an1n16x5 FILLER_191_1004 ();
 b15zdnd11an1n04x5 FILLER_191_1020 ();
 b15zdnd11an1n64x5 FILLER_191_1027 ();
 b15zdnd11an1n64x5 FILLER_191_1091 ();
 b15zdnd11an1n64x5 FILLER_191_1155 ();
 b15zdnd11an1n64x5 FILLER_191_1219 ();
 b15zdnd11an1n64x5 FILLER_191_1283 ();
 b15zdnd11an1n16x5 FILLER_191_1347 ();
 b15zdnd11an1n04x5 FILLER_191_1363 ();
 b15zdnd00an1n02x5 FILLER_191_1367 ();
 b15zdnd00an1n01x5 FILLER_191_1369 ();
 b15zdnd11an1n16x5 FILLER_191_1374 ();
 b15zdnd11an1n04x5 FILLER_191_1393 ();
 b15zdnd11an1n04x5 FILLER_191_1400 ();
 b15zdnd11an1n64x5 FILLER_191_1407 ();
 b15zdnd11an1n32x5 FILLER_191_1471 ();
 b15zdnd11an1n16x5 FILLER_191_1503 ();
 b15zdnd11an1n04x5 FILLER_191_1519 ();
 b15zdnd00an1n02x5 FILLER_191_1523 ();
 b15zdnd11an1n04x5 FILLER_191_1528 ();
 b15zdnd11an1n04x5 FILLER_191_1535 ();
 b15zdnd11an1n64x5 FILLER_191_1542 ();
 b15zdnd11an1n64x5 FILLER_191_1606 ();
 b15zdnd11an1n64x5 FILLER_191_1670 ();
 b15zdnd11an1n64x5 FILLER_191_1734 ();
 b15zdnd11an1n64x5 FILLER_191_1798 ();
 b15zdnd11an1n04x5 FILLER_191_1902 ();
 b15zdnd11an1n64x5 FILLER_191_1909 ();
 b15zdnd11an1n64x5 FILLER_191_1973 ();
 b15zdnd11an1n64x5 FILLER_191_2037 ();
 b15zdnd11an1n64x5 FILLER_191_2101 ();
 b15zdnd11an1n64x5 FILLER_191_2165 ();
 b15zdnd11an1n32x5 FILLER_191_2229 ();
 b15zdnd11an1n16x5 FILLER_191_2261 ();
 b15zdnd11an1n04x5 FILLER_191_2277 ();
 b15zdnd00an1n02x5 FILLER_191_2281 ();
 b15zdnd00an1n01x5 FILLER_191_2283 ();
 b15zdnd11an1n64x5 FILLER_192_8 ();
 b15zdnd11an1n64x5 FILLER_192_103 ();
 b15zdnd11an1n64x5 FILLER_192_167 ();
 b15zdnd11an1n64x5 FILLER_192_231 ();
 b15zdnd11an1n08x5 FILLER_192_295 ();
 b15zdnd00an1n02x5 FILLER_192_303 ();
 b15zdnd00an1n01x5 FILLER_192_305 ();
 b15zdnd11an1n32x5 FILLER_192_348 ();
 b15zdnd11an1n16x5 FILLER_192_380 ();
 b15zdnd11an1n04x5 FILLER_192_396 ();
 b15zdnd00an1n02x5 FILLER_192_400 ();
 b15zdnd00an1n01x5 FILLER_192_402 ();
 b15zdnd11an1n08x5 FILLER_192_419 ();
 b15zdnd00an1n02x5 FILLER_192_427 ();
 b15zdnd11an1n64x5 FILLER_192_440 ();
 b15zdnd11an1n64x5 FILLER_192_504 ();
 b15zdnd11an1n64x5 FILLER_192_568 ();
 b15zdnd11an1n16x5 FILLER_192_632 ();
 b15zdnd11an1n08x5 FILLER_192_648 ();
 b15zdnd11an1n04x5 FILLER_192_656 ();
 b15zdnd00an1n02x5 FILLER_192_660 ();
 b15zdnd11an1n32x5 FILLER_192_665 ();
 b15zdnd11an1n16x5 FILLER_192_697 ();
 b15zdnd11an1n04x5 FILLER_192_713 ();
 b15zdnd00an1n01x5 FILLER_192_717 ();
 b15zdnd11an1n32x5 FILLER_192_726 ();
 b15zdnd11an1n16x5 FILLER_192_758 ();
 b15zdnd11an1n04x5 FILLER_192_774 ();
 b15zdnd11an1n04x5 FILLER_192_782 ();
 b15zdnd00an1n01x5 FILLER_192_786 ();
 b15zdnd11an1n16x5 FILLER_192_793 ();
 b15zdnd11an1n08x5 FILLER_192_809 ();
 b15zdnd11an1n04x5 FILLER_192_817 ();
 b15zdnd11an1n08x5 FILLER_192_833 ();
 b15zdnd11an1n04x5 FILLER_192_841 ();
 b15zdnd00an1n01x5 FILLER_192_845 ();
 b15zdnd11an1n64x5 FILLER_192_877 ();
 b15zdnd11an1n08x5 FILLER_192_941 ();
 b15zdnd11an1n04x5 FILLER_192_949 ();
 b15zdnd11an1n64x5 FILLER_192_958 ();
 b15zdnd11an1n64x5 FILLER_192_1022 ();
 b15zdnd11an1n64x5 FILLER_192_1086 ();
 b15zdnd11an1n64x5 FILLER_192_1150 ();
 b15zdnd11an1n64x5 FILLER_192_1214 ();
 b15zdnd11an1n64x5 FILLER_192_1278 ();
 b15zdnd11an1n16x5 FILLER_192_1342 ();
 b15zdnd11an1n08x5 FILLER_192_1358 ();
 b15zdnd11an1n04x5 FILLER_192_1366 ();
 b15zdnd00an1n02x5 FILLER_192_1370 ();
 b15zdnd11an1n64x5 FILLER_192_1424 ();
 b15zdnd11an1n32x5 FILLER_192_1488 ();
 b15zdnd11an1n04x5 FILLER_192_1520 ();
 b15zdnd00an1n02x5 FILLER_192_1524 ();
 b15zdnd00an1n01x5 FILLER_192_1526 ();
 b15zdnd11an1n64x5 FILLER_192_1530 ();
 b15zdnd11an1n64x5 FILLER_192_1594 ();
 b15zdnd11an1n64x5 FILLER_192_1658 ();
 b15zdnd11an1n32x5 FILLER_192_1722 ();
 b15zdnd11an1n08x5 FILLER_192_1754 ();
 b15zdnd11an1n04x5 FILLER_192_1762 ();
 b15zdnd00an1n02x5 FILLER_192_1766 ();
 b15zdnd00an1n01x5 FILLER_192_1768 ();
 b15zdnd11an1n64x5 FILLER_192_1775 ();
 b15zdnd11an1n32x5 FILLER_192_1839 ();
 b15zdnd11an1n16x5 FILLER_192_1871 ();
 b15zdnd11an1n04x5 FILLER_192_1887 ();
 b15zdnd00an1n02x5 FILLER_192_1891 ();
 b15zdnd11an1n32x5 FILLER_192_1896 ();
 b15zdnd11an1n16x5 FILLER_192_1928 ();
 b15zdnd11an1n08x5 FILLER_192_1944 ();
 b15zdnd00an1n02x5 FILLER_192_1952 ();
 b15zdnd11an1n16x5 FILLER_192_1959 ();
 b15zdnd11an1n04x5 FILLER_192_1975 ();
 b15zdnd00an1n02x5 FILLER_192_1979 ();
 b15zdnd11an1n64x5 FILLER_192_1988 ();
 b15zdnd11an1n32x5 FILLER_192_2052 ();
 b15zdnd11an1n08x5 FILLER_192_2084 ();
 b15zdnd11an1n32x5 FILLER_192_2096 ();
 b15zdnd11an1n16x5 FILLER_192_2128 ();
 b15zdnd11an1n08x5 FILLER_192_2144 ();
 b15zdnd00an1n02x5 FILLER_192_2152 ();
 b15zdnd11an1n32x5 FILLER_192_2162 ();
 b15zdnd11an1n16x5 FILLER_192_2194 ();
 b15zdnd11an1n08x5 FILLER_192_2210 ();
 b15zdnd00an1n02x5 FILLER_192_2218 ();
 b15zdnd00an1n01x5 FILLER_192_2220 ();
 b15zdnd11an1n08x5 FILLER_192_2263 ();
 b15zdnd11an1n04x5 FILLER_192_2271 ();
 b15zdnd00an1n01x5 FILLER_192_2275 ();
 b15zdnd11an1n64x5 FILLER_193_0 ();
 b15zdnd11an1n64x5 FILLER_193_64 ();
 b15zdnd11an1n64x5 FILLER_193_128 ();
 b15zdnd11an1n64x5 FILLER_193_192 ();
 b15zdnd11an1n32x5 FILLER_193_256 ();
 b15zdnd11an1n08x5 FILLER_193_288 ();
 b15zdnd11an1n04x5 FILLER_193_296 ();
 b15zdnd00an1n02x5 FILLER_193_300 ();
 b15zdnd00an1n01x5 FILLER_193_302 ();
 b15zdnd11an1n04x5 FILLER_193_308 ();
 b15zdnd00an1n02x5 FILLER_193_312 ();
 b15zdnd00an1n01x5 FILLER_193_314 ();
 b15zdnd11an1n64x5 FILLER_193_357 ();
 b15zdnd11an1n04x5 FILLER_193_421 ();
 b15zdnd11an1n08x5 FILLER_193_435 ();
 b15zdnd11an1n04x5 FILLER_193_443 ();
 b15zdnd11an1n32x5 FILLER_193_453 ();
 b15zdnd11an1n16x5 FILLER_193_507 ();
 b15zdnd11an1n04x5 FILLER_193_523 ();
 b15zdnd00an1n01x5 FILLER_193_527 ();
 b15zdnd11an1n16x5 FILLER_193_540 ();
 b15zdnd11an1n08x5 FILLER_193_556 ();
 b15zdnd11an1n16x5 FILLER_193_570 ();
 b15zdnd11an1n08x5 FILLER_193_586 ();
 b15zdnd00an1n02x5 FILLER_193_594 ();
 b15zdnd11an1n64x5 FILLER_193_600 ();
 b15zdnd11an1n08x5 FILLER_193_664 ();
 b15zdnd11an1n04x5 FILLER_193_672 ();
 b15zdnd00an1n02x5 FILLER_193_676 ();
 b15zdnd11an1n64x5 FILLER_193_686 ();
 b15zdnd11an1n16x5 FILLER_193_750 ();
 b15zdnd11an1n08x5 FILLER_193_766 ();
 b15zdnd11an1n04x5 FILLER_193_774 ();
 b15zdnd00an1n02x5 FILLER_193_778 ();
 b15zdnd00an1n01x5 FILLER_193_780 ();
 b15zdnd11an1n64x5 FILLER_193_798 ();
 b15zdnd11an1n16x5 FILLER_193_862 ();
 b15zdnd11an1n08x5 FILLER_193_878 ();
 b15zdnd11an1n04x5 FILLER_193_886 ();
 b15zdnd00an1n02x5 FILLER_193_890 ();
 b15zdnd00an1n01x5 FILLER_193_892 ();
 b15zdnd11an1n16x5 FILLER_193_913 ();
 b15zdnd11an1n08x5 FILLER_193_929 ();
 b15zdnd11an1n04x5 FILLER_193_937 ();
 b15zdnd11an1n64x5 FILLER_193_961 ();
 b15zdnd11an1n64x5 FILLER_193_1025 ();
 b15zdnd11an1n64x5 FILLER_193_1089 ();
 b15zdnd11an1n64x5 FILLER_193_1153 ();
 b15zdnd11an1n64x5 FILLER_193_1217 ();
 b15zdnd11an1n32x5 FILLER_193_1281 ();
 b15zdnd11an1n16x5 FILLER_193_1313 ();
 b15zdnd11an1n08x5 FILLER_193_1329 ();
 b15zdnd11an1n32x5 FILLER_193_1342 ();
 b15zdnd00an1n02x5 FILLER_193_1374 ();
 b15zdnd00an1n01x5 FILLER_193_1376 ();
 b15zdnd11an1n16x5 FILLER_193_1381 ();
 b15zdnd11an1n64x5 FILLER_193_1400 ();
 b15zdnd11an1n64x5 FILLER_193_1464 ();
 b15zdnd11an1n64x5 FILLER_193_1528 ();
 b15zdnd11an1n64x5 FILLER_193_1592 ();
 b15zdnd11an1n64x5 FILLER_193_1656 ();
 b15zdnd11an1n32x5 FILLER_193_1720 ();
 b15zdnd11an1n08x5 FILLER_193_1752 ();
 b15zdnd11an1n04x5 FILLER_193_1760 ();
 b15zdnd11an1n64x5 FILLER_193_1768 ();
 b15zdnd11an1n64x5 FILLER_193_1832 ();
 b15zdnd11an1n64x5 FILLER_193_1896 ();
 b15zdnd11an1n16x5 FILLER_193_1960 ();
 b15zdnd11an1n08x5 FILLER_193_1976 ();
 b15zdnd00an1n01x5 FILLER_193_1984 ();
 b15zdnd11an1n16x5 FILLER_193_2002 ();
 b15zdnd11an1n08x5 FILLER_193_2018 ();
 b15zdnd11an1n04x5 FILLER_193_2026 ();
 b15zdnd00an1n01x5 FILLER_193_2030 ();
 b15zdnd11an1n64x5 FILLER_193_2039 ();
 b15zdnd11an1n64x5 FILLER_193_2103 ();
 b15zdnd11an1n32x5 FILLER_193_2167 ();
 b15zdnd11an1n08x5 FILLER_193_2199 ();
 b15zdnd11an1n04x5 FILLER_193_2220 ();
 b15zdnd11an1n32x5 FILLER_193_2238 ();
 b15zdnd11an1n08x5 FILLER_193_2270 ();
 b15zdnd11an1n04x5 FILLER_193_2278 ();
 b15zdnd00an1n02x5 FILLER_193_2282 ();
 b15zdnd11an1n64x5 FILLER_194_8 ();
 b15zdnd11an1n64x5 FILLER_194_72 ();
 b15zdnd11an1n64x5 FILLER_194_136 ();
 b15zdnd11an1n16x5 FILLER_194_200 ();
 b15zdnd11an1n08x5 FILLER_194_216 ();
 b15zdnd11an1n04x5 FILLER_194_224 ();
 b15zdnd00an1n02x5 FILLER_194_228 ();
 b15zdnd00an1n01x5 FILLER_194_230 ();
 b15zdnd11an1n16x5 FILLER_194_273 ();
 b15zdnd11an1n08x5 FILLER_194_289 ();
 b15zdnd11an1n04x5 FILLER_194_297 ();
 b15zdnd00an1n02x5 FILLER_194_301 ();
 b15zdnd00an1n01x5 FILLER_194_303 ();
 b15zdnd11an1n64x5 FILLER_194_356 ();
 b15zdnd11an1n08x5 FILLER_194_420 ();
 b15zdnd11an1n04x5 FILLER_194_428 ();
 b15zdnd11an1n16x5 FILLER_194_454 ();
 b15zdnd11an1n04x5 FILLER_194_470 ();
 b15zdnd00an1n02x5 FILLER_194_474 ();
 b15zdnd00an1n01x5 FILLER_194_476 ();
 b15zdnd11an1n16x5 FILLER_194_491 ();
 b15zdnd11an1n08x5 FILLER_194_507 ();
 b15zdnd11an1n04x5 FILLER_194_515 ();
 b15zdnd11an1n64x5 FILLER_194_545 ();
 b15zdnd11an1n64x5 FILLER_194_609 ();
 b15zdnd11an1n32x5 FILLER_194_673 ();
 b15zdnd11an1n08x5 FILLER_194_705 ();
 b15zdnd11an1n04x5 FILLER_194_713 ();
 b15zdnd00an1n01x5 FILLER_194_717 ();
 b15zdnd11an1n64x5 FILLER_194_726 ();
 b15zdnd11an1n64x5 FILLER_194_790 ();
 b15zdnd11an1n64x5 FILLER_194_854 ();
 b15zdnd11an1n08x5 FILLER_194_918 ();
 b15zdnd00an1n02x5 FILLER_194_926 ();
 b15zdnd11an1n64x5 FILLER_194_940 ();
 b15zdnd11an1n64x5 FILLER_194_1004 ();
 b15zdnd11an1n32x5 FILLER_194_1068 ();
 b15zdnd11an1n08x5 FILLER_194_1100 ();
 b15zdnd11an1n64x5 FILLER_194_1113 ();
 b15zdnd11an1n64x5 FILLER_194_1177 ();
 b15zdnd11an1n64x5 FILLER_194_1241 ();
 b15zdnd11an1n64x5 FILLER_194_1305 ();
 b15zdnd11an1n64x5 FILLER_194_1369 ();
 b15zdnd11an1n64x5 FILLER_194_1433 ();
 b15zdnd11an1n64x5 FILLER_194_1497 ();
 b15zdnd11an1n64x5 FILLER_194_1561 ();
 b15zdnd11an1n64x5 FILLER_194_1625 ();
 b15zdnd11an1n64x5 FILLER_194_1689 ();
 b15zdnd11an1n64x5 FILLER_194_1753 ();
 b15zdnd11an1n64x5 FILLER_194_1817 ();
 b15zdnd11an1n64x5 FILLER_194_1881 ();
 b15zdnd11an1n64x5 FILLER_194_1945 ();
 b15zdnd11an1n64x5 FILLER_194_2009 ();
 b15zdnd11an1n64x5 FILLER_194_2073 ();
 b15zdnd11an1n16x5 FILLER_194_2137 ();
 b15zdnd00an1n01x5 FILLER_194_2153 ();
 b15zdnd11an1n64x5 FILLER_194_2162 ();
 b15zdnd11an1n32x5 FILLER_194_2226 ();
 b15zdnd11an1n16x5 FILLER_194_2258 ();
 b15zdnd00an1n02x5 FILLER_194_2274 ();
 b15zdnd00an1n02x5 FILLER_195_0 ();
 b15zdnd11an1n08x5 FILLER_195_6 ();
 b15zdnd00an1n02x5 FILLER_195_14 ();
 b15zdnd00an1n01x5 FILLER_195_16 ();
 b15zdnd11an1n64x5 FILLER_195_21 ();
 b15zdnd11an1n64x5 FILLER_195_85 ();
 b15zdnd11an1n64x5 FILLER_195_149 ();
 b15zdnd11an1n08x5 FILLER_195_213 ();
 b15zdnd11an1n04x5 FILLER_195_221 ();
 b15zdnd00an1n02x5 FILLER_195_225 ();
 b15zdnd00an1n01x5 FILLER_195_227 ();
 b15zdnd11an1n32x5 FILLER_195_270 ();
 b15zdnd11an1n08x5 FILLER_195_302 ();
 b15zdnd11an1n64x5 FILLER_195_341 ();
 b15zdnd11an1n64x5 FILLER_195_405 ();
 b15zdnd11an1n08x5 FILLER_195_469 ();
 b15zdnd11an1n04x5 FILLER_195_477 ();
 b15zdnd00an1n02x5 FILLER_195_481 ();
 b15zdnd00an1n01x5 FILLER_195_483 ();
 b15zdnd11an1n04x5 FILLER_195_504 ();
 b15zdnd11an1n64x5 FILLER_195_528 ();
 b15zdnd11an1n64x5 FILLER_195_592 ();
 b15zdnd11an1n64x5 FILLER_195_656 ();
 b15zdnd11an1n32x5 FILLER_195_720 ();
 b15zdnd11an1n16x5 FILLER_195_752 ();
 b15zdnd11an1n04x5 FILLER_195_768 ();
 b15zdnd00an1n02x5 FILLER_195_772 ();
 b15zdnd11an1n64x5 FILLER_195_780 ();
 b15zdnd11an1n64x5 FILLER_195_844 ();
 b15zdnd11an1n16x5 FILLER_195_908 ();
 b15zdnd11an1n08x5 FILLER_195_924 ();
 b15zdnd00an1n01x5 FILLER_195_932 ();
 b15zdnd11an1n64x5 FILLER_195_937 ();
 b15zdnd11an1n16x5 FILLER_195_1001 ();
 b15zdnd11an1n04x5 FILLER_195_1017 ();
 b15zdnd00an1n02x5 FILLER_195_1021 ();
 b15zdnd11an1n08x5 FILLER_195_1040 ();
 b15zdnd11an1n04x5 FILLER_195_1048 ();
 b15zdnd00an1n01x5 FILLER_195_1052 ();
 b15zdnd11an1n64x5 FILLER_195_1058 ();
 b15zdnd11an1n64x5 FILLER_195_1122 ();
 b15zdnd11an1n32x5 FILLER_195_1186 ();
 b15zdnd11an1n04x5 FILLER_195_1218 ();
 b15zdnd00an1n02x5 FILLER_195_1222 ();
 b15zdnd11an1n04x5 FILLER_195_1227 ();
 b15zdnd11an1n64x5 FILLER_195_1234 ();
 b15zdnd11an1n64x5 FILLER_195_1298 ();
 b15zdnd11an1n08x5 FILLER_195_1362 ();
 b15zdnd11an1n04x5 FILLER_195_1370 ();
 b15zdnd00an1n02x5 FILLER_195_1374 ();
 b15zdnd00an1n01x5 FILLER_195_1376 ();
 b15zdnd11an1n64x5 FILLER_195_1388 ();
 b15zdnd11an1n64x5 FILLER_195_1452 ();
 b15zdnd11an1n64x5 FILLER_195_1516 ();
 b15zdnd11an1n64x5 FILLER_195_1580 ();
 b15zdnd11an1n64x5 FILLER_195_1644 ();
 b15zdnd11an1n64x5 FILLER_195_1708 ();
 b15zdnd11an1n64x5 FILLER_195_1772 ();
 b15zdnd11an1n64x5 FILLER_195_1836 ();
 b15zdnd11an1n64x5 FILLER_195_1900 ();
 b15zdnd11an1n64x5 FILLER_195_1964 ();
 b15zdnd11an1n64x5 FILLER_195_2028 ();
 b15zdnd11an1n64x5 FILLER_195_2092 ();
 b15zdnd11an1n64x5 FILLER_195_2156 ();
 b15zdnd11an1n64x5 FILLER_195_2220 ();
 b15zdnd11an1n32x5 FILLER_196_8 ();
 b15zdnd11an1n16x5 FILLER_196_40 ();
 b15zdnd11an1n04x5 FILLER_196_56 ();
 b15zdnd00an1n02x5 FILLER_196_60 ();
 b15zdnd11an1n64x5 FILLER_196_65 ();
 b15zdnd11an1n64x5 FILLER_196_129 ();
 b15zdnd11an1n64x5 FILLER_196_193 ();
 b15zdnd11an1n64x5 FILLER_196_257 ();
 b15zdnd11an1n08x5 FILLER_196_321 ();
 b15zdnd00an1n01x5 FILLER_196_329 ();
 b15zdnd11an1n32x5 FILLER_196_333 ();
 b15zdnd11an1n08x5 FILLER_196_365 ();
 b15zdnd11an1n08x5 FILLER_196_377 ();
 b15zdnd11an1n04x5 FILLER_196_385 ();
 b15zdnd00an1n01x5 FILLER_196_389 ();
 b15zdnd11an1n04x5 FILLER_196_402 ();
 b15zdnd11an1n32x5 FILLER_196_422 ();
 b15zdnd11an1n04x5 FILLER_196_454 ();
 b15zdnd00an1n02x5 FILLER_196_458 ();
 b15zdnd11an1n32x5 FILLER_196_472 ();
 b15zdnd11an1n04x5 FILLER_196_504 ();
 b15zdnd11an1n04x5 FILLER_196_532 ();
 b15zdnd00an1n02x5 FILLER_196_536 ();
 b15zdnd00an1n01x5 FILLER_196_538 ();
 b15zdnd11an1n64x5 FILLER_196_558 ();
 b15zdnd11an1n64x5 FILLER_196_622 ();
 b15zdnd11an1n32x5 FILLER_196_686 ();
 b15zdnd11an1n64x5 FILLER_196_726 ();
 b15zdnd11an1n64x5 FILLER_196_790 ();
 b15zdnd11an1n64x5 FILLER_196_854 ();
 b15zdnd11an1n64x5 FILLER_196_918 ();
 b15zdnd11an1n32x5 FILLER_196_982 ();
 b15zdnd11an1n32x5 FILLER_196_1040 ();
 b15zdnd11an1n08x5 FILLER_196_1072 ();
 b15zdnd11an1n04x5 FILLER_196_1080 ();
 b15zdnd00an1n02x5 FILLER_196_1084 ();
 b15zdnd00an1n01x5 FILLER_196_1086 ();
 b15zdnd11an1n64x5 FILLER_196_1092 ();
 b15zdnd11an1n32x5 FILLER_196_1156 ();
 b15zdnd11an1n08x5 FILLER_196_1188 ();
 b15zdnd11an1n04x5 FILLER_196_1196 ();
 b15zdnd00an1n02x5 FILLER_196_1200 ();
 b15zdnd00an1n01x5 FILLER_196_1202 ();
 b15zdnd11an1n64x5 FILLER_196_1255 ();
 b15zdnd11an1n64x5 FILLER_196_1319 ();
 b15zdnd11an1n64x5 FILLER_196_1383 ();
 b15zdnd11an1n64x5 FILLER_196_1447 ();
 b15zdnd11an1n64x5 FILLER_196_1511 ();
 b15zdnd11an1n64x5 FILLER_196_1575 ();
 b15zdnd11an1n64x5 FILLER_196_1639 ();
 b15zdnd11an1n64x5 FILLER_196_1703 ();
 b15zdnd11an1n64x5 FILLER_196_1767 ();
 b15zdnd11an1n64x5 FILLER_196_1831 ();
 b15zdnd11an1n32x5 FILLER_196_1895 ();
 b15zdnd11an1n04x5 FILLER_196_1927 ();
 b15zdnd00an1n02x5 FILLER_196_1931 ();
 b15zdnd00an1n01x5 FILLER_196_1933 ();
 b15zdnd11an1n64x5 FILLER_196_1986 ();
 b15zdnd11an1n32x5 FILLER_196_2050 ();
 b15zdnd11an1n08x5 FILLER_196_2082 ();
 b15zdnd11an1n32x5 FILLER_196_2111 ();
 b15zdnd11an1n08x5 FILLER_196_2143 ();
 b15zdnd00an1n02x5 FILLER_196_2151 ();
 b15zdnd00an1n01x5 FILLER_196_2153 ();
 b15zdnd11an1n64x5 FILLER_196_2162 ();
 b15zdnd11an1n32x5 FILLER_196_2226 ();
 b15zdnd11an1n16x5 FILLER_196_2258 ();
 b15zdnd00an1n02x5 FILLER_196_2274 ();
 b15zdnd11an1n32x5 FILLER_197_0 ();
 b15zdnd00an1n02x5 FILLER_197_32 ();
 b15zdnd00an1n01x5 FILLER_197_34 ();
 b15zdnd11an1n64x5 FILLER_197_87 ();
 b15zdnd11an1n64x5 FILLER_197_151 ();
 b15zdnd11an1n64x5 FILLER_197_215 ();
 b15zdnd11an1n32x5 FILLER_197_279 ();
 b15zdnd11an1n16x5 FILLER_197_311 ();
 b15zdnd00an1n02x5 FILLER_197_327 ();
 b15zdnd11an1n32x5 FILLER_197_332 ();
 b15zdnd11an1n16x5 FILLER_197_364 ();
 b15zdnd00an1n02x5 FILLER_197_380 ();
 b15zdnd00an1n01x5 FILLER_197_382 ();
 b15zdnd11an1n32x5 FILLER_197_399 ();
 b15zdnd11an1n04x5 FILLER_197_431 ();
 b15zdnd00an1n01x5 FILLER_197_435 ();
 b15zdnd11an1n32x5 FILLER_197_443 ();
 b15zdnd11an1n04x5 FILLER_197_475 ();
 b15zdnd00an1n02x5 FILLER_197_479 ();
 b15zdnd00an1n01x5 FILLER_197_481 ();
 b15zdnd11an1n64x5 FILLER_197_492 ();
 b15zdnd11an1n64x5 FILLER_197_556 ();
 b15zdnd11an1n64x5 FILLER_197_620 ();
 b15zdnd11an1n64x5 FILLER_197_684 ();
 b15zdnd11an1n16x5 FILLER_197_748 ();
 b15zdnd11an1n08x5 FILLER_197_764 ();
 b15zdnd11an1n04x5 FILLER_197_772 ();
 b15zdnd11an1n64x5 FILLER_197_780 ();
 b15zdnd11an1n64x5 FILLER_197_844 ();
 b15zdnd11an1n32x5 FILLER_197_908 ();
 b15zdnd11an1n08x5 FILLER_197_940 ();
 b15zdnd00an1n01x5 FILLER_197_948 ();
 b15zdnd11an1n64x5 FILLER_197_957 ();
 b15zdnd11an1n32x5 FILLER_197_1021 ();
 b15zdnd11an1n16x5 FILLER_197_1053 ();
 b15zdnd11an1n08x5 FILLER_197_1069 ();
 b15zdnd11an1n04x5 FILLER_197_1077 ();
 b15zdnd11an1n04x5 FILLER_197_1084 ();
 b15zdnd00an1n02x5 FILLER_197_1088 ();
 b15zdnd11an1n64x5 FILLER_197_1107 ();
 b15zdnd11an1n16x5 FILLER_197_1171 ();
 b15zdnd11an1n08x5 FILLER_197_1187 ();
 b15zdnd00an1n02x5 FILLER_197_1195 ();
 b15zdnd11an1n64x5 FILLER_197_1249 ();
 b15zdnd11an1n64x5 FILLER_197_1313 ();
 b15zdnd11an1n64x5 FILLER_197_1377 ();
 b15zdnd11an1n64x5 FILLER_197_1441 ();
 b15zdnd11an1n64x5 FILLER_197_1505 ();
 b15zdnd11an1n64x5 FILLER_197_1569 ();
 b15zdnd11an1n64x5 FILLER_197_1633 ();
 b15zdnd11an1n32x5 FILLER_197_1697 ();
 b15zdnd11an1n16x5 FILLER_197_1729 ();
 b15zdnd11an1n04x5 FILLER_197_1745 ();
 b15zdnd00an1n02x5 FILLER_197_1749 ();
 b15zdnd00an1n01x5 FILLER_197_1751 ();
 b15zdnd11an1n64x5 FILLER_197_1756 ();
 b15zdnd11an1n64x5 FILLER_197_1820 ();
 b15zdnd11an1n64x5 FILLER_197_1884 ();
 b15zdnd11an1n04x5 FILLER_197_1948 ();
 b15zdnd11an1n04x5 FILLER_197_1955 ();
 b15zdnd11an1n04x5 FILLER_197_1962 ();
 b15zdnd11an1n08x5 FILLER_197_1969 ();
 b15zdnd11an1n04x5 FILLER_197_1977 ();
 b15zdnd11an1n64x5 FILLER_197_2023 ();
 b15zdnd11an1n16x5 FILLER_197_2087 ();
 b15zdnd11an1n04x5 FILLER_197_2103 ();
 b15zdnd11an1n64x5 FILLER_197_2115 ();
 b15zdnd11an1n64x5 FILLER_197_2179 ();
 b15zdnd11an1n32x5 FILLER_197_2243 ();
 b15zdnd11an1n08x5 FILLER_197_2275 ();
 b15zdnd00an1n01x5 FILLER_197_2283 ();
 b15zdnd11an1n32x5 FILLER_198_8 ();
 b15zdnd11an1n08x5 FILLER_198_40 ();
 b15zdnd11an1n04x5 FILLER_198_53 ();
 b15zdnd11an1n64x5 FILLER_198_60 ();
 b15zdnd11an1n16x5 FILLER_198_124 ();
 b15zdnd11an1n04x5 FILLER_198_140 ();
 b15zdnd00an1n01x5 FILLER_198_144 ();
 b15zdnd11an1n64x5 FILLER_198_177 ();
 b15zdnd11an1n64x5 FILLER_198_241 ();
 b15zdnd11an1n64x5 FILLER_198_305 ();
 b15zdnd00an1n02x5 FILLER_198_369 ();
 b15zdnd11an1n64x5 FILLER_198_389 ();
 b15zdnd11an1n08x5 FILLER_198_453 ();
 b15zdnd11an1n04x5 FILLER_198_461 ();
 b15zdnd00an1n01x5 FILLER_198_465 ();
 b15zdnd11an1n16x5 FILLER_198_482 ();
 b15zdnd11an1n08x5 FILLER_198_498 ();
 b15zdnd11an1n04x5 FILLER_198_506 ();
 b15zdnd11an1n16x5 FILLER_198_521 ();
 b15zdnd00an1n02x5 FILLER_198_537 ();
 b15zdnd00an1n01x5 FILLER_198_539 ();
 b15zdnd11an1n64x5 FILLER_198_554 ();
 b15zdnd11an1n64x5 FILLER_198_618 ();
 b15zdnd11an1n32x5 FILLER_198_682 ();
 b15zdnd11an1n04x5 FILLER_198_714 ();
 b15zdnd11an1n64x5 FILLER_198_726 ();
 b15zdnd11an1n64x5 FILLER_198_790 ();
 b15zdnd11an1n64x5 FILLER_198_854 ();
 b15zdnd11an1n08x5 FILLER_198_918 ();
 b15zdnd00an1n02x5 FILLER_198_926 ();
 b15zdnd11an1n08x5 FILLER_198_932 ();
 b15zdnd11an1n04x5 FILLER_198_940 ();
 b15zdnd00an1n02x5 FILLER_198_944 ();
 b15zdnd00an1n01x5 FILLER_198_946 ();
 b15zdnd11an1n04x5 FILLER_198_957 ();
 b15zdnd11an1n64x5 FILLER_198_973 ();
 b15zdnd11an1n16x5 FILLER_198_1037 ();
 b15zdnd11an1n04x5 FILLER_198_1053 ();
 b15zdnd11an1n04x5 FILLER_198_1101 ();
 b15zdnd11an1n64x5 FILLER_198_1136 ();
 b15zdnd11an1n16x5 FILLER_198_1200 ();
 b15zdnd11an1n04x5 FILLER_198_1219 ();
 b15zdnd11an1n04x5 FILLER_198_1226 ();
 b15zdnd11an1n64x5 FILLER_198_1233 ();
 b15zdnd11an1n64x5 FILLER_198_1297 ();
 b15zdnd11an1n64x5 FILLER_198_1361 ();
 b15zdnd11an1n64x5 FILLER_198_1425 ();
 b15zdnd11an1n64x5 FILLER_198_1489 ();
 b15zdnd11an1n64x5 FILLER_198_1553 ();
 b15zdnd11an1n64x5 FILLER_198_1617 ();
 b15zdnd11an1n64x5 FILLER_198_1681 ();
 b15zdnd11an1n64x5 FILLER_198_1745 ();
 b15zdnd11an1n64x5 FILLER_198_1809 ();
 b15zdnd11an1n64x5 FILLER_198_1873 ();
 b15zdnd11an1n16x5 FILLER_198_1937 ();
 b15zdnd11an1n04x5 FILLER_198_1953 ();
 b15zdnd00an1n02x5 FILLER_198_1957 ();
 b15zdnd11an1n64x5 FILLER_198_1984 ();
 b15zdnd11an1n32x5 FILLER_198_2048 ();
 b15zdnd11an1n08x5 FILLER_198_2080 ();
 b15zdnd11an1n32x5 FILLER_198_2096 ();
 b15zdnd11an1n16x5 FILLER_198_2128 ();
 b15zdnd11an1n08x5 FILLER_198_2144 ();
 b15zdnd00an1n02x5 FILLER_198_2152 ();
 b15zdnd11an1n64x5 FILLER_198_2162 ();
 b15zdnd11an1n32x5 FILLER_198_2226 ();
 b15zdnd11an1n16x5 FILLER_198_2258 ();
 b15zdnd00an1n02x5 FILLER_198_2274 ();
 b15zdnd11an1n32x5 FILLER_199_0 ();
 b15zdnd11an1n16x5 FILLER_199_32 ();
 b15zdnd11an1n08x5 FILLER_199_48 ();
 b15zdnd00an1n02x5 FILLER_199_56 ();
 b15zdnd00an1n01x5 FILLER_199_58 ();
 b15zdnd11an1n64x5 FILLER_199_62 ();
 b15zdnd11an1n64x5 FILLER_199_126 ();
 b15zdnd11an1n64x5 FILLER_199_190 ();
 b15zdnd11an1n16x5 FILLER_199_254 ();
 b15zdnd11an1n08x5 FILLER_199_270 ();
 b15zdnd11an1n04x5 FILLER_199_278 ();
 b15zdnd00an1n02x5 FILLER_199_282 ();
 b15zdnd11an1n64x5 FILLER_199_326 ();
 b15zdnd11an1n64x5 FILLER_199_390 ();
 b15zdnd11an1n32x5 FILLER_199_454 ();
 b15zdnd11an1n16x5 FILLER_199_486 ();
 b15zdnd11an1n08x5 FILLER_199_502 ();
 b15zdnd00an1n02x5 FILLER_199_510 ();
 b15zdnd00an1n01x5 FILLER_199_512 ();
 b15zdnd11an1n32x5 FILLER_199_539 ();
 b15zdnd00an1n02x5 FILLER_199_571 ();
 b15zdnd00an1n01x5 FILLER_199_573 ();
 b15zdnd11an1n64x5 FILLER_199_594 ();
 b15zdnd11an1n64x5 FILLER_199_658 ();
 b15zdnd11an1n64x5 FILLER_199_722 ();
 b15zdnd11an1n64x5 FILLER_199_786 ();
 b15zdnd11an1n64x5 FILLER_199_850 ();
 b15zdnd11an1n64x5 FILLER_199_914 ();
 b15zdnd11an1n64x5 FILLER_199_978 ();
 b15zdnd11an1n16x5 FILLER_199_1042 ();
 b15zdnd11an1n08x5 FILLER_199_1058 ();
 b15zdnd11an1n04x5 FILLER_199_1066 ();
 b15zdnd00an1n02x5 FILLER_199_1070 ();
 b15zdnd00an1n01x5 FILLER_199_1072 ();
 b15zdnd11an1n04x5 FILLER_199_1076 ();
 b15zdnd11an1n64x5 FILLER_199_1083 ();
 b15zdnd11an1n64x5 FILLER_199_1147 ();
 b15zdnd11an1n16x5 FILLER_199_1211 ();
 b15zdnd00an1n01x5 FILLER_199_1227 ();
 b15zdnd11an1n64x5 FILLER_199_1231 ();
 b15zdnd11an1n64x5 FILLER_199_1295 ();
 b15zdnd11an1n64x5 FILLER_199_1359 ();
 b15zdnd11an1n64x5 FILLER_199_1423 ();
 b15zdnd11an1n64x5 FILLER_199_1487 ();
 b15zdnd11an1n64x5 FILLER_199_1551 ();
 b15zdnd11an1n64x5 FILLER_199_1615 ();
 b15zdnd11an1n64x5 FILLER_199_1679 ();
 b15zdnd11an1n64x5 FILLER_199_1743 ();
 b15zdnd11an1n64x5 FILLER_199_1807 ();
 b15zdnd11an1n64x5 FILLER_199_1871 ();
 b15zdnd11an1n64x5 FILLER_199_1935 ();
 b15zdnd11an1n64x5 FILLER_199_1999 ();
 b15zdnd11an1n64x5 FILLER_199_2063 ();
 b15zdnd11an1n64x5 FILLER_199_2127 ();
 b15zdnd11an1n64x5 FILLER_199_2191 ();
 b15zdnd11an1n16x5 FILLER_199_2255 ();
 b15zdnd11an1n08x5 FILLER_199_2271 ();
 b15zdnd11an1n04x5 FILLER_199_2279 ();
 b15zdnd00an1n01x5 FILLER_199_2283 ();
 b15zdnd11an1n64x5 FILLER_200_8 ();
 b15zdnd00an1n02x5 FILLER_200_72 ();
 b15zdnd00an1n01x5 FILLER_200_74 ();
 b15zdnd11an1n64x5 FILLER_200_89 ();
 b15zdnd11an1n64x5 FILLER_200_153 ();
 b15zdnd11an1n08x5 FILLER_200_217 ();
 b15zdnd11an1n04x5 FILLER_200_225 ();
 b15zdnd00an1n02x5 FILLER_200_229 ();
 b15zdnd00an1n01x5 FILLER_200_231 ();
 b15zdnd11an1n64x5 FILLER_200_235 ();
 b15zdnd11an1n64x5 FILLER_200_299 ();
 b15zdnd11an1n32x5 FILLER_200_363 ();
 b15zdnd11an1n16x5 FILLER_200_395 ();
 b15zdnd00an1n02x5 FILLER_200_411 ();
 b15zdnd11an1n64x5 FILLER_200_429 ();
 b15zdnd11an1n64x5 FILLER_200_493 ();
 b15zdnd11an1n64x5 FILLER_200_557 ();
 b15zdnd11an1n64x5 FILLER_200_621 ();
 b15zdnd11an1n32x5 FILLER_200_685 ();
 b15zdnd00an1n01x5 FILLER_200_717 ();
 b15zdnd11an1n64x5 FILLER_200_726 ();
 b15zdnd11an1n64x5 FILLER_200_790 ();
 b15zdnd11an1n64x5 FILLER_200_854 ();
 b15zdnd11an1n64x5 FILLER_200_918 ();
 b15zdnd11an1n64x5 FILLER_200_982 ();
 b15zdnd11an1n64x5 FILLER_200_1046 ();
 b15zdnd11an1n64x5 FILLER_200_1110 ();
 b15zdnd11an1n64x5 FILLER_200_1174 ();
 b15zdnd11an1n64x5 FILLER_200_1238 ();
 b15zdnd11an1n16x5 FILLER_200_1302 ();
 b15zdnd11an1n04x5 FILLER_200_1318 ();
 b15zdnd11an1n64x5 FILLER_200_1342 ();
 b15zdnd11an1n64x5 FILLER_200_1406 ();
 b15zdnd11an1n64x5 FILLER_200_1470 ();
 b15zdnd11an1n64x5 FILLER_200_1534 ();
 b15zdnd11an1n64x5 FILLER_200_1598 ();
 b15zdnd11an1n64x5 FILLER_200_1662 ();
 b15zdnd11an1n32x5 FILLER_200_1726 ();
 b15zdnd11an1n08x5 FILLER_200_1758 ();
 b15zdnd11an1n64x5 FILLER_200_1770 ();
 b15zdnd11an1n64x5 FILLER_200_1834 ();
 b15zdnd11an1n64x5 FILLER_200_1898 ();
 b15zdnd11an1n64x5 FILLER_200_1962 ();
 b15zdnd11an1n64x5 FILLER_200_2026 ();
 b15zdnd11an1n64x5 FILLER_200_2090 ();
 b15zdnd11an1n32x5 FILLER_200_2162 ();
 b15zdnd11an1n04x5 FILLER_200_2194 ();
 b15zdnd00an1n02x5 FILLER_200_2198 ();
 b15zdnd00an1n01x5 FILLER_200_2200 ();
 b15zdnd11an1n04x5 FILLER_200_2204 ();
 b15zdnd11an1n64x5 FILLER_200_2211 ();
 b15zdnd00an1n01x5 FILLER_200_2275 ();
 b15zdnd11an1n64x5 FILLER_201_0 ();
 b15zdnd11an1n32x5 FILLER_201_64 ();
 b15zdnd11an1n64x5 FILLER_201_116 ();
 b15zdnd11an1n16x5 FILLER_201_180 ();
 b15zdnd11an1n08x5 FILLER_201_196 ();
 b15zdnd00an1n01x5 FILLER_201_204 ();
 b15zdnd11an1n64x5 FILLER_201_257 ();
 b15zdnd11an1n64x5 FILLER_201_321 ();
 b15zdnd11an1n64x5 FILLER_201_385 ();
 b15zdnd11an1n64x5 FILLER_201_449 ();
 b15zdnd11an1n64x5 FILLER_201_513 ();
 b15zdnd11an1n16x5 FILLER_201_577 ();
 b15zdnd11an1n04x5 FILLER_201_593 ();
 b15zdnd00an1n02x5 FILLER_201_597 ();
 b15zdnd00an1n01x5 FILLER_201_599 ();
 b15zdnd11an1n64x5 FILLER_201_611 ();
 b15zdnd11an1n64x5 FILLER_201_675 ();
 b15zdnd11an1n64x5 FILLER_201_739 ();
 b15zdnd11an1n64x5 FILLER_201_803 ();
 b15zdnd11an1n64x5 FILLER_201_867 ();
 b15zdnd11an1n64x5 FILLER_201_931 ();
 b15zdnd11an1n64x5 FILLER_201_995 ();
 b15zdnd11an1n64x5 FILLER_201_1059 ();
 b15zdnd11an1n64x5 FILLER_201_1123 ();
 b15zdnd11an1n64x5 FILLER_201_1187 ();
 b15zdnd11an1n64x5 FILLER_201_1251 ();
 b15zdnd11an1n64x5 FILLER_201_1315 ();
 b15zdnd11an1n64x5 FILLER_201_1379 ();
 b15zdnd11an1n64x5 FILLER_201_1443 ();
 b15zdnd11an1n64x5 FILLER_201_1507 ();
 b15zdnd11an1n64x5 FILLER_201_1571 ();
 b15zdnd11an1n64x5 FILLER_201_1635 ();
 b15zdnd11an1n64x5 FILLER_201_1699 ();
 b15zdnd11an1n64x5 FILLER_201_1763 ();
 b15zdnd11an1n64x5 FILLER_201_1827 ();
 b15zdnd11an1n32x5 FILLER_201_1891 ();
 b15zdnd11an1n16x5 FILLER_201_1923 ();
 b15zdnd11an1n04x5 FILLER_201_1939 ();
 b15zdnd00an1n02x5 FILLER_201_1943 ();
 b15zdnd11an1n64x5 FILLER_201_1987 ();
 b15zdnd11an1n64x5 FILLER_201_2051 ();
 b15zdnd11an1n32x5 FILLER_201_2115 ();
 b15zdnd11an1n16x5 FILLER_201_2147 ();
 b15zdnd11an1n08x5 FILLER_201_2163 ();
 b15zdnd11an1n04x5 FILLER_201_2171 ();
 b15zdnd00an1n01x5 FILLER_201_2175 ();
 b15zdnd11an1n32x5 FILLER_201_2228 ();
 b15zdnd11an1n16x5 FILLER_201_2260 ();
 b15zdnd11an1n08x5 FILLER_201_2276 ();
 b15zdnd11an1n64x5 FILLER_202_8 ();
 b15zdnd00an1n02x5 FILLER_202_72 ();
 b15zdnd00an1n01x5 FILLER_202_74 ();
 b15zdnd11an1n04x5 FILLER_202_120 ();
 b15zdnd11an1n64x5 FILLER_202_144 ();
 b15zdnd11an1n08x5 FILLER_202_208 ();
 b15zdnd00an1n01x5 FILLER_202_216 ();
 b15zdnd11an1n16x5 FILLER_202_269 ();
 b15zdnd11an1n08x5 FILLER_202_285 ();
 b15zdnd11an1n64x5 FILLER_202_300 ();
 b15zdnd11an1n08x5 FILLER_202_364 ();
 b15zdnd00an1n02x5 FILLER_202_372 ();
 b15zdnd00an1n01x5 FILLER_202_374 ();
 b15zdnd11an1n64x5 FILLER_202_386 ();
 b15zdnd11an1n64x5 FILLER_202_450 ();
 b15zdnd11an1n32x5 FILLER_202_514 ();
 b15zdnd00an1n02x5 FILLER_202_546 ();
 b15zdnd11an1n16x5 FILLER_202_570 ();
 b15zdnd11an1n08x5 FILLER_202_586 ();
 b15zdnd11an1n04x5 FILLER_202_594 ();
 b15zdnd11an1n64x5 FILLER_202_612 ();
 b15zdnd11an1n32x5 FILLER_202_676 ();
 b15zdnd11an1n08x5 FILLER_202_708 ();
 b15zdnd00an1n02x5 FILLER_202_716 ();
 b15zdnd11an1n64x5 FILLER_202_726 ();
 b15zdnd11an1n64x5 FILLER_202_790 ();
 b15zdnd11an1n64x5 FILLER_202_854 ();
 b15zdnd11an1n16x5 FILLER_202_918 ();
 b15zdnd00an1n02x5 FILLER_202_934 ();
 b15zdnd00an1n01x5 FILLER_202_936 ();
 b15zdnd11an1n64x5 FILLER_202_941 ();
 b15zdnd11an1n64x5 FILLER_202_1005 ();
 b15zdnd11an1n64x5 FILLER_202_1069 ();
 b15zdnd11an1n64x5 FILLER_202_1133 ();
 b15zdnd11an1n64x5 FILLER_202_1197 ();
 b15zdnd11an1n64x5 FILLER_202_1261 ();
 b15zdnd11an1n64x5 FILLER_202_1325 ();
 b15zdnd00an1n01x5 FILLER_202_1389 ();
 b15zdnd11an1n64x5 FILLER_202_1394 ();
 b15zdnd11an1n64x5 FILLER_202_1458 ();
 b15zdnd11an1n08x5 FILLER_202_1522 ();
 b15zdnd00an1n02x5 FILLER_202_1530 ();
 b15zdnd00an1n01x5 FILLER_202_1532 ();
 b15zdnd11an1n64x5 FILLER_202_1537 ();
 b15zdnd11an1n64x5 FILLER_202_1601 ();
 b15zdnd11an1n64x5 FILLER_202_1665 ();
 b15zdnd11an1n64x5 FILLER_202_1729 ();
 b15zdnd11an1n64x5 FILLER_202_1793 ();
 b15zdnd11an1n64x5 FILLER_202_1857 ();
 b15zdnd11an1n64x5 FILLER_202_1921 ();
 b15zdnd11an1n64x5 FILLER_202_1985 ();
 b15zdnd11an1n08x5 FILLER_202_2049 ();
 b15zdnd11an1n04x5 FILLER_202_2060 ();
 b15zdnd11an1n64x5 FILLER_202_2067 ();
 b15zdnd11an1n16x5 FILLER_202_2131 ();
 b15zdnd11an1n04x5 FILLER_202_2147 ();
 b15zdnd00an1n02x5 FILLER_202_2151 ();
 b15zdnd00an1n01x5 FILLER_202_2153 ();
 b15zdnd11an1n32x5 FILLER_202_2162 ();
 b15zdnd11an1n08x5 FILLER_202_2194 ();
 b15zdnd11an1n64x5 FILLER_202_2205 ();
 b15zdnd11an1n04x5 FILLER_202_2269 ();
 b15zdnd00an1n02x5 FILLER_202_2273 ();
 b15zdnd00an1n01x5 FILLER_202_2275 ();
 b15zdnd11an1n64x5 FILLER_203_0 ();
 b15zdnd11an1n64x5 FILLER_203_64 ();
 b15zdnd11an1n64x5 FILLER_203_128 ();
 b15zdnd11an1n16x5 FILLER_203_192 ();
 b15zdnd11an1n08x5 FILLER_203_208 ();
 b15zdnd11an1n04x5 FILLER_203_216 ();
 b15zdnd11an1n04x5 FILLER_203_223 ();
 b15zdnd00an1n02x5 FILLER_203_227 ();
 b15zdnd00an1n01x5 FILLER_203_229 ();
 b15zdnd11an1n04x5 FILLER_203_233 ();
 b15zdnd00an1n01x5 FILLER_203_237 ();
 b15zdnd11an1n04x5 FILLER_203_241 ();
 b15zdnd11an1n08x5 FILLER_203_248 ();
 b15zdnd00an1n02x5 FILLER_203_256 ();
 b15zdnd00an1n01x5 FILLER_203_258 ();
 b15zdnd11an1n64x5 FILLER_203_265 ();
 b15zdnd11an1n64x5 FILLER_203_329 ();
 b15zdnd11an1n32x5 FILLER_203_393 ();
 b15zdnd11an1n04x5 FILLER_203_425 ();
 b15zdnd00an1n01x5 FILLER_203_429 ();
 b15zdnd11an1n64x5 FILLER_203_450 ();
 b15zdnd11an1n64x5 FILLER_203_514 ();
 b15zdnd11an1n32x5 FILLER_203_578 ();
 b15zdnd11an1n16x5 FILLER_203_610 ();
 b15zdnd11an1n04x5 FILLER_203_626 ();
 b15zdnd11an1n64x5 FILLER_203_634 ();
 b15zdnd11an1n64x5 FILLER_203_698 ();
 b15zdnd11an1n64x5 FILLER_203_762 ();
 b15zdnd11an1n16x5 FILLER_203_826 ();
 b15zdnd11an1n08x5 FILLER_203_842 ();
 b15zdnd00an1n01x5 FILLER_203_850 ();
 b15zdnd11an1n64x5 FILLER_203_859 ();
 b15zdnd11an1n64x5 FILLER_203_923 ();
 b15zdnd11an1n64x5 FILLER_203_987 ();
 b15zdnd11an1n64x5 FILLER_203_1051 ();
 b15zdnd11an1n64x5 FILLER_203_1115 ();
 b15zdnd11an1n64x5 FILLER_203_1179 ();
 b15zdnd11an1n64x5 FILLER_203_1243 ();
 b15zdnd11an1n64x5 FILLER_203_1307 ();
 b15zdnd11an1n64x5 FILLER_203_1371 ();
 b15zdnd11an1n64x5 FILLER_203_1435 ();
 b15zdnd11an1n64x5 FILLER_203_1499 ();
 b15zdnd11an1n16x5 FILLER_203_1563 ();
 b15zdnd11an1n08x5 FILLER_203_1579 ();
 b15zdnd11an1n04x5 FILLER_203_1587 ();
 b15zdnd11an1n16x5 FILLER_203_1598 ();
 b15zdnd11an1n04x5 FILLER_203_1614 ();
 b15zdnd00an1n01x5 FILLER_203_1618 ();
 b15zdnd11an1n64x5 FILLER_203_1622 ();
 b15zdnd11an1n64x5 FILLER_203_1686 ();
 b15zdnd11an1n16x5 FILLER_203_1750 ();
 b15zdnd11an1n08x5 FILLER_203_1766 ();
 b15zdnd00an1n02x5 FILLER_203_1774 ();
 b15zdnd11an1n64x5 FILLER_203_1780 ();
 b15zdnd11an1n64x5 FILLER_203_1844 ();
 b15zdnd11an1n16x5 FILLER_203_1908 ();
 b15zdnd11an1n64x5 FILLER_203_1930 ();
 b15zdnd11an1n16x5 FILLER_203_1994 ();
 b15zdnd11an1n08x5 FILLER_203_2013 ();
 b15zdnd00an1n02x5 FILLER_203_2021 ();
 b15zdnd11an1n08x5 FILLER_203_2026 ();
 b15zdnd11an1n04x5 FILLER_203_2034 ();
 b15zdnd00an1n01x5 FILLER_203_2038 ();
 b15zdnd11an1n32x5 FILLER_203_2091 ();
 b15zdnd11an1n08x5 FILLER_203_2123 ();
 b15zdnd00an1n01x5 FILLER_203_2131 ();
 b15zdnd11an1n64x5 FILLER_203_2174 ();
 b15zdnd11an1n32x5 FILLER_203_2238 ();
 b15zdnd11an1n08x5 FILLER_203_2270 ();
 b15zdnd11an1n04x5 FILLER_203_2278 ();
 b15zdnd00an1n02x5 FILLER_203_2282 ();
 b15zdnd11an1n64x5 FILLER_204_8 ();
 b15zdnd11an1n64x5 FILLER_204_72 ();
 b15zdnd11an1n16x5 FILLER_204_136 ();
 b15zdnd11an1n08x5 FILLER_204_152 ();
 b15zdnd00an1n02x5 FILLER_204_160 ();
 b15zdnd11an1n32x5 FILLER_204_176 ();
 b15zdnd11an1n16x5 FILLER_204_208 ();
 b15zdnd11an1n08x5 FILLER_204_224 ();
 b15zdnd11an1n04x5 FILLER_204_232 ();
 b15zdnd00an1n02x5 FILLER_204_236 ();
 b15zdnd00an1n01x5 FILLER_204_238 ();
 b15zdnd11an1n04x5 FILLER_204_242 ();
 b15zdnd11an1n64x5 FILLER_204_253 ();
 b15zdnd11an1n32x5 FILLER_204_317 ();
 b15zdnd11an1n16x5 FILLER_204_349 ();
 b15zdnd11an1n08x5 FILLER_204_365 ();
 b15zdnd00an1n02x5 FILLER_204_373 ();
 b15zdnd11an1n04x5 FILLER_204_395 ();
 b15zdnd11an1n64x5 FILLER_204_413 ();
 b15zdnd11an1n64x5 FILLER_204_477 ();
 b15zdnd11an1n08x5 FILLER_204_541 ();
 b15zdnd11an1n04x5 FILLER_204_549 ();
 b15zdnd00an1n01x5 FILLER_204_553 ();
 b15zdnd11an1n64x5 FILLER_204_576 ();
 b15zdnd11an1n64x5 FILLER_204_640 ();
 b15zdnd11an1n08x5 FILLER_204_704 ();
 b15zdnd11an1n04x5 FILLER_204_712 ();
 b15zdnd00an1n02x5 FILLER_204_716 ();
 b15zdnd11an1n64x5 FILLER_204_726 ();
 b15zdnd11an1n64x5 FILLER_204_790 ();
 b15zdnd11an1n64x5 FILLER_204_854 ();
 b15zdnd11an1n64x5 FILLER_204_918 ();
 b15zdnd11an1n64x5 FILLER_204_982 ();
 b15zdnd11an1n64x5 FILLER_204_1046 ();
 b15zdnd11an1n64x5 FILLER_204_1110 ();
 b15zdnd11an1n64x5 FILLER_204_1174 ();
 b15zdnd11an1n64x5 FILLER_204_1238 ();
 b15zdnd11an1n64x5 FILLER_204_1302 ();
 b15zdnd11an1n64x5 FILLER_204_1366 ();
 b15zdnd11an1n64x5 FILLER_204_1430 ();
 b15zdnd11an1n64x5 FILLER_204_1494 ();
 b15zdnd11an1n32x5 FILLER_204_1558 ();
 b15zdnd11an1n16x5 FILLER_204_1590 ();
 b15zdnd11an1n08x5 FILLER_204_1606 ();
 b15zdnd00an1n02x5 FILLER_204_1614 ();
 b15zdnd00an1n01x5 FILLER_204_1616 ();
 b15zdnd11an1n04x5 FILLER_204_1620 ();
 b15zdnd11an1n64x5 FILLER_204_1627 ();
 b15zdnd11an1n64x5 FILLER_204_1691 ();
 b15zdnd11an1n64x5 FILLER_204_1755 ();
 b15zdnd11an1n64x5 FILLER_204_1819 ();
 b15zdnd11an1n32x5 FILLER_204_1883 ();
 b15zdnd11an1n08x5 FILLER_204_1915 ();
 b15zdnd00an1n02x5 FILLER_204_1923 ();
 b15zdnd00an1n01x5 FILLER_204_1925 ();
 b15zdnd11an1n32x5 FILLER_204_1939 ();
 b15zdnd11an1n16x5 FILLER_204_1971 ();
 b15zdnd00an1n01x5 FILLER_204_1987 ();
 b15zdnd11an1n16x5 FILLER_204_2040 ();
 b15zdnd11an1n08x5 FILLER_204_2056 ();
 b15zdnd00an1n01x5 FILLER_204_2064 ();
 b15zdnd11an1n64x5 FILLER_204_2068 ();
 b15zdnd11an1n16x5 FILLER_204_2132 ();
 b15zdnd11an1n04x5 FILLER_204_2148 ();
 b15zdnd00an1n02x5 FILLER_204_2152 ();
 b15zdnd11an1n32x5 FILLER_204_2162 ();
 b15zdnd11an1n08x5 FILLER_204_2194 ();
 b15zdnd11an1n04x5 FILLER_204_2207 ();
 b15zdnd11an1n32x5 FILLER_204_2217 ();
 b15zdnd11an1n16x5 FILLER_204_2249 ();
 b15zdnd11an1n08x5 FILLER_204_2265 ();
 b15zdnd00an1n02x5 FILLER_204_2273 ();
 b15zdnd00an1n01x5 FILLER_204_2275 ();
 b15zdnd11an1n64x5 FILLER_205_0 ();
 b15zdnd11an1n04x5 FILLER_205_64 ();
 b15zdnd00an1n02x5 FILLER_205_68 ();
 b15zdnd11an1n16x5 FILLER_205_91 ();
 b15zdnd11an1n04x5 FILLER_205_107 ();
 b15zdnd00an1n02x5 FILLER_205_111 ();
 b15zdnd11an1n64x5 FILLER_205_119 ();
 b15zdnd11an1n64x5 FILLER_205_183 ();
 b15zdnd11an1n64x5 FILLER_205_247 ();
 b15zdnd11an1n64x5 FILLER_205_311 ();
 b15zdnd11an1n64x5 FILLER_205_375 ();
 b15zdnd00an1n02x5 FILLER_205_439 ();
 b15zdnd00an1n01x5 FILLER_205_441 ();
 b15zdnd11an1n64x5 FILLER_205_456 ();
 b15zdnd11an1n32x5 FILLER_205_520 ();
 b15zdnd11an1n08x5 FILLER_205_552 ();
 b15zdnd11an1n04x5 FILLER_205_560 ();
 b15zdnd00an1n02x5 FILLER_205_564 ();
 b15zdnd00an1n01x5 FILLER_205_566 ();
 b15zdnd11an1n32x5 FILLER_205_587 ();
 b15zdnd11an1n16x5 FILLER_205_619 ();
 b15zdnd11an1n08x5 FILLER_205_635 ();
 b15zdnd11an1n04x5 FILLER_205_643 ();
 b15zdnd00an1n01x5 FILLER_205_647 ();
 b15zdnd11an1n64x5 FILLER_205_652 ();
 b15zdnd11an1n64x5 FILLER_205_716 ();
 b15zdnd11an1n32x5 FILLER_205_780 ();
 b15zdnd11an1n04x5 FILLER_205_812 ();
 b15zdnd00an1n02x5 FILLER_205_816 ();
 b15zdnd00an1n01x5 FILLER_205_818 ();
 b15zdnd11an1n32x5 FILLER_205_861 ();
 b15zdnd11an1n16x5 FILLER_205_893 ();
 b15zdnd00an1n02x5 FILLER_205_909 ();
 b15zdnd00an1n01x5 FILLER_205_911 ();
 b15zdnd11an1n08x5 FILLER_205_921 ();
 b15zdnd11an1n04x5 FILLER_205_929 ();
 b15zdnd00an1n02x5 FILLER_205_933 ();
 b15zdnd00an1n01x5 FILLER_205_935 ();
 b15zdnd11an1n64x5 FILLER_205_940 ();
 b15zdnd11an1n64x5 FILLER_205_1004 ();
 b15zdnd11an1n64x5 FILLER_205_1068 ();
 b15zdnd11an1n64x5 FILLER_205_1132 ();
 b15zdnd11an1n64x5 FILLER_205_1196 ();
 b15zdnd11an1n64x5 FILLER_205_1260 ();
 b15zdnd11an1n64x5 FILLER_205_1324 ();
 b15zdnd11an1n64x5 FILLER_205_1388 ();
 b15zdnd11an1n64x5 FILLER_205_1452 ();
 b15zdnd11an1n64x5 FILLER_205_1516 ();
 b15zdnd11an1n16x5 FILLER_205_1580 ();
 b15zdnd00an1n02x5 FILLER_205_1596 ();
 b15zdnd00an1n01x5 FILLER_205_1598 ();
 b15zdnd11an1n64x5 FILLER_205_1651 ();
 b15zdnd11an1n64x5 FILLER_205_1715 ();
 b15zdnd11an1n64x5 FILLER_205_1779 ();
 b15zdnd11an1n64x5 FILLER_205_1843 ();
 b15zdnd11an1n08x5 FILLER_205_1907 ();
 b15zdnd00an1n02x5 FILLER_205_1915 ();
 b15zdnd11an1n16x5 FILLER_205_1922 ();
 b15zdnd11an1n04x5 FILLER_205_1938 ();
 b15zdnd11an1n16x5 FILLER_205_1984 ();
 b15zdnd00an1n02x5 FILLER_205_2000 ();
 b15zdnd00an1n01x5 FILLER_205_2002 ();
 b15zdnd11an1n64x5 FILLER_205_2045 ();
 b15zdnd11an1n64x5 FILLER_205_2109 ();
 b15zdnd11an1n32x5 FILLER_205_2173 ();
 b15zdnd11an1n04x5 FILLER_205_2205 ();
 b15zdnd00an1n02x5 FILLER_205_2209 ();
 b15zdnd11an1n16x5 FILLER_205_2253 ();
 b15zdnd11an1n08x5 FILLER_205_2269 ();
 b15zdnd11an1n04x5 FILLER_205_2277 ();
 b15zdnd00an1n02x5 FILLER_205_2281 ();
 b15zdnd00an1n01x5 FILLER_205_2283 ();
 b15zdnd11an1n64x5 FILLER_206_8 ();
 b15zdnd11an1n64x5 FILLER_206_72 ();
 b15zdnd11an1n04x5 FILLER_206_136 ();
 b15zdnd00an1n02x5 FILLER_206_140 ();
 b15zdnd11an1n64x5 FILLER_206_149 ();
 b15zdnd11an1n64x5 FILLER_206_213 ();
 b15zdnd11an1n64x5 FILLER_206_277 ();
 b15zdnd11an1n64x5 FILLER_206_341 ();
 b15zdnd11an1n64x5 FILLER_206_405 ();
 b15zdnd11an1n64x5 FILLER_206_469 ();
 b15zdnd11an1n16x5 FILLER_206_533 ();
 b15zdnd11an1n08x5 FILLER_206_549 ();
 b15zdnd11an1n64x5 FILLER_206_581 ();
 b15zdnd11an1n64x5 FILLER_206_645 ();
 b15zdnd11an1n08x5 FILLER_206_709 ();
 b15zdnd00an1n01x5 FILLER_206_717 ();
 b15zdnd11an1n64x5 FILLER_206_726 ();
 b15zdnd11an1n32x5 FILLER_206_790 ();
 b15zdnd11an1n04x5 FILLER_206_822 ();
 b15zdnd00an1n01x5 FILLER_206_826 ();
 b15zdnd11an1n64x5 FILLER_206_869 ();
 b15zdnd11an1n64x5 FILLER_206_933 ();
 b15zdnd11an1n64x5 FILLER_206_997 ();
 b15zdnd11an1n64x5 FILLER_206_1061 ();
 b15zdnd11an1n64x5 FILLER_206_1125 ();
 b15zdnd11an1n64x5 FILLER_206_1189 ();
 b15zdnd11an1n64x5 FILLER_206_1253 ();
 b15zdnd11an1n64x5 FILLER_206_1317 ();
 b15zdnd11an1n64x5 FILLER_206_1381 ();
 b15zdnd11an1n64x5 FILLER_206_1445 ();
 b15zdnd11an1n08x5 FILLER_206_1509 ();
 b15zdnd11an1n04x5 FILLER_206_1517 ();
 b15zdnd00an1n02x5 FILLER_206_1521 ();
 b15zdnd00an1n01x5 FILLER_206_1523 ();
 b15zdnd11an1n32x5 FILLER_206_1528 ();
 b15zdnd11an1n16x5 FILLER_206_1560 ();
 b15zdnd11an1n08x5 FILLER_206_1576 ();
 b15zdnd11an1n08x5 FILLER_206_1590 ();
 b15zdnd00an1n01x5 FILLER_206_1598 ();
 b15zdnd11an1n64x5 FILLER_206_1651 ();
 b15zdnd11an1n64x5 FILLER_206_1715 ();
 b15zdnd11an1n64x5 FILLER_206_1779 ();
 b15zdnd11an1n64x5 FILLER_206_1843 ();
 b15zdnd11an1n08x5 FILLER_206_1907 ();
 b15zdnd11an1n04x5 FILLER_206_1915 ();
 b15zdnd00an1n02x5 FILLER_206_1919 ();
 b15zdnd11an1n04x5 FILLER_206_1924 ();
 b15zdnd11an1n04x5 FILLER_206_1938 ();
 b15zdnd11an1n04x5 FILLER_206_1954 ();
 b15zdnd11an1n04x5 FILLER_206_1963 ();
 b15zdnd00an1n02x5 FILLER_206_1967 ();
 b15zdnd00an1n01x5 FILLER_206_1969 ();
 b15zdnd11an1n04x5 FILLER_206_2012 ();
 b15zdnd11an1n64x5 FILLER_206_2019 ();
 b15zdnd11an1n64x5 FILLER_206_2083 ();
 b15zdnd11an1n04x5 FILLER_206_2147 ();
 b15zdnd00an1n02x5 FILLER_206_2151 ();
 b15zdnd00an1n01x5 FILLER_206_2153 ();
 b15zdnd11an1n32x5 FILLER_206_2162 ();
 b15zdnd11an1n08x5 FILLER_206_2194 ();
 b15zdnd00an1n02x5 FILLER_206_2202 ();
 b15zdnd00an1n01x5 FILLER_206_2204 ();
 b15zdnd11an1n64x5 FILLER_206_2210 ();
 b15zdnd00an1n02x5 FILLER_206_2274 ();
 b15zdnd11an1n64x5 FILLER_207_0 ();
 b15zdnd11an1n64x5 FILLER_207_64 ();
 b15zdnd11an1n32x5 FILLER_207_128 ();
 b15zdnd11an1n04x5 FILLER_207_160 ();
 b15zdnd00an1n02x5 FILLER_207_164 ();
 b15zdnd00an1n01x5 FILLER_207_166 ();
 b15zdnd11an1n64x5 FILLER_207_170 ();
 b15zdnd11an1n64x5 FILLER_207_234 ();
 b15zdnd11an1n64x5 FILLER_207_298 ();
 b15zdnd11an1n64x5 FILLER_207_362 ();
 b15zdnd11an1n64x5 FILLER_207_426 ();
 b15zdnd11an1n32x5 FILLER_207_490 ();
 b15zdnd00an1n02x5 FILLER_207_522 ();
 b15zdnd00an1n01x5 FILLER_207_524 ();
 b15zdnd11an1n64x5 FILLER_207_551 ();
 b15zdnd11an1n64x5 FILLER_207_615 ();
 b15zdnd11an1n64x5 FILLER_207_679 ();
 b15zdnd11an1n64x5 FILLER_207_743 ();
 b15zdnd11an1n64x5 FILLER_207_807 ();
 b15zdnd11an1n64x5 FILLER_207_871 ();
 b15zdnd11an1n64x5 FILLER_207_935 ();
 b15zdnd11an1n64x5 FILLER_207_999 ();
 b15zdnd11an1n64x5 FILLER_207_1063 ();
 b15zdnd11an1n64x5 FILLER_207_1127 ();
 b15zdnd11an1n64x5 FILLER_207_1191 ();
 b15zdnd11an1n64x5 FILLER_207_1255 ();
 b15zdnd11an1n64x5 FILLER_207_1319 ();
 b15zdnd11an1n64x5 FILLER_207_1383 ();
 b15zdnd11an1n32x5 FILLER_207_1447 ();
 b15zdnd11an1n08x5 FILLER_207_1479 ();
 b15zdnd11an1n04x5 FILLER_207_1487 ();
 b15zdnd00an1n01x5 FILLER_207_1491 ();
 b15zdnd11an1n08x5 FILLER_207_1512 ();
 b15zdnd11an1n04x5 FILLER_207_1520 ();
 b15zdnd11an1n64x5 FILLER_207_1528 ();
 b15zdnd11an1n16x5 FILLER_207_1592 ();
 b15zdnd11an1n08x5 FILLER_207_1608 ();
 b15zdnd00an1n01x5 FILLER_207_1616 ();
 b15zdnd11an1n04x5 FILLER_207_1620 ();
 b15zdnd11an1n16x5 FILLER_207_1627 ();
 b15zdnd11an1n04x5 FILLER_207_1643 ();
 b15zdnd00an1n01x5 FILLER_207_1647 ();
 b15zdnd11an1n64x5 FILLER_207_1655 ();
 b15zdnd11an1n32x5 FILLER_207_1719 ();
 b15zdnd11an1n08x5 FILLER_207_1751 ();
 b15zdnd00an1n02x5 FILLER_207_1759 ();
 b15zdnd00an1n01x5 FILLER_207_1761 ();
 b15zdnd11an1n04x5 FILLER_207_1765 ();
 b15zdnd11an1n08x5 FILLER_207_1772 ();
 b15zdnd11an1n04x5 FILLER_207_1780 ();
 b15zdnd00an1n02x5 FILLER_207_1784 ();
 b15zdnd00an1n01x5 FILLER_207_1786 ();
 b15zdnd11an1n64x5 FILLER_207_1791 ();
 b15zdnd11an1n64x5 FILLER_207_1855 ();
 b15zdnd00an1n01x5 FILLER_207_1919 ();
 b15zdnd11an1n04x5 FILLER_207_1930 ();
 b15zdnd11an1n04x5 FILLER_207_1940 ();
 b15zdnd00an1n02x5 FILLER_207_1944 ();
 b15zdnd00an1n01x5 FILLER_207_1946 ();
 b15zdnd11an1n08x5 FILLER_207_1951 ();
 b15zdnd11an1n04x5 FILLER_207_1959 ();
 b15zdnd00an1n02x5 FILLER_207_1963 ();
 b15zdnd00an1n01x5 FILLER_207_1965 ();
 b15zdnd11an1n04x5 FILLER_207_1969 ();
 b15zdnd00an1n02x5 FILLER_207_1973 ();
 b15zdnd00an1n01x5 FILLER_207_1975 ();
 b15zdnd11an1n64x5 FILLER_207_1982 ();
 b15zdnd11an1n64x5 FILLER_207_2046 ();
 b15zdnd11an1n64x5 FILLER_207_2110 ();
 b15zdnd11an1n64x5 FILLER_207_2174 ();
 b15zdnd11an1n32x5 FILLER_207_2238 ();
 b15zdnd11an1n08x5 FILLER_207_2270 ();
 b15zdnd11an1n04x5 FILLER_207_2278 ();
 b15zdnd00an1n02x5 FILLER_207_2282 ();
 b15zdnd11an1n64x5 FILLER_208_8 ();
 b15zdnd11an1n64x5 FILLER_208_72 ();
 b15zdnd11an1n04x5 FILLER_208_136 ();
 b15zdnd11an1n64x5 FILLER_208_192 ();
 b15zdnd11an1n64x5 FILLER_208_256 ();
 b15zdnd11an1n64x5 FILLER_208_320 ();
 b15zdnd11an1n64x5 FILLER_208_384 ();
 b15zdnd11an1n64x5 FILLER_208_448 ();
 b15zdnd11an1n64x5 FILLER_208_512 ();
 b15zdnd11an1n08x5 FILLER_208_576 ();
 b15zdnd11an1n04x5 FILLER_208_584 ();
 b15zdnd00an1n01x5 FILLER_208_588 ();
 b15zdnd11an1n64x5 FILLER_208_609 ();
 b15zdnd11an1n32x5 FILLER_208_673 ();
 b15zdnd11an1n08x5 FILLER_208_705 ();
 b15zdnd11an1n04x5 FILLER_208_713 ();
 b15zdnd00an1n01x5 FILLER_208_717 ();
 b15zdnd11an1n64x5 FILLER_208_726 ();
 b15zdnd11an1n64x5 FILLER_208_790 ();
 b15zdnd11an1n64x5 FILLER_208_854 ();
 b15zdnd11an1n64x5 FILLER_208_918 ();
 b15zdnd11an1n64x5 FILLER_208_982 ();
 b15zdnd11an1n08x5 FILLER_208_1046 ();
 b15zdnd11an1n04x5 FILLER_208_1054 ();
 b15zdnd00an1n02x5 FILLER_208_1058 ();
 b15zdnd11an1n64x5 FILLER_208_1063 ();
 b15zdnd11an1n64x5 FILLER_208_1127 ();
 b15zdnd11an1n64x5 FILLER_208_1191 ();
 b15zdnd11an1n64x5 FILLER_208_1255 ();
 b15zdnd11an1n32x5 FILLER_208_1319 ();
 b15zdnd11an1n08x5 FILLER_208_1351 ();
 b15zdnd00an1n02x5 FILLER_208_1359 ();
 b15zdnd00an1n01x5 FILLER_208_1361 ();
 b15zdnd11an1n04x5 FILLER_208_1365 ();
 b15zdnd11an1n32x5 FILLER_208_1372 ();
 b15zdnd11an1n08x5 FILLER_208_1404 ();
 b15zdnd00an1n02x5 FILLER_208_1412 ();
 b15zdnd00an1n01x5 FILLER_208_1414 ();
 b15zdnd11an1n64x5 FILLER_208_1419 ();
 b15zdnd11an1n32x5 FILLER_208_1483 ();
 b15zdnd11an1n08x5 FILLER_208_1515 ();
 b15zdnd11an1n04x5 FILLER_208_1523 ();
 b15zdnd00an1n02x5 FILLER_208_1527 ();
 b15zdnd00an1n01x5 FILLER_208_1529 ();
 b15zdnd11an1n64x5 FILLER_208_1550 ();
 b15zdnd11an1n08x5 FILLER_208_1614 ();
 b15zdnd00an1n01x5 FILLER_208_1622 ();
 b15zdnd11an1n64x5 FILLER_208_1626 ();
 b15zdnd11an1n16x5 FILLER_208_1690 ();
 b15zdnd11an1n08x5 FILLER_208_1706 ();
 b15zdnd00an1n01x5 FILLER_208_1714 ();
 b15zdnd11an1n08x5 FILLER_208_1722 ();
 b15zdnd11an1n04x5 FILLER_208_1730 ();
 b15zdnd00an1n02x5 FILLER_208_1734 ();
 b15zdnd00an1n01x5 FILLER_208_1736 ();
 b15zdnd11an1n16x5 FILLER_208_1789 ();
 b15zdnd11an1n08x5 FILLER_208_1805 ();
 b15zdnd11an1n04x5 FILLER_208_1813 ();
 b15zdnd00an1n01x5 FILLER_208_1817 ();
 b15zdnd11an1n64x5 FILLER_208_1826 ();
 b15zdnd11an1n64x5 FILLER_208_1890 ();
 b15zdnd11an1n64x5 FILLER_208_1954 ();
 b15zdnd11an1n64x5 FILLER_208_2018 ();
 b15zdnd11an1n32x5 FILLER_208_2082 ();
 b15zdnd11an1n04x5 FILLER_208_2114 ();
 b15zdnd00an1n01x5 FILLER_208_2118 ();
 b15zdnd11an1n04x5 FILLER_208_2122 ();
 b15zdnd11an1n16x5 FILLER_208_2129 ();
 b15zdnd11an1n08x5 FILLER_208_2145 ();
 b15zdnd00an1n01x5 FILLER_208_2153 ();
 b15zdnd11an1n64x5 FILLER_208_2162 ();
 b15zdnd11an1n32x5 FILLER_208_2226 ();
 b15zdnd11an1n16x5 FILLER_208_2258 ();
 b15zdnd00an1n02x5 FILLER_208_2274 ();
 b15zdnd11an1n64x5 FILLER_209_0 ();
 b15zdnd11an1n64x5 FILLER_209_64 ();
 b15zdnd11an1n08x5 FILLER_209_128 ();
 b15zdnd11an1n04x5 FILLER_209_136 ();
 b15zdnd00an1n02x5 FILLER_209_140 ();
 b15zdnd11an1n08x5 FILLER_209_149 ();
 b15zdnd00an1n01x5 FILLER_209_157 ();
 b15zdnd11an1n04x5 FILLER_209_161 ();
 b15zdnd11an1n64x5 FILLER_209_168 ();
 b15zdnd11an1n64x5 FILLER_209_232 ();
 b15zdnd11an1n64x5 FILLER_209_296 ();
 b15zdnd11an1n64x5 FILLER_209_360 ();
 b15zdnd11an1n64x5 FILLER_209_424 ();
 b15zdnd11an1n64x5 FILLER_209_488 ();
 b15zdnd11an1n08x5 FILLER_209_552 ();
 b15zdnd00an1n02x5 FILLER_209_560 ();
 b15zdnd11an1n64x5 FILLER_209_582 ();
 b15zdnd11an1n04x5 FILLER_209_646 ();
 b15zdnd00an1n02x5 FILLER_209_650 ();
 b15zdnd00an1n01x5 FILLER_209_652 ();
 b15zdnd11an1n64x5 FILLER_209_667 ();
 b15zdnd11an1n64x5 FILLER_209_731 ();
 b15zdnd11an1n08x5 FILLER_209_795 ();
 b15zdnd00an1n02x5 FILLER_209_803 ();
 b15zdnd11an1n64x5 FILLER_209_836 ();
 b15zdnd11an1n64x5 FILLER_209_900 ();
 b15zdnd11an1n16x5 FILLER_209_964 ();
 b15zdnd11an1n08x5 FILLER_209_980 ();
 b15zdnd00an1n02x5 FILLER_209_988 ();
 b15zdnd00an1n01x5 FILLER_209_990 ();
 b15zdnd11an1n32x5 FILLER_209_995 ();
 b15zdnd11an1n04x5 FILLER_209_1027 ();
 b15zdnd00an1n02x5 FILLER_209_1031 ();
 b15zdnd11an1n64x5 FILLER_209_1085 ();
 b15zdnd11an1n64x5 FILLER_209_1149 ();
 b15zdnd11an1n64x5 FILLER_209_1213 ();
 b15zdnd11an1n32x5 FILLER_209_1277 ();
 b15zdnd11an1n08x5 FILLER_209_1309 ();
 b15zdnd11an1n04x5 FILLER_209_1317 ();
 b15zdnd11an1n16x5 FILLER_209_1324 ();
 b15zdnd11an1n04x5 FILLER_209_1340 ();
 b15zdnd11an1n64x5 FILLER_209_1396 ();
 b15zdnd11an1n64x5 FILLER_209_1460 ();
 b15zdnd11an1n64x5 FILLER_209_1524 ();
 b15zdnd11an1n64x5 FILLER_209_1588 ();
 b15zdnd11an1n64x5 FILLER_209_1652 ();
 b15zdnd11an1n16x5 FILLER_209_1716 ();
 b15zdnd11an1n08x5 FILLER_209_1732 ();
 b15zdnd11an1n04x5 FILLER_209_1740 ();
 b15zdnd00an1n01x5 FILLER_209_1744 ();
 b15zdnd11an1n04x5 FILLER_209_1748 ();
 b15zdnd11an1n04x5 FILLER_209_1755 ();
 b15zdnd00an1n02x5 FILLER_209_1759 ();
 b15zdnd00an1n01x5 FILLER_209_1761 ();
 b15zdnd11an1n64x5 FILLER_209_1765 ();
 b15zdnd11an1n64x5 FILLER_209_1829 ();
 b15zdnd11an1n64x5 FILLER_209_1893 ();
 b15zdnd11an1n64x5 FILLER_209_1957 ();
 b15zdnd11an1n64x5 FILLER_209_2021 ();
 b15zdnd11an1n16x5 FILLER_209_2085 ();
 b15zdnd11an1n64x5 FILLER_209_2153 ();
 b15zdnd11an1n64x5 FILLER_209_2217 ();
 b15zdnd00an1n02x5 FILLER_209_2281 ();
 b15zdnd00an1n01x5 FILLER_209_2283 ();
 b15zdnd11an1n64x5 FILLER_210_8 ();
 b15zdnd11an1n64x5 FILLER_210_72 ();
 b15zdnd11an1n64x5 FILLER_210_136 ();
 b15zdnd11an1n64x5 FILLER_210_200 ();
 b15zdnd11an1n64x5 FILLER_210_264 ();
 b15zdnd11an1n64x5 FILLER_210_328 ();
 b15zdnd11an1n64x5 FILLER_210_392 ();
 b15zdnd11an1n64x5 FILLER_210_456 ();
 b15zdnd11an1n32x5 FILLER_210_520 ();
 b15zdnd11an1n16x5 FILLER_210_552 ();
 b15zdnd11an1n04x5 FILLER_210_568 ();
 b15zdnd11an1n64x5 FILLER_210_614 ();
 b15zdnd11an1n08x5 FILLER_210_678 ();
 b15zdnd11an1n04x5 FILLER_210_686 ();
 b15zdnd00an1n02x5 FILLER_210_690 ();
 b15zdnd00an1n01x5 FILLER_210_692 ();
 b15zdnd11an1n04x5 FILLER_210_713 ();
 b15zdnd00an1n01x5 FILLER_210_717 ();
 b15zdnd11an1n16x5 FILLER_210_726 ();
 b15zdnd11an1n08x5 FILLER_210_742 ();
 b15zdnd11an1n04x5 FILLER_210_750 ();
 b15zdnd00an1n02x5 FILLER_210_754 ();
 b15zdnd11an1n08x5 FILLER_210_763 ();
 b15zdnd11an1n04x5 FILLER_210_771 ();
 b15zdnd00an1n01x5 FILLER_210_775 ();
 b15zdnd11an1n64x5 FILLER_210_779 ();
 b15zdnd11an1n64x5 FILLER_210_843 ();
 b15zdnd11an1n64x5 FILLER_210_907 ();
 b15zdnd11an1n64x5 FILLER_210_971 ();
 b15zdnd11an1n16x5 FILLER_210_1035 ();
 b15zdnd11an1n04x5 FILLER_210_1054 ();
 b15zdnd11an1n16x5 FILLER_210_1061 ();
 b15zdnd11an1n04x5 FILLER_210_1077 ();
 b15zdnd11an1n64x5 FILLER_210_1112 ();
 b15zdnd11an1n04x5 FILLER_210_1176 ();
 b15zdnd00an1n02x5 FILLER_210_1180 ();
 b15zdnd11an1n64x5 FILLER_210_1190 ();
 b15zdnd11an1n32x5 FILLER_210_1254 ();
 b15zdnd00an1n01x5 FILLER_210_1286 ();
 b15zdnd11an1n32x5 FILLER_210_1327 ();
 b15zdnd11an1n08x5 FILLER_210_1359 ();
 b15zdnd00an1n02x5 FILLER_210_1367 ();
 b15zdnd00an1n01x5 FILLER_210_1369 ();
 b15zdnd11an1n64x5 FILLER_210_1373 ();
 b15zdnd11an1n64x5 FILLER_210_1437 ();
 b15zdnd11an1n64x5 FILLER_210_1501 ();
 b15zdnd11an1n32x5 FILLER_210_1565 ();
 b15zdnd11an1n16x5 FILLER_210_1597 ();
 b15zdnd00an1n02x5 FILLER_210_1613 ();
 b15zdnd11an1n64x5 FILLER_210_1623 ();
 b15zdnd11an1n32x5 FILLER_210_1687 ();
 b15zdnd00an1n01x5 FILLER_210_1719 ();
 b15zdnd11an1n64x5 FILLER_210_1772 ();
 b15zdnd11an1n64x5 FILLER_210_1836 ();
 b15zdnd11an1n64x5 FILLER_210_1900 ();
 b15zdnd11an1n64x5 FILLER_210_1964 ();
 b15zdnd11an1n64x5 FILLER_210_2028 ();
 b15zdnd11an1n32x5 FILLER_210_2092 ();
 b15zdnd00an1n02x5 FILLER_210_2124 ();
 b15zdnd11an1n16x5 FILLER_210_2129 ();
 b15zdnd11an1n08x5 FILLER_210_2145 ();
 b15zdnd00an1n01x5 FILLER_210_2153 ();
 b15zdnd11an1n64x5 FILLER_210_2162 ();
 b15zdnd11an1n32x5 FILLER_210_2226 ();
 b15zdnd11an1n16x5 FILLER_210_2258 ();
 b15zdnd00an1n02x5 FILLER_210_2274 ();
 b15zdnd11an1n64x5 FILLER_211_0 ();
 b15zdnd11an1n64x5 FILLER_211_64 ();
 b15zdnd11an1n64x5 FILLER_211_128 ();
 b15zdnd11an1n64x5 FILLER_211_192 ();
 b15zdnd11an1n64x5 FILLER_211_256 ();
 b15zdnd11an1n64x5 FILLER_211_320 ();
 b15zdnd11an1n64x5 FILLER_211_384 ();
 b15zdnd11an1n16x5 FILLER_211_448 ();
 b15zdnd11an1n08x5 FILLER_211_464 ();
 b15zdnd11an1n64x5 FILLER_211_482 ();
 b15zdnd11an1n16x5 FILLER_211_546 ();
 b15zdnd11an1n08x5 FILLER_211_562 ();
 b15zdnd11an1n16x5 FILLER_211_601 ();
 b15zdnd11an1n08x5 FILLER_211_617 ();
 b15zdnd00an1n02x5 FILLER_211_625 ();
 b15zdnd11an1n08x5 FILLER_211_638 ();
 b15zdnd11an1n04x5 FILLER_211_646 ();
 b15zdnd00an1n01x5 FILLER_211_650 ();
 b15zdnd11an1n04x5 FILLER_211_675 ();
 b15zdnd11an1n32x5 FILLER_211_705 ();
 b15zdnd11an1n08x5 FILLER_211_737 ();
 b15zdnd11an1n04x5 FILLER_211_745 ();
 b15zdnd00an1n02x5 FILLER_211_749 ();
 b15zdnd11an1n64x5 FILLER_211_803 ();
 b15zdnd11an1n64x5 FILLER_211_867 ();
 b15zdnd11an1n64x5 FILLER_211_931 ();
 b15zdnd11an1n64x5 FILLER_211_995 ();
 b15zdnd11an1n64x5 FILLER_211_1059 ();
 b15zdnd11an1n16x5 FILLER_211_1123 ();
 b15zdnd11an1n08x5 FILLER_211_1139 ();
 b15zdnd11an1n04x5 FILLER_211_1147 ();
 b15zdnd00an1n01x5 FILLER_211_1151 ();
 b15zdnd11an1n32x5 FILLER_211_1191 ();
 b15zdnd11an1n08x5 FILLER_211_1223 ();
 b15zdnd11an1n04x5 FILLER_211_1231 ();
 b15zdnd00an1n02x5 FILLER_211_1235 ();
 b15zdnd11an1n32x5 FILLER_211_1279 ();
 b15zdnd11an1n08x5 FILLER_211_1311 ();
 b15zdnd11an1n04x5 FILLER_211_1319 ();
 b15zdnd11an1n64x5 FILLER_211_1326 ();
 b15zdnd11an1n64x5 FILLER_211_1390 ();
 b15zdnd11an1n32x5 FILLER_211_1454 ();
 b15zdnd11an1n16x5 FILLER_211_1486 ();
 b15zdnd11an1n04x5 FILLER_211_1529 ();
 b15zdnd11an1n64x5 FILLER_211_1539 ();
 b15zdnd00an1n02x5 FILLER_211_1603 ();
 b15zdnd00an1n01x5 FILLER_211_1605 ();
 b15zdnd11an1n04x5 FILLER_211_1609 ();
 b15zdnd11an1n08x5 FILLER_211_1640 ();
 b15zdnd11an1n04x5 FILLER_211_1648 ();
 b15zdnd00an1n02x5 FILLER_211_1652 ();
 b15zdnd00an1n01x5 FILLER_211_1654 ();
 b15zdnd11an1n32x5 FILLER_211_1664 ();
 b15zdnd11an1n08x5 FILLER_211_1696 ();
 b15zdnd11an1n04x5 FILLER_211_1704 ();
 b15zdnd00an1n02x5 FILLER_211_1708 ();
 b15zdnd11an1n16x5 FILLER_211_1719 ();
 b15zdnd11an1n08x5 FILLER_211_1735 ();
 b15zdnd00an1n02x5 FILLER_211_1743 ();
 b15zdnd00an1n01x5 FILLER_211_1745 ();
 b15zdnd11an1n64x5 FILLER_211_1749 ();
 b15zdnd11an1n64x5 FILLER_211_1813 ();
 b15zdnd11an1n64x5 FILLER_211_1877 ();
 b15zdnd11an1n64x5 FILLER_211_1941 ();
 b15zdnd11an1n64x5 FILLER_211_2005 ();
 b15zdnd11an1n64x5 FILLER_211_2069 ();
 b15zdnd11an1n64x5 FILLER_211_2133 ();
 b15zdnd11an1n64x5 FILLER_211_2197 ();
 b15zdnd11an1n16x5 FILLER_211_2261 ();
 b15zdnd11an1n04x5 FILLER_211_2277 ();
 b15zdnd00an1n02x5 FILLER_211_2281 ();
 b15zdnd00an1n01x5 FILLER_211_2283 ();
 b15zdnd11an1n64x5 FILLER_212_8 ();
 b15zdnd11an1n64x5 FILLER_212_72 ();
 b15zdnd11an1n64x5 FILLER_212_136 ();
 b15zdnd11an1n32x5 FILLER_212_200 ();
 b15zdnd11an1n16x5 FILLER_212_232 ();
 b15zdnd00an1n02x5 FILLER_212_248 ();
 b15zdnd11an1n64x5 FILLER_212_257 ();
 b15zdnd11an1n64x5 FILLER_212_321 ();
 b15zdnd11an1n64x5 FILLER_212_385 ();
 b15zdnd11an1n64x5 FILLER_212_449 ();
 b15zdnd11an1n64x5 FILLER_212_513 ();
 b15zdnd00an1n02x5 FILLER_212_577 ();
 b15zdnd11an1n16x5 FILLER_212_593 ();
 b15zdnd11an1n32x5 FILLER_212_612 ();
 b15zdnd11an1n16x5 FILLER_212_644 ();
 b15zdnd11an1n08x5 FILLER_212_660 ();
 b15zdnd11an1n04x5 FILLER_212_668 ();
 b15zdnd00an1n02x5 FILLER_212_672 ();
 b15zdnd00an1n01x5 FILLER_212_674 ();
 b15zdnd11an1n32x5 FILLER_212_686 ();
 b15zdnd11an1n32x5 FILLER_212_726 ();
 b15zdnd11an1n08x5 FILLER_212_758 ();
 b15zdnd00an1n02x5 FILLER_212_766 ();
 b15zdnd00an1n01x5 FILLER_212_768 ();
 b15zdnd11an1n04x5 FILLER_212_772 ();
 b15zdnd11an1n64x5 FILLER_212_779 ();
 b15zdnd11an1n64x5 FILLER_212_843 ();
 b15zdnd11an1n64x5 FILLER_212_907 ();
 b15zdnd11an1n64x5 FILLER_212_971 ();
 b15zdnd11an1n64x5 FILLER_212_1035 ();
 b15zdnd11an1n64x5 FILLER_212_1099 ();
 b15zdnd11an1n32x5 FILLER_212_1163 ();
 b15zdnd11an1n16x5 FILLER_212_1195 ();
 b15zdnd11an1n04x5 FILLER_212_1211 ();
 b15zdnd00an1n01x5 FILLER_212_1215 ();
 b15zdnd11an1n64x5 FILLER_212_1220 ();
 b15zdnd11an1n64x5 FILLER_212_1284 ();
 b15zdnd11an1n64x5 FILLER_212_1348 ();
 b15zdnd11an1n64x5 FILLER_212_1412 ();
 b15zdnd11an1n32x5 FILLER_212_1476 ();
 b15zdnd11an1n08x5 FILLER_212_1508 ();
 b15zdnd00an1n02x5 FILLER_212_1516 ();
 b15zdnd11an1n64x5 FILLER_212_1526 ();
 b15zdnd11an1n32x5 FILLER_212_1590 ();
 b15zdnd11an1n64x5 FILLER_212_1625 ();
 b15zdnd11an1n64x5 FILLER_212_1689 ();
 b15zdnd11an1n64x5 FILLER_212_1753 ();
 b15zdnd11an1n64x5 FILLER_212_1817 ();
 b15zdnd11an1n64x5 FILLER_212_1881 ();
 b15zdnd11an1n64x5 FILLER_212_1945 ();
 b15zdnd11an1n64x5 FILLER_212_2009 ();
 b15zdnd11an1n64x5 FILLER_212_2073 ();
 b15zdnd11an1n16x5 FILLER_212_2137 ();
 b15zdnd00an1n01x5 FILLER_212_2153 ();
 b15zdnd11an1n64x5 FILLER_212_2162 ();
 b15zdnd11an1n32x5 FILLER_212_2226 ();
 b15zdnd11an1n16x5 FILLER_212_2258 ();
 b15zdnd00an1n02x5 FILLER_212_2274 ();
 b15zdnd11an1n64x5 FILLER_213_0 ();
 b15zdnd11an1n64x5 FILLER_213_64 ();
 b15zdnd11an1n16x5 FILLER_213_128 ();
 b15zdnd11an1n16x5 FILLER_213_158 ();
 b15zdnd00an1n01x5 FILLER_213_174 ();
 b15zdnd11an1n64x5 FILLER_213_192 ();
 b15zdnd11an1n64x5 FILLER_213_256 ();
 b15zdnd11an1n64x5 FILLER_213_320 ();
 b15zdnd11an1n16x5 FILLER_213_384 ();
 b15zdnd11an1n08x5 FILLER_213_400 ();
 b15zdnd11an1n04x5 FILLER_213_408 ();
 b15zdnd00an1n02x5 FILLER_213_412 ();
 b15zdnd11an1n64x5 FILLER_213_418 ();
 b15zdnd11an1n64x5 FILLER_213_482 ();
 b15zdnd11an1n32x5 FILLER_213_546 ();
 b15zdnd11an1n04x5 FILLER_213_578 ();
 b15zdnd11an1n04x5 FILLER_213_634 ();
 b15zdnd11an1n64x5 FILLER_213_644 ();
 b15zdnd11an1n64x5 FILLER_213_708 ();
 b15zdnd11an1n64x5 FILLER_213_772 ();
 b15zdnd11an1n64x5 FILLER_213_836 ();
 b15zdnd11an1n64x5 FILLER_213_900 ();
 b15zdnd11an1n64x5 FILLER_213_964 ();
 b15zdnd11an1n64x5 FILLER_213_1028 ();
 b15zdnd11an1n08x5 FILLER_213_1092 ();
 b15zdnd00an1n01x5 FILLER_213_1100 ();
 b15zdnd11an1n32x5 FILLER_213_1108 ();
 b15zdnd11an1n08x5 FILLER_213_1140 ();
 b15zdnd00an1n01x5 FILLER_213_1148 ();
 b15zdnd11an1n64x5 FILLER_213_1201 ();
 b15zdnd11an1n64x5 FILLER_213_1265 ();
 b15zdnd11an1n32x5 FILLER_213_1329 ();
 b15zdnd11an1n16x5 FILLER_213_1361 ();
 b15zdnd11an1n04x5 FILLER_213_1377 ();
 b15zdnd11an1n64x5 FILLER_213_1384 ();
 b15zdnd11an1n64x5 FILLER_213_1448 ();
 b15zdnd11an1n64x5 FILLER_213_1512 ();
 b15zdnd11an1n32x5 FILLER_213_1576 ();
 b15zdnd11an1n08x5 FILLER_213_1608 ();
 b15zdnd11an1n04x5 FILLER_213_1616 ();
 b15zdnd00an1n02x5 FILLER_213_1620 ();
 b15zdnd00an1n01x5 FILLER_213_1622 ();
 b15zdnd11an1n64x5 FILLER_213_1626 ();
 b15zdnd11an1n08x5 FILLER_213_1690 ();
 b15zdnd11an1n04x5 FILLER_213_1698 ();
 b15zdnd11an1n16x5 FILLER_213_1711 ();
 b15zdnd11an1n08x5 FILLER_213_1727 ();
 b15zdnd11an1n04x5 FILLER_213_1735 ();
 b15zdnd00an1n02x5 FILLER_213_1739 ();
 b15zdnd00an1n01x5 FILLER_213_1741 ();
 b15zdnd11an1n64x5 FILLER_213_1794 ();
 b15zdnd11an1n64x5 FILLER_213_1858 ();
 b15zdnd11an1n64x5 FILLER_213_1922 ();
 b15zdnd11an1n64x5 FILLER_213_1986 ();
 b15zdnd11an1n64x5 FILLER_213_2050 ();
 b15zdnd11an1n64x5 FILLER_213_2114 ();
 b15zdnd11an1n64x5 FILLER_213_2178 ();
 b15zdnd11an1n32x5 FILLER_213_2242 ();
 b15zdnd11an1n08x5 FILLER_213_2274 ();
 b15zdnd00an1n02x5 FILLER_213_2282 ();
 b15zdnd11an1n64x5 FILLER_214_8 ();
 b15zdnd11an1n64x5 FILLER_214_72 ();
 b15zdnd11an1n08x5 FILLER_214_136 ();
 b15zdnd11an1n04x5 FILLER_214_144 ();
 b15zdnd00an1n02x5 FILLER_214_148 ();
 b15zdnd00an1n01x5 FILLER_214_150 ();
 b15zdnd11an1n64x5 FILLER_214_158 ();
 b15zdnd11an1n64x5 FILLER_214_222 ();
 b15zdnd11an1n64x5 FILLER_214_286 ();
 b15zdnd11an1n32x5 FILLER_214_350 ();
 b15zdnd11an1n08x5 FILLER_214_382 ();
 b15zdnd11an1n08x5 FILLER_214_401 ();
 b15zdnd00an1n01x5 FILLER_214_409 ();
 b15zdnd11an1n64x5 FILLER_214_417 ();
 b15zdnd11an1n32x5 FILLER_214_481 ();
 b15zdnd11an1n16x5 FILLER_214_513 ();
 b15zdnd11an1n08x5 FILLER_214_529 ();
 b15zdnd11an1n04x5 FILLER_214_537 ();
 b15zdnd11an1n32x5 FILLER_214_568 ();
 b15zdnd11an1n04x5 FILLER_214_603 ();
 b15zdnd11an1n64x5 FILLER_214_610 ();
 b15zdnd11an1n32x5 FILLER_214_674 ();
 b15zdnd11an1n08x5 FILLER_214_706 ();
 b15zdnd11an1n04x5 FILLER_214_714 ();
 b15zdnd11an1n64x5 FILLER_214_726 ();
 b15zdnd11an1n64x5 FILLER_214_790 ();
 b15zdnd11an1n64x5 FILLER_214_854 ();
 b15zdnd11an1n16x5 FILLER_214_918 ();
 b15zdnd11an1n64x5 FILLER_214_937 ();
 b15zdnd11an1n64x5 FILLER_214_1001 ();
 b15zdnd11an1n64x5 FILLER_214_1065 ();
 b15zdnd11an1n32x5 FILLER_214_1129 ();
 b15zdnd11an1n04x5 FILLER_214_1161 ();
 b15zdnd00an1n02x5 FILLER_214_1165 ();
 b15zdnd11an1n04x5 FILLER_214_1170 ();
 b15zdnd11an1n04x5 FILLER_214_1177 ();
 b15zdnd11an1n32x5 FILLER_214_1184 ();
 b15zdnd11an1n16x5 FILLER_214_1216 ();
 b15zdnd00an1n01x5 FILLER_214_1232 ();
 b15zdnd11an1n64x5 FILLER_214_1264 ();
 b15zdnd11an1n16x5 FILLER_214_1328 ();
 b15zdnd11an1n08x5 FILLER_214_1344 ();
 b15zdnd11an1n04x5 FILLER_214_1352 ();
 b15zdnd11an1n64x5 FILLER_214_1384 ();
 b15zdnd11an1n64x5 FILLER_214_1448 ();
 b15zdnd11an1n64x5 FILLER_214_1512 ();
 b15zdnd00an1n02x5 FILLER_214_1576 ();
 b15zdnd11an1n08x5 FILLER_214_1585 ();
 b15zdnd11an1n04x5 FILLER_214_1593 ();
 b15zdnd00an1n01x5 FILLER_214_1597 ();
 b15zdnd11an1n64x5 FILLER_214_1650 ();
 b15zdnd11an1n32x5 FILLER_214_1714 ();
 b15zdnd11an1n16x5 FILLER_214_1746 ();
 b15zdnd00an1n02x5 FILLER_214_1762 ();
 b15zdnd00an1n01x5 FILLER_214_1764 ();
 b15zdnd11an1n04x5 FILLER_214_1768 ();
 b15zdnd11an1n64x5 FILLER_214_1775 ();
 b15zdnd11an1n64x5 FILLER_214_1839 ();
 b15zdnd11an1n64x5 FILLER_214_1903 ();
 b15zdnd11an1n64x5 FILLER_214_1967 ();
 b15zdnd11an1n64x5 FILLER_214_2031 ();
 b15zdnd11an1n32x5 FILLER_214_2095 ();
 b15zdnd11an1n16x5 FILLER_214_2127 ();
 b15zdnd11an1n08x5 FILLER_214_2143 ();
 b15zdnd00an1n02x5 FILLER_214_2151 ();
 b15zdnd00an1n01x5 FILLER_214_2153 ();
 b15zdnd11an1n64x5 FILLER_214_2162 ();
 b15zdnd11an1n32x5 FILLER_214_2226 ();
 b15zdnd11an1n16x5 FILLER_214_2258 ();
 b15zdnd00an1n02x5 FILLER_214_2274 ();
 b15zdnd11an1n64x5 FILLER_215_0 ();
 b15zdnd11an1n16x5 FILLER_215_64 ();
 b15zdnd11an1n04x5 FILLER_215_80 ();
 b15zdnd00an1n01x5 FILLER_215_84 ();
 b15zdnd11an1n32x5 FILLER_215_127 ();
 b15zdnd11an1n04x5 FILLER_215_159 ();
 b15zdnd00an1n01x5 FILLER_215_163 ();
 b15zdnd11an1n16x5 FILLER_215_209 ();
 b15zdnd11an1n08x5 FILLER_215_225 ();
 b15zdnd00an1n01x5 FILLER_215_233 ();
 b15zdnd11an1n64x5 FILLER_215_248 ();
 b15zdnd11an1n64x5 FILLER_215_312 ();
 b15zdnd11an1n16x5 FILLER_215_376 ();
 b15zdnd00an1n02x5 FILLER_215_392 ();
 b15zdnd00an1n01x5 FILLER_215_394 ();
 b15zdnd11an1n64x5 FILLER_215_411 ();
 b15zdnd11an1n16x5 FILLER_215_475 ();
 b15zdnd11an1n04x5 FILLER_215_491 ();
 b15zdnd00an1n02x5 FILLER_215_495 ();
 b15zdnd11an1n16x5 FILLER_215_515 ();
 b15zdnd11an1n08x5 FILLER_215_531 ();
 b15zdnd11an1n04x5 FILLER_215_539 ();
 b15zdnd00an1n02x5 FILLER_215_543 ();
 b15zdnd00an1n01x5 FILLER_215_545 ();
 b15zdnd11an1n04x5 FILLER_215_557 ();
 b15zdnd11an1n64x5 FILLER_215_569 ();
 b15zdnd11an1n32x5 FILLER_215_633 ();
 b15zdnd11an1n04x5 FILLER_215_665 ();
 b15zdnd11an1n64x5 FILLER_215_673 ();
 b15zdnd11an1n16x5 FILLER_215_737 ();
 b15zdnd11an1n08x5 FILLER_215_753 ();
 b15zdnd00an1n01x5 FILLER_215_761 ();
 b15zdnd11an1n04x5 FILLER_215_765 ();
 b15zdnd11an1n04x5 FILLER_215_772 ();
 b15zdnd11an1n04x5 FILLER_215_779 ();
 b15zdnd11an1n64x5 FILLER_215_786 ();
 b15zdnd11an1n32x5 FILLER_215_850 ();
 b15zdnd11an1n16x5 FILLER_215_882 ();
 b15zdnd11an1n08x5 FILLER_215_898 ();
 b15zdnd11an1n04x5 FILLER_215_906 ();
 b15zdnd00an1n01x5 FILLER_215_910 ();
 b15zdnd11an1n04x5 FILLER_215_918 ();
 b15zdnd00an1n01x5 FILLER_215_922 ();
 b15zdnd11an1n04x5 FILLER_215_926 ();
 b15zdnd11an1n04x5 FILLER_215_933 ();
 b15zdnd11an1n04x5 FILLER_215_940 ();
 b15zdnd11an1n64x5 FILLER_215_947 ();
 b15zdnd11an1n64x5 FILLER_215_1011 ();
 b15zdnd11an1n64x5 FILLER_215_1075 ();
 b15zdnd11an1n64x5 FILLER_215_1139 ();
 b15zdnd11an1n64x5 FILLER_215_1203 ();
 b15zdnd11an1n64x5 FILLER_215_1267 ();
 b15zdnd11an1n32x5 FILLER_215_1331 ();
 b15zdnd11an1n08x5 FILLER_215_1363 ();
 b15zdnd11an1n04x5 FILLER_215_1371 ();
 b15zdnd00an1n02x5 FILLER_215_1375 ();
 b15zdnd00an1n01x5 FILLER_215_1377 ();
 b15zdnd11an1n64x5 FILLER_215_1381 ();
 b15zdnd11an1n64x5 FILLER_215_1445 ();
 b15zdnd11an1n64x5 FILLER_215_1509 ();
 b15zdnd11an1n32x5 FILLER_215_1573 ();
 b15zdnd11an1n08x5 FILLER_215_1605 ();
 b15zdnd11an1n04x5 FILLER_215_1613 ();
 b15zdnd00an1n02x5 FILLER_215_1617 ();
 b15zdnd00an1n01x5 FILLER_215_1619 ();
 b15zdnd11an1n64x5 FILLER_215_1627 ();
 b15zdnd11an1n64x5 FILLER_215_1691 ();
 b15zdnd11an1n08x5 FILLER_215_1755 ();
 b15zdnd00an1n02x5 FILLER_215_1763 ();
 b15zdnd11an1n64x5 FILLER_215_1768 ();
 b15zdnd11an1n64x5 FILLER_215_1832 ();
 b15zdnd11an1n64x5 FILLER_215_1896 ();
 b15zdnd11an1n64x5 FILLER_215_1960 ();
 b15zdnd11an1n64x5 FILLER_215_2024 ();
 b15zdnd11an1n64x5 FILLER_215_2088 ();
 b15zdnd11an1n64x5 FILLER_215_2152 ();
 b15zdnd11an1n64x5 FILLER_215_2216 ();
 b15zdnd11an1n04x5 FILLER_215_2280 ();
 b15zdnd11an1n64x5 FILLER_216_8 ();
 b15zdnd11an1n64x5 FILLER_216_72 ();
 b15zdnd11an1n64x5 FILLER_216_136 ();
 b15zdnd11an1n08x5 FILLER_216_200 ();
 b15zdnd11an1n64x5 FILLER_216_228 ();
 b15zdnd11an1n16x5 FILLER_216_292 ();
 b15zdnd11an1n04x5 FILLER_216_308 ();
 b15zdnd00an1n02x5 FILLER_216_312 ();
 b15zdnd11an1n32x5 FILLER_216_325 ();
 b15zdnd11an1n16x5 FILLER_216_357 ();
 b15zdnd11an1n04x5 FILLER_216_373 ();
 b15zdnd11an1n04x5 FILLER_216_382 ();
 b15zdnd11an1n08x5 FILLER_216_391 ();
 b15zdnd00an1n02x5 FILLER_216_399 ();
 b15zdnd11an1n64x5 FILLER_216_443 ();
 b15zdnd11an1n64x5 FILLER_216_507 ();
 b15zdnd11an1n64x5 FILLER_216_571 ();
 b15zdnd11an1n64x5 FILLER_216_635 ();
 b15zdnd11an1n16x5 FILLER_216_699 ();
 b15zdnd00an1n02x5 FILLER_216_715 ();
 b15zdnd00an1n01x5 FILLER_216_717 ();
 b15zdnd11an1n08x5 FILLER_216_726 ();
 b15zdnd11an1n08x5 FILLER_216_741 ();
 b15zdnd11an1n16x5 FILLER_216_801 ();
 b15zdnd11an1n04x5 FILLER_216_817 ();
 b15zdnd11an1n32x5 FILLER_216_830 ();
 b15zdnd11an1n08x5 FILLER_216_862 ();
 b15zdnd11an1n04x5 FILLER_216_870 ();
 b15zdnd00an1n02x5 FILLER_216_874 ();
 b15zdnd00an1n01x5 FILLER_216_876 ();
 b15zdnd11an1n08x5 FILLER_216_886 ();
 b15zdnd11an1n04x5 FILLER_216_894 ();
 b15zdnd00an1n01x5 FILLER_216_898 ();
 b15zdnd11an1n04x5 FILLER_216_906 ();
 b15zdnd11an1n64x5 FILLER_216_962 ();
 b15zdnd11an1n64x5 FILLER_216_1026 ();
 b15zdnd11an1n64x5 FILLER_216_1090 ();
 b15zdnd11an1n32x5 FILLER_216_1154 ();
 b15zdnd11an1n08x5 FILLER_216_1186 ();
 b15zdnd00an1n02x5 FILLER_216_1194 ();
 b15zdnd11an1n04x5 FILLER_216_1199 ();
 b15zdnd11an1n64x5 FILLER_216_1206 ();
 b15zdnd11an1n64x5 FILLER_216_1270 ();
 b15zdnd11an1n64x5 FILLER_216_1334 ();
 b15zdnd11an1n64x5 FILLER_216_1398 ();
 b15zdnd11an1n64x5 FILLER_216_1462 ();
 b15zdnd11an1n04x5 FILLER_216_1526 ();
 b15zdnd00an1n01x5 FILLER_216_1530 ();
 b15zdnd11an1n64x5 FILLER_216_1535 ();
 b15zdnd11an1n16x5 FILLER_216_1599 ();
 b15zdnd11an1n04x5 FILLER_216_1615 ();
 b15zdnd00an1n01x5 FILLER_216_1619 ();
 b15zdnd11an1n08x5 FILLER_216_1623 ();
 b15zdnd11an1n04x5 FILLER_216_1631 ();
 b15zdnd00an1n01x5 FILLER_216_1635 ();
 b15zdnd11an1n64x5 FILLER_216_1643 ();
 b15zdnd11an1n64x5 FILLER_216_1707 ();
 b15zdnd11an1n32x5 FILLER_216_1771 ();
 b15zdnd11an1n08x5 FILLER_216_1803 ();
 b15zdnd11an1n04x5 FILLER_216_1811 ();
 b15zdnd00an1n02x5 FILLER_216_1815 ();
 b15zdnd11an1n64x5 FILLER_216_1824 ();
 b15zdnd11an1n64x5 FILLER_216_1888 ();
 b15zdnd11an1n64x5 FILLER_216_1952 ();
 b15zdnd11an1n64x5 FILLER_216_2016 ();
 b15zdnd11an1n64x5 FILLER_216_2080 ();
 b15zdnd11an1n08x5 FILLER_216_2144 ();
 b15zdnd00an1n02x5 FILLER_216_2152 ();
 b15zdnd11an1n64x5 FILLER_216_2162 ();
 b15zdnd11an1n32x5 FILLER_216_2226 ();
 b15zdnd11an1n16x5 FILLER_216_2258 ();
 b15zdnd00an1n02x5 FILLER_216_2274 ();
 b15zdnd11an1n64x5 FILLER_217_0 ();
 b15zdnd11an1n64x5 FILLER_217_64 ();
 b15zdnd11an1n04x5 FILLER_217_128 ();
 b15zdnd00an1n02x5 FILLER_217_132 ();
 b15zdnd00an1n01x5 FILLER_217_134 ();
 b15zdnd11an1n64x5 FILLER_217_157 ();
 b15zdnd11an1n64x5 FILLER_217_221 ();
 b15zdnd11an1n16x5 FILLER_217_285 ();
 b15zdnd00an1n02x5 FILLER_217_301 ();
 b15zdnd11an1n32x5 FILLER_217_313 ();
 b15zdnd11an1n04x5 FILLER_217_345 ();
 b15zdnd00an1n02x5 FILLER_217_349 ();
 b15zdnd00an1n01x5 FILLER_217_351 ();
 b15zdnd11an1n04x5 FILLER_217_404 ();
 b15zdnd11an1n64x5 FILLER_217_417 ();
 b15zdnd11an1n32x5 FILLER_217_481 ();
 b15zdnd11an1n16x5 FILLER_217_513 ();
 b15zdnd00an1n02x5 FILLER_217_529 ();
 b15zdnd11an1n64x5 FILLER_217_535 ();
 b15zdnd11an1n64x5 FILLER_217_599 ();
 b15zdnd11an1n64x5 FILLER_217_663 ();
 b15zdnd11an1n08x5 FILLER_217_727 ();
 b15zdnd11an1n04x5 FILLER_217_735 ();
 b15zdnd11an1n04x5 FILLER_217_745 ();
 b15zdnd11an1n08x5 FILLER_217_791 ();
 b15zdnd00an1n01x5 FILLER_217_799 ();
 b15zdnd11an1n16x5 FILLER_217_842 ();
 b15zdnd00an1n02x5 FILLER_217_858 ();
 b15zdnd00an1n01x5 FILLER_217_860 ();
 b15zdnd11an1n32x5 FILLER_217_870 ();
 b15zdnd11an1n04x5 FILLER_217_902 ();
 b15zdnd00an1n02x5 FILLER_217_906 ();
 b15zdnd00an1n01x5 FILLER_217_908 ();
 b15zdnd11an1n04x5 FILLER_217_961 ();
 b15zdnd11an1n32x5 FILLER_217_972 ();
 b15zdnd11an1n16x5 FILLER_217_1004 ();
 b15zdnd11an1n04x5 FILLER_217_1020 ();
 b15zdnd11an1n64x5 FILLER_217_1066 ();
 b15zdnd11an1n32x5 FILLER_217_1130 ();
 b15zdnd11an1n16x5 FILLER_217_1162 ();
 b15zdnd11an1n64x5 FILLER_217_1230 ();
 b15zdnd11an1n64x5 FILLER_217_1294 ();
 b15zdnd11an1n64x5 FILLER_217_1358 ();
 b15zdnd11an1n64x5 FILLER_217_1422 ();
 b15zdnd11an1n64x5 FILLER_217_1486 ();
 b15zdnd11an1n64x5 FILLER_217_1550 ();
 b15zdnd11an1n04x5 FILLER_217_1614 ();
 b15zdnd00an1n02x5 FILLER_217_1618 ();
 b15zdnd11an1n04x5 FILLER_217_1623 ();
 b15zdnd11an1n64x5 FILLER_217_1630 ();
 b15zdnd11an1n64x5 FILLER_217_1694 ();
 b15zdnd11an1n64x5 FILLER_217_1758 ();
 b15zdnd11an1n64x5 FILLER_217_1822 ();
 b15zdnd11an1n64x5 FILLER_217_1886 ();
 b15zdnd11an1n64x5 FILLER_217_1950 ();
 b15zdnd11an1n64x5 FILLER_217_2014 ();
 b15zdnd11an1n64x5 FILLER_217_2078 ();
 b15zdnd11an1n64x5 FILLER_217_2142 ();
 b15zdnd11an1n64x5 FILLER_217_2206 ();
 b15zdnd11an1n08x5 FILLER_217_2270 ();
 b15zdnd11an1n04x5 FILLER_217_2278 ();
 b15zdnd00an1n02x5 FILLER_217_2282 ();
 b15zdnd11an1n64x5 FILLER_218_8 ();
 b15zdnd11an1n64x5 FILLER_218_72 ();
 b15zdnd11an1n64x5 FILLER_218_136 ();
 b15zdnd11an1n64x5 FILLER_218_200 ();
 b15zdnd11an1n64x5 FILLER_218_264 ();
 b15zdnd11an1n32x5 FILLER_218_328 ();
 b15zdnd11an1n08x5 FILLER_218_360 ();
 b15zdnd00an1n01x5 FILLER_218_368 ();
 b15zdnd11an1n04x5 FILLER_218_372 ();
 b15zdnd11an1n04x5 FILLER_218_379 ();
 b15zdnd11an1n04x5 FILLER_218_390 ();
 b15zdnd11an1n64x5 FILLER_218_436 ();
 b15zdnd11an1n64x5 FILLER_218_500 ();
 b15zdnd11an1n64x5 FILLER_218_564 ();
 b15zdnd11an1n32x5 FILLER_218_628 ();
 b15zdnd11an1n08x5 FILLER_218_660 ();
 b15zdnd00an1n01x5 FILLER_218_668 ();
 b15zdnd11an1n32x5 FILLER_218_673 ();
 b15zdnd11an1n08x5 FILLER_218_705 ();
 b15zdnd11an1n04x5 FILLER_218_713 ();
 b15zdnd00an1n01x5 FILLER_218_717 ();
 b15zdnd11an1n16x5 FILLER_218_726 ();
 b15zdnd00an1n01x5 FILLER_218_742 ();
 b15zdnd11an1n04x5 FILLER_218_785 ();
 b15zdnd11an1n04x5 FILLER_218_792 ();
 b15zdnd00an1n02x5 FILLER_218_796 ();
 b15zdnd00an1n01x5 FILLER_218_798 ();
 b15zdnd11an1n04x5 FILLER_218_806 ();
 b15zdnd11an1n64x5 FILLER_218_813 ();
 b15zdnd11an1n16x5 FILLER_218_877 ();
 b15zdnd11an1n08x5 FILLER_218_893 ();
 b15zdnd11an1n04x5 FILLER_218_901 ();
 b15zdnd00an1n01x5 FILLER_218_905 ();
 b15zdnd11an1n64x5 FILLER_218_958 ();
 b15zdnd11an1n64x5 FILLER_218_1022 ();
 b15zdnd11an1n64x5 FILLER_218_1086 ();
 b15zdnd11an1n32x5 FILLER_218_1150 ();
 b15zdnd11an1n16x5 FILLER_218_1182 ();
 b15zdnd11an1n04x5 FILLER_218_1198 ();
 b15zdnd00an1n01x5 FILLER_218_1202 ();
 b15zdnd11an1n64x5 FILLER_218_1206 ();
 b15zdnd11an1n64x5 FILLER_218_1270 ();
 b15zdnd11an1n64x5 FILLER_218_1334 ();
 b15zdnd11an1n64x5 FILLER_218_1398 ();
 b15zdnd11an1n64x5 FILLER_218_1462 ();
 b15zdnd11an1n64x5 FILLER_218_1526 ();
 b15zdnd11an1n08x5 FILLER_218_1590 ();
 b15zdnd11an1n04x5 FILLER_218_1598 ();
 b15zdnd11an1n64x5 FILLER_218_1654 ();
 b15zdnd11an1n08x5 FILLER_218_1718 ();
 b15zdnd00an1n02x5 FILLER_218_1726 ();
 b15zdnd00an1n01x5 FILLER_218_1728 ();
 b15zdnd11an1n08x5 FILLER_218_1735 ();
 b15zdnd11an1n04x5 FILLER_218_1743 ();
 b15zdnd00an1n02x5 FILLER_218_1747 ();
 b15zdnd11an1n04x5 FILLER_218_1752 ();
 b15zdnd00an1n01x5 FILLER_218_1756 ();
 b15zdnd11an1n64x5 FILLER_218_1760 ();
 b15zdnd11an1n64x5 FILLER_218_1824 ();
 b15zdnd11an1n08x5 FILLER_218_1888 ();
 b15zdnd11an1n04x5 FILLER_218_1896 ();
 b15zdnd11an1n64x5 FILLER_218_1903 ();
 b15zdnd11an1n64x5 FILLER_218_1967 ();
 b15zdnd11an1n64x5 FILLER_218_2031 ();
 b15zdnd11an1n32x5 FILLER_218_2095 ();
 b15zdnd11an1n16x5 FILLER_218_2127 ();
 b15zdnd11an1n08x5 FILLER_218_2143 ();
 b15zdnd00an1n02x5 FILLER_218_2151 ();
 b15zdnd00an1n01x5 FILLER_218_2153 ();
 b15zdnd11an1n64x5 FILLER_218_2162 ();
 b15zdnd11an1n32x5 FILLER_218_2226 ();
 b15zdnd11an1n16x5 FILLER_218_2258 ();
 b15zdnd00an1n02x5 FILLER_218_2274 ();
 b15zdnd11an1n64x5 FILLER_219_0 ();
 b15zdnd11an1n64x5 FILLER_219_64 ();
 b15zdnd11an1n64x5 FILLER_219_128 ();
 b15zdnd11an1n32x5 FILLER_219_192 ();
 b15zdnd11an1n16x5 FILLER_219_224 ();
 b15zdnd11an1n08x5 FILLER_219_240 ();
 b15zdnd11an1n64x5 FILLER_219_255 ();
 b15zdnd11an1n32x5 FILLER_219_319 ();
 b15zdnd11an1n16x5 FILLER_219_351 ();
 b15zdnd00an1n02x5 FILLER_219_367 ();
 b15zdnd00an1n01x5 FILLER_219_369 ();
 b15zdnd11an1n04x5 FILLER_219_373 ();
 b15zdnd11an1n04x5 FILLER_219_381 ();
 b15zdnd11an1n64x5 FILLER_219_427 ();
 b15zdnd11an1n16x5 FILLER_219_491 ();
 b15zdnd00an1n02x5 FILLER_219_507 ();
 b15zdnd00an1n01x5 FILLER_219_509 ();
 b15zdnd11an1n64x5 FILLER_219_513 ();
 b15zdnd11an1n64x5 FILLER_219_577 ();
 b15zdnd11an1n64x5 FILLER_219_641 ();
 b15zdnd11an1n32x5 FILLER_219_705 ();
 b15zdnd11an1n16x5 FILLER_219_737 ();
 b15zdnd11an1n04x5 FILLER_219_753 ();
 b15zdnd00an1n02x5 FILLER_219_757 ();
 b15zdnd00an1n01x5 FILLER_219_759 ();
 b15zdnd11an1n04x5 FILLER_219_812 ();
 b15zdnd11an1n64x5 FILLER_219_822 ();
 b15zdnd11an1n16x5 FILLER_219_886 ();
 b15zdnd11an1n04x5 FILLER_219_902 ();
 b15zdnd00an1n02x5 FILLER_219_906 ();
 b15zdnd00an1n01x5 FILLER_219_908 ();
 b15zdnd11an1n04x5 FILLER_219_936 ();
 b15zdnd11an1n04x5 FILLER_219_943 ();
 b15zdnd11an1n64x5 FILLER_219_950 ();
 b15zdnd11an1n64x5 FILLER_219_1014 ();
 b15zdnd11an1n64x5 FILLER_219_1078 ();
 b15zdnd11an1n64x5 FILLER_219_1142 ();
 b15zdnd11an1n64x5 FILLER_219_1206 ();
 b15zdnd11an1n64x5 FILLER_219_1270 ();
 b15zdnd11an1n16x5 FILLER_219_1334 ();
 b15zdnd11an1n08x5 FILLER_219_1350 ();
 b15zdnd00an1n02x5 FILLER_219_1358 ();
 b15zdnd00an1n01x5 FILLER_219_1360 ();
 b15zdnd11an1n32x5 FILLER_219_1403 ();
 b15zdnd11an1n16x5 FILLER_219_1435 ();
 b15zdnd11an1n04x5 FILLER_219_1451 ();
 b15zdnd00an1n02x5 FILLER_219_1455 ();
 b15zdnd00an1n01x5 FILLER_219_1457 ();
 b15zdnd11an1n04x5 FILLER_219_1461 ();
 b15zdnd11an1n04x5 FILLER_219_1468 ();
 b15zdnd11an1n16x5 FILLER_219_1475 ();
 b15zdnd11an1n08x5 FILLER_219_1491 ();
 b15zdnd11an1n04x5 FILLER_219_1499 ();
 b15zdnd00an1n02x5 FILLER_219_1503 ();
 b15zdnd00an1n01x5 FILLER_219_1505 ();
 b15zdnd11an1n64x5 FILLER_219_1548 ();
 b15zdnd11an1n08x5 FILLER_219_1612 ();
 b15zdnd11an1n04x5 FILLER_219_1620 ();
 b15zdnd00an1n02x5 FILLER_219_1624 ();
 b15zdnd00an1n01x5 FILLER_219_1626 ();
 b15zdnd11an1n64x5 FILLER_219_1630 ();
 b15zdnd11an1n16x5 FILLER_219_1694 ();
 b15zdnd11an1n08x5 FILLER_219_1710 ();
 b15zdnd11an1n04x5 FILLER_219_1718 ();
 b15zdnd00an1n02x5 FILLER_219_1722 ();
 b15zdnd00an1n01x5 FILLER_219_1724 ();
 b15zdnd11an1n64x5 FILLER_219_1777 ();
 b15zdnd11an1n32x5 FILLER_219_1841 ();
 b15zdnd11an1n16x5 FILLER_219_1873 ();
 b15zdnd11an1n08x5 FILLER_219_1889 ();
 b15zdnd00an1n02x5 FILLER_219_1897 ();
 b15zdnd11an1n64x5 FILLER_219_1902 ();
 b15zdnd11an1n64x5 FILLER_219_1966 ();
 b15zdnd11an1n64x5 FILLER_219_2030 ();
 b15zdnd11an1n64x5 FILLER_219_2094 ();
 b15zdnd11an1n32x5 FILLER_219_2158 ();
 b15zdnd11an1n16x5 FILLER_219_2190 ();
 b15zdnd11an1n04x5 FILLER_219_2206 ();
 b15zdnd00an1n02x5 FILLER_219_2210 ();
 b15zdnd00an1n01x5 FILLER_219_2212 ();
 b15zdnd11an1n16x5 FILLER_219_2216 ();
 b15zdnd11an1n08x5 FILLER_219_2232 ();
 b15zdnd11an1n04x5 FILLER_219_2240 ();
 b15zdnd00an1n02x5 FILLER_219_2244 ();
 b15zdnd11an1n32x5 FILLER_219_2250 ();
 b15zdnd00an1n02x5 FILLER_219_2282 ();
 b15zdnd11an1n16x5 FILLER_220_8 ();
 b15zdnd00an1n01x5 FILLER_220_24 ();
 b15zdnd11an1n64x5 FILLER_220_29 ();
 b15zdnd11an1n64x5 FILLER_220_93 ();
 b15zdnd11an1n32x5 FILLER_220_157 ();
 b15zdnd11an1n16x5 FILLER_220_189 ();
 b15zdnd11an1n04x5 FILLER_220_205 ();
 b15zdnd00an1n02x5 FILLER_220_209 ();
 b15zdnd00an1n01x5 FILLER_220_211 ();
 b15zdnd11an1n64x5 FILLER_220_220 ();
 b15zdnd11an1n64x5 FILLER_220_284 ();
 b15zdnd11an1n32x5 FILLER_220_348 ();
 b15zdnd11an1n08x5 FILLER_220_380 ();
 b15zdnd11an1n64x5 FILLER_220_391 ();
 b15zdnd11an1n16x5 FILLER_220_455 ();
 b15zdnd11an1n08x5 FILLER_220_471 ();
 b15zdnd11an1n04x5 FILLER_220_479 ();
 b15zdnd11an1n64x5 FILLER_220_535 ();
 b15zdnd11an1n64x5 FILLER_220_599 ();
 b15zdnd11an1n32x5 FILLER_220_663 ();
 b15zdnd11an1n16x5 FILLER_220_695 ();
 b15zdnd11an1n04x5 FILLER_220_711 ();
 b15zdnd00an1n02x5 FILLER_220_715 ();
 b15zdnd00an1n01x5 FILLER_220_717 ();
 b15zdnd11an1n16x5 FILLER_220_726 ();
 b15zdnd11an1n04x5 FILLER_220_742 ();
 b15zdnd00an1n01x5 FILLER_220_746 ();
 b15zdnd11an1n08x5 FILLER_220_799 ();
 b15zdnd11an1n04x5 FILLER_220_807 ();
 b15zdnd11an1n32x5 FILLER_220_853 ();
 b15zdnd11an1n16x5 FILLER_220_885 ();
 b15zdnd11an1n04x5 FILLER_220_901 ();
 b15zdnd00an1n02x5 FILLER_220_905 ();
 b15zdnd00an1n01x5 FILLER_220_907 ();
 b15zdnd11an1n16x5 FILLER_220_911 ();
 b15zdnd00an1n01x5 FILLER_220_927 ();
 b15zdnd11an1n04x5 FILLER_220_931 ();
 b15zdnd11an1n64x5 FILLER_220_938 ();
 b15zdnd11an1n64x5 FILLER_220_1002 ();
 b15zdnd11an1n64x5 FILLER_220_1066 ();
 b15zdnd11an1n64x5 FILLER_220_1130 ();
 b15zdnd11an1n64x5 FILLER_220_1194 ();
 b15zdnd11an1n64x5 FILLER_220_1258 ();
 b15zdnd11an1n64x5 FILLER_220_1322 ();
 b15zdnd11an1n32x5 FILLER_220_1386 ();
 b15zdnd11an1n16x5 FILLER_220_1418 ();
 b15zdnd11an1n04x5 FILLER_220_1434 ();
 b15zdnd00an1n01x5 FILLER_220_1438 ();
 b15zdnd11an1n64x5 FILLER_220_1491 ();
 b15zdnd11an1n32x5 FILLER_220_1555 ();
 b15zdnd11an1n16x5 FILLER_220_1587 ();
 b15zdnd00an1n01x5 FILLER_220_1603 ();
 b15zdnd11an1n64x5 FILLER_220_1611 ();
 b15zdnd11an1n64x5 FILLER_220_1675 ();
 b15zdnd11an1n08x5 FILLER_220_1739 ();
 b15zdnd00an1n02x5 FILLER_220_1747 ();
 b15zdnd00an1n01x5 FILLER_220_1749 ();
 b15zdnd11an1n32x5 FILLER_220_1753 ();
 b15zdnd11an1n04x5 FILLER_220_1785 ();
 b15zdnd00an1n02x5 FILLER_220_1789 ();
 b15zdnd00an1n01x5 FILLER_220_1791 ();
 b15zdnd11an1n64x5 FILLER_220_1799 ();
 b15zdnd11an1n08x5 FILLER_220_1863 ();
 b15zdnd00an1n02x5 FILLER_220_1871 ();
 b15zdnd00an1n01x5 FILLER_220_1873 ();
 b15zdnd11an1n64x5 FILLER_220_1926 ();
 b15zdnd11an1n64x5 FILLER_220_1990 ();
 b15zdnd11an1n64x5 FILLER_220_2054 ();
 b15zdnd11an1n32x5 FILLER_220_2118 ();
 b15zdnd11an1n04x5 FILLER_220_2150 ();
 b15zdnd11an1n64x5 FILLER_220_2162 ();
 b15zdnd11an1n08x5 FILLER_220_2226 ();
 b15zdnd11an1n04x5 FILLER_220_2234 ();
 b15zdnd11an1n32x5 FILLER_220_2242 ();
 b15zdnd00an1n02x5 FILLER_220_2274 ();
 b15zdnd11an1n64x5 FILLER_221_0 ();
 b15zdnd11an1n64x5 FILLER_221_64 ();
 b15zdnd11an1n64x5 FILLER_221_128 ();
 b15zdnd11an1n64x5 FILLER_221_192 ();
 b15zdnd11an1n32x5 FILLER_221_256 ();
 b15zdnd11an1n16x5 FILLER_221_288 ();
 b15zdnd11an1n08x5 FILLER_221_304 ();
 b15zdnd11an1n04x5 FILLER_221_312 ();
 b15zdnd00an1n02x5 FILLER_221_316 ();
 b15zdnd11an1n64x5 FILLER_221_358 ();
 b15zdnd11an1n64x5 FILLER_221_422 ();
 b15zdnd11an1n08x5 FILLER_221_486 ();
 b15zdnd11an1n04x5 FILLER_221_494 ();
 b15zdnd00an1n02x5 FILLER_221_498 ();
 b15zdnd00an1n01x5 FILLER_221_500 ();
 b15zdnd11an1n04x5 FILLER_221_504 ();
 b15zdnd11an1n64x5 FILLER_221_511 ();
 b15zdnd11an1n64x5 FILLER_221_575 ();
 b15zdnd11an1n64x5 FILLER_221_639 ();
 b15zdnd11an1n32x5 FILLER_221_703 ();
 b15zdnd11an1n16x5 FILLER_221_735 ();
 b15zdnd11an1n08x5 FILLER_221_751 ();
 b15zdnd00an1n02x5 FILLER_221_759 ();
 b15zdnd00an1n01x5 FILLER_221_761 ();
 b15zdnd11an1n04x5 FILLER_221_769 ();
 b15zdnd11an1n08x5 FILLER_221_776 ();
 b15zdnd00an1n01x5 FILLER_221_784 ();
 b15zdnd11an1n64x5 FILLER_221_837 ();
 b15zdnd11an1n64x5 FILLER_221_901 ();
 b15zdnd11an1n64x5 FILLER_221_965 ();
 b15zdnd11an1n64x5 FILLER_221_1029 ();
 b15zdnd11an1n64x5 FILLER_221_1093 ();
 b15zdnd11an1n64x5 FILLER_221_1157 ();
 b15zdnd11an1n64x5 FILLER_221_1221 ();
 b15zdnd11an1n64x5 FILLER_221_1285 ();
 b15zdnd11an1n64x5 FILLER_221_1349 ();
 b15zdnd11an1n64x5 FILLER_221_1413 ();
 b15zdnd11an1n64x5 FILLER_221_1477 ();
 b15zdnd11an1n64x5 FILLER_221_1541 ();
 b15zdnd11an1n64x5 FILLER_221_1605 ();
 b15zdnd11an1n64x5 FILLER_221_1669 ();
 b15zdnd11an1n64x5 FILLER_221_1733 ();
 b15zdnd11an1n64x5 FILLER_221_1797 ();
 b15zdnd11an1n32x5 FILLER_221_1861 ();
 b15zdnd11an1n04x5 FILLER_221_1893 ();
 b15zdnd00an1n02x5 FILLER_221_1897 ();
 b15zdnd00an1n01x5 FILLER_221_1899 ();
 b15zdnd11an1n64x5 FILLER_221_1903 ();
 b15zdnd11an1n64x5 FILLER_221_1967 ();
 b15zdnd11an1n64x5 FILLER_221_2031 ();
 b15zdnd11an1n64x5 FILLER_221_2095 ();
 b15zdnd00an1n02x5 FILLER_221_2159 ();
 b15zdnd00an1n01x5 FILLER_221_2161 ();
 b15zdnd11an1n16x5 FILLER_221_2168 ();
 b15zdnd11an1n08x5 FILLER_221_2184 ();
 b15zdnd00an1n02x5 FILLER_221_2192 ();
 b15zdnd00an1n01x5 FILLER_221_2194 ();
 b15zdnd11an1n16x5 FILLER_221_2198 ();
 b15zdnd11an1n04x5 FILLER_221_2214 ();
 b15zdnd11an1n16x5 FILLER_221_2221 ();
 b15zdnd11an1n04x5 FILLER_221_2237 ();
 b15zdnd00an1n01x5 FILLER_221_2241 ();
 b15zdnd11an1n16x5 FILLER_221_2254 ();
 b15zdnd11an1n08x5 FILLER_221_2270 ();
 b15zdnd11an1n04x5 FILLER_221_2278 ();
 b15zdnd00an1n02x5 FILLER_221_2282 ();
 b15zdnd11an1n64x5 FILLER_222_8 ();
 b15zdnd11an1n64x5 FILLER_222_72 ();
 b15zdnd11an1n64x5 FILLER_222_136 ();
 b15zdnd11an1n64x5 FILLER_222_200 ();
 b15zdnd11an1n64x5 FILLER_222_264 ();
 b15zdnd11an1n16x5 FILLER_222_328 ();
 b15zdnd11an1n04x5 FILLER_222_344 ();
 b15zdnd00an1n02x5 FILLER_222_348 ();
 b15zdnd11an1n04x5 FILLER_222_353 ();
 b15zdnd11an1n16x5 FILLER_222_360 ();
 b15zdnd11an1n08x5 FILLER_222_376 ();
 b15zdnd11an1n04x5 FILLER_222_384 ();
 b15zdnd00an1n02x5 FILLER_222_388 ();
 b15zdnd00an1n01x5 FILLER_222_390 ();
 b15zdnd11an1n64x5 FILLER_222_399 ();
 b15zdnd11an1n64x5 FILLER_222_463 ();
 b15zdnd11an1n64x5 FILLER_222_527 ();
 b15zdnd11an1n32x5 FILLER_222_591 ();
 b15zdnd11an1n08x5 FILLER_222_623 ();
 b15zdnd00an1n02x5 FILLER_222_631 ();
 b15zdnd00an1n01x5 FILLER_222_633 ();
 b15zdnd11an1n32x5 FILLER_222_661 ();
 b15zdnd11an1n16x5 FILLER_222_693 ();
 b15zdnd11an1n08x5 FILLER_222_709 ();
 b15zdnd00an1n01x5 FILLER_222_717 ();
 b15zdnd11an1n32x5 FILLER_222_726 ();
 b15zdnd11an1n04x5 FILLER_222_758 ();
 b15zdnd00an1n01x5 FILLER_222_762 ();
 b15zdnd11an1n04x5 FILLER_222_805 ();
 b15zdnd00an1n01x5 FILLER_222_809 ();
 b15zdnd11an1n64x5 FILLER_222_852 ();
 b15zdnd11an1n64x5 FILLER_222_916 ();
 b15zdnd11an1n64x5 FILLER_222_980 ();
 b15zdnd11an1n64x5 FILLER_222_1044 ();
 b15zdnd11an1n64x5 FILLER_222_1108 ();
 b15zdnd11an1n64x5 FILLER_222_1172 ();
 b15zdnd11an1n64x5 FILLER_222_1236 ();
 b15zdnd11an1n64x5 FILLER_222_1300 ();
 b15zdnd11an1n04x5 FILLER_222_1364 ();
 b15zdnd00an1n01x5 FILLER_222_1368 ();
 b15zdnd11an1n32x5 FILLER_222_1372 ();
 b15zdnd11an1n16x5 FILLER_222_1404 ();
 b15zdnd11an1n08x5 FILLER_222_1420 ();
 b15zdnd00an1n02x5 FILLER_222_1428 ();
 b15zdnd00an1n01x5 FILLER_222_1430 ();
 b15zdnd11an1n64x5 FILLER_222_1473 ();
 b15zdnd11an1n64x5 FILLER_222_1537 ();
 b15zdnd11an1n64x5 FILLER_222_1601 ();
 b15zdnd11an1n64x5 FILLER_222_1665 ();
 b15zdnd11an1n64x5 FILLER_222_1729 ();
 b15zdnd11an1n64x5 FILLER_222_1793 ();
 b15zdnd11an1n64x5 FILLER_222_1857 ();
 b15zdnd11an1n64x5 FILLER_222_1921 ();
 b15zdnd11an1n64x5 FILLER_222_1985 ();
 b15zdnd11an1n32x5 FILLER_222_2049 ();
 b15zdnd11an1n16x5 FILLER_222_2081 ();
 b15zdnd11an1n04x5 FILLER_222_2097 ();
 b15zdnd00an1n01x5 FILLER_222_2101 ();
 b15zdnd11an1n32x5 FILLER_222_2106 ();
 b15zdnd11an1n16x5 FILLER_222_2138 ();
 b15zdnd11an1n16x5 FILLER_222_2162 ();
 b15zdnd11an1n08x5 FILLER_222_2178 ();
 b15zdnd00an1n02x5 FILLER_222_2186 ();
 b15zdnd11an1n04x5 FILLER_222_2240 ();
 b15zdnd11an1n04x5 FILLER_222_2258 ();
 b15zdnd11an1n04x5 FILLER_222_2270 ();
 b15zdnd00an1n02x5 FILLER_222_2274 ();
 b15zdnd11an1n64x5 FILLER_223_0 ();
 b15zdnd11an1n64x5 FILLER_223_64 ();
 b15zdnd11an1n64x5 FILLER_223_128 ();
 b15zdnd11an1n08x5 FILLER_223_192 ();
 b15zdnd00an1n01x5 FILLER_223_200 ();
 b15zdnd11an1n64x5 FILLER_223_204 ();
 b15zdnd11an1n64x5 FILLER_223_268 ();
 b15zdnd11an1n64x5 FILLER_223_332 ();
 b15zdnd11an1n64x5 FILLER_223_396 ();
 b15zdnd11an1n64x5 FILLER_223_460 ();
 b15zdnd11an1n64x5 FILLER_223_524 ();
 b15zdnd11an1n64x5 FILLER_223_588 ();
 b15zdnd11an1n64x5 FILLER_223_652 ();
 b15zdnd11an1n32x5 FILLER_223_716 ();
 b15zdnd11an1n16x5 FILLER_223_748 ();
 b15zdnd00an1n01x5 FILLER_223_764 ();
 b15zdnd11an1n04x5 FILLER_223_768 ();
 b15zdnd11an1n08x5 FILLER_223_775 ();
 b15zdnd11an1n04x5 FILLER_223_783 ();
 b15zdnd11an1n04x5 FILLER_223_795 ();
 b15zdnd00an1n02x5 FILLER_223_799 ();
 b15zdnd11an1n04x5 FILLER_223_804 ();
 b15zdnd11an1n08x5 FILLER_223_811 ();
 b15zdnd00an1n02x5 FILLER_223_819 ();
 b15zdnd11an1n04x5 FILLER_223_828 ();
 b15zdnd00an1n02x5 FILLER_223_832 ();
 b15zdnd00an1n01x5 FILLER_223_834 ();
 b15zdnd11an1n64x5 FILLER_223_842 ();
 b15zdnd11an1n64x5 FILLER_223_906 ();
 b15zdnd11an1n64x5 FILLER_223_970 ();
 b15zdnd11an1n64x5 FILLER_223_1034 ();
 b15zdnd11an1n64x5 FILLER_223_1098 ();
 b15zdnd11an1n32x5 FILLER_223_1162 ();
 b15zdnd11an1n16x5 FILLER_223_1194 ();
 b15zdnd11an1n04x5 FILLER_223_1210 ();
 b15zdnd00an1n01x5 FILLER_223_1214 ();
 b15zdnd11an1n64x5 FILLER_223_1227 ();
 b15zdnd11an1n64x5 FILLER_223_1291 ();
 b15zdnd11an1n08x5 FILLER_223_1355 ();
 b15zdnd00an1n02x5 FILLER_223_1363 ();
 b15zdnd00an1n01x5 FILLER_223_1365 ();
 b15zdnd11an1n64x5 FILLER_223_1405 ();
 b15zdnd11an1n64x5 FILLER_223_1469 ();
 b15zdnd11an1n64x5 FILLER_223_1533 ();
 b15zdnd11an1n64x5 FILLER_223_1597 ();
 b15zdnd11an1n64x5 FILLER_223_1661 ();
 b15zdnd11an1n64x5 FILLER_223_1725 ();
 b15zdnd11an1n64x5 FILLER_223_1789 ();
 b15zdnd11an1n64x5 FILLER_223_1853 ();
 b15zdnd11an1n64x5 FILLER_223_1917 ();
 b15zdnd11an1n64x5 FILLER_223_1981 ();
 b15zdnd11an1n64x5 FILLER_223_2045 ();
 b15zdnd11an1n64x5 FILLER_223_2109 ();
 b15zdnd11an1n32x5 FILLER_223_2173 ();
 b15zdnd11an1n04x5 FILLER_223_2205 ();
 b15zdnd00an1n01x5 FILLER_223_2209 ();
 b15zdnd11an1n64x5 FILLER_223_2214 ();
 b15zdnd11an1n04x5 FILLER_223_2278 ();
 b15zdnd00an1n02x5 FILLER_223_2282 ();
 b15zdnd11an1n64x5 FILLER_224_8 ();
 b15zdnd11an1n64x5 FILLER_224_72 ();
 b15zdnd11an1n64x5 FILLER_224_136 ();
 b15zdnd11an1n04x5 FILLER_224_200 ();
 b15zdnd00an1n02x5 FILLER_224_204 ();
 b15zdnd00an1n01x5 FILLER_224_206 ();
 b15zdnd11an1n04x5 FILLER_224_210 ();
 b15zdnd11an1n32x5 FILLER_224_266 ();
 b15zdnd11an1n08x5 FILLER_224_298 ();
 b15zdnd11an1n04x5 FILLER_224_306 ();
 b15zdnd00an1n02x5 FILLER_224_310 ();
 b15zdnd00an1n01x5 FILLER_224_312 ();
 b15zdnd11an1n64x5 FILLER_224_322 ();
 b15zdnd11an1n64x5 FILLER_224_386 ();
 b15zdnd11an1n32x5 FILLER_224_450 ();
 b15zdnd11an1n16x5 FILLER_224_482 ();
 b15zdnd11an1n04x5 FILLER_224_498 ();
 b15zdnd00an1n01x5 FILLER_224_502 ();
 b15zdnd11an1n64x5 FILLER_224_545 ();
 b15zdnd11an1n32x5 FILLER_224_609 ();
 b15zdnd11an1n04x5 FILLER_224_641 ();
 b15zdnd00an1n02x5 FILLER_224_645 ();
 b15zdnd00an1n01x5 FILLER_224_647 ();
 b15zdnd11an1n32x5 FILLER_224_656 ();
 b15zdnd11an1n16x5 FILLER_224_688 ();
 b15zdnd11an1n08x5 FILLER_224_704 ();
 b15zdnd11an1n04x5 FILLER_224_712 ();
 b15zdnd00an1n02x5 FILLER_224_716 ();
 b15zdnd11an1n64x5 FILLER_224_726 ();
 b15zdnd11an1n16x5 FILLER_224_790 ();
 b15zdnd11an1n04x5 FILLER_224_806 ();
 b15zdnd00an1n01x5 FILLER_224_810 ();
 b15zdnd11an1n64x5 FILLER_224_814 ();
 b15zdnd11an1n64x5 FILLER_224_878 ();
 b15zdnd11an1n64x5 FILLER_224_942 ();
 b15zdnd11an1n32x5 FILLER_224_1006 ();
 b15zdnd11an1n16x5 FILLER_224_1038 ();
 b15zdnd11an1n04x5 FILLER_224_1054 ();
 b15zdnd00an1n02x5 FILLER_224_1058 ();
 b15zdnd11an1n08x5 FILLER_224_1063 ();
 b15zdnd11an1n64x5 FILLER_224_1098 ();
 b15zdnd11an1n64x5 FILLER_224_1162 ();
 b15zdnd11an1n64x5 FILLER_224_1226 ();
 b15zdnd11an1n32x5 FILLER_224_1290 ();
 b15zdnd11an1n16x5 FILLER_224_1322 ();
 b15zdnd11an1n04x5 FILLER_224_1338 ();
 b15zdnd11an1n64x5 FILLER_224_1394 ();
 b15zdnd11an1n64x5 FILLER_224_1458 ();
 b15zdnd11an1n32x5 FILLER_224_1522 ();
 b15zdnd11an1n16x5 FILLER_224_1554 ();
 b15zdnd11an1n08x5 FILLER_224_1570 ();
 b15zdnd00an1n02x5 FILLER_224_1578 ();
 b15zdnd00an1n01x5 FILLER_224_1580 ();
 b15zdnd11an1n64x5 FILLER_224_1585 ();
 b15zdnd11an1n64x5 FILLER_224_1649 ();
 b15zdnd11an1n64x5 FILLER_224_1713 ();
 b15zdnd11an1n64x5 FILLER_224_1777 ();
 b15zdnd11an1n64x5 FILLER_224_1841 ();
 b15zdnd11an1n64x5 FILLER_224_1905 ();
 b15zdnd11an1n16x5 FILLER_224_1969 ();
 b15zdnd11an1n08x5 FILLER_224_1985 ();
 b15zdnd11an1n04x5 FILLER_224_1993 ();
 b15zdnd00an1n01x5 FILLER_224_1997 ();
 b15zdnd11an1n04x5 FILLER_224_2001 ();
 b15zdnd11an1n04x5 FILLER_224_2008 ();
 b15zdnd11an1n64x5 FILLER_224_2018 ();
 b15zdnd11an1n16x5 FILLER_224_2082 ();
 b15zdnd11an1n04x5 FILLER_224_2098 ();
 b15zdnd11an1n32x5 FILLER_224_2116 ();
 b15zdnd11an1n04x5 FILLER_224_2148 ();
 b15zdnd00an1n02x5 FILLER_224_2152 ();
 b15zdnd11an1n32x5 FILLER_224_2162 ();
 b15zdnd11an1n04x5 FILLER_224_2194 ();
 b15zdnd00an1n02x5 FILLER_224_2198 ();
 b15zdnd00an1n01x5 FILLER_224_2200 ();
 b15zdnd11an1n04x5 FILLER_224_2208 ();
 b15zdnd11an1n16x5 FILLER_224_2221 ();
 b15zdnd11an1n08x5 FILLER_224_2237 ();
 b15zdnd11an1n04x5 FILLER_224_2245 ();
 b15zdnd00an1n02x5 FILLER_224_2249 ();
 b15zdnd11an1n16x5 FILLER_224_2256 ();
 b15zdnd11an1n04x5 FILLER_224_2272 ();
 b15zdnd11an1n64x5 FILLER_225_0 ();
 b15zdnd11an1n64x5 FILLER_225_64 ();
 b15zdnd11an1n64x5 FILLER_225_128 ();
 b15zdnd11an1n16x5 FILLER_225_192 ();
 b15zdnd11an1n04x5 FILLER_225_208 ();
 b15zdnd00an1n01x5 FILLER_225_212 ();
 b15zdnd11an1n64x5 FILLER_225_216 ();
 b15zdnd11an1n64x5 FILLER_225_280 ();
 b15zdnd11an1n64x5 FILLER_225_344 ();
 b15zdnd11an1n64x5 FILLER_225_408 ();
 b15zdnd11an1n32x5 FILLER_225_472 ();
 b15zdnd00an1n02x5 FILLER_225_504 ();
 b15zdnd00an1n01x5 FILLER_225_506 ();
 b15zdnd11an1n64x5 FILLER_225_549 ();
 b15zdnd11an1n64x5 FILLER_225_613 ();
 b15zdnd11an1n64x5 FILLER_225_677 ();
 b15zdnd11an1n64x5 FILLER_225_741 ();
 b15zdnd11an1n16x5 FILLER_225_805 ();
 b15zdnd11an1n08x5 FILLER_225_821 ();
 b15zdnd11an1n64x5 FILLER_225_860 ();
 b15zdnd11an1n64x5 FILLER_225_924 ();
 b15zdnd11an1n32x5 FILLER_225_988 ();
 b15zdnd11an1n08x5 FILLER_225_1020 ();
 b15zdnd11an1n04x5 FILLER_225_1028 ();
 b15zdnd00an1n01x5 FILLER_225_1032 ();
 b15zdnd11an1n64x5 FILLER_225_1085 ();
 b15zdnd11an1n32x5 FILLER_225_1149 ();
 b15zdnd00an1n02x5 FILLER_225_1181 ();
 b15zdnd11an1n64x5 FILLER_225_1225 ();
 b15zdnd11an1n64x5 FILLER_225_1289 ();
 b15zdnd11an1n08x5 FILLER_225_1353 ();
 b15zdnd00an1n01x5 FILLER_225_1361 ();
 b15zdnd11an1n04x5 FILLER_225_1365 ();
 b15zdnd11an1n04x5 FILLER_225_1372 ();
 b15zdnd11an1n04x5 FILLER_225_1379 ();
 b15zdnd00an1n02x5 FILLER_225_1383 ();
 b15zdnd00an1n01x5 FILLER_225_1385 ();
 b15zdnd11an1n64x5 FILLER_225_1393 ();
 b15zdnd11an1n32x5 FILLER_225_1457 ();
 b15zdnd11an1n16x5 FILLER_225_1489 ();
 b15zdnd11an1n08x5 FILLER_225_1505 ();
 b15zdnd00an1n02x5 FILLER_225_1513 ();
 b15zdnd11an1n04x5 FILLER_225_1518 ();
 b15zdnd11an1n64x5 FILLER_225_1525 ();
 b15zdnd11an1n64x5 FILLER_225_1589 ();
 b15zdnd11an1n64x5 FILLER_225_1653 ();
 b15zdnd11an1n64x5 FILLER_225_1717 ();
 b15zdnd11an1n64x5 FILLER_225_1781 ();
 b15zdnd11an1n64x5 FILLER_225_1845 ();
 b15zdnd11an1n32x5 FILLER_225_1909 ();
 b15zdnd11an1n16x5 FILLER_225_1941 ();
 b15zdnd11an1n08x5 FILLER_225_1957 ();
 b15zdnd11an1n04x5 FILLER_225_1965 ();
 b15zdnd00an1n02x5 FILLER_225_1969 ();
 b15zdnd00an1n01x5 FILLER_225_1971 ();
 b15zdnd11an1n08x5 FILLER_225_2006 ();
 b15zdnd11an1n04x5 FILLER_225_2014 ();
 b15zdnd11an1n04x5 FILLER_225_2045 ();
 b15zdnd11an1n32x5 FILLER_225_2055 ();
 b15zdnd11an1n08x5 FILLER_225_2087 ();
 b15zdnd00an1n02x5 FILLER_225_2095 ();
 b15zdnd11an1n16x5 FILLER_225_2109 ();
 b15zdnd11an1n32x5 FILLER_225_2129 ();
 b15zdnd11an1n16x5 FILLER_225_2161 ();
 b15zdnd00an1n01x5 FILLER_225_2177 ();
 b15zdnd11an1n04x5 FILLER_225_2184 ();
 b15zdnd00an1n01x5 FILLER_225_2188 ();
 b15zdnd11an1n08x5 FILLER_225_2199 ();
 b15zdnd00an1n02x5 FILLER_225_2207 ();
 b15zdnd00an1n01x5 FILLER_225_2209 ();
 b15zdnd11an1n16x5 FILLER_225_2216 ();
 b15zdnd11an1n08x5 FILLER_225_2232 ();
 b15zdnd00an1n02x5 FILLER_225_2240 ();
 b15zdnd11an1n32x5 FILLER_225_2246 ();
 b15zdnd11an1n04x5 FILLER_225_2278 ();
 b15zdnd00an1n02x5 FILLER_225_2282 ();
 b15zdnd11an1n64x5 FILLER_226_8 ();
 b15zdnd11an1n64x5 FILLER_226_72 ();
 b15zdnd11an1n64x5 FILLER_226_136 ();
 b15zdnd11an1n64x5 FILLER_226_200 ();
 b15zdnd11an1n64x5 FILLER_226_264 ();
 b15zdnd11an1n64x5 FILLER_226_328 ();
 b15zdnd11an1n64x5 FILLER_226_392 ();
 b15zdnd11an1n32x5 FILLER_226_456 ();
 b15zdnd11an1n04x5 FILLER_226_488 ();
 b15zdnd00an1n01x5 FILLER_226_492 ();
 b15zdnd11an1n64x5 FILLER_226_535 ();
 b15zdnd11an1n64x5 FILLER_226_599 ();
 b15zdnd11an1n32x5 FILLER_226_663 ();
 b15zdnd11an1n16x5 FILLER_226_695 ();
 b15zdnd11an1n04x5 FILLER_226_711 ();
 b15zdnd00an1n02x5 FILLER_226_715 ();
 b15zdnd00an1n01x5 FILLER_226_717 ();
 b15zdnd11an1n64x5 FILLER_226_726 ();
 b15zdnd11an1n64x5 FILLER_226_790 ();
 b15zdnd11an1n64x5 FILLER_226_854 ();
 b15zdnd11an1n64x5 FILLER_226_918 ();
 b15zdnd11an1n64x5 FILLER_226_982 ();
 b15zdnd11an1n04x5 FILLER_226_1046 ();
 b15zdnd00an1n01x5 FILLER_226_1050 ();
 b15zdnd11an1n04x5 FILLER_226_1054 ();
 b15zdnd11an1n08x5 FILLER_226_1061 ();
 b15zdnd11an1n04x5 FILLER_226_1069 ();
 b15zdnd11an1n64x5 FILLER_226_1076 ();
 b15zdnd11an1n64x5 FILLER_226_1140 ();
 b15zdnd11an1n64x5 FILLER_226_1204 ();
 b15zdnd11an1n64x5 FILLER_226_1268 ();
 b15zdnd11an1n32x5 FILLER_226_1332 ();
 b15zdnd00an1n01x5 FILLER_226_1364 ();
 b15zdnd11an1n64x5 FILLER_226_1368 ();
 b15zdnd11an1n32x5 FILLER_226_1432 ();
 b15zdnd11an1n16x5 FILLER_226_1464 ();
 b15zdnd11an1n04x5 FILLER_226_1480 ();
 b15zdnd11an1n64x5 FILLER_226_1524 ();
 b15zdnd11an1n64x5 FILLER_226_1588 ();
 b15zdnd11an1n64x5 FILLER_226_1652 ();
 b15zdnd11an1n64x5 FILLER_226_1716 ();
 b15zdnd11an1n64x5 FILLER_226_1780 ();
 b15zdnd11an1n64x5 FILLER_226_1844 ();
 b15zdnd11an1n64x5 FILLER_226_1908 ();
 b15zdnd11an1n64x5 FILLER_226_1972 ();
 b15zdnd11an1n04x5 FILLER_226_2036 ();
 b15zdnd00an1n01x5 FILLER_226_2040 ();
 b15zdnd11an1n32x5 FILLER_226_2049 ();
 b15zdnd11an1n08x5 FILLER_226_2081 ();
 b15zdnd00an1n02x5 FILLER_226_2089 ();
 b15zdnd00an1n01x5 FILLER_226_2091 ();
 b15zdnd11an1n04x5 FILLER_226_2097 ();
 b15zdnd11an1n04x5 FILLER_226_2107 ();
 b15zdnd00an1n02x5 FILLER_226_2111 ();
 b15zdnd11an1n04x5 FILLER_226_2116 ();
 b15zdnd11an1n16x5 FILLER_226_2134 ();
 b15zdnd11an1n04x5 FILLER_226_2150 ();
 b15zdnd11an1n04x5 FILLER_226_2162 ();
 b15zdnd00an1n02x5 FILLER_226_2166 ();
 b15zdnd00an1n01x5 FILLER_226_2168 ();
 b15zdnd11an1n16x5 FILLER_226_2178 ();
 b15zdnd11an1n08x5 FILLER_226_2194 ();
 b15zdnd00an1n02x5 FILLER_226_2202 ();
 b15zdnd00an1n01x5 FILLER_226_2204 ();
 b15zdnd11an1n04x5 FILLER_226_2210 ();
 b15zdnd11an1n32x5 FILLER_226_2218 ();
 b15zdnd11an1n08x5 FILLER_226_2250 ();
 b15zdnd00an1n02x5 FILLER_226_2258 ();
 b15zdnd00an1n01x5 FILLER_226_2260 ();
 b15zdnd11an1n08x5 FILLER_226_2265 ();
 b15zdnd00an1n02x5 FILLER_226_2273 ();
 b15zdnd00an1n01x5 FILLER_226_2275 ();
 b15zdnd11an1n32x5 FILLER_227_0 ();
 b15zdnd11an1n16x5 FILLER_227_32 ();
 b15zdnd11an1n04x5 FILLER_227_48 ();
 b15zdnd00an1n02x5 FILLER_227_52 ();
 b15zdnd11an1n16x5 FILLER_227_57 ();
 b15zdnd00an1n02x5 FILLER_227_73 ();
 b15zdnd00an1n01x5 FILLER_227_75 ();
 b15zdnd11an1n64x5 FILLER_227_90 ();
 b15zdnd11an1n64x5 FILLER_227_154 ();
 b15zdnd11an1n32x5 FILLER_227_218 ();
 b15zdnd11an1n08x5 FILLER_227_250 ();
 b15zdnd00an1n01x5 FILLER_227_258 ();
 b15zdnd11an1n64x5 FILLER_227_301 ();
 b15zdnd11an1n64x5 FILLER_227_365 ();
 b15zdnd11an1n64x5 FILLER_227_429 ();
 b15zdnd11an1n64x5 FILLER_227_535 ();
 b15zdnd11an1n64x5 FILLER_227_599 ();
 b15zdnd11an1n64x5 FILLER_227_663 ();
 b15zdnd11an1n64x5 FILLER_227_727 ();
 b15zdnd11an1n64x5 FILLER_227_791 ();
 b15zdnd11an1n64x5 FILLER_227_855 ();
 b15zdnd11an1n64x5 FILLER_227_919 ();
 b15zdnd11an1n64x5 FILLER_227_983 ();
 b15zdnd11an1n64x5 FILLER_227_1047 ();
 b15zdnd11an1n64x5 FILLER_227_1111 ();
 b15zdnd11an1n64x5 FILLER_227_1175 ();
 b15zdnd11an1n64x5 FILLER_227_1239 ();
 b15zdnd11an1n08x5 FILLER_227_1303 ();
 b15zdnd11an1n04x5 FILLER_227_1311 ();
 b15zdnd00an1n02x5 FILLER_227_1315 ();
 b15zdnd00an1n01x5 FILLER_227_1317 ();
 b15zdnd11an1n32x5 FILLER_227_1334 ();
 b15zdnd11an1n08x5 FILLER_227_1366 ();
 b15zdnd11an1n04x5 FILLER_227_1374 ();
 b15zdnd11an1n64x5 FILLER_227_1390 ();
 b15zdnd11an1n32x5 FILLER_227_1454 ();
 b15zdnd11an1n08x5 FILLER_227_1486 ();
 b15zdnd11an1n04x5 FILLER_227_1494 ();
 b15zdnd00an1n02x5 FILLER_227_1498 ();
 b15zdnd11an1n64x5 FILLER_227_1505 ();
 b15zdnd11an1n64x5 FILLER_227_1569 ();
 b15zdnd11an1n64x5 FILLER_227_1633 ();
 b15zdnd11an1n64x5 FILLER_227_1697 ();
 b15zdnd11an1n64x5 FILLER_227_1761 ();
 b15zdnd11an1n64x5 FILLER_227_1825 ();
 b15zdnd11an1n64x5 FILLER_227_1889 ();
 b15zdnd11an1n32x5 FILLER_227_1953 ();
 b15zdnd11an1n16x5 FILLER_227_1985 ();
 b15zdnd11an1n08x5 FILLER_227_2001 ();
 b15zdnd11an1n04x5 FILLER_227_2009 ();
 b15zdnd00an1n02x5 FILLER_227_2013 ();
 b15zdnd00an1n01x5 FILLER_227_2015 ();
 b15zdnd11an1n32x5 FILLER_227_2021 ();
 b15zdnd11an1n16x5 FILLER_227_2053 ();
 b15zdnd11an1n04x5 FILLER_227_2069 ();
 b15zdnd00an1n02x5 FILLER_227_2073 ();
 b15zdnd00an1n01x5 FILLER_227_2075 ();
 b15zdnd11an1n04x5 FILLER_227_2082 ();
 b15zdnd11an1n04x5 FILLER_227_2101 ();
 b15zdnd11an1n64x5 FILLER_227_2114 ();
 b15zdnd11an1n64x5 FILLER_227_2178 ();
 b15zdnd00an1n02x5 FILLER_227_2242 ();
 b15zdnd11an1n16x5 FILLER_227_2258 ();
 b15zdnd00an1n02x5 FILLER_227_2282 ();
 b15zdnd11an1n32x5 FILLER_228_8 ();
 b15zdnd11an1n08x5 FILLER_228_40 ();
 b15zdnd11an1n04x5 FILLER_228_48 ();
 b15zdnd00an1n01x5 FILLER_228_52 ();
 b15zdnd11an1n04x5 FILLER_228_56 ();
 b15zdnd11an1n64x5 FILLER_228_63 ();
 b15zdnd11an1n64x5 FILLER_228_127 ();
 b15zdnd11an1n16x5 FILLER_228_191 ();
 b15zdnd00an1n01x5 FILLER_228_207 ();
 b15zdnd11an1n64x5 FILLER_228_250 ();
 b15zdnd11an1n64x5 FILLER_228_314 ();
 b15zdnd11an1n64x5 FILLER_228_378 ();
 b15zdnd11an1n32x5 FILLER_228_442 ();
 b15zdnd11an1n08x5 FILLER_228_474 ();
 b15zdnd11an1n04x5 FILLER_228_482 ();
 b15zdnd00an1n02x5 FILLER_228_486 ();
 b15zdnd00an1n01x5 FILLER_228_488 ();
 b15zdnd11an1n04x5 FILLER_228_493 ();
 b15zdnd11an1n64x5 FILLER_228_536 ();
 b15zdnd11an1n64x5 FILLER_228_600 ();
 b15zdnd11an1n32x5 FILLER_228_664 ();
 b15zdnd11an1n16x5 FILLER_228_696 ();
 b15zdnd11an1n04x5 FILLER_228_712 ();
 b15zdnd00an1n02x5 FILLER_228_716 ();
 b15zdnd11an1n64x5 FILLER_228_726 ();
 b15zdnd11an1n64x5 FILLER_228_790 ();
 b15zdnd11an1n64x5 FILLER_228_854 ();
 b15zdnd11an1n64x5 FILLER_228_918 ();
 b15zdnd11an1n64x5 FILLER_228_982 ();
 b15zdnd11an1n64x5 FILLER_228_1046 ();
 b15zdnd11an1n64x5 FILLER_228_1110 ();
 b15zdnd11an1n64x5 FILLER_228_1174 ();
 b15zdnd11an1n64x5 FILLER_228_1238 ();
 b15zdnd11an1n32x5 FILLER_228_1302 ();
 b15zdnd00an1n02x5 FILLER_228_1334 ();
 b15zdnd11an1n16x5 FILLER_228_1344 ();
 b15zdnd11an1n64x5 FILLER_228_1399 ();
 b15zdnd11an1n64x5 FILLER_228_1463 ();
 b15zdnd11an1n64x5 FILLER_228_1527 ();
 b15zdnd11an1n64x5 FILLER_228_1591 ();
 b15zdnd11an1n64x5 FILLER_228_1655 ();
 b15zdnd11an1n64x5 FILLER_228_1719 ();
 b15zdnd11an1n64x5 FILLER_228_1783 ();
 b15zdnd11an1n16x5 FILLER_228_1847 ();
 b15zdnd11an1n08x5 FILLER_228_1863 ();
 b15zdnd11an1n04x5 FILLER_228_1871 ();
 b15zdnd11an1n64x5 FILLER_228_1896 ();
 b15zdnd11an1n16x5 FILLER_228_1960 ();
 b15zdnd00an1n02x5 FILLER_228_1976 ();
 b15zdnd11an1n64x5 FILLER_228_2030 ();
 b15zdnd11an1n32x5 FILLER_228_2094 ();
 b15zdnd11an1n16x5 FILLER_228_2126 ();
 b15zdnd11an1n08x5 FILLER_228_2142 ();
 b15zdnd11an1n04x5 FILLER_228_2150 ();
 b15zdnd11an1n64x5 FILLER_228_2162 ();
 b15zdnd11an1n16x5 FILLER_228_2226 ();
 b15zdnd11an1n08x5 FILLER_228_2256 ();
 b15zdnd00an1n01x5 FILLER_228_2264 ();
 b15zdnd00an1n02x5 FILLER_228_2273 ();
 b15zdnd00an1n01x5 FILLER_228_2275 ();
 b15zdnd11an1n16x5 FILLER_229_0 ();
 b15zdnd00an1n02x5 FILLER_229_16 ();
 b15zdnd00an1n01x5 FILLER_229_18 ();
 b15zdnd11an1n08x5 FILLER_229_23 ();
 b15zdnd00an1n02x5 FILLER_229_31 ();
 b15zdnd11an1n64x5 FILLER_229_85 ();
 b15zdnd11an1n64x5 FILLER_229_149 ();
 b15zdnd11an1n64x5 FILLER_229_213 ();
 b15zdnd11an1n64x5 FILLER_229_277 ();
 b15zdnd11an1n64x5 FILLER_229_341 ();
 b15zdnd11an1n64x5 FILLER_229_405 ();
 b15zdnd11an1n16x5 FILLER_229_469 ();
 b15zdnd11an1n08x5 FILLER_229_485 ();
 b15zdnd00an1n02x5 FILLER_229_493 ();
 b15zdnd00an1n01x5 FILLER_229_495 ();
 b15zdnd11an1n08x5 FILLER_229_507 ();
 b15zdnd00an1n02x5 FILLER_229_515 ();
 b15zdnd11an1n64x5 FILLER_229_524 ();
 b15zdnd11an1n32x5 FILLER_229_588 ();
 b15zdnd11an1n16x5 FILLER_229_620 ();
 b15zdnd11an1n64x5 FILLER_229_640 ();
 b15zdnd11an1n64x5 FILLER_229_704 ();
 b15zdnd11an1n64x5 FILLER_229_768 ();
 b15zdnd11an1n64x5 FILLER_229_832 ();
 b15zdnd11an1n64x5 FILLER_229_896 ();
 b15zdnd11an1n64x5 FILLER_229_960 ();
 b15zdnd11an1n64x5 FILLER_229_1024 ();
 b15zdnd11an1n64x5 FILLER_229_1088 ();
 b15zdnd11an1n04x5 FILLER_229_1152 ();
 b15zdnd00an1n01x5 FILLER_229_1156 ();
 b15zdnd11an1n64x5 FILLER_229_1172 ();
 b15zdnd11an1n64x5 FILLER_229_1236 ();
 b15zdnd11an1n32x5 FILLER_229_1300 ();
 b15zdnd00an1n02x5 FILLER_229_1332 ();
 b15zdnd00an1n01x5 FILLER_229_1334 ();
 b15zdnd11an1n64x5 FILLER_229_1342 ();
 b15zdnd11an1n64x5 FILLER_229_1406 ();
 b15zdnd11an1n64x5 FILLER_229_1470 ();
 b15zdnd11an1n64x5 FILLER_229_1534 ();
 b15zdnd11an1n64x5 FILLER_229_1598 ();
 b15zdnd11an1n64x5 FILLER_229_1662 ();
 b15zdnd11an1n64x5 FILLER_229_1726 ();
 b15zdnd11an1n08x5 FILLER_229_1790 ();
 b15zdnd11an1n04x5 FILLER_229_1798 ();
 b15zdnd00an1n02x5 FILLER_229_1802 ();
 b15zdnd00an1n01x5 FILLER_229_1804 ();
 b15zdnd11an1n16x5 FILLER_229_1813 ();
 b15zdnd11an1n04x5 FILLER_229_1881 ();
 b15zdnd00an1n01x5 FILLER_229_1885 ();
 b15zdnd11an1n64x5 FILLER_229_1890 ();
 b15zdnd11an1n32x5 FILLER_229_1954 ();
 b15zdnd11an1n08x5 FILLER_229_1986 ();
 b15zdnd00an1n02x5 FILLER_229_1994 ();
 b15zdnd11an1n04x5 FILLER_229_1999 ();
 b15zdnd00an1n01x5 FILLER_229_2003 ();
 b15zdnd11an1n32x5 FILLER_229_2007 ();
 b15zdnd11an1n08x5 FILLER_229_2039 ();
 b15zdnd00an1n01x5 FILLER_229_2047 ();
 b15zdnd11an1n64x5 FILLER_229_2055 ();
 b15zdnd11an1n64x5 FILLER_229_2119 ();
 b15zdnd11an1n64x5 FILLER_229_2183 ();
 b15zdnd11an1n32x5 FILLER_229_2247 ();
 b15zdnd11an1n04x5 FILLER_229_2279 ();
 b15zdnd00an1n01x5 FILLER_229_2283 ();
 b15zdnd11an1n32x5 FILLER_230_8 ();
 b15zdnd11an1n08x5 FILLER_230_40 ();
 b15zdnd11an1n04x5 FILLER_230_48 ();
 b15zdnd00an1n01x5 FILLER_230_52 ();
 b15zdnd11an1n04x5 FILLER_230_84 ();
 b15zdnd11an1n64x5 FILLER_230_114 ();
 b15zdnd11an1n64x5 FILLER_230_178 ();
 b15zdnd11an1n08x5 FILLER_230_242 ();
 b15zdnd00an1n02x5 FILLER_230_250 ();
 b15zdnd00an1n01x5 FILLER_230_252 ();
 b15zdnd11an1n64x5 FILLER_230_271 ();
 b15zdnd11an1n64x5 FILLER_230_335 ();
 b15zdnd11an1n64x5 FILLER_230_399 ();
 b15zdnd11an1n32x5 FILLER_230_463 ();
 b15zdnd11an1n04x5 FILLER_230_495 ();
 b15zdnd11an1n64x5 FILLER_230_506 ();
 b15zdnd11an1n64x5 FILLER_230_570 ();
 b15zdnd11an1n04x5 FILLER_230_634 ();
 b15zdnd00an1n01x5 FILLER_230_638 ();
 b15zdnd11an1n32x5 FILLER_230_681 ();
 b15zdnd11an1n04x5 FILLER_230_713 ();
 b15zdnd00an1n01x5 FILLER_230_717 ();
 b15zdnd11an1n64x5 FILLER_230_726 ();
 b15zdnd11an1n64x5 FILLER_230_790 ();
 b15zdnd11an1n64x5 FILLER_230_854 ();
 b15zdnd11an1n64x5 FILLER_230_918 ();
 b15zdnd11an1n64x5 FILLER_230_982 ();
 b15zdnd11an1n64x5 FILLER_230_1046 ();
 b15zdnd11an1n16x5 FILLER_230_1110 ();
 b15zdnd00an1n02x5 FILLER_230_1126 ();
 b15zdnd11an1n04x5 FILLER_230_1131 ();
 b15zdnd11an1n16x5 FILLER_230_1138 ();
 b15zdnd11an1n04x5 FILLER_230_1154 ();
 b15zdnd00an1n02x5 FILLER_230_1158 ();
 b15zdnd00an1n01x5 FILLER_230_1160 ();
 b15zdnd11an1n64x5 FILLER_230_1165 ();
 b15zdnd11an1n64x5 FILLER_230_1229 ();
 b15zdnd11an1n64x5 FILLER_230_1293 ();
 b15zdnd00an1n02x5 FILLER_230_1357 ();
 b15zdnd00an1n01x5 FILLER_230_1359 ();
 b15zdnd11an1n64x5 FILLER_230_1364 ();
 b15zdnd11an1n64x5 FILLER_230_1428 ();
 b15zdnd11an1n64x5 FILLER_230_1492 ();
 b15zdnd11an1n64x5 FILLER_230_1556 ();
 b15zdnd11an1n64x5 FILLER_230_1620 ();
 b15zdnd11an1n64x5 FILLER_230_1684 ();
 b15zdnd11an1n64x5 FILLER_230_1748 ();
 b15zdnd11an1n32x5 FILLER_230_1812 ();
 b15zdnd00an1n02x5 FILLER_230_1844 ();
 b15zdnd00an1n01x5 FILLER_230_1846 ();
 b15zdnd11an1n04x5 FILLER_230_1850 ();
 b15zdnd11an1n04x5 FILLER_230_1857 ();
 b15zdnd11an1n16x5 FILLER_230_1864 ();
 b15zdnd11an1n64x5 FILLER_230_1907 ();
 b15zdnd11an1n16x5 FILLER_230_1971 ();
 b15zdnd11an1n08x5 FILLER_230_1987 ();
 b15zdnd11an1n04x5 FILLER_230_1995 ();
 b15zdnd00an1n02x5 FILLER_230_1999 ();
 b15zdnd00an1n01x5 FILLER_230_2001 ();
 b15zdnd11an1n32x5 FILLER_230_2005 ();
 b15zdnd11an1n16x5 FILLER_230_2037 ();
 b15zdnd11an1n32x5 FILLER_230_2095 ();
 b15zdnd11an1n16x5 FILLER_230_2127 ();
 b15zdnd11an1n08x5 FILLER_230_2143 ();
 b15zdnd00an1n02x5 FILLER_230_2151 ();
 b15zdnd00an1n01x5 FILLER_230_2153 ();
 b15zdnd11an1n64x5 FILLER_230_2162 ();
 b15zdnd11an1n32x5 FILLER_230_2226 ();
 b15zdnd11an1n16x5 FILLER_230_2258 ();
 b15zdnd00an1n02x5 FILLER_230_2274 ();
 b15zdnd11an1n64x5 FILLER_231_0 ();
 b15zdnd00an1n01x5 FILLER_231_64 ();
 b15zdnd11an1n16x5 FILLER_231_110 ();
 b15zdnd11an1n08x5 FILLER_231_126 ();
 b15zdnd11an1n64x5 FILLER_231_145 ();
 b15zdnd11an1n32x5 FILLER_231_209 ();
 b15zdnd00an1n02x5 FILLER_231_241 ();
 b15zdnd00an1n01x5 FILLER_231_243 ();
 b15zdnd11an1n04x5 FILLER_231_247 ();
 b15zdnd11an1n64x5 FILLER_231_293 ();
 b15zdnd11an1n64x5 FILLER_231_357 ();
 b15zdnd11an1n64x5 FILLER_231_421 ();
 b15zdnd11an1n08x5 FILLER_231_485 ();
 b15zdnd11an1n04x5 FILLER_231_493 ();
 b15zdnd00an1n02x5 FILLER_231_497 ();
 b15zdnd11an1n04x5 FILLER_231_504 ();
 b15zdnd11an1n64x5 FILLER_231_513 ();
 b15zdnd11an1n64x5 FILLER_231_577 ();
 b15zdnd11an1n64x5 FILLER_231_641 ();
 b15zdnd11an1n64x5 FILLER_231_705 ();
 b15zdnd11an1n64x5 FILLER_231_769 ();
 b15zdnd11an1n64x5 FILLER_231_833 ();
 b15zdnd11an1n64x5 FILLER_231_897 ();
 b15zdnd11an1n64x5 FILLER_231_961 ();
 b15zdnd11an1n64x5 FILLER_231_1025 ();
 b15zdnd11an1n16x5 FILLER_231_1089 ();
 b15zdnd00an1n02x5 FILLER_231_1105 ();
 b15zdnd00an1n01x5 FILLER_231_1107 ();
 b15zdnd11an1n64x5 FILLER_231_1160 ();
 b15zdnd11an1n32x5 FILLER_231_1224 ();
 b15zdnd11an1n04x5 FILLER_231_1256 ();
 b15zdnd00an1n01x5 FILLER_231_1260 ();
 b15zdnd11an1n04x5 FILLER_231_1264 ();
 b15zdnd11an1n64x5 FILLER_231_1271 ();
 b15zdnd11an1n64x5 FILLER_231_1335 ();
 b15zdnd11an1n32x5 FILLER_231_1399 ();
 b15zdnd11an1n04x5 FILLER_231_1431 ();
 b15zdnd00an1n02x5 FILLER_231_1435 ();
 b15zdnd00an1n01x5 FILLER_231_1437 ();
 b15zdnd11an1n04x5 FILLER_231_1469 ();
 b15zdnd00an1n01x5 FILLER_231_1473 ();
 b15zdnd11an1n64x5 FILLER_231_1489 ();
 b15zdnd11an1n64x5 FILLER_231_1553 ();
 b15zdnd11an1n64x5 FILLER_231_1617 ();
 b15zdnd11an1n64x5 FILLER_231_1681 ();
 b15zdnd11an1n64x5 FILLER_231_1745 ();
 b15zdnd11an1n32x5 FILLER_231_1809 ();
 b15zdnd11an1n08x5 FILLER_231_1841 ();
 b15zdnd11an1n04x5 FILLER_231_1849 ();
 b15zdnd00an1n02x5 FILLER_231_1853 ();
 b15zdnd00an1n01x5 FILLER_231_1855 ();
 b15zdnd11an1n16x5 FILLER_231_1864 ();
 b15zdnd00an1n02x5 FILLER_231_1880 ();
 b15zdnd00an1n01x5 FILLER_231_1882 ();
 b15zdnd11an1n32x5 FILLER_231_1889 ();
 b15zdnd11an1n04x5 FILLER_231_1921 ();
 b15zdnd11an1n64x5 FILLER_231_1930 ();
 b15zdnd11an1n16x5 FILLER_231_1994 ();
 b15zdnd11an1n08x5 FILLER_231_2010 ();
 b15zdnd11an1n04x5 FILLER_231_2018 ();
 b15zdnd00an1n02x5 FILLER_231_2022 ();
 b15zdnd00an1n01x5 FILLER_231_2024 ();
 b15zdnd11an1n32x5 FILLER_231_2029 ();
 b15zdnd11an1n08x5 FILLER_231_2061 ();
 b15zdnd11an1n04x5 FILLER_231_2069 ();
 b15zdnd00an1n02x5 FILLER_231_2073 ();
 b15zdnd11an1n64x5 FILLER_231_2085 ();
 b15zdnd11an1n64x5 FILLER_231_2149 ();
 b15zdnd11an1n64x5 FILLER_231_2213 ();
 b15zdnd11an1n04x5 FILLER_231_2277 ();
 b15zdnd00an1n02x5 FILLER_231_2281 ();
 b15zdnd00an1n01x5 FILLER_231_2283 ();
 b15zdnd11an1n16x5 FILLER_232_8 ();
 b15zdnd11an1n04x5 FILLER_232_24 ();
 b15zdnd11an1n16x5 FILLER_232_42 ();
 b15zdnd11an1n04x5 FILLER_232_58 ();
 b15zdnd00an1n01x5 FILLER_232_62 ();
 b15zdnd11an1n64x5 FILLER_232_77 ();
 b15zdnd11an1n64x5 FILLER_232_141 ();
 b15zdnd11an1n16x5 FILLER_232_205 ();
 b15zdnd11an1n04x5 FILLER_232_221 ();
 b15zdnd00an1n01x5 FILLER_232_225 ();
 b15zdnd11an1n64x5 FILLER_232_278 ();
 b15zdnd11an1n64x5 FILLER_232_342 ();
 b15zdnd11an1n64x5 FILLER_232_406 ();
 b15zdnd11an1n16x5 FILLER_232_470 ();
 b15zdnd11an1n08x5 FILLER_232_486 ();
 b15zdnd11an1n04x5 FILLER_232_494 ();
 b15zdnd00an1n02x5 FILLER_232_498 ();
 b15zdnd11an1n64x5 FILLER_232_510 ();
 b15zdnd11an1n64x5 FILLER_232_574 ();
 b15zdnd11an1n16x5 FILLER_232_638 ();
 b15zdnd11an1n08x5 FILLER_232_654 ();
 b15zdnd00an1n01x5 FILLER_232_662 ();
 b15zdnd00an1n02x5 FILLER_232_715 ();
 b15zdnd00an1n01x5 FILLER_232_717 ();
 b15zdnd11an1n16x5 FILLER_232_726 ();
 b15zdnd11an1n08x5 FILLER_232_742 ();
 b15zdnd00an1n02x5 FILLER_232_750 ();
 b15zdnd00an1n01x5 FILLER_232_752 ();
 b15zdnd11an1n64x5 FILLER_232_761 ();
 b15zdnd11an1n64x5 FILLER_232_825 ();
 b15zdnd11an1n64x5 FILLER_232_889 ();
 b15zdnd11an1n64x5 FILLER_232_953 ();
 b15zdnd11an1n64x5 FILLER_232_1017 ();
 b15zdnd11an1n32x5 FILLER_232_1081 ();
 b15zdnd11an1n08x5 FILLER_232_1113 ();
 b15zdnd00an1n02x5 FILLER_232_1121 ();
 b15zdnd00an1n01x5 FILLER_232_1123 ();
 b15zdnd11an1n04x5 FILLER_232_1127 ();
 b15zdnd11an1n04x5 FILLER_232_1134 ();
 b15zdnd11an1n64x5 FILLER_232_1141 ();
 b15zdnd11an1n16x5 FILLER_232_1205 ();
 b15zdnd11an1n08x5 FILLER_232_1221 ();
 b15zdnd00an1n01x5 FILLER_232_1229 ();
 b15zdnd11an1n64x5 FILLER_232_1270 ();
 b15zdnd11an1n64x5 FILLER_232_1334 ();
 b15zdnd11an1n64x5 FILLER_232_1398 ();
 b15zdnd11an1n64x5 FILLER_232_1462 ();
 b15zdnd11an1n64x5 FILLER_232_1526 ();
 b15zdnd11an1n64x5 FILLER_232_1590 ();
 b15zdnd11an1n64x5 FILLER_232_1654 ();
 b15zdnd11an1n64x5 FILLER_232_1718 ();
 b15zdnd11an1n64x5 FILLER_232_1782 ();
 b15zdnd11an1n04x5 FILLER_232_1846 ();
 b15zdnd00an1n02x5 FILLER_232_1850 ();
 b15zdnd00an1n01x5 FILLER_232_1852 ();
 b15zdnd11an1n64x5 FILLER_232_1895 ();
 b15zdnd11an1n64x5 FILLER_232_1959 ();
 b15zdnd11an1n64x5 FILLER_232_2023 ();
 b15zdnd11an1n64x5 FILLER_232_2087 ();
 b15zdnd00an1n02x5 FILLER_232_2151 ();
 b15zdnd00an1n01x5 FILLER_232_2153 ();
 b15zdnd11an1n64x5 FILLER_232_2162 ();
 b15zdnd11an1n32x5 FILLER_232_2226 ();
 b15zdnd11an1n16x5 FILLER_232_2258 ();
 b15zdnd00an1n02x5 FILLER_232_2274 ();
 b15zdnd11an1n08x5 FILLER_233_0 ();
 b15zdnd11an1n04x5 FILLER_233_8 ();
 b15zdnd00an1n02x5 FILLER_233_12 ();
 b15zdnd11an1n04x5 FILLER_233_22 ();
 b15zdnd00an1n02x5 FILLER_233_26 ();
 b15zdnd11an1n64x5 FILLER_233_42 ();
 b15zdnd11an1n64x5 FILLER_233_106 ();
 b15zdnd11an1n64x5 FILLER_233_170 ();
 b15zdnd11an1n08x5 FILLER_233_234 ();
 b15zdnd00an1n02x5 FILLER_233_242 ();
 b15zdnd11an1n04x5 FILLER_233_247 ();
 b15zdnd11an1n64x5 FILLER_233_254 ();
 b15zdnd11an1n64x5 FILLER_233_318 ();
 b15zdnd11an1n64x5 FILLER_233_382 ();
 b15zdnd11an1n32x5 FILLER_233_446 ();
 b15zdnd11an1n16x5 FILLER_233_478 ();
 b15zdnd11an1n04x5 FILLER_233_494 ();
 b15zdnd11an1n04x5 FILLER_233_502 ();
 b15zdnd11an1n64x5 FILLER_233_510 ();
 b15zdnd11an1n64x5 FILLER_233_574 ();
 b15zdnd11an1n32x5 FILLER_233_638 ();
 b15zdnd11an1n04x5 FILLER_233_670 ();
 b15zdnd00an1n02x5 FILLER_233_674 ();
 b15zdnd00an1n01x5 FILLER_233_676 ();
 b15zdnd11an1n04x5 FILLER_233_680 ();
 b15zdnd00an1n02x5 FILLER_233_684 ();
 b15zdnd00an1n01x5 FILLER_233_686 ();
 b15zdnd11an1n08x5 FILLER_233_690 ();
 b15zdnd11an1n04x5 FILLER_233_698 ();
 b15zdnd11an1n64x5 FILLER_233_706 ();
 b15zdnd11an1n64x5 FILLER_233_770 ();
 b15zdnd11an1n32x5 FILLER_233_834 ();
 b15zdnd11an1n16x5 FILLER_233_866 ();
 b15zdnd11an1n04x5 FILLER_233_882 ();
 b15zdnd11an1n64x5 FILLER_233_901 ();
 b15zdnd11an1n64x5 FILLER_233_965 ();
 b15zdnd11an1n64x5 FILLER_233_1029 ();
 b15zdnd11an1n64x5 FILLER_233_1093 ();
 b15zdnd11an1n64x5 FILLER_233_1157 ();
 b15zdnd11an1n64x5 FILLER_233_1221 ();
 b15zdnd11an1n08x5 FILLER_233_1285 ();
 b15zdnd00an1n02x5 FILLER_233_1293 ();
 b15zdnd11an1n04x5 FILLER_233_1298 ();
 b15zdnd11an1n64x5 FILLER_233_1305 ();
 b15zdnd11an1n64x5 FILLER_233_1369 ();
 b15zdnd11an1n64x5 FILLER_233_1433 ();
 b15zdnd11an1n64x5 FILLER_233_1497 ();
 b15zdnd11an1n64x5 FILLER_233_1561 ();
 b15zdnd11an1n64x5 FILLER_233_1625 ();
 b15zdnd11an1n64x5 FILLER_233_1689 ();
 b15zdnd11an1n64x5 FILLER_233_1753 ();
 b15zdnd11an1n16x5 FILLER_233_1817 ();
 b15zdnd00an1n01x5 FILLER_233_1833 ();
 b15zdnd11an1n64x5 FILLER_233_1837 ();
 b15zdnd11an1n64x5 FILLER_233_1901 ();
 b15zdnd11an1n64x5 FILLER_233_1965 ();
 b15zdnd11an1n32x5 FILLER_233_2029 ();
 b15zdnd11an1n16x5 FILLER_233_2061 ();
 b15zdnd11an1n64x5 FILLER_233_2119 ();
 b15zdnd11an1n64x5 FILLER_233_2183 ();
 b15zdnd11an1n04x5 FILLER_233_2247 ();
 b15zdnd00an1n01x5 FILLER_233_2251 ();
 b15zdnd11an1n16x5 FILLER_233_2256 ();
 b15zdnd11an1n08x5 FILLER_233_2272 ();
 b15zdnd11an1n04x5 FILLER_233_2280 ();
 b15zdnd11an1n16x5 FILLER_234_8 ();
 b15zdnd11an1n64x5 FILLER_234_28 ();
 b15zdnd11an1n64x5 FILLER_234_92 ();
 b15zdnd11an1n64x5 FILLER_234_156 ();
 b15zdnd11an1n64x5 FILLER_234_220 ();
 b15zdnd11an1n64x5 FILLER_234_284 ();
 b15zdnd11an1n32x5 FILLER_234_348 ();
 b15zdnd11an1n08x5 FILLER_234_380 ();
 b15zdnd11an1n64x5 FILLER_234_393 ();
 b15zdnd11an1n32x5 FILLER_234_457 ();
 b15zdnd11an1n08x5 FILLER_234_489 ();
 b15zdnd11an1n04x5 FILLER_234_497 ();
 b15zdnd00an1n02x5 FILLER_234_501 ();
 b15zdnd11an1n32x5 FILLER_234_509 ();
 b15zdnd11an1n08x5 FILLER_234_541 ();
 b15zdnd11an1n04x5 FILLER_234_549 ();
 b15zdnd00an1n02x5 FILLER_234_553 ();
 b15zdnd00an1n01x5 FILLER_234_555 ();
 b15zdnd11an1n64x5 FILLER_234_560 ();
 b15zdnd11an1n16x5 FILLER_234_624 ();
 b15zdnd00an1n02x5 FILLER_234_640 ();
 b15zdnd11an1n16x5 FILLER_234_662 ();
 b15zdnd00an1n02x5 FILLER_234_678 ();
 b15zdnd00an1n01x5 FILLER_234_680 ();
 b15zdnd11an1n32x5 FILLER_234_684 ();
 b15zdnd00an1n02x5 FILLER_234_716 ();
 b15zdnd11an1n64x5 FILLER_234_726 ();
 b15zdnd11an1n64x5 FILLER_234_790 ();
 b15zdnd11an1n64x5 FILLER_234_854 ();
 b15zdnd11an1n64x5 FILLER_234_918 ();
 b15zdnd11an1n64x5 FILLER_234_982 ();
 b15zdnd11an1n64x5 FILLER_234_1046 ();
 b15zdnd11an1n64x5 FILLER_234_1110 ();
 b15zdnd11an1n64x5 FILLER_234_1174 ();
 b15zdnd11an1n32x5 FILLER_234_1238 ();
 b15zdnd11an1n64x5 FILLER_234_1322 ();
 b15zdnd11an1n64x5 FILLER_234_1386 ();
 b15zdnd11an1n64x5 FILLER_234_1450 ();
 b15zdnd11an1n64x5 FILLER_234_1514 ();
 b15zdnd11an1n16x5 FILLER_234_1578 ();
 b15zdnd11an1n08x5 FILLER_234_1594 ();
 b15zdnd00an1n02x5 FILLER_234_1602 ();
 b15zdnd11an1n64x5 FILLER_234_1643 ();
 b15zdnd11an1n64x5 FILLER_234_1707 ();
 b15zdnd11an1n32x5 FILLER_234_1771 ();
 b15zdnd11an1n16x5 FILLER_234_1803 ();
 b15zdnd11an1n04x5 FILLER_234_1819 ();
 b15zdnd00an1n02x5 FILLER_234_1823 ();
 b15zdnd00an1n01x5 FILLER_234_1825 ();
 b15zdnd11an1n04x5 FILLER_234_1829 ();
 b15zdnd11an1n64x5 FILLER_234_1836 ();
 b15zdnd11an1n64x5 FILLER_234_1900 ();
 b15zdnd11an1n64x5 FILLER_234_1964 ();
 b15zdnd11an1n64x5 FILLER_234_2028 ();
 b15zdnd11an1n32x5 FILLER_234_2092 ();
 b15zdnd11an1n16x5 FILLER_234_2124 ();
 b15zdnd11an1n08x5 FILLER_234_2140 ();
 b15zdnd11an1n04x5 FILLER_234_2148 ();
 b15zdnd00an1n02x5 FILLER_234_2152 ();
 b15zdnd11an1n64x5 FILLER_234_2162 ();
 b15zdnd11an1n32x5 FILLER_234_2226 ();
 b15zdnd11an1n16x5 FILLER_234_2258 ();
 b15zdnd00an1n02x5 FILLER_234_2274 ();
 b15zdnd11an1n64x5 FILLER_235_0 ();
 b15zdnd11an1n32x5 FILLER_235_64 ();
 b15zdnd11an1n16x5 FILLER_235_96 ();
 b15zdnd00an1n01x5 FILLER_235_112 ();
 b15zdnd11an1n64x5 FILLER_235_116 ();
 b15zdnd11an1n64x5 FILLER_235_180 ();
 b15zdnd11an1n64x5 FILLER_235_244 ();
 b15zdnd11an1n64x5 FILLER_235_308 ();
 b15zdnd11an1n64x5 FILLER_235_372 ();
 b15zdnd11an1n64x5 FILLER_235_436 ();
 b15zdnd11an1n64x5 FILLER_235_500 ();
 b15zdnd11an1n32x5 FILLER_235_564 ();
 b15zdnd11an1n16x5 FILLER_235_596 ();
 b15zdnd11an1n08x5 FILLER_235_612 ();
 b15zdnd11an1n04x5 FILLER_235_620 ();
 b15zdnd00an1n01x5 FILLER_235_624 ();
 b15zdnd11an1n04x5 FILLER_235_665 ();
 b15zdnd11an1n64x5 FILLER_235_672 ();
 b15zdnd11an1n64x5 FILLER_235_736 ();
 b15zdnd11an1n64x5 FILLER_235_800 ();
 b15zdnd11an1n64x5 FILLER_235_864 ();
 b15zdnd11an1n32x5 FILLER_235_928 ();
 b15zdnd11an1n04x5 FILLER_235_960 ();
 b15zdnd00an1n02x5 FILLER_235_964 ();
 b15zdnd11an1n64x5 FILLER_235_973 ();
 b15zdnd11an1n32x5 FILLER_235_1037 ();
 b15zdnd11an1n16x5 FILLER_235_1069 ();
 b15zdnd11an1n64x5 FILLER_235_1124 ();
 b15zdnd11an1n64x5 FILLER_235_1188 ();
 b15zdnd11an1n32x5 FILLER_235_1252 ();
 b15zdnd11an1n08x5 FILLER_235_1284 ();
 b15zdnd11an1n04x5 FILLER_235_1292 ();
 b15zdnd11an1n64x5 FILLER_235_1299 ();
 b15zdnd11an1n64x5 FILLER_235_1363 ();
 b15zdnd11an1n64x5 FILLER_235_1427 ();
 b15zdnd11an1n64x5 FILLER_235_1491 ();
 b15zdnd11an1n32x5 FILLER_235_1555 ();
 b15zdnd11an1n16x5 FILLER_235_1587 ();
 b15zdnd11an1n08x5 FILLER_235_1603 ();
 b15zdnd00an1n02x5 FILLER_235_1611 ();
 b15zdnd00an1n01x5 FILLER_235_1613 ();
 b15zdnd11an1n08x5 FILLER_235_1621 ();
 b15zdnd11an1n04x5 FILLER_235_1629 ();
 b15zdnd11an1n64x5 FILLER_235_1644 ();
 b15zdnd11an1n16x5 FILLER_235_1708 ();
 b15zdnd00an1n02x5 FILLER_235_1724 ();
 b15zdnd00an1n01x5 FILLER_235_1726 ();
 b15zdnd11an1n32x5 FILLER_235_1754 ();
 b15zdnd11an1n16x5 FILLER_235_1786 ();
 b15zdnd11an1n04x5 FILLER_235_1802 ();
 b15zdnd11an1n64x5 FILLER_235_1858 ();
 b15zdnd11an1n64x5 FILLER_235_1922 ();
 b15zdnd11an1n64x5 FILLER_235_1986 ();
 b15zdnd11an1n64x5 FILLER_235_2050 ();
 b15zdnd11an1n64x5 FILLER_235_2114 ();
 b15zdnd11an1n64x5 FILLER_235_2178 ();
 b15zdnd11an1n32x5 FILLER_235_2242 ();
 b15zdnd11an1n08x5 FILLER_235_2274 ();
 b15zdnd00an1n02x5 FILLER_235_2282 ();
 b15zdnd11an1n16x5 FILLER_236_8 ();
 b15zdnd00an1n01x5 FILLER_236_24 ();
 b15zdnd11an1n64x5 FILLER_236_29 ();
 b15zdnd11an1n64x5 FILLER_236_93 ();
 b15zdnd11an1n64x5 FILLER_236_157 ();
 b15zdnd11an1n32x5 FILLER_236_221 ();
 b15zdnd11an1n16x5 FILLER_236_253 ();
 b15zdnd11an1n08x5 FILLER_236_269 ();
 b15zdnd11an1n04x5 FILLER_236_277 ();
 b15zdnd11an1n64x5 FILLER_236_323 ();
 b15zdnd11an1n64x5 FILLER_236_387 ();
 b15zdnd11an1n64x5 FILLER_236_451 ();
 b15zdnd11an1n64x5 FILLER_236_515 ();
 b15zdnd11an1n08x5 FILLER_236_579 ();
 b15zdnd00an1n02x5 FILLER_236_587 ();
 b15zdnd11an1n04x5 FILLER_236_629 ();
 b15zdnd11an1n16x5 FILLER_236_636 ();
 b15zdnd11an1n08x5 FILLER_236_652 ();
 b15zdnd00an1n01x5 FILLER_236_660 ();
 b15zdnd11an1n08x5 FILLER_236_664 ();
 b15zdnd00an1n02x5 FILLER_236_672 ();
 b15zdnd00an1n01x5 FILLER_236_674 ();
 b15zdnd11an1n32x5 FILLER_236_679 ();
 b15zdnd11an1n04x5 FILLER_236_711 ();
 b15zdnd00an1n02x5 FILLER_236_715 ();
 b15zdnd00an1n01x5 FILLER_236_717 ();
 b15zdnd11an1n64x5 FILLER_236_726 ();
 b15zdnd11an1n64x5 FILLER_236_790 ();
 b15zdnd11an1n16x5 FILLER_236_854 ();
 b15zdnd11an1n08x5 FILLER_236_870 ();
 b15zdnd11an1n04x5 FILLER_236_878 ();
 b15zdnd00an1n02x5 FILLER_236_882 ();
 b15zdnd11an1n32x5 FILLER_236_896 ();
 b15zdnd11an1n16x5 FILLER_236_928 ();
 b15zdnd00an1n02x5 FILLER_236_944 ();
 b15zdnd11an1n64x5 FILLER_236_985 ();
 b15zdnd11an1n64x5 FILLER_236_1052 ();
 b15zdnd11an1n64x5 FILLER_236_1116 ();
 b15zdnd11an1n64x5 FILLER_236_1180 ();
 b15zdnd11an1n64x5 FILLER_236_1244 ();
 b15zdnd11an1n64x5 FILLER_236_1308 ();
 b15zdnd11an1n64x5 FILLER_236_1372 ();
 b15zdnd11an1n08x5 FILLER_236_1436 ();
 b15zdnd11an1n04x5 FILLER_236_1444 ();
 b15zdnd00an1n02x5 FILLER_236_1448 ();
 b15zdnd00an1n01x5 FILLER_236_1450 ();
 b15zdnd11an1n08x5 FILLER_236_1456 ();
 b15zdnd00an1n01x5 FILLER_236_1464 ();
 b15zdnd11an1n64x5 FILLER_236_1468 ();
 b15zdnd11an1n32x5 FILLER_236_1532 ();
 b15zdnd11an1n08x5 FILLER_236_1564 ();
 b15zdnd00an1n02x5 FILLER_236_1572 ();
 b15zdnd00an1n01x5 FILLER_236_1574 ();
 b15zdnd11an1n08x5 FILLER_236_1586 ();
 b15zdnd11an1n04x5 FILLER_236_1594 ();
 b15zdnd11an1n64x5 FILLER_236_1608 ();
 b15zdnd11an1n16x5 FILLER_236_1672 ();
 b15zdnd00an1n02x5 FILLER_236_1688 ();
 b15zdnd00an1n01x5 FILLER_236_1690 ();
 b15zdnd11an1n16x5 FILLER_236_1743 ();
 b15zdnd11an1n04x5 FILLER_236_1759 ();
 b15zdnd00an1n02x5 FILLER_236_1763 ();
 b15zdnd11an1n16x5 FILLER_236_1807 ();
 b15zdnd11an1n08x5 FILLER_236_1823 ();
 b15zdnd11an1n04x5 FILLER_236_1834 ();
 b15zdnd11an1n64x5 FILLER_236_1841 ();
 b15zdnd11an1n64x5 FILLER_236_1905 ();
 b15zdnd11an1n64x5 FILLER_236_1969 ();
 b15zdnd11an1n64x5 FILLER_236_2033 ();
 b15zdnd11an1n32x5 FILLER_236_2097 ();
 b15zdnd11an1n16x5 FILLER_236_2129 ();
 b15zdnd11an1n08x5 FILLER_236_2145 ();
 b15zdnd00an1n01x5 FILLER_236_2153 ();
 b15zdnd11an1n32x5 FILLER_236_2162 ();
 b15zdnd11an1n08x5 FILLER_236_2194 ();
 b15zdnd11an1n04x5 FILLER_236_2205 ();
 b15zdnd11an1n64x5 FILLER_236_2212 ();
 b15zdnd11an1n64x5 FILLER_237_0 ();
 b15zdnd11an1n64x5 FILLER_237_64 ();
 b15zdnd11an1n16x5 FILLER_237_128 ();
 b15zdnd11an1n04x5 FILLER_237_144 ();
 b15zdnd00an1n02x5 FILLER_237_148 ();
 b15zdnd00an1n01x5 FILLER_237_150 ();
 b15zdnd11an1n64x5 FILLER_237_154 ();
 b15zdnd11an1n32x5 FILLER_237_218 ();
 b15zdnd11an1n08x5 FILLER_237_250 ();
 b15zdnd11an1n04x5 FILLER_237_258 ();
 b15zdnd00an1n01x5 FILLER_237_262 ();
 b15zdnd11an1n16x5 FILLER_237_269 ();
 b15zdnd11an1n04x5 FILLER_237_285 ();
 b15zdnd00an1n02x5 FILLER_237_289 ();
 b15zdnd11an1n32x5 FILLER_237_333 ();
 b15zdnd11an1n16x5 FILLER_237_365 ();
 b15zdnd11an1n64x5 FILLER_237_385 ();
 b15zdnd11an1n32x5 FILLER_237_449 ();
 b15zdnd11an1n16x5 FILLER_237_481 ();
 b15zdnd11an1n04x5 FILLER_237_497 ();
 b15zdnd00an1n02x5 FILLER_237_501 ();
 b15zdnd00an1n01x5 FILLER_237_503 ();
 b15zdnd11an1n64x5 FILLER_237_510 ();
 b15zdnd11an1n32x5 FILLER_237_574 ();
 b15zdnd11an1n16x5 FILLER_237_606 ();
 b15zdnd00an1n02x5 FILLER_237_622 ();
 b15zdnd00an1n01x5 FILLER_237_624 ();
 b15zdnd11an1n32x5 FILLER_237_628 ();
 b15zdnd11an1n16x5 FILLER_237_660 ();
 b15zdnd11an1n08x5 FILLER_237_676 ();
 b15zdnd11an1n04x5 FILLER_237_684 ();
 b15zdnd11an1n64x5 FILLER_237_730 ();
 b15zdnd11an1n64x5 FILLER_237_794 ();
 b15zdnd11an1n32x5 FILLER_237_858 ();
 b15zdnd00an1n02x5 FILLER_237_890 ();
 b15zdnd00an1n01x5 FILLER_237_892 ();
 b15zdnd11an1n16x5 FILLER_237_900 ();
 b15zdnd11an1n08x5 FILLER_237_916 ();
 b15zdnd11an1n04x5 FILLER_237_924 ();
 b15zdnd00an1n01x5 FILLER_237_928 ();
 b15zdnd11an1n04x5 FILLER_237_940 ();
 b15zdnd11an1n32x5 FILLER_237_949 ();
 b15zdnd11an1n16x5 FILLER_237_981 ();
 b15zdnd11an1n08x5 FILLER_237_997 ();
 b15zdnd11an1n04x5 FILLER_237_1005 ();
 b15zdnd00an1n01x5 FILLER_237_1009 ();
 b15zdnd11an1n04x5 FILLER_237_1018 ();
 b15zdnd11an1n64x5 FILLER_237_1074 ();
 b15zdnd11an1n16x5 FILLER_237_1138 ();
 b15zdnd11an1n08x5 FILLER_237_1154 ();
 b15zdnd00an1n01x5 FILLER_237_1162 ();
 b15zdnd11an1n64x5 FILLER_237_1205 ();
 b15zdnd11an1n64x5 FILLER_237_1269 ();
 b15zdnd11an1n64x5 FILLER_237_1333 ();
 b15zdnd11an1n32x5 FILLER_237_1397 ();
 b15zdnd11an1n16x5 FILLER_237_1429 ();
 b15zdnd00an1n01x5 FILLER_237_1445 ();
 b15zdnd11an1n04x5 FILLER_237_1459 ();
 b15zdnd00an1n01x5 FILLER_237_1463 ();
 b15zdnd11an1n04x5 FILLER_237_1474 ();
 b15zdnd11an1n32x5 FILLER_237_1484 ();
 b15zdnd11an1n08x5 FILLER_237_1516 ();
 b15zdnd00an1n02x5 FILLER_237_1524 ();
 b15zdnd00an1n01x5 FILLER_237_1526 ();
 b15zdnd11an1n08x5 FILLER_237_1569 ();
 b15zdnd00an1n02x5 FILLER_237_1577 ();
 b15zdnd11an1n16x5 FILLER_237_1582 ();
 b15zdnd11an1n04x5 FILLER_237_1598 ();
 b15zdnd00an1n02x5 FILLER_237_1602 ();
 b15zdnd11an1n64x5 FILLER_237_1608 ();
 b15zdnd11an1n32x5 FILLER_237_1672 ();
 b15zdnd00an1n02x5 FILLER_237_1704 ();
 b15zdnd00an1n01x5 FILLER_237_1706 ();
 b15zdnd11an1n04x5 FILLER_237_1710 ();
 b15zdnd11an1n04x5 FILLER_237_1717 ();
 b15zdnd00an1n01x5 FILLER_237_1721 ();
 b15zdnd11an1n04x5 FILLER_237_1726 ();
 b15zdnd00an1n02x5 FILLER_237_1730 ();
 b15zdnd00an1n01x5 FILLER_237_1732 ();
 b15zdnd11an1n64x5 FILLER_237_1741 ();
 b15zdnd11an1n64x5 FILLER_237_1805 ();
 b15zdnd11an1n64x5 FILLER_237_1869 ();
 b15zdnd11an1n64x5 FILLER_237_1933 ();
 b15zdnd11an1n64x5 FILLER_237_1997 ();
 b15zdnd11an1n64x5 FILLER_237_2061 ();
 b15zdnd11an1n32x5 FILLER_237_2125 ();
 b15zdnd11an1n08x5 FILLER_237_2157 ();
 b15zdnd11an1n04x5 FILLER_237_2165 ();
 b15zdnd00an1n01x5 FILLER_237_2169 ();
 b15zdnd11an1n64x5 FILLER_237_2210 ();
 b15zdnd11an1n08x5 FILLER_237_2274 ();
 b15zdnd00an1n02x5 FILLER_237_2282 ();
 b15zdnd11an1n64x5 FILLER_238_8 ();
 b15zdnd11an1n32x5 FILLER_238_72 ();
 b15zdnd11an1n08x5 FILLER_238_104 ();
 b15zdnd11an1n16x5 FILLER_238_118 ();
 b15zdnd11an1n08x5 FILLER_238_134 ();
 b15zdnd11an1n04x5 FILLER_238_142 ();
 b15zdnd00an1n02x5 FILLER_238_146 ();
 b15zdnd00an1n01x5 FILLER_238_148 ();
 b15zdnd11an1n08x5 FILLER_238_152 ();
 b15zdnd00an1n02x5 FILLER_238_160 ();
 b15zdnd11an1n64x5 FILLER_238_165 ();
 b15zdnd11an1n64x5 FILLER_238_229 ();
 b15zdnd11an1n64x5 FILLER_238_293 ();
 b15zdnd11an1n32x5 FILLER_238_357 ();
 b15zdnd00an1n02x5 FILLER_238_389 ();
 b15zdnd00an1n01x5 FILLER_238_391 ();
 b15zdnd11an1n16x5 FILLER_238_395 ();
 b15zdnd00an1n02x5 FILLER_238_411 ();
 b15zdnd11an1n64x5 FILLER_238_444 ();
 b15zdnd11an1n64x5 FILLER_238_508 ();
 b15zdnd11an1n64x5 FILLER_238_572 ();
 b15zdnd11an1n64x5 FILLER_238_636 ();
 b15zdnd11an1n16x5 FILLER_238_700 ();
 b15zdnd00an1n02x5 FILLER_238_716 ();
 b15zdnd11an1n64x5 FILLER_238_726 ();
 b15zdnd11an1n64x5 FILLER_238_790 ();
 b15zdnd11an1n64x5 FILLER_238_854 ();
 b15zdnd11an1n08x5 FILLER_238_918 ();
 b15zdnd11an1n04x5 FILLER_238_926 ();
 b15zdnd00an1n02x5 FILLER_238_930 ();
 b15zdnd00an1n01x5 FILLER_238_932 ();
 b15zdnd11an1n16x5 FILLER_238_936 ();
 b15zdnd11an1n08x5 FILLER_238_952 ();
 b15zdnd00an1n01x5 FILLER_238_960 ();
 b15zdnd11an1n08x5 FILLER_238_972 ();
 b15zdnd11an1n04x5 FILLER_238_985 ();
 b15zdnd11an1n08x5 FILLER_238_1028 ();
 b15zdnd11an1n04x5 FILLER_238_1036 ();
 b15zdnd11an1n04x5 FILLER_238_1043 ();
 b15zdnd11an1n64x5 FILLER_238_1050 ();
 b15zdnd11an1n64x5 FILLER_238_1114 ();
 b15zdnd11an1n64x5 FILLER_238_1178 ();
 b15zdnd11an1n64x5 FILLER_238_1242 ();
 b15zdnd11an1n64x5 FILLER_238_1306 ();
 b15zdnd11an1n64x5 FILLER_238_1370 ();
 b15zdnd11an1n64x5 FILLER_238_1434 ();
 b15zdnd11an1n32x5 FILLER_238_1498 ();
 b15zdnd11an1n16x5 FILLER_238_1530 ();
 b15zdnd11an1n08x5 FILLER_238_1546 ();
 b15zdnd11an1n64x5 FILLER_238_1606 ();
 b15zdnd11an1n32x5 FILLER_238_1670 ();
 b15zdnd11an1n08x5 FILLER_238_1702 ();
 b15zdnd11an1n04x5 FILLER_238_1710 ();
 b15zdnd00an1n02x5 FILLER_238_1714 ();
 b15zdnd11an1n64x5 FILLER_238_1719 ();
 b15zdnd11an1n64x5 FILLER_238_1783 ();
 b15zdnd11an1n64x5 FILLER_238_1847 ();
 b15zdnd11an1n64x5 FILLER_238_1911 ();
 b15zdnd11an1n64x5 FILLER_238_1975 ();
 b15zdnd11an1n64x5 FILLER_238_2039 ();
 b15zdnd11an1n32x5 FILLER_238_2103 ();
 b15zdnd11an1n16x5 FILLER_238_2135 ();
 b15zdnd00an1n02x5 FILLER_238_2151 ();
 b15zdnd00an1n01x5 FILLER_238_2153 ();
 b15zdnd11an1n64x5 FILLER_238_2162 ();
 b15zdnd11an1n32x5 FILLER_238_2226 ();
 b15zdnd11an1n16x5 FILLER_238_2258 ();
 b15zdnd00an1n02x5 FILLER_238_2274 ();
 b15zdnd00an1n02x5 FILLER_239_0 ();
 b15zdnd11an1n04x5 FILLER_239_6 ();
 b15zdnd11an1n16x5 FILLER_239_18 ();
 b15zdnd11an1n04x5 FILLER_239_34 ();
 b15zdnd11an1n32x5 FILLER_239_52 ();
 b15zdnd11an1n16x5 FILLER_239_84 ();
 b15zdnd11an1n08x5 FILLER_239_100 ();
 b15zdnd00an1n02x5 FILLER_239_108 ();
 b15zdnd11an1n04x5 FILLER_239_114 ();
 b15zdnd11an1n04x5 FILLER_239_122 ();
 b15zdnd11an1n64x5 FILLER_239_178 ();
 b15zdnd11an1n64x5 FILLER_239_242 ();
 b15zdnd11an1n64x5 FILLER_239_306 ();
 b15zdnd11an1n08x5 FILLER_239_370 ();
 b15zdnd11an1n64x5 FILLER_239_420 ();
 b15zdnd11an1n64x5 FILLER_239_484 ();
 b15zdnd11an1n64x5 FILLER_239_548 ();
 b15zdnd11an1n64x5 FILLER_239_612 ();
 b15zdnd11an1n64x5 FILLER_239_676 ();
 b15zdnd11an1n64x5 FILLER_239_740 ();
 b15zdnd11an1n64x5 FILLER_239_804 ();
 b15zdnd11an1n16x5 FILLER_239_868 ();
 b15zdnd11an1n08x5 FILLER_239_884 ();
 b15zdnd00an1n02x5 FILLER_239_892 ();
 b15zdnd00an1n01x5 FILLER_239_894 ();
 b15zdnd11an1n16x5 FILLER_239_935 ();
 b15zdnd11an1n04x5 FILLER_239_951 ();
 b15zdnd00an1n01x5 FILLER_239_955 ();
 b15zdnd11an1n64x5 FILLER_239_977 ();
 b15zdnd11an1n32x5 FILLER_239_1041 ();
 b15zdnd11an1n04x5 FILLER_239_1073 ();
 b15zdnd11an1n64x5 FILLER_239_1081 ();
 b15zdnd11an1n64x5 FILLER_239_1145 ();
 b15zdnd11an1n64x5 FILLER_239_1209 ();
 b15zdnd11an1n64x5 FILLER_239_1273 ();
 b15zdnd11an1n64x5 FILLER_239_1337 ();
 b15zdnd11an1n32x5 FILLER_239_1401 ();
 b15zdnd11an1n16x5 FILLER_239_1433 ();
 b15zdnd11an1n64x5 FILLER_239_1458 ();
 b15zdnd11an1n32x5 FILLER_239_1522 ();
 b15zdnd11an1n16x5 FILLER_239_1554 ();
 b15zdnd11an1n08x5 FILLER_239_1570 ();
 b15zdnd00an1n01x5 FILLER_239_1578 ();
 b15zdnd11an1n04x5 FILLER_239_1582 ();
 b15zdnd11an1n32x5 FILLER_239_1589 ();
 b15zdnd11an1n08x5 FILLER_239_1621 ();
 b15zdnd00an1n02x5 FILLER_239_1629 ();
 b15zdnd11an1n64x5 FILLER_239_1634 ();
 b15zdnd11an1n64x5 FILLER_239_1698 ();
 b15zdnd11an1n64x5 FILLER_239_1762 ();
 b15zdnd11an1n16x5 FILLER_239_1826 ();
 b15zdnd11an1n08x5 FILLER_239_1842 ();
 b15zdnd11an1n04x5 FILLER_239_1850 ();
 b15zdnd11an1n64x5 FILLER_239_1896 ();
 b15zdnd11an1n64x5 FILLER_239_1960 ();
 b15zdnd11an1n64x5 FILLER_239_2024 ();
 b15zdnd11an1n64x5 FILLER_239_2088 ();
 b15zdnd11an1n64x5 FILLER_239_2152 ();
 b15zdnd11an1n64x5 FILLER_239_2216 ();
 b15zdnd11an1n04x5 FILLER_239_2280 ();
 b15zdnd11an1n16x5 FILLER_240_8 ();
 b15zdnd11an1n04x5 FILLER_240_24 ();
 b15zdnd11an1n64x5 FILLER_240_42 ();
 b15zdnd11an1n64x5 FILLER_240_106 ();
 b15zdnd11an1n64x5 FILLER_240_170 ();
 b15zdnd11an1n64x5 FILLER_240_234 ();
 b15zdnd11an1n64x5 FILLER_240_298 ();
 b15zdnd11an1n08x5 FILLER_240_362 ();
 b15zdnd00an1n02x5 FILLER_240_370 ();
 b15zdnd11an1n08x5 FILLER_240_424 ();
 b15zdnd11an1n04x5 FILLER_240_432 ();
 b15zdnd00an1n02x5 FILLER_240_436 ();
 b15zdnd11an1n64x5 FILLER_240_444 ();
 b15zdnd11an1n16x5 FILLER_240_508 ();
 b15zdnd00an1n02x5 FILLER_240_524 ();
 b15zdnd11an1n64x5 FILLER_240_568 ();
 b15zdnd11an1n64x5 FILLER_240_632 ();
 b15zdnd11an1n16x5 FILLER_240_696 ();
 b15zdnd11an1n04x5 FILLER_240_712 ();
 b15zdnd00an1n02x5 FILLER_240_716 ();
 b15zdnd11an1n64x5 FILLER_240_726 ();
 b15zdnd11an1n64x5 FILLER_240_790 ();
 b15zdnd11an1n64x5 FILLER_240_854 ();
 b15zdnd11an1n08x5 FILLER_240_918 ();
 b15zdnd11an1n04x5 FILLER_240_926 ();
 b15zdnd00an1n01x5 FILLER_240_930 ();
 b15zdnd11an1n16x5 FILLER_240_934 ();
 b15zdnd11an1n04x5 FILLER_240_950 ();
 b15zdnd11an1n64x5 FILLER_240_958 ();
 b15zdnd11an1n64x5 FILLER_240_1022 ();
 b15zdnd11an1n64x5 FILLER_240_1086 ();
 b15zdnd11an1n64x5 FILLER_240_1150 ();
 b15zdnd11an1n64x5 FILLER_240_1214 ();
 b15zdnd11an1n64x5 FILLER_240_1278 ();
 b15zdnd11an1n64x5 FILLER_240_1342 ();
 b15zdnd11an1n32x5 FILLER_240_1406 ();
 b15zdnd11an1n08x5 FILLER_240_1438 ();
 b15zdnd11an1n04x5 FILLER_240_1446 ();
 b15zdnd00an1n01x5 FILLER_240_1450 ();
 b15zdnd11an1n64x5 FILLER_240_1465 ();
 b15zdnd11an1n32x5 FILLER_240_1529 ();
 b15zdnd11an1n16x5 FILLER_240_1561 ();
 b15zdnd11an1n64x5 FILLER_240_1616 ();
 b15zdnd11an1n64x5 FILLER_240_1680 ();
 b15zdnd11an1n64x5 FILLER_240_1744 ();
 b15zdnd11an1n64x5 FILLER_240_1808 ();
 b15zdnd11an1n64x5 FILLER_240_1872 ();
 b15zdnd11an1n64x5 FILLER_240_1936 ();
 b15zdnd11an1n64x5 FILLER_240_2000 ();
 b15zdnd11an1n64x5 FILLER_240_2064 ();
 b15zdnd11an1n16x5 FILLER_240_2128 ();
 b15zdnd11an1n08x5 FILLER_240_2144 ();
 b15zdnd00an1n02x5 FILLER_240_2152 ();
 b15zdnd11an1n64x5 FILLER_240_2162 ();
 b15zdnd11an1n32x5 FILLER_240_2226 ();
 b15zdnd11an1n16x5 FILLER_240_2258 ();
 b15zdnd00an1n02x5 FILLER_240_2274 ();
 b15zdnd11an1n16x5 FILLER_241_0 ();
 b15zdnd11an1n04x5 FILLER_241_16 ();
 b15zdnd00an1n02x5 FILLER_241_20 ();
 b15zdnd11an1n64x5 FILLER_241_30 ();
 b15zdnd11an1n64x5 FILLER_241_94 ();
 b15zdnd11an1n64x5 FILLER_241_158 ();
 b15zdnd11an1n64x5 FILLER_241_222 ();
 b15zdnd11an1n08x5 FILLER_241_286 ();
 b15zdnd11an1n04x5 FILLER_241_294 ();
 b15zdnd00an1n02x5 FILLER_241_298 ();
 b15zdnd00an1n01x5 FILLER_241_300 ();
 b15zdnd11an1n64x5 FILLER_241_310 ();
 b15zdnd11an1n16x5 FILLER_241_374 ();
 b15zdnd00an1n02x5 FILLER_241_390 ();
 b15zdnd11an1n04x5 FILLER_241_395 ();
 b15zdnd11an1n64x5 FILLER_241_402 ();
 b15zdnd11an1n32x5 FILLER_241_466 ();
 b15zdnd11an1n08x5 FILLER_241_498 ();
 b15zdnd11an1n04x5 FILLER_241_506 ();
 b15zdnd11an1n64x5 FILLER_241_513 ();
 b15zdnd11an1n64x5 FILLER_241_577 ();
 b15zdnd11an1n64x5 FILLER_241_641 ();
 b15zdnd11an1n16x5 FILLER_241_705 ();
 b15zdnd11an1n08x5 FILLER_241_721 ();
 b15zdnd11an1n04x5 FILLER_241_729 ();
 b15zdnd00an1n01x5 FILLER_241_733 ();
 b15zdnd11an1n64x5 FILLER_241_752 ();
 b15zdnd11an1n64x5 FILLER_241_816 ();
 b15zdnd11an1n64x5 FILLER_241_880 ();
 b15zdnd11an1n64x5 FILLER_241_944 ();
 b15zdnd11an1n64x5 FILLER_241_1008 ();
 b15zdnd11an1n64x5 FILLER_241_1072 ();
 b15zdnd11an1n32x5 FILLER_241_1136 ();
 b15zdnd11an1n16x5 FILLER_241_1168 ();
 b15zdnd00an1n02x5 FILLER_241_1184 ();
 b15zdnd11an1n04x5 FILLER_241_1197 ();
 b15zdnd11an1n64x5 FILLER_241_1211 ();
 b15zdnd11an1n64x5 FILLER_241_1275 ();
 b15zdnd11an1n64x5 FILLER_241_1339 ();
 b15zdnd11an1n32x5 FILLER_241_1403 ();
 b15zdnd11an1n16x5 FILLER_241_1435 ();
 b15zdnd00an1n02x5 FILLER_241_1451 ();
 b15zdnd11an1n04x5 FILLER_241_1458 ();
 b15zdnd00an1n02x5 FILLER_241_1462 ();
 b15zdnd00an1n01x5 FILLER_241_1464 ();
 b15zdnd11an1n64x5 FILLER_241_1469 ();
 b15zdnd11an1n32x5 FILLER_241_1533 ();
 b15zdnd11an1n16x5 FILLER_241_1565 ();
 b15zdnd11an1n08x5 FILLER_241_1581 ();
 b15zdnd11an1n04x5 FILLER_241_1589 ();
 b15zdnd11an1n64x5 FILLER_241_1635 ();
 b15zdnd11an1n64x5 FILLER_241_1699 ();
 b15zdnd11an1n64x5 FILLER_241_1763 ();
 b15zdnd11an1n64x5 FILLER_241_1827 ();
 b15zdnd11an1n64x5 FILLER_241_1891 ();
 b15zdnd11an1n64x5 FILLER_241_1955 ();
 b15zdnd11an1n64x5 FILLER_241_2019 ();
 b15zdnd11an1n64x5 FILLER_241_2083 ();
 b15zdnd11an1n64x5 FILLER_241_2147 ();
 b15zdnd11an1n64x5 FILLER_241_2211 ();
 b15zdnd11an1n08x5 FILLER_241_2275 ();
 b15zdnd00an1n01x5 FILLER_241_2283 ();
 b15zdnd11an1n64x5 FILLER_242_8 ();
 b15zdnd11an1n32x5 FILLER_242_72 ();
 b15zdnd11an1n04x5 FILLER_242_104 ();
 b15zdnd00an1n02x5 FILLER_242_108 ();
 b15zdnd00an1n01x5 FILLER_242_110 ();
 b15zdnd11an1n64x5 FILLER_242_114 ();
 b15zdnd11an1n64x5 FILLER_242_178 ();
 b15zdnd11an1n32x5 FILLER_242_242 ();
 b15zdnd11an1n16x5 FILLER_242_274 ();
 b15zdnd11an1n04x5 FILLER_242_290 ();
 b15zdnd00an1n02x5 FILLER_242_294 ();
 b15zdnd11an1n04x5 FILLER_242_300 ();
 b15zdnd11an1n64x5 FILLER_242_307 ();
 b15zdnd11an1n64x5 FILLER_242_371 ();
 b15zdnd11an1n64x5 FILLER_242_435 ();
 b15zdnd11an1n04x5 FILLER_242_499 ();
 b15zdnd00an1n01x5 FILLER_242_503 ();
 b15zdnd11an1n64x5 FILLER_242_546 ();
 b15zdnd11an1n64x5 FILLER_242_610 ();
 b15zdnd11an1n32x5 FILLER_242_674 ();
 b15zdnd11an1n08x5 FILLER_242_706 ();
 b15zdnd11an1n04x5 FILLER_242_714 ();
 b15zdnd11an1n32x5 FILLER_242_726 ();
 b15zdnd11an1n16x5 FILLER_242_758 ();
 b15zdnd11an1n08x5 FILLER_242_774 ();
 b15zdnd11an1n64x5 FILLER_242_788 ();
 b15zdnd11an1n64x5 FILLER_242_852 ();
 b15zdnd11an1n64x5 FILLER_242_916 ();
 b15zdnd11an1n64x5 FILLER_242_980 ();
 b15zdnd11an1n64x5 FILLER_242_1044 ();
 b15zdnd11an1n32x5 FILLER_242_1108 ();
 b15zdnd11an1n16x5 FILLER_242_1140 ();
 b15zdnd11an1n04x5 FILLER_242_1156 ();
 b15zdnd11an1n04x5 FILLER_242_1200 ();
 b15zdnd00an1n02x5 FILLER_242_1204 ();
 b15zdnd00an1n01x5 FILLER_242_1206 ();
 b15zdnd11an1n64x5 FILLER_242_1211 ();
 b15zdnd11an1n64x5 FILLER_242_1275 ();
 b15zdnd11an1n64x5 FILLER_242_1339 ();
 b15zdnd11an1n64x5 FILLER_242_1403 ();
 b15zdnd11an1n64x5 FILLER_242_1467 ();
 b15zdnd11an1n32x5 FILLER_242_1531 ();
 b15zdnd11an1n16x5 FILLER_242_1563 ();
 b15zdnd11an1n04x5 FILLER_242_1579 ();
 b15zdnd11an1n04x5 FILLER_242_1608 ();
 b15zdnd11an1n64x5 FILLER_242_1643 ();
 b15zdnd11an1n64x5 FILLER_242_1707 ();
 b15zdnd11an1n64x5 FILLER_242_1771 ();
 b15zdnd11an1n64x5 FILLER_242_1835 ();
 b15zdnd11an1n64x5 FILLER_242_1899 ();
 b15zdnd11an1n64x5 FILLER_242_1963 ();
 b15zdnd11an1n64x5 FILLER_242_2027 ();
 b15zdnd11an1n32x5 FILLER_242_2091 ();
 b15zdnd11an1n16x5 FILLER_242_2123 ();
 b15zdnd11an1n08x5 FILLER_242_2139 ();
 b15zdnd11an1n04x5 FILLER_242_2147 ();
 b15zdnd00an1n02x5 FILLER_242_2151 ();
 b15zdnd00an1n01x5 FILLER_242_2153 ();
 b15zdnd11an1n64x5 FILLER_242_2162 ();
 b15zdnd11an1n32x5 FILLER_242_2226 ();
 b15zdnd11an1n16x5 FILLER_242_2258 ();
 b15zdnd00an1n02x5 FILLER_242_2274 ();
 b15zdnd11an1n64x5 FILLER_243_0 ();
 b15zdnd11an1n64x5 FILLER_243_64 ();
 b15zdnd11an1n16x5 FILLER_243_128 ();
 b15zdnd11an1n04x5 FILLER_243_144 ();
 b15zdnd11an1n64x5 FILLER_243_190 ();
 b15zdnd11an1n64x5 FILLER_243_254 ();
 b15zdnd11an1n64x5 FILLER_243_318 ();
 b15zdnd11an1n64x5 FILLER_243_382 ();
 b15zdnd11an1n64x5 FILLER_243_446 ();
 b15zdnd11an1n64x5 FILLER_243_515 ();
 b15zdnd11an1n64x5 FILLER_243_579 ();
 b15zdnd11an1n32x5 FILLER_243_643 ();
 b15zdnd11an1n08x5 FILLER_243_675 ();
 b15zdnd11an1n04x5 FILLER_243_683 ();
 b15zdnd00an1n02x5 FILLER_243_687 ();
 b15zdnd00an1n01x5 FILLER_243_689 ();
 b15zdnd11an1n64x5 FILLER_243_695 ();
 b15zdnd11an1n64x5 FILLER_243_759 ();
 b15zdnd11an1n64x5 FILLER_243_823 ();
 b15zdnd11an1n64x5 FILLER_243_887 ();
 b15zdnd11an1n04x5 FILLER_243_951 ();
 b15zdnd00an1n01x5 FILLER_243_955 ();
 b15zdnd11an1n64x5 FILLER_243_998 ();
 b15zdnd11an1n64x5 FILLER_243_1062 ();
 b15zdnd11an1n32x5 FILLER_243_1126 ();
 b15zdnd11an1n08x5 FILLER_243_1158 ();
 b15zdnd11an1n04x5 FILLER_243_1166 ();
 b15zdnd11an1n04x5 FILLER_243_1184 ();
 b15zdnd11an1n04x5 FILLER_243_1191 ();
 b15zdnd00an1n01x5 FILLER_243_1195 ();
 b15zdnd11an1n64x5 FILLER_243_1199 ();
 b15zdnd11an1n64x5 FILLER_243_1263 ();
 b15zdnd11an1n64x5 FILLER_243_1327 ();
 b15zdnd11an1n64x5 FILLER_243_1391 ();
 b15zdnd11an1n64x5 FILLER_243_1455 ();
 b15zdnd11an1n64x5 FILLER_243_1519 ();
 b15zdnd11an1n64x5 FILLER_243_1583 ();
 b15zdnd11an1n64x5 FILLER_243_1647 ();
 b15zdnd11an1n64x5 FILLER_243_1711 ();
 b15zdnd11an1n08x5 FILLER_243_1775 ();
 b15zdnd11an1n64x5 FILLER_243_1810 ();
 b15zdnd11an1n64x5 FILLER_243_1874 ();
 b15zdnd11an1n16x5 FILLER_243_1938 ();
 b15zdnd11an1n04x5 FILLER_243_1954 ();
 b15zdnd00an1n01x5 FILLER_243_1958 ();
 b15zdnd11an1n64x5 FILLER_243_1974 ();
 b15zdnd11an1n64x5 FILLER_243_2038 ();
 b15zdnd11an1n64x5 FILLER_243_2102 ();
 b15zdnd11an1n64x5 FILLER_243_2166 ();
 b15zdnd11an1n32x5 FILLER_243_2230 ();
 b15zdnd11an1n16x5 FILLER_243_2262 ();
 b15zdnd11an1n04x5 FILLER_243_2278 ();
 b15zdnd00an1n02x5 FILLER_243_2282 ();
 b15zdnd11an1n64x5 FILLER_244_8 ();
 b15zdnd11an1n64x5 FILLER_244_72 ();
 b15zdnd11an1n64x5 FILLER_244_136 ();
 b15zdnd11an1n64x5 FILLER_244_200 ();
 b15zdnd11an1n64x5 FILLER_244_264 ();
 b15zdnd11an1n64x5 FILLER_244_328 ();
 b15zdnd11an1n64x5 FILLER_244_392 ();
 b15zdnd11an1n32x5 FILLER_244_456 ();
 b15zdnd11an1n16x5 FILLER_244_488 ();
 b15zdnd11an1n04x5 FILLER_244_504 ();
 b15zdnd11an1n16x5 FILLER_244_512 ();
 b15zdnd00an1n01x5 FILLER_244_528 ();
 b15zdnd11an1n64x5 FILLER_244_571 ();
 b15zdnd11an1n64x5 FILLER_244_635 ();
 b15zdnd11an1n16x5 FILLER_244_699 ();
 b15zdnd00an1n02x5 FILLER_244_715 ();
 b15zdnd00an1n01x5 FILLER_244_717 ();
 b15zdnd11an1n64x5 FILLER_244_726 ();
 b15zdnd11an1n64x5 FILLER_244_790 ();
 b15zdnd11an1n64x5 FILLER_244_854 ();
 b15zdnd11an1n64x5 FILLER_244_918 ();
 b15zdnd11an1n64x5 FILLER_244_982 ();
 b15zdnd11an1n64x5 FILLER_244_1046 ();
 b15zdnd11an1n64x5 FILLER_244_1110 ();
 b15zdnd11an1n08x5 FILLER_244_1174 ();
 b15zdnd11an1n04x5 FILLER_244_1182 ();
 b15zdnd11an1n64x5 FILLER_244_1206 ();
 b15zdnd11an1n64x5 FILLER_244_1270 ();
 b15zdnd11an1n32x5 FILLER_244_1334 ();
 b15zdnd11an1n16x5 FILLER_244_1366 ();
 b15zdnd11an1n04x5 FILLER_244_1382 ();
 b15zdnd11an1n32x5 FILLER_244_1395 ();
 b15zdnd11an1n16x5 FILLER_244_1427 ();
 b15zdnd11an1n08x5 FILLER_244_1443 ();
 b15zdnd11an1n04x5 FILLER_244_1451 ();
 b15zdnd11an1n04x5 FILLER_244_1461 ();
 b15zdnd11an1n04x5 FILLER_244_1470 ();
 b15zdnd11an1n64x5 FILLER_244_1477 ();
 b15zdnd11an1n64x5 FILLER_244_1541 ();
 b15zdnd11an1n64x5 FILLER_244_1605 ();
 b15zdnd11an1n32x5 FILLER_244_1669 ();
 b15zdnd11an1n08x5 FILLER_244_1701 ();
 b15zdnd11an1n04x5 FILLER_244_1709 ();
 b15zdnd00an1n02x5 FILLER_244_1713 ();
 b15zdnd11an1n16x5 FILLER_244_1757 ();
 b15zdnd11an1n08x5 FILLER_244_1773 ();
 b15zdnd11an1n04x5 FILLER_244_1781 ();
 b15zdnd00an1n01x5 FILLER_244_1785 ();
 b15zdnd11an1n64x5 FILLER_244_1790 ();
 b15zdnd11an1n64x5 FILLER_244_1854 ();
 b15zdnd11an1n64x5 FILLER_244_1918 ();
 b15zdnd11an1n64x5 FILLER_244_1982 ();
 b15zdnd11an1n64x5 FILLER_244_2046 ();
 b15zdnd11an1n32x5 FILLER_244_2110 ();
 b15zdnd11an1n08x5 FILLER_244_2142 ();
 b15zdnd11an1n04x5 FILLER_244_2150 ();
 b15zdnd11an1n64x5 FILLER_244_2162 ();
 b15zdnd11an1n32x5 FILLER_244_2226 ();
 b15zdnd11an1n16x5 FILLER_244_2258 ();
 b15zdnd00an1n02x5 FILLER_244_2274 ();
 b15zdnd11an1n64x5 FILLER_245_0 ();
 b15zdnd11an1n64x5 FILLER_245_64 ();
 b15zdnd11an1n64x5 FILLER_245_128 ();
 b15zdnd11an1n64x5 FILLER_245_192 ();
 b15zdnd11an1n32x5 FILLER_245_256 ();
 b15zdnd11an1n08x5 FILLER_245_288 ();
 b15zdnd11an1n04x5 FILLER_245_296 ();
 b15zdnd00an1n02x5 FILLER_245_300 ();
 b15zdnd11an1n64x5 FILLER_245_314 ();
 b15zdnd11an1n64x5 FILLER_245_378 ();
 b15zdnd11an1n32x5 FILLER_245_442 ();
 b15zdnd11an1n16x5 FILLER_245_474 ();
 b15zdnd11an1n04x5 FILLER_245_490 ();
 b15zdnd00an1n02x5 FILLER_245_494 ();
 b15zdnd00an1n01x5 FILLER_245_496 ();
 b15zdnd11an1n64x5 FILLER_245_549 ();
 b15zdnd11an1n64x5 FILLER_245_613 ();
 b15zdnd11an1n64x5 FILLER_245_677 ();
 b15zdnd11an1n64x5 FILLER_245_741 ();
 b15zdnd11an1n64x5 FILLER_245_805 ();
 b15zdnd11an1n64x5 FILLER_245_869 ();
 b15zdnd11an1n64x5 FILLER_245_933 ();
 b15zdnd11an1n64x5 FILLER_245_997 ();
 b15zdnd11an1n64x5 FILLER_245_1061 ();
 b15zdnd11an1n64x5 FILLER_245_1125 ();
 b15zdnd11an1n64x5 FILLER_245_1189 ();
 b15zdnd11an1n64x5 FILLER_245_1253 ();
 b15zdnd11an1n64x5 FILLER_245_1317 ();
 b15zdnd11an1n64x5 FILLER_245_1381 ();
 b15zdnd11an1n08x5 FILLER_245_1445 ();
 b15zdnd11an1n04x5 FILLER_245_1453 ();
 b15zdnd00an1n02x5 FILLER_245_1457 ();
 b15zdnd00an1n01x5 FILLER_245_1459 ();
 b15zdnd11an1n64x5 FILLER_245_1502 ();
 b15zdnd11an1n16x5 FILLER_245_1566 ();
 b15zdnd11an1n04x5 FILLER_245_1582 ();
 b15zdnd00an1n02x5 FILLER_245_1586 ();
 b15zdnd11an1n64x5 FILLER_245_1627 ();
 b15zdnd11an1n64x5 FILLER_245_1691 ();
 b15zdnd11an1n32x5 FILLER_245_1755 ();
 b15zdnd11an1n04x5 FILLER_245_1787 ();
 b15zdnd00an1n02x5 FILLER_245_1791 ();
 b15zdnd11an1n64x5 FILLER_245_1809 ();
 b15zdnd11an1n64x5 FILLER_245_1873 ();
 b15zdnd11an1n64x5 FILLER_245_1937 ();
 b15zdnd11an1n16x5 FILLER_245_2001 ();
 b15zdnd11an1n08x5 FILLER_245_2017 ();
 b15zdnd11an1n04x5 FILLER_245_2025 ();
 b15zdnd11an1n64x5 FILLER_245_2038 ();
 b15zdnd11an1n64x5 FILLER_245_2102 ();
 b15zdnd11an1n64x5 FILLER_245_2166 ();
 b15zdnd11an1n32x5 FILLER_245_2230 ();
 b15zdnd11an1n16x5 FILLER_245_2262 ();
 b15zdnd11an1n04x5 FILLER_245_2278 ();
 b15zdnd00an1n02x5 FILLER_245_2282 ();
 b15zdnd11an1n64x5 FILLER_246_8 ();
 b15zdnd11an1n16x5 FILLER_246_72 ();
 b15zdnd11an1n04x5 FILLER_246_88 ();
 b15zdnd11an1n04x5 FILLER_246_95 ();
 b15zdnd11an1n04x5 FILLER_246_109 ();
 b15zdnd11an1n04x5 FILLER_246_120 ();
 b15zdnd11an1n64x5 FILLER_246_166 ();
 b15zdnd11an1n64x5 FILLER_246_230 ();
 b15zdnd11an1n08x5 FILLER_246_294 ();
 b15zdnd00an1n01x5 FILLER_246_302 ();
 b15zdnd11an1n04x5 FILLER_246_312 ();
 b15zdnd11an1n64x5 FILLER_246_323 ();
 b15zdnd11an1n32x5 FILLER_246_387 ();
 b15zdnd11an1n16x5 FILLER_246_419 ();
 b15zdnd11an1n08x5 FILLER_246_435 ();
 b15zdnd11an1n04x5 FILLER_246_443 ();
 b15zdnd11an1n64x5 FILLER_246_450 ();
 b15zdnd11an1n04x5 FILLER_246_514 ();
 b15zdnd00an1n02x5 FILLER_246_518 ();
 b15zdnd11an1n04x5 FILLER_246_523 ();
 b15zdnd11an1n64x5 FILLER_246_530 ();
 b15zdnd11an1n64x5 FILLER_246_594 ();
 b15zdnd11an1n32x5 FILLER_246_658 ();
 b15zdnd11an1n16x5 FILLER_246_690 ();
 b15zdnd11an1n08x5 FILLER_246_706 ();
 b15zdnd11an1n04x5 FILLER_246_714 ();
 b15zdnd11an1n64x5 FILLER_246_726 ();
 b15zdnd11an1n64x5 FILLER_246_790 ();
 b15zdnd11an1n64x5 FILLER_246_854 ();
 b15zdnd11an1n64x5 FILLER_246_918 ();
 b15zdnd11an1n64x5 FILLER_246_982 ();
 b15zdnd11an1n64x5 FILLER_246_1046 ();
 b15zdnd11an1n64x5 FILLER_246_1110 ();
 b15zdnd11an1n64x5 FILLER_246_1174 ();
 b15zdnd11an1n64x5 FILLER_246_1238 ();
 b15zdnd11an1n32x5 FILLER_246_1302 ();
 b15zdnd11an1n16x5 FILLER_246_1334 ();
 b15zdnd11an1n64x5 FILLER_246_1353 ();
 b15zdnd11an1n32x5 FILLER_246_1417 ();
 b15zdnd11an1n08x5 FILLER_246_1449 ();
 b15zdnd11an1n04x5 FILLER_246_1457 ();
 b15zdnd00an1n02x5 FILLER_246_1461 ();
 b15zdnd11an1n64x5 FILLER_246_1505 ();
 b15zdnd11an1n32x5 FILLER_246_1569 ();
 b15zdnd11an1n16x5 FILLER_246_1601 ();
 b15zdnd00an1n02x5 FILLER_246_1617 ();
 b15zdnd11an1n64x5 FILLER_246_1627 ();
 b15zdnd11an1n64x5 FILLER_246_1691 ();
 b15zdnd11an1n64x5 FILLER_246_1755 ();
 b15zdnd11an1n16x5 FILLER_246_1819 ();
 b15zdnd11an1n04x5 FILLER_246_1835 ();
 b15zdnd00an1n02x5 FILLER_246_1839 ();
 b15zdnd00an1n01x5 FILLER_246_1841 ();
 b15zdnd11an1n64x5 FILLER_246_1882 ();
 b15zdnd11an1n08x5 FILLER_246_1946 ();
 b15zdnd00an1n02x5 FILLER_246_1954 ();
 b15zdnd00an1n01x5 FILLER_246_1956 ();
 b15zdnd11an1n04x5 FILLER_246_1960 ();
 b15zdnd11an1n08x5 FILLER_246_1967 ();
 b15zdnd00an1n02x5 FILLER_246_1975 ();
 b15zdnd00an1n01x5 FILLER_246_1977 ();
 b15zdnd11an1n64x5 FILLER_246_2020 ();
 b15zdnd11an1n08x5 FILLER_246_2084 ();
 b15zdnd00an1n02x5 FILLER_246_2092 ();
 b15zdnd00an1n01x5 FILLER_246_2094 ();
 b15zdnd11an1n32x5 FILLER_246_2098 ();
 b15zdnd11an1n16x5 FILLER_246_2130 ();
 b15zdnd11an1n08x5 FILLER_246_2146 ();
 b15zdnd11an1n64x5 FILLER_246_2162 ();
 b15zdnd11an1n32x5 FILLER_246_2226 ();
 b15zdnd11an1n16x5 FILLER_246_2258 ();
 b15zdnd00an1n02x5 FILLER_246_2274 ();
 b15zdnd11an1n64x5 FILLER_247_0 ();
 b15zdnd11an1n64x5 FILLER_247_64 ();
 b15zdnd11an1n64x5 FILLER_247_128 ();
 b15zdnd11an1n64x5 FILLER_247_192 ();
 b15zdnd11an1n32x5 FILLER_247_256 ();
 b15zdnd00an1n02x5 FILLER_247_288 ();
 b15zdnd00an1n01x5 FILLER_247_290 ();
 b15zdnd11an1n04x5 FILLER_247_298 ();
 b15zdnd11an1n64x5 FILLER_247_344 ();
 b15zdnd00an1n02x5 FILLER_247_408 ();
 b15zdnd11an1n64x5 FILLER_247_450 ();
 b15zdnd11an1n04x5 FILLER_247_514 ();
 b15zdnd00an1n02x5 FILLER_247_518 ();
 b15zdnd11an1n64x5 FILLER_247_523 ();
 b15zdnd11an1n64x5 FILLER_247_587 ();
 b15zdnd11an1n64x5 FILLER_247_651 ();
 b15zdnd11an1n64x5 FILLER_247_715 ();
 b15zdnd11an1n64x5 FILLER_247_779 ();
 b15zdnd11an1n16x5 FILLER_247_843 ();
 b15zdnd11an1n08x5 FILLER_247_859 ();
 b15zdnd00an1n02x5 FILLER_247_867 ();
 b15zdnd11an1n64x5 FILLER_247_908 ();
 b15zdnd11an1n64x5 FILLER_247_972 ();
 b15zdnd11an1n64x5 FILLER_247_1036 ();
 b15zdnd11an1n64x5 FILLER_247_1100 ();
 b15zdnd11an1n64x5 FILLER_247_1164 ();
 b15zdnd11an1n64x5 FILLER_247_1228 ();
 b15zdnd11an1n32x5 FILLER_247_1292 ();
 b15zdnd11an1n16x5 FILLER_247_1324 ();
 b15zdnd00an1n02x5 FILLER_247_1340 ();
 b15zdnd11an1n04x5 FILLER_247_1345 ();
 b15zdnd11an1n64x5 FILLER_247_1352 ();
 b15zdnd11an1n32x5 FILLER_247_1416 ();
 b15zdnd11an1n08x5 FILLER_247_1448 ();
 b15zdnd11an1n04x5 FILLER_247_1456 ();
 b15zdnd00an1n02x5 FILLER_247_1460 ();
 b15zdnd11an1n64x5 FILLER_247_1504 ();
 b15zdnd11an1n64x5 FILLER_247_1568 ();
 b15zdnd11an1n64x5 FILLER_247_1632 ();
 b15zdnd11an1n64x5 FILLER_247_1696 ();
 b15zdnd11an1n64x5 FILLER_247_1760 ();
 b15zdnd11an1n32x5 FILLER_247_1824 ();
 b15zdnd11an1n08x5 FILLER_247_1856 ();
 b15zdnd11an1n04x5 FILLER_247_1864 ();
 b15zdnd00an1n02x5 FILLER_247_1868 ();
 b15zdnd11an1n04x5 FILLER_247_1873 ();
 b15zdnd00an1n02x5 FILLER_247_1877 ();
 b15zdnd11an1n32x5 FILLER_247_1882 ();
 b15zdnd11an1n16x5 FILLER_247_1914 ();
 b15zdnd11an1n08x5 FILLER_247_1930 ();
 b15zdnd00an1n01x5 FILLER_247_1938 ();
 b15zdnd11an1n64x5 FILLER_247_1991 ();
 b15zdnd11an1n04x5 FILLER_247_2055 ();
 b15zdnd00an1n02x5 FILLER_247_2059 ();
 b15zdnd11an1n64x5 FILLER_247_2101 ();
 b15zdnd11an1n16x5 FILLER_247_2165 ();
 b15zdnd00an1n02x5 FILLER_247_2181 ();
 b15zdnd00an1n01x5 FILLER_247_2183 ();
 b15zdnd11an1n32x5 FILLER_247_2236 ();
 b15zdnd11an1n16x5 FILLER_247_2268 ();
 b15zdnd11an1n64x5 FILLER_248_8 ();
 b15zdnd11an1n64x5 FILLER_248_72 ();
 b15zdnd11an1n64x5 FILLER_248_136 ();
 b15zdnd11an1n64x5 FILLER_248_200 ();
 b15zdnd11an1n16x5 FILLER_248_264 ();
 b15zdnd11an1n08x5 FILLER_248_280 ();
 b15zdnd11an1n04x5 FILLER_248_288 ();
 b15zdnd00an1n01x5 FILLER_248_292 ();
 b15zdnd11an1n04x5 FILLER_248_298 ();
 b15zdnd11an1n04x5 FILLER_248_306 ();
 b15zdnd00an1n02x5 FILLER_248_310 ();
 b15zdnd11an1n64x5 FILLER_248_316 ();
 b15zdnd11an1n32x5 FILLER_248_380 ();
 b15zdnd11an1n16x5 FILLER_248_412 ();
 b15zdnd00an1n02x5 FILLER_248_428 ();
 b15zdnd11an1n08x5 FILLER_248_436 ();
 b15zdnd00an1n02x5 FILLER_248_444 ();
 b15zdnd11an1n64x5 FILLER_248_449 ();
 b15zdnd11an1n64x5 FILLER_248_513 ();
 b15zdnd11an1n64x5 FILLER_248_577 ();
 b15zdnd11an1n64x5 FILLER_248_641 ();
 b15zdnd11an1n08x5 FILLER_248_705 ();
 b15zdnd11an1n04x5 FILLER_248_713 ();
 b15zdnd00an1n01x5 FILLER_248_717 ();
 b15zdnd11an1n16x5 FILLER_248_726 ();
 b15zdnd11an1n04x5 FILLER_248_742 ();
 b15zdnd00an1n01x5 FILLER_248_746 ();
 b15zdnd11an1n16x5 FILLER_248_756 ();
 b15zdnd11an1n04x5 FILLER_248_772 ();
 b15zdnd00an1n02x5 FILLER_248_776 ();
 b15zdnd00an1n01x5 FILLER_248_778 ();
 b15zdnd11an1n04x5 FILLER_248_782 ();
 b15zdnd11an1n64x5 FILLER_248_789 ();
 b15zdnd11an1n32x5 FILLER_248_853 ();
 b15zdnd11an1n04x5 FILLER_248_885 ();
 b15zdnd11an1n64x5 FILLER_248_896 ();
 b15zdnd11an1n64x5 FILLER_248_960 ();
 b15zdnd11an1n64x5 FILLER_248_1024 ();
 b15zdnd11an1n64x5 FILLER_248_1088 ();
 b15zdnd11an1n64x5 FILLER_248_1152 ();
 b15zdnd00an1n01x5 FILLER_248_1216 ();
 b15zdnd11an1n64x5 FILLER_248_1220 ();
 b15zdnd11an1n32x5 FILLER_248_1284 ();
 b15zdnd11an1n04x5 FILLER_248_1316 ();
 b15zdnd00an1n02x5 FILLER_248_1320 ();
 b15zdnd11an1n64x5 FILLER_248_1374 ();
 b15zdnd11an1n64x5 FILLER_248_1438 ();
 b15zdnd11an1n64x5 FILLER_248_1502 ();
 b15zdnd11an1n32x5 FILLER_248_1566 ();
 b15zdnd11an1n08x5 FILLER_248_1598 ();
 b15zdnd11an1n04x5 FILLER_248_1606 ();
 b15zdnd11an1n64x5 FILLER_248_1617 ();
 b15zdnd11an1n32x5 FILLER_248_1681 ();
 b15zdnd11an1n04x5 FILLER_248_1713 ();
 b15zdnd11an1n64x5 FILLER_248_1737 ();
 b15zdnd11an1n64x5 FILLER_248_1801 ();
 b15zdnd11an1n64x5 FILLER_248_1865 ();
 b15zdnd11an1n32x5 FILLER_248_1929 ();
 b15zdnd11an1n04x5 FILLER_248_1961 ();
 b15zdnd11an1n16x5 FILLER_248_1968 ();
 b15zdnd11an1n04x5 FILLER_248_1984 ();
 b15zdnd00an1n01x5 FILLER_248_1988 ();
 b15zdnd11an1n64x5 FILLER_248_2009 ();
 b15zdnd11an1n16x5 FILLER_248_2073 ();
 b15zdnd11an1n04x5 FILLER_248_2089 ();
 b15zdnd00an1n02x5 FILLER_248_2093 ();
 b15zdnd00an1n01x5 FILLER_248_2095 ();
 b15zdnd11an1n32x5 FILLER_248_2099 ();
 b15zdnd11an1n16x5 FILLER_248_2131 ();
 b15zdnd11an1n04x5 FILLER_248_2147 ();
 b15zdnd00an1n02x5 FILLER_248_2151 ();
 b15zdnd00an1n01x5 FILLER_248_2153 ();
 b15zdnd11an1n32x5 FILLER_248_2162 ();
 b15zdnd11an1n08x5 FILLER_248_2194 ();
 b15zdnd11an1n04x5 FILLER_248_2205 ();
 b15zdnd11an1n04x5 FILLER_248_2212 ();
 b15zdnd11an1n32x5 FILLER_248_2219 ();
 b15zdnd11an1n16x5 FILLER_248_2251 ();
 b15zdnd11an1n08x5 FILLER_248_2267 ();
 b15zdnd00an1n01x5 FILLER_248_2275 ();
 b15zdnd11an1n64x5 FILLER_249_0 ();
 b15zdnd11an1n32x5 FILLER_249_64 ();
 b15zdnd11an1n04x5 FILLER_249_96 ();
 b15zdnd00an1n02x5 FILLER_249_100 ();
 b15zdnd11an1n64x5 FILLER_249_144 ();
 b15zdnd11an1n64x5 FILLER_249_208 ();
 b15zdnd11an1n64x5 FILLER_249_272 ();
 b15zdnd11an1n64x5 FILLER_249_336 ();
 b15zdnd11an1n64x5 FILLER_249_400 ();
 b15zdnd11an1n64x5 FILLER_249_464 ();
 b15zdnd11an1n64x5 FILLER_249_528 ();
 b15zdnd11an1n64x5 FILLER_249_592 ();
 b15zdnd11an1n32x5 FILLER_249_656 ();
 b15zdnd11an1n08x5 FILLER_249_688 ();
 b15zdnd11an1n32x5 FILLER_249_738 ();
 b15zdnd11an1n08x5 FILLER_249_770 ();
 b15zdnd00an1n02x5 FILLER_249_778 ();
 b15zdnd11an1n64x5 FILLER_249_822 ();
 b15zdnd11an1n04x5 FILLER_249_886 ();
 b15zdnd00an1n01x5 FILLER_249_890 ();
 b15zdnd11an1n64x5 FILLER_249_902 ();
 b15zdnd11an1n64x5 FILLER_249_966 ();
 b15zdnd11an1n64x5 FILLER_249_1030 ();
 b15zdnd11an1n64x5 FILLER_249_1094 ();
 b15zdnd11an1n32x5 FILLER_249_1158 ();
 b15zdnd11an1n16x5 FILLER_249_1190 ();
 b15zdnd11an1n08x5 FILLER_249_1206 ();
 b15zdnd00an1n02x5 FILLER_249_1214 ();
 b15zdnd11an1n04x5 FILLER_249_1219 ();
 b15zdnd00an1n02x5 FILLER_249_1223 ();
 b15zdnd11an1n64x5 FILLER_249_1228 ();
 b15zdnd11an1n32x5 FILLER_249_1292 ();
 b15zdnd11an1n16x5 FILLER_249_1324 ();
 b15zdnd11an1n04x5 FILLER_249_1343 ();
 b15zdnd11an1n64x5 FILLER_249_1350 ();
 b15zdnd11an1n64x5 FILLER_249_1414 ();
 b15zdnd11an1n64x5 FILLER_249_1478 ();
 b15zdnd11an1n64x5 FILLER_249_1542 ();
 b15zdnd11an1n32x5 FILLER_249_1637 ();
 b15zdnd11an1n16x5 FILLER_249_1669 ();
 b15zdnd00an1n02x5 FILLER_249_1685 ();
 b15zdnd00an1n01x5 FILLER_249_1687 ();
 b15zdnd11an1n04x5 FILLER_249_1728 ();
 b15zdnd11an1n64x5 FILLER_249_1735 ();
 b15zdnd11an1n64x5 FILLER_249_1799 ();
 b15zdnd11an1n64x5 FILLER_249_1863 ();
 b15zdnd11an1n64x5 FILLER_249_1927 ();
 b15zdnd11an1n64x5 FILLER_249_1991 ();
 b15zdnd11an1n16x5 FILLER_249_2055 ();
 b15zdnd11an1n04x5 FILLER_249_2071 ();
 b15zdnd00an1n01x5 FILLER_249_2075 ();
 b15zdnd11an1n04x5 FILLER_249_2089 ();
 b15zdnd11an1n64x5 FILLER_249_2113 ();
 b15zdnd11an1n32x5 FILLER_249_2177 ();
 b15zdnd11an1n04x5 FILLER_249_2209 ();
 b15zdnd00an1n02x5 FILLER_249_2213 ();
 b15zdnd00an1n01x5 FILLER_249_2215 ();
 b15zdnd11an1n64x5 FILLER_249_2219 ();
 b15zdnd00an1n01x5 FILLER_249_2283 ();
 b15zdnd11an1n64x5 FILLER_250_8 ();
 b15zdnd11an1n64x5 FILLER_250_72 ();
 b15zdnd11an1n64x5 FILLER_250_136 ();
 b15zdnd11an1n64x5 FILLER_250_200 ();
 b15zdnd11an1n64x5 FILLER_250_264 ();
 b15zdnd11an1n64x5 FILLER_250_328 ();
 b15zdnd11an1n64x5 FILLER_250_392 ();
 b15zdnd11an1n64x5 FILLER_250_456 ();
 b15zdnd11an1n64x5 FILLER_250_520 ();
 b15zdnd11an1n32x5 FILLER_250_584 ();
 b15zdnd11an1n16x5 FILLER_250_616 ();
 b15zdnd11an1n08x5 FILLER_250_632 ();
 b15zdnd00an1n02x5 FILLER_250_640 ();
 b15zdnd11an1n32x5 FILLER_250_673 ();
 b15zdnd11an1n08x5 FILLER_250_705 ();
 b15zdnd11an1n04x5 FILLER_250_713 ();
 b15zdnd00an1n01x5 FILLER_250_717 ();
 b15zdnd11an1n08x5 FILLER_250_726 ();
 b15zdnd11an1n04x5 FILLER_250_734 ();
 b15zdnd00an1n02x5 FILLER_250_738 ();
 b15zdnd00an1n01x5 FILLER_250_740 ();
 b15zdnd11an1n08x5 FILLER_250_747 ();
 b15zdnd00an1n01x5 FILLER_250_755 ();
 b15zdnd11an1n64x5 FILLER_250_808 ();
 b15zdnd11an1n64x5 FILLER_250_872 ();
 b15zdnd11an1n64x5 FILLER_250_936 ();
 b15zdnd11an1n64x5 FILLER_250_1000 ();
 b15zdnd11an1n64x5 FILLER_250_1064 ();
 b15zdnd11an1n32x5 FILLER_250_1128 ();
 b15zdnd00an1n01x5 FILLER_250_1160 ();
 b15zdnd11an1n16x5 FILLER_250_1167 ();
 b15zdnd11an1n08x5 FILLER_250_1183 ();
 b15zdnd00an1n02x5 FILLER_250_1191 ();
 b15zdnd00an1n01x5 FILLER_250_1193 ();
 b15zdnd11an1n64x5 FILLER_250_1246 ();
 b15zdnd11an1n64x5 FILLER_250_1310 ();
 b15zdnd11an1n32x5 FILLER_250_1374 ();
 b15zdnd11an1n08x5 FILLER_250_1406 ();
 b15zdnd00an1n02x5 FILLER_250_1414 ();
 b15zdnd11an1n64x5 FILLER_250_1468 ();
 b15zdnd11an1n64x5 FILLER_250_1532 ();
 b15zdnd11an1n64x5 FILLER_250_1596 ();
 b15zdnd11an1n32x5 FILLER_250_1660 ();
 b15zdnd11an1n16x5 FILLER_250_1692 ();
 b15zdnd11an1n08x5 FILLER_250_1708 ();
 b15zdnd11an1n04x5 FILLER_250_1716 ();
 b15zdnd11an1n64x5 FILLER_250_1723 ();
 b15zdnd11an1n64x5 FILLER_250_1787 ();
 b15zdnd11an1n64x5 FILLER_250_1851 ();
 b15zdnd11an1n64x5 FILLER_250_1915 ();
 b15zdnd11an1n64x5 FILLER_250_1979 ();
 b15zdnd11an1n32x5 FILLER_250_2043 ();
 b15zdnd00an1n02x5 FILLER_250_2075 ();
 b15zdnd00an1n01x5 FILLER_250_2077 ();
 b15zdnd11an1n64x5 FILLER_250_2081 ();
 b15zdnd11an1n08x5 FILLER_250_2145 ();
 b15zdnd00an1n01x5 FILLER_250_2153 ();
 b15zdnd11an1n32x5 FILLER_250_2162 ();
 b15zdnd11an1n16x5 FILLER_250_2194 ();
 b15zdnd11an1n08x5 FILLER_250_2215 ();
 b15zdnd11an1n04x5 FILLER_250_2223 ();
 b15zdnd00an1n02x5 FILLER_250_2227 ();
 b15zdnd11an1n04x5 FILLER_250_2271 ();
 b15zdnd00an1n01x5 FILLER_250_2275 ();
 b15zdnd11an1n64x5 FILLER_251_0 ();
 b15zdnd11an1n08x5 FILLER_251_64 ();
 b15zdnd11an1n04x5 FILLER_251_72 ();
 b15zdnd00an1n01x5 FILLER_251_76 ();
 b15zdnd11an1n04x5 FILLER_251_80 ();
 b15zdnd00an1n02x5 FILLER_251_84 ();
 b15zdnd11an1n04x5 FILLER_251_96 ();
 b15zdnd00an1n02x5 FILLER_251_100 ();
 b15zdnd00an1n01x5 FILLER_251_102 ();
 b15zdnd11an1n64x5 FILLER_251_119 ();
 b15zdnd11an1n64x5 FILLER_251_183 ();
 b15zdnd11an1n64x5 FILLER_251_247 ();
 b15zdnd11an1n64x5 FILLER_251_311 ();
 b15zdnd11an1n64x5 FILLER_251_375 ();
 b15zdnd11an1n64x5 FILLER_251_439 ();
 b15zdnd11an1n64x5 FILLER_251_503 ();
 b15zdnd11an1n64x5 FILLER_251_567 ();
 b15zdnd11an1n32x5 FILLER_251_631 ();
 b15zdnd11an1n16x5 FILLER_251_663 ();
 b15zdnd11an1n08x5 FILLER_251_679 ();
 b15zdnd11an1n04x5 FILLER_251_694 ();
 b15zdnd00an1n01x5 FILLER_251_698 ();
 b15zdnd11an1n32x5 FILLER_251_741 ();
 b15zdnd11an1n16x5 FILLER_251_773 ();
 b15zdnd11an1n64x5 FILLER_251_792 ();
 b15zdnd11an1n64x5 FILLER_251_856 ();
 b15zdnd11an1n64x5 FILLER_251_920 ();
 b15zdnd11an1n64x5 FILLER_251_984 ();
 b15zdnd11an1n64x5 FILLER_251_1048 ();
 b15zdnd11an1n64x5 FILLER_251_1112 ();
 b15zdnd11an1n32x5 FILLER_251_1176 ();
 b15zdnd11an1n16x5 FILLER_251_1208 ();
 b15zdnd11an1n08x5 FILLER_251_1224 ();
 b15zdnd11an1n04x5 FILLER_251_1236 ();
 b15zdnd11an1n32x5 FILLER_251_1282 ();
 b15zdnd11an1n16x5 FILLER_251_1314 ();
 b15zdnd00an1n01x5 FILLER_251_1330 ();
 b15zdnd11an1n32x5 FILLER_251_1373 ();
 b15zdnd11an1n08x5 FILLER_251_1405 ();
 b15zdnd00an1n01x5 FILLER_251_1413 ();
 b15zdnd11an1n08x5 FILLER_251_1428 ();
 b15zdnd11an1n64x5 FILLER_251_1439 ();
 b15zdnd11an1n64x5 FILLER_251_1503 ();
 b15zdnd11an1n64x5 FILLER_251_1567 ();
 b15zdnd11an1n64x5 FILLER_251_1631 ();
 b15zdnd11an1n64x5 FILLER_251_1695 ();
 b15zdnd11an1n64x5 FILLER_251_1759 ();
 b15zdnd11an1n64x5 FILLER_251_1823 ();
 b15zdnd11an1n64x5 FILLER_251_1887 ();
 b15zdnd11an1n64x5 FILLER_251_1951 ();
 b15zdnd11an1n64x5 FILLER_251_2015 ();
 b15zdnd11an1n64x5 FILLER_251_2079 ();
 b15zdnd11an1n64x5 FILLER_251_2143 ();
 b15zdnd00an1n02x5 FILLER_251_2207 ();
 b15zdnd00an1n01x5 FILLER_251_2209 ();
 b15zdnd11an1n04x5 FILLER_251_2213 ();
 b15zdnd11an1n32x5 FILLER_251_2224 ();
 b15zdnd11an1n16x5 FILLER_251_2256 ();
 b15zdnd11an1n08x5 FILLER_251_2272 ();
 b15zdnd11an1n04x5 FILLER_251_2280 ();
 b15zdnd11an1n64x5 FILLER_252_8 ();
 b15zdnd11an1n64x5 FILLER_252_72 ();
 b15zdnd11an1n32x5 FILLER_252_136 ();
 b15zdnd11an1n08x5 FILLER_252_168 ();
 b15zdnd00an1n01x5 FILLER_252_176 ();
 b15zdnd11an1n16x5 FILLER_252_182 ();
 b15zdnd11an1n08x5 FILLER_252_198 ();
 b15zdnd11an1n64x5 FILLER_252_209 ();
 b15zdnd11an1n16x5 FILLER_252_273 ();
 b15zdnd11an1n08x5 FILLER_252_289 ();
 b15zdnd11an1n04x5 FILLER_252_297 ();
 b15zdnd11an1n32x5 FILLER_252_343 ();
 b15zdnd11an1n04x5 FILLER_252_375 ();
 b15zdnd11an1n64x5 FILLER_252_388 ();
 b15zdnd11an1n64x5 FILLER_252_452 ();
 b15zdnd11an1n64x5 FILLER_252_516 ();
 b15zdnd11an1n64x5 FILLER_252_580 ();
 b15zdnd11an1n32x5 FILLER_252_644 ();
 b15zdnd00an1n02x5 FILLER_252_676 ();
 b15zdnd00an1n01x5 FILLER_252_678 ();
 b15zdnd11an1n04x5 FILLER_252_684 ();
 b15zdnd11an1n04x5 FILLER_252_701 ();
 b15zdnd00an1n02x5 FILLER_252_716 ();
 b15zdnd11an1n64x5 FILLER_252_726 ();
 b15zdnd11an1n08x5 FILLER_252_790 ();
 b15zdnd00an1n01x5 FILLER_252_798 ();
 b15zdnd11an1n64x5 FILLER_252_802 ();
 b15zdnd11an1n32x5 FILLER_252_866 ();
 b15zdnd00an1n01x5 FILLER_252_898 ();
 b15zdnd11an1n64x5 FILLER_252_941 ();
 b15zdnd11an1n32x5 FILLER_252_1005 ();
 b15zdnd00an1n02x5 FILLER_252_1037 ();
 b15zdnd11an1n64x5 FILLER_252_1091 ();
 b15zdnd11an1n64x5 FILLER_252_1155 ();
 b15zdnd11an1n64x5 FILLER_252_1219 ();
 b15zdnd11an1n64x5 FILLER_252_1283 ();
 b15zdnd11an1n64x5 FILLER_252_1347 ();
 b15zdnd11an1n16x5 FILLER_252_1411 ();
 b15zdnd11an1n08x5 FILLER_252_1427 ();
 b15zdnd11an1n04x5 FILLER_252_1438 ();
 b15zdnd11an1n16x5 FILLER_252_1445 ();
 b15zdnd11an1n08x5 FILLER_252_1461 ();
 b15zdnd00an1n02x5 FILLER_252_1469 ();
 b15zdnd11an1n64x5 FILLER_252_1513 ();
 b15zdnd11an1n64x5 FILLER_252_1577 ();
 b15zdnd11an1n64x5 FILLER_252_1641 ();
 b15zdnd11an1n64x5 FILLER_252_1705 ();
 b15zdnd11an1n64x5 FILLER_252_1769 ();
 b15zdnd11an1n64x5 FILLER_252_1833 ();
 b15zdnd11an1n64x5 FILLER_252_1897 ();
 b15zdnd11an1n64x5 FILLER_252_1961 ();
 b15zdnd11an1n64x5 FILLER_252_2025 ();
 b15zdnd11an1n64x5 FILLER_252_2089 ();
 b15zdnd00an1n01x5 FILLER_252_2153 ();
 b15zdnd11an1n32x5 FILLER_252_2162 ();
 b15zdnd11an1n16x5 FILLER_252_2194 ();
 b15zdnd00an1n02x5 FILLER_252_2210 ();
 b15zdnd11an1n04x5 FILLER_252_2217 ();
 b15zdnd11an1n32x5 FILLER_252_2225 ();
 b15zdnd11an1n16x5 FILLER_252_2257 ();
 b15zdnd00an1n02x5 FILLER_252_2273 ();
 b15zdnd00an1n01x5 FILLER_252_2275 ();
 b15zdnd11an1n64x5 FILLER_253_0 ();
 b15zdnd11an1n64x5 FILLER_253_64 ();
 b15zdnd11an1n64x5 FILLER_253_128 ();
 b15zdnd00an1n02x5 FILLER_253_192 ();
 b15zdnd00an1n01x5 FILLER_253_194 ();
 b15zdnd11an1n64x5 FILLER_253_237 ();
 b15zdnd11an1n64x5 FILLER_253_301 ();
 b15zdnd11an1n64x5 FILLER_253_365 ();
 b15zdnd11an1n64x5 FILLER_253_429 ();
 b15zdnd11an1n64x5 FILLER_253_493 ();
 b15zdnd11an1n32x5 FILLER_253_557 ();
 b15zdnd11an1n16x5 FILLER_253_589 ();
 b15zdnd11an1n08x5 FILLER_253_605 ();
 b15zdnd11an1n32x5 FILLER_253_631 ();
 b15zdnd11an1n04x5 FILLER_253_663 ();
 b15zdnd00an1n02x5 FILLER_253_667 ();
 b15zdnd11an1n04x5 FILLER_253_673 ();
 b15zdnd11an1n04x5 FILLER_253_719 ();
 b15zdnd11an1n04x5 FILLER_253_765 ();
 b15zdnd00an1n02x5 FILLER_253_769 ();
 b15zdnd00an1n01x5 FILLER_253_771 ();
 b15zdnd11an1n64x5 FILLER_253_824 ();
 b15zdnd11an1n32x5 FILLER_253_888 ();
 b15zdnd11an1n08x5 FILLER_253_920 ();
 b15zdnd11an1n04x5 FILLER_253_928 ();
 b15zdnd00an1n01x5 FILLER_253_932 ();
 b15zdnd11an1n64x5 FILLER_253_936 ();
 b15zdnd11an1n32x5 FILLER_253_1000 ();
 b15zdnd11an1n16x5 FILLER_253_1032 ();
 b15zdnd11an1n08x5 FILLER_253_1048 ();
 b15zdnd00an1n02x5 FILLER_253_1056 ();
 b15zdnd00an1n01x5 FILLER_253_1058 ();
 b15zdnd11an1n04x5 FILLER_253_1062 ();
 b15zdnd11an1n64x5 FILLER_253_1069 ();
 b15zdnd11an1n64x5 FILLER_253_1133 ();
 b15zdnd11an1n64x5 FILLER_253_1197 ();
 b15zdnd11an1n32x5 FILLER_253_1261 ();
 b15zdnd00an1n02x5 FILLER_253_1293 ();
 b15zdnd11an1n04x5 FILLER_253_1337 ();
 b15zdnd11an1n04x5 FILLER_253_1344 ();
 b15zdnd11an1n64x5 FILLER_253_1351 ();
 b15zdnd11an1n64x5 FILLER_253_1415 ();
 b15zdnd11an1n64x5 FILLER_253_1479 ();
 b15zdnd11an1n64x5 FILLER_253_1543 ();
 b15zdnd11an1n64x5 FILLER_253_1607 ();
 b15zdnd11an1n64x5 FILLER_253_1671 ();
 b15zdnd11an1n64x5 FILLER_253_1735 ();
 b15zdnd11an1n64x5 FILLER_253_1799 ();
 b15zdnd11an1n64x5 FILLER_253_1863 ();
 b15zdnd11an1n64x5 FILLER_253_1927 ();
 b15zdnd11an1n64x5 FILLER_253_1991 ();
 b15zdnd11an1n16x5 FILLER_253_2055 ();
 b15zdnd11an1n08x5 FILLER_253_2071 ();
 b15zdnd00an1n02x5 FILLER_253_2079 ();
 b15zdnd00an1n01x5 FILLER_253_2081 ();
 b15zdnd11an1n64x5 FILLER_253_2088 ();
 b15zdnd11an1n32x5 FILLER_253_2152 ();
 b15zdnd11an1n16x5 FILLER_253_2184 ();
 b15zdnd11an1n08x5 FILLER_253_2200 ();
 b15zdnd11an1n04x5 FILLER_253_2208 ();
 b15zdnd00an1n01x5 FILLER_253_2212 ();
 b15zdnd11an1n32x5 FILLER_253_2226 ();
 b15zdnd11an1n16x5 FILLER_253_2258 ();
 b15zdnd11an1n08x5 FILLER_253_2274 ();
 b15zdnd00an1n02x5 FILLER_253_2282 ();
 b15zdnd11an1n64x5 FILLER_254_8 ();
 b15zdnd11an1n08x5 FILLER_254_72 ();
 b15zdnd11an1n04x5 FILLER_254_80 ();
 b15zdnd00an1n01x5 FILLER_254_84 ();
 b15zdnd11an1n08x5 FILLER_254_91 ();
 b15zdnd11an1n04x5 FILLER_254_99 ();
 b15zdnd00an1n02x5 FILLER_254_103 ();
 b15zdnd11an1n64x5 FILLER_254_113 ();
 b15zdnd00an1n02x5 FILLER_254_177 ();
 b15zdnd11an1n64x5 FILLER_254_231 ();
 b15zdnd11an1n32x5 FILLER_254_295 ();
 b15zdnd11an1n04x5 FILLER_254_327 ();
 b15zdnd11an1n64x5 FILLER_254_334 ();
 b15zdnd11an1n64x5 FILLER_254_398 ();
 b15zdnd11an1n64x5 FILLER_254_462 ();
 b15zdnd11an1n64x5 FILLER_254_526 ();
 b15zdnd11an1n64x5 FILLER_254_590 ();
 b15zdnd11an1n16x5 FILLER_254_654 ();
 b15zdnd11an1n04x5 FILLER_254_670 ();
 b15zdnd00an1n02x5 FILLER_254_716 ();
 b15zdnd11an1n64x5 FILLER_254_726 ();
 b15zdnd11an1n04x5 FILLER_254_790 ();
 b15zdnd00an1n02x5 FILLER_254_794 ();
 b15zdnd00an1n01x5 FILLER_254_796 ();
 b15zdnd11an1n64x5 FILLER_254_800 ();
 b15zdnd11an1n32x5 FILLER_254_864 ();
 b15zdnd00an1n01x5 FILLER_254_896 ();
 b15zdnd11an1n04x5 FILLER_254_937 ();
 b15zdnd11an1n04x5 FILLER_254_944 ();
 b15zdnd00an1n02x5 FILLER_254_948 ();
 b15zdnd11an1n04x5 FILLER_254_955 ();
 b15zdnd11an1n64x5 FILLER_254_977 ();
 b15zdnd11an1n16x5 FILLER_254_1041 ();
 b15zdnd11an1n08x5 FILLER_254_1057 ();
 b15zdnd00an1n01x5 FILLER_254_1065 ();
 b15zdnd11an1n64x5 FILLER_254_1069 ();
 b15zdnd11an1n64x5 FILLER_254_1133 ();
 b15zdnd11an1n64x5 FILLER_254_1197 ();
 b15zdnd11an1n16x5 FILLER_254_1261 ();
 b15zdnd00an1n02x5 FILLER_254_1277 ();
 b15zdnd00an1n01x5 FILLER_254_1279 ();
 b15zdnd11an1n08x5 FILLER_254_1298 ();
 b15zdnd00an1n01x5 FILLER_254_1306 ();
 b15zdnd11an1n64x5 FILLER_254_1359 ();
 b15zdnd11an1n64x5 FILLER_254_1423 ();
 b15zdnd11an1n64x5 FILLER_254_1487 ();
 b15zdnd11an1n64x5 FILLER_254_1551 ();
 b15zdnd11an1n32x5 FILLER_254_1615 ();
 b15zdnd11an1n16x5 FILLER_254_1647 ();
 b15zdnd11an1n08x5 FILLER_254_1663 ();
 b15zdnd00an1n01x5 FILLER_254_1671 ();
 b15zdnd11an1n64x5 FILLER_254_1680 ();
 b15zdnd11an1n64x5 FILLER_254_1744 ();
 b15zdnd11an1n64x5 FILLER_254_1808 ();
 b15zdnd11an1n64x5 FILLER_254_1872 ();
 b15zdnd11an1n64x5 FILLER_254_1936 ();
 b15zdnd11an1n64x5 FILLER_254_2000 ();
 b15zdnd11an1n08x5 FILLER_254_2064 ();
 b15zdnd11an1n04x5 FILLER_254_2072 ();
 b15zdnd00an1n02x5 FILLER_254_2076 ();
 b15zdnd00an1n01x5 FILLER_254_2078 ();
 b15zdnd11an1n04x5 FILLER_254_2097 ();
 b15zdnd11an1n32x5 FILLER_254_2106 ();
 b15zdnd11an1n16x5 FILLER_254_2138 ();
 b15zdnd11an1n32x5 FILLER_254_2162 ();
 b15zdnd11an1n08x5 FILLER_254_2194 ();
 b15zdnd11an1n04x5 FILLER_254_2202 ();
 b15zdnd11an1n04x5 FILLER_254_2210 ();
 b15zdnd11an1n04x5 FILLER_254_2220 ();
 b15zdnd11an1n32x5 FILLER_254_2227 ();
 b15zdnd11an1n16x5 FILLER_254_2259 ();
 b15zdnd00an1n01x5 FILLER_254_2275 ();
 b15zdnd11an1n64x5 FILLER_255_0 ();
 b15zdnd11an1n64x5 FILLER_255_64 ();
 b15zdnd11an1n64x5 FILLER_255_128 ();
 b15zdnd11an1n04x5 FILLER_255_192 ();
 b15zdnd00an1n01x5 FILLER_255_196 ();
 b15zdnd11an1n04x5 FILLER_255_200 ();
 b15zdnd11an1n64x5 FILLER_255_207 ();
 b15zdnd11an1n32x5 FILLER_255_271 ();
 b15zdnd00an1n01x5 FILLER_255_303 ();
 b15zdnd11an1n64x5 FILLER_255_356 ();
 b15zdnd11an1n64x5 FILLER_255_420 ();
 b15zdnd11an1n64x5 FILLER_255_484 ();
 b15zdnd11an1n16x5 FILLER_255_548 ();
 b15zdnd11an1n08x5 FILLER_255_564 ();
 b15zdnd00an1n02x5 FILLER_255_572 ();
 b15zdnd00an1n01x5 FILLER_255_574 ();
 b15zdnd11an1n64x5 FILLER_255_581 ();
 b15zdnd11an1n08x5 FILLER_255_645 ();
 b15zdnd11an1n04x5 FILLER_255_653 ();
 b15zdnd00an1n02x5 FILLER_255_657 ();
 b15zdnd00an1n01x5 FILLER_255_659 ();
 b15zdnd11an1n04x5 FILLER_255_702 ();
 b15zdnd11an1n32x5 FILLER_255_748 ();
 b15zdnd11an1n16x5 FILLER_255_780 ();
 b15zdnd00an1n01x5 FILLER_255_796 ();
 b15zdnd11an1n64x5 FILLER_255_800 ();
 b15zdnd11an1n32x5 FILLER_255_864 ();
 b15zdnd11an1n16x5 FILLER_255_896 ();
 b15zdnd11an1n08x5 FILLER_255_912 ();
 b15zdnd11an1n04x5 FILLER_255_920 ();
 b15zdnd00an1n02x5 FILLER_255_924 ();
 b15zdnd11an1n64x5 FILLER_255_968 ();
 b15zdnd11an1n32x5 FILLER_255_1032 ();
 b15zdnd11an1n04x5 FILLER_255_1064 ();
 b15zdnd00an1n02x5 FILLER_255_1068 ();
 b15zdnd11an1n64x5 FILLER_255_1074 ();
 b15zdnd11an1n64x5 FILLER_255_1138 ();
 b15zdnd11an1n08x5 FILLER_255_1202 ();
 b15zdnd11an1n04x5 FILLER_255_1210 ();
 b15zdnd00an1n02x5 FILLER_255_1214 ();
 b15zdnd00an1n01x5 FILLER_255_1216 ();
 b15zdnd11an1n64x5 FILLER_255_1221 ();
 b15zdnd11an1n32x5 FILLER_255_1285 ();
 b15zdnd11an1n08x5 FILLER_255_1317 ();
 b15zdnd11an1n04x5 FILLER_255_1325 ();
 b15zdnd00an1n02x5 FILLER_255_1329 ();
 b15zdnd00an1n01x5 FILLER_255_1331 ();
 b15zdnd11an1n64x5 FILLER_255_1335 ();
 b15zdnd11an1n64x5 FILLER_255_1399 ();
 b15zdnd11an1n64x5 FILLER_255_1463 ();
 b15zdnd11an1n32x5 FILLER_255_1527 ();
 b15zdnd11an1n16x5 FILLER_255_1559 ();
 b15zdnd00an1n02x5 FILLER_255_1575 ();
 b15zdnd11an1n64x5 FILLER_255_1588 ();
 b15zdnd11an1n32x5 FILLER_255_1652 ();
 b15zdnd11an1n08x5 FILLER_255_1684 ();
 b15zdnd11an1n04x5 FILLER_255_1692 ();
 b15zdnd11an1n04x5 FILLER_255_1699 ();
 b15zdnd11an1n64x5 FILLER_255_1706 ();
 b15zdnd11an1n64x5 FILLER_255_1770 ();
 b15zdnd11an1n32x5 FILLER_255_1834 ();
 b15zdnd11an1n16x5 FILLER_255_1866 ();
 b15zdnd00an1n02x5 FILLER_255_1882 ();
 b15zdnd11an1n64x5 FILLER_255_1887 ();
 b15zdnd00an1n02x5 FILLER_255_1951 ();
 b15zdnd00an1n01x5 FILLER_255_1953 ();
 b15zdnd11an1n04x5 FILLER_255_1959 ();
 b15zdnd11an1n64x5 FILLER_255_1966 ();
 b15zdnd11an1n32x5 FILLER_255_2030 ();
 b15zdnd11an1n16x5 FILLER_255_2062 ();
 b15zdnd11an1n64x5 FILLER_255_2120 ();
 b15zdnd11an1n16x5 FILLER_255_2184 ();
 b15zdnd11an1n08x5 FILLER_255_2200 ();
 b15zdnd11an1n04x5 FILLER_255_2208 ();
 b15zdnd00an1n02x5 FILLER_255_2212 ();
 b15zdnd00an1n01x5 FILLER_255_2214 ();
 b15zdnd11an1n64x5 FILLER_255_2218 ();
 b15zdnd00an1n02x5 FILLER_255_2282 ();
 b15zdnd11an1n64x5 FILLER_256_8 ();
 b15zdnd11an1n32x5 FILLER_256_72 ();
 b15zdnd11an1n16x5 FILLER_256_104 ();
 b15zdnd00an1n01x5 FILLER_256_120 ();
 b15zdnd11an1n64x5 FILLER_256_127 ();
 b15zdnd11an1n64x5 FILLER_256_191 ();
 b15zdnd11an1n64x5 FILLER_256_255 ();
 b15zdnd11an1n08x5 FILLER_256_319 ();
 b15zdnd00an1n02x5 FILLER_256_327 ();
 b15zdnd11an1n04x5 FILLER_256_332 ();
 b15zdnd11an1n64x5 FILLER_256_339 ();
 b15zdnd11an1n64x5 FILLER_256_403 ();
 b15zdnd11an1n64x5 FILLER_256_467 ();
 b15zdnd11an1n64x5 FILLER_256_531 ();
 b15zdnd11an1n32x5 FILLER_256_595 ();
 b15zdnd11an1n16x5 FILLER_256_627 ();
 b15zdnd11an1n08x5 FILLER_256_643 ();
 b15zdnd00an1n02x5 FILLER_256_651 ();
 b15zdnd00an1n01x5 FILLER_256_653 ();
 b15zdnd11an1n04x5 FILLER_256_706 ();
 b15zdnd00an1n02x5 FILLER_256_715 ();
 b15zdnd00an1n01x5 FILLER_256_717 ();
 b15zdnd11an1n64x5 FILLER_256_726 ();
 b15zdnd11an1n64x5 FILLER_256_790 ();
 b15zdnd11an1n64x5 FILLER_256_854 ();
 b15zdnd00an1n02x5 FILLER_256_918 ();
 b15zdnd00an1n01x5 FILLER_256_920 ();
 b15zdnd11an1n04x5 FILLER_256_973 ();
 b15zdnd11an1n32x5 FILLER_256_1019 ();
 b15zdnd11an1n08x5 FILLER_256_1051 ();
 b15zdnd00an1n02x5 FILLER_256_1059 ();
 b15zdnd11an1n04x5 FILLER_256_1064 ();
 b15zdnd11an1n64x5 FILLER_256_1074 ();
 b15zdnd11an1n64x5 FILLER_256_1138 ();
 b15zdnd00an1n01x5 FILLER_256_1202 ();
 b15zdnd11an1n04x5 FILLER_256_1206 ();
 b15zdnd11an1n64x5 FILLER_256_1215 ();
 b15zdnd11an1n64x5 FILLER_256_1279 ();
 b15zdnd11an1n64x5 FILLER_256_1343 ();
 b15zdnd11an1n64x5 FILLER_256_1407 ();
 b15zdnd11an1n64x5 FILLER_256_1471 ();
 b15zdnd11an1n32x5 FILLER_256_1535 ();
 b15zdnd11an1n08x5 FILLER_256_1567 ();
 b15zdnd11an1n04x5 FILLER_256_1575 ();
 b15zdnd11an1n04x5 FILLER_256_1589 ();
 b15zdnd11an1n32x5 FILLER_256_1597 ();
 b15zdnd11an1n08x5 FILLER_256_1629 ();
 b15zdnd11an1n04x5 FILLER_256_1637 ();
 b15zdnd00an1n02x5 FILLER_256_1641 ();
 b15zdnd11an1n04x5 FILLER_256_1674 ();
 b15zdnd11an1n64x5 FILLER_256_1730 ();
 b15zdnd11an1n32x5 FILLER_256_1794 ();
 b15zdnd11an1n16x5 FILLER_256_1826 ();
 b15zdnd11an1n08x5 FILLER_256_1842 ();
 b15zdnd00an1n02x5 FILLER_256_1850 ();
 b15zdnd00an1n01x5 FILLER_256_1852 ();
 b15zdnd11an1n04x5 FILLER_256_1893 ();
 b15zdnd11an1n32x5 FILLER_256_1900 ();
 b15zdnd11an1n08x5 FILLER_256_1932 ();
 b15zdnd00an1n02x5 FILLER_256_1940 ();
 b15zdnd00an1n01x5 FILLER_256_1942 ();
 b15zdnd11an1n08x5 FILLER_256_1947 ();
 b15zdnd11an1n64x5 FILLER_256_1958 ();
 b15zdnd11an1n16x5 FILLER_256_2022 ();
 b15zdnd11an1n08x5 FILLER_256_2038 ();
 b15zdnd11an1n04x5 FILLER_256_2046 ();
 b15zdnd11an1n04x5 FILLER_256_2053 ();
 b15zdnd11an1n04x5 FILLER_256_2060 ();
 b15zdnd11an1n04x5 FILLER_256_2067 ();
 b15zdnd11an1n32x5 FILLER_256_2111 ();
 b15zdnd11an1n08x5 FILLER_256_2143 ();
 b15zdnd00an1n02x5 FILLER_256_2151 ();
 b15zdnd00an1n01x5 FILLER_256_2153 ();
 b15zdnd11an1n32x5 FILLER_256_2162 ();
 b15zdnd11an1n16x5 FILLER_256_2194 ();
 b15zdnd11an1n32x5 FILLER_256_2214 ();
 b15zdnd11an1n16x5 FILLER_256_2246 ();
 b15zdnd11an1n08x5 FILLER_256_2262 ();
 b15zdnd11an1n04x5 FILLER_256_2270 ();
 b15zdnd00an1n02x5 FILLER_256_2274 ();
 b15zdnd11an1n64x5 FILLER_257_0 ();
 b15zdnd00an1n01x5 FILLER_257_64 ();
 b15zdnd11an1n64x5 FILLER_257_75 ();
 b15zdnd11an1n64x5 FILLER_257_139 ();
 b15zdnd11an1n64x5 FILLER_257_203 ();
 b15zdnd11an1n64x5 FILLER_257_267 ();
 b15zdnd11an1n64x5 FILLER_257_331 ();
 b15zdnd11an1n64x5 FILLER_257_395 ();
 b15zdnd11an1n64x5 FILLER_257_459 ();
 b15zdnd11an1n64x5 FILLER_257_523 ();
 b15zdnd11an1n64x5 FILLER_257_587 ();
 b15zdnd11an1n16x5 FILLER_257_651 ();
 b15zdnd11an1n04x5 FILLER_257_667 ();
 b15zdnd11an1n04x5 FILLER_257_674 ();
 b15zdnd11an1n64x5 FILLER_257_720 ();
 b15zdnd11an1n64x5 FILLER_257_784 ();
 b15zdnd11an1n64x5 FILLER_257_848 ();
 b15zdnd11an1n16x5 FILLER_257_912 ();
 b15zdnd11an1n04x5 FILLER_257_928 ();
 b15zdnd00an1n02x5 FILLER_257_932 ();
 b15zdnd11an1n04x5 FILLER_257_937 ();
 b15zdnd11an1n04x5 FILLER_257_944 ();
 b15zdnd11an1n64x5 FILLER_257_951 ();
 b15zdnd11an1n32x5 FILLER_257_1015 ();
 b15zdnd11an1n16x5 FILLER_257_1047 ();
 b15zdnd11an1n04x5 FILLER_257_1063 ();
 b15zdnd11an1n64x5 FILLER_257_1071 ();
 b15zdnd11an1n32x5 FILLER_257_1135 ();
 b15zdnd11an1n16x5 FILLER_257_1167 ();
 b15zdnd11an1n08x5 FILLER_257_1183 ();
 b15zdnd11an1n04x5 FILLER_257_1191 ();
 b15zdnd00an1n01x5 FILLER_257_1195 ();
 b15zdnd11an1n64x5 FILLER_257_1207 ();
 b15zdnd11an1n64x5 FILLER_257_1271 ();
 b15zdnd11an1n64x5 FILLER_257_1335 ();
 b15zdnd11an1n64x5 FILLER_257_1399 ();
 b15zdnd11an1n08x5 FILLER_257_1463 ();
 b15zdnd11an1n04x5 FILLER_257_1474 ();
 b15zdnd11an1n64x5 FILLER_257_1481 ();
 b15zdnd11an1n64x5 FILLER_257_1545 ();
 b15zdnd11an1n32x5 FILLER_257_1609 ();
 b15zdnd11an1n16x5 FILLER_257_1641 ();
 b15zdnd11an1n08x5 FILLER_257_1657 ();
 b15zdnd11an1n04x5 FILLER_257_1665 ();
 b15zdnd00an1n02x5 FILLER_257_1669 ();
 b15zdnd11an1n04x5 FILLER_257_1713 ();
 b15zdnd11an1n64x5 FILLER_257_1759 ();
 b15zdnd11an1n64x5 FILLER_257_1823 ();
 b15zdnd11an1n64x5 FILLER_257_1887 ();
 b15zdnd11an1n04x5 FILLER_257_1951 ();
 b15zdnd00an1n01x5 FILLER_257_1955 ();
 b15zdnd11an1n64x5 FILLER_257_1966 ();
 b15zdnd11an1n16x5 FILLER_257_2082 ();
 b15zdnd11an1n08x5 FILLER_257_2098 ();
 b15zdnd11an1n64x5 FILLER_257_2109 ();
 b15zdnd11an1n64x5 FILLER_257_2173 ();
 b15zdnd11an1n32x5 FILLER_257_2237 ();
 b15zdnd11an1n08x5 FILLER_257_2269 ();
 b15zdnd11an1n04x5 FILLER_257_2277 ();
 b15zdnd00an1n02x5 FILLER_257_2281 ();
 b15zdnd00an1n01x5 FILLER_257_2283 ();
 b15zdnd11an1n64x5 FILLER_258_8 ();
 b15zdnd11an1n64x5 FILLER_258_72 ();
 b15zdnd11an1n64x5 FILLER_258_136 ();
 b15zdnd11an1n64x5 FILLER_258_200 ();
 b15zdnd11an1n64x5 FILLER_258_264 ();
 b15zdnd11an1n64x5 FILLER_258_328 ();
 b15zdnd11an1n64x5 FILLER_258_392 ();
 b15zdnd11an1n64x5 FILLER_258_456 ();
 b15zdnd11an1n64x5 FILLER_258_520 ();
 b15zdnd11an1n64x5 FILLER_258_584 ();
 b15zdnd11an1n32x5 FILLER_258_648 ();
 b15zdnd00an1n01x5 FILLER_258_680 ();
 b15zdnd11an1n04x5 FILLER_258_684 ();
 b15zdnd00an1n02x5 FILLER_258_688 ();
 b15zdnd00an1n01x5 FILLER_258_690 ();
 b15zdnd11an1n16x5 FILLER_258_694 ();
 b15zdnd11an1n08x5 FILLER_258_710 ();
 b15zdnd11an1n64x5 FILLER_258_726 ();
 b15zdnd11an1n64x5 FILLER_258_790 ();
 b15zdnd11an1n64x5 FILLER_258_854 ();
 b15zdnd11an1n32x5 FILLER_258_918 ();
 b15zdnd11an1n08x5 FILLER_258_950 ();
 b15zdnd11an1n64x5 FILLER_258_962 ();
 b15zdnd11an1n04x5 FILLER_258_1026 ();
 b15zdnd00an1n02x5 FILLER_258_1030 ();
 b15zdnd00an1n01x5 FILLER_258_1032 ();
 b15zdnd11an1n08x5 FILLER_258_1039 ();
 b15zdnd00an1n02x5 FILLER_258_1047 ();
 b15zdnd00an1n01x5 FILLER_258_1049 ();
 b15zdnd11an1n64x5 FILLER_258_1063 ();
 b15zdnd11an1n64x5 FILLER_258_1127 ();
 b15zdnd11an1n64x5 FILLER_258_1191 ();
 b15zdnd11an1n64x5 FILLER_258_1255 ();
 b15zdnd11an1n64x5 FILLER_258_1319 ();
 b15zdnd11an1n64x5 FILLER_258_1383 ();
 b15zdnd11an1n04x5 FILLER_258_1447 ();
 b15zdnd00an1n02x5 FILLER_258_1451 ();
 b15zdnd11an1n16x5 FILLER_258_1505 ();
 b15zdnd11an1n04x5 FILLER_258_1521 ();
 b15zdnd00an1n02x5 FILLER_258_1525 ();
 b15zdnd11an1n32x5 FILLER_258_1552 ();
 b15zdnd11an1n04x5 FILLER_258_1584 ();
 b15zdnd00an1n02x5 FILLER_258_1588 ();
 b15zdnd00an1n01x5 FILLER_258_1590 ();
 b15zdnd11an1n64x5 FILLER_258_1594 ();
 b15zdnd11an1n16x5 FILLER_258_1658 ();
 b15zdnd00an1n01x5 FILLER_258_1674 ();
 b15zdnd11an1n16x5 FILLER_258_1678 ();
 b15zdnd11an1n08x5 FILLER_258_1694 ();
 b15zdnd00an1n02x5 FILLER_258_1702 ();
 b15zdnd11an1n64x5 FILLER_258_1707 ();
 b15zdnd11an1n32x5 FILLER_258_1771 ();
 b15zdnd11an1n08x5 FILLER_258_1803 ();
 b15zdnd00an1n02x5 FILLER_258_1811 ();
 b15zdnd00an1n01x5 FILLER_258_1813 ();
 b15zdnd11an1n64x5 FILLER_258_1866 ();
 b15zdnd11an1n08x5 FILLER_258_1930 ();
 b15zdnd11an1n04x5 FILLER_258_1938 ();
 b15zdnd11an1n04x5 FILLER_258_1947 ();
 b15zdnd00an1n02x5 FILLER_258_1951 ();
 b15zdnd11an1n64x5 FILLER_258_1957 ();
 b15zdnd11an1n16x5 FILLER_258_2021 ();
 b15zdnd11an1n08x5 FILLER_258_2037 ();
 b15zdnd00an1n02x5 FILLER_258_2045 ();
 b15zdnd00an1n01x5 FILLER_258_2047 ();
 b15zdnd11an1n04x5 FILLER_258_2051 ();
 b15zdnd11an1n32x5 FILLER_258_2058 ();
 b15zdnd11an1n16x5 FILLER_258_2090 ();
 b15zdnd00an1n02x5 FILLER_258_2106 ();
 b15zdnd00an1n01x5 FILLER_258_2108 ();
 b15zdnd11an1n32x5 FILLER_258_2112 ();
 b15zdnd11an1n08x5 FILLER_258_2144 ();
 b15zdnd00an1n02x5 FILLER_258_2152 ();
 b15zdnd11an1n64x5 FILLER_258_2162 ();
 b15zdnd11an1n32x5 FILLER_258_2226 ();
 b15zdnd11an1n16x5 FILLER_258_2258 ();
 b15zdnd00an1n02x5 FILLER_258_2274 ();
 b15zdnd11an1n08x5 FILLER_259_0 ();
 b15zdnd11an1n04x5 FILLER_259_8 ();
 b15zdnd00an1n02x5 FILLER_259_12 ();
 b15zdnd11an1n64x5 FILLER_259_25 ();
 b15zdnd11an1n32x5 FILLER_259_89 ();
 b15zdnd11an1n08x5 FILLER_259_121 ();
 b15zdnd00an1n02x5 FILLER_259_129 ();
 b15zdnd00an1n01x5 FILLER_259_131 ();
 b15zdnd11an1n04x5 FILLER_259_174 ();
 b15zdnd11an1n64x5 FILLER_259_203 ();
 b15zdnd11an1n64x5 FILLER_259_267 ();
 b15zdnd11an1n64x5 FILLER_259_331 ();
 b15zdnd11an1n64x5 FILLER_259_395 ();
 b15zdnd11an1n64x5 FILLER_259_459 ();
 b15zdnd11an1n04x5 FILLER_259_523 ();
 b15zdnd00an1n02x5 FILLER_259_527 ();
 b15zdnd00an1n01x5 FILLER_259_529 ();
 b15zdnd11an1n64x5 FILLER_259_534 ();
 b15zdnd11an1n64x5 FILLER_259_598 ();
 b15zdnd11an1n16x5 FILLER_259_662 ();
 b15zdnd11an1n08x5 FILLER_259_678 ();
 b15zdnd11an1n64x5 FILLER_259_689 ();
 b15zdnd11an1n16x5 FILLER_259_753 ();
 b15zdnd11an1n08x5 FILLER_259_769 ();
 b15zdnd00an1n01x5 FILLER_259_777 ();
 b15zdnd11an1n64x5 FILLER_259_820 ();
 b15zdnd11an1n64x5 FILLER_259_884 ();
 b15zdnd11an1n64x5 FILLER_259_948 ();
 b15zdnd11an1n32x5 FILLER_259_1012 ();
 b15zdnd11an1n08x5 FILLER_259_1044 ();
 b15zdnd00an1n02x5 FILLER_259_1052 ();
 b15zdnd00an1n01x5 FILLER_259_1054 ();
 b15zdnd11an1n64x5 FILLER_259_1060 ();
 b15zdnd11an1n64x5 FILLER_259_1124 ();
 b15zdnd11an1n08x5 FILLER_259_1188 ();
 b15zdnd11an1n64x5 FILLER_259_1202 ();
 b15zdnd11an1n64x5 FILLER_259_1266 ();
 b15zdnd11an1n64x5 FILLER_259_1330 ();
 b15zdnd11an1n64x5 FILLER_259_1394 ();
 b15zdnd11an1n16x5 FILLER_259_1458 ();
 b15zdnd11an1n04x5 FILLER_259_1474 ();
 b15zdnd00an1n01x5 FILLER_259_1478 ();
 b15zdnd11an1n32x5 FILLER_259_1482 ();
 b15zdnd00an1n02x5 FILLER_259_1514 ();
 b15zdnd11an1n64x5 FILLER_259_1558 ();
 b15zdnd11an1n16x5 FILLER_259_1622 ();
 b15zdnd00an1n02x5 FILLER_259_1638 ();
 b15zdnd11an1n64x5 FILLER_259_1680 ();
 b15zdnd11an1n16x5 FILLER_259_1744 ();
 b15zdnd11an1n08x5 FILLER_259_1760 ();
 b15zdnd11an1n04x5 FILLER_259_1768 ();
 b15zdnd00an1n02x5 FILLER_259_1772 ();
 b15zdnd00an1n01x5 FILLER_259_1774 ();
 b15zdnd11an1n16x5 FILLER_259_1815 ();
 b15zdnd00an1n01x5 FILLER_259_1831 ();
 b15zdnd11an1n04x5 FILLER_259_1835 ();
 b15zdnd11an1n04x5 FILLER_259_1842 ();
 b15zdnd11an1n64x5 FILLER_259_1849 ();
 b15zdnd11an1n32x5 FILLER_259_1913 ();
 b15zdnd11an1n04x5 FILLER_259_1945 ();
 b15zdnd00an1n02x5 FILLER_259_1949 ();
 b15zdnd11an1n64x5 FILLER_259_1961 ();
 b15zdnd11an1n64x5 FILLER_259_2025 ();
 b15zdnd11an1n64x5 FILLER_259_2089 ();
 b15zdnd11an1n64x5 FILLER_259_2153 ();
 b15zdnd11an1n64x5 FILLER_259_2217 ();
 b15zdnd00an1n02x5 FILLER_259_2281 ();
 b15zdnd00an1n01x5 FILLER_259_2283 ();
 b15zdnd11an1n16x5 FILLER_260_8 ();
 b15zdnd00an1n02x5 FILLER_260_24 ();
 b15zdnd00an1n01x5 FILLER_260_26 ();
 b15zdnd11an1n64x5 FILLER_260_41 ();
 b15zdnd11an1n32x5 FILLER_260_105 ();
 b15zdnd11an1n16x5 FILLER_260_137 ();
 b15zdnd11an1n08x5 FILLER_260_153 ();
 b15zdnd11an1n04x5 FILLER_260_161 ();
 b15zdnd00an1n01x5 FILLER_260_165 ();
 b15zdnd11an1n08x5 FILLER_260_169 ();
 b15zdnd11an1n04x5 FILLER_260_177 ();
 b15zdnd00an1n01x5 FILLER_260_181 ();
 b15zdnd11an1n64x5 FILLER_260_224 ();
 b15zdnd11an1n64x5 FILLER_260_288 ();
 b15zdnd11an1n64x5 FILLER_260_352 ();
 b15zdnd11an1n64x5 FILLER_260_416 ();
 b15zdnd11an1n32x5 FILLER_260_480 ();
 b15zdnd11an1n16x5 FILLER_260_512 ();
 b15zdnd00an1n01x5 FILLER_260_528 ();
 b15zdnd11an1n32x5 FILLER_260_535 ();
 b15zdnd11an1n08x5 FILLER_260_567 ();
 b15zdnd11an1n04x5 FILLER_260_575 ();
 b15zdnd00an1n02x5 FILLER_260_579 ();
 b15zdnd11an1n04x5 FILLER_260_592 ();
 b15zdnd11an1n04x5 FILLER_260_599 ();
 b15zdnd00an1n02x5 FILLER_260_603 ();
 b15zdnd00an1n01x5 FILLER_260_605 ();
 b15zdnd11an1n64x5 FILLER_260_609 ();
 b15zdnd11an1n32x5 FILLER_260_673 ();
 b15zdnd11an1n08x5 FILLER_260_705 ();
 b15zdnd11an1n04x5 FILLER_260_713 ();
 b15zdnd00an1n01x5 FILLER_260_717 ();
 b15zdnd11an1n64x5 FILLER_260_726 ();
 b15zdnd11an1n64x5 FILLER_260_790 ();
 b15zdnd11an1n64x5 FILLER_260_854 ();
 b15zdnd11an1n64x5 FILLER_260_918 ();
 b15zdnd11an1n64x5 FILLER_260_982 ();
 b15zdnd11an1n64x5 FILLER_260_1046 ();
 b15zdnd11an1n64x5 FILLER_260_1110 ();
 b15zdnd11an1n08x5 FILLER_260_1174 ();
 b15zdnd00an1n02x5 FILLER_260_1182 ();
 b15zdnd11an1n04x5 FILLER_260_1189 ();
 b15zdnd11an1n64x5 FILLER_260_1206 ();
 b15zdnd11an1n64x5 FILLER_260_1270 ();
 b15zdnd11an1n32x5 FILLER_260_1334 ();
 b15zdnd11an1n16x5 FILLER_260_1366 ();
 b15zdnd00an1n02x5 FILLER_260_1382 ();
 b15zdnd00an1n01x5 FILLER_260_1384 ();
 b15zdnd11an1n64x5 FILLER_260_1389 ();
 b15zdnd11an1n64x5 FILLER_260_1453 ();
 b15zdnd11an1n64x5 FILLER_260_1517 ();
 b15zdnd11an1n64x5 FILLER_260_1581 ();
 b15zdnd11an1n32x5 FILLER_260_1645 ();
 b15zdnd11an1n64x5 FILLER_260_1680 ();
 b15zdnd11an1n32x5 FILLER_260_1744 ();
 b15zdnd11an1n16x5 FILLER_260_1776 ();
 b15zdnd11an1n08x5 FILLER_260_1792 ();
 b15zdnd11an1n04x5 FILLER_260_1800 ();
 b15zdnd00an1n02x5 FILLER_260_1804 ();
 b15zdnd11an1n04x5 FILLER_260_1809 ();
 b15zdnd00an1n02x5 FILLER_260_1813 ();
 b15zdnd11an1n64x5 FILLER_260_1818 ();
 b15zdnd11an1n64x5 FILLER_260_1882 ();
 b15zdnd11an1n08x5 FILLER_260_1946 ();
 b15zdnd11an1n04x5 FILLER_260_1954 ();
 b15zdnd11an1n64x5 FILLER_260_1964 ();
 b15zdnd11an1n64x5 FILLER_260_2028 ();
 b15zdnd11an1n32x5 FILLER_260_2092 ();
 b15zdnd11an1n16x5 FILLER_260_2124 ();
 b15zdnd11an1n08x5 FILLER_260_2140 ();
 b15zdnd11an1n04x5 FILLER_260_2148 ();
 b15zdnd00an1n02x5 FILLER_260_2152 ();
 b15zdnd11an1n64x5 FILLER_260_2162 ();
 b15zdnd11an1n32x5 FILLER_260_2226 ();
 b15zdnd11an1n16x5 FILLER_260_2258 ();
 b15zdnd00an1n02x5 FILLER_260_2274 ();
 b15zdnd11an1n64x5 FILLER_261_0 ();
 b15zdnd11an1n64x5 FILLER_261_64 ();
 b15zdnd11an1n08x5 FILLER_261_128 ();
 b15zdnd00an1n02x5 FILLER_261_136 ();
 b15zdnd00an1n01x5 FILLER_261_138 ();
 b15zdnd11an1n64x5 FILLER_261_191 ();
 b15zdnd11an1n64x5 FILLER_261_255 ();
 b15zdnd11an1n64x5 FILLER_261_319 ();
 b15zdnd11an1n64x5 FILLER_261_383 ();
 b15zdnd11an1n64x5 FILLER_261_447 ();
 b15zdnd11an1n16x5 FILLER_261_511 ();
 b15zdnd00an1n02x5 FILLER_261_527 ();
 b15zdnd00an1n01x5 FILLER_261_529 ();
 b15zdnd11an1n32x5 FILLER_261_536 ();
 b15zdnd11an1n16x5 FILLER_261_568 ();
 b15zdnd11an1n08x5 FILLER_261_584 ();
 b15zdnd11an1n64x5 FILLER_261_634 ();
 b15zdnd11an1n64x5 FILLER_261_698 ();
 b15zdnd11an1n64x5 FILLER_261_762 ();
 b15zdnd11an1n64x5 FILLER_261_826 ();
 b15zdnd11an1n64x5 FILLER_261_890 ();
 b15zdnd11an1n64x5 FILLER_261_954 ();
 b15zdnd11an1n32x5 FILLER_261_1018 ();
 b15zdnd11an1n08x5 FILLER_261_1050 ();
 b15zdnd00an1n02x5 FILLER_261_1058 ();
 b15zdnd00an1n01x5 FILLER_261_1060 ();
 b15zdnd11an1n08x5 FILLER_261_1071 ();
 b15zdnd00an1n02x5 FILLER_261_1079 ();
 b15zdnd00an1n01x5 FILLER_261_1081 ();
 b15zdnd11an1n64x5 FILLER_261_1086 ();
 b15zdnd11an1n16x5 FILLER_261_1150 ();
 b15zdnd11an1n08x5 FILLER_261_1166 ();
 b15zdnd11an1n04x5 FILLER_261_1174 ();
 b15zdnd00an1n02x5 FILLER_261_1178 ();
 b15zdnd11an1n04x5 FILLER_261_1191 ();
 b15zdnd11an1n64x5 FILLER_261_1211 ();
 b15zdnd11an1n64x5 FILLER_261_1275 ();
 b15zdnd11an1n64x5 FILLER_261_1339 ();
 b15zdnd11an1n64x5 FILLER_261_1403 ();
 b15zdnd11an1n64x5 FILLER_261_1467 ();
 b15zdnd11an1n64x5 FILLER_261_1531 ();
 b15zdnd11an1n64x5 FILLER_261_1595 ();
 b15zdnd11an1n64x5 FILLER_261_1659 ();
 b15zdnd11an1n64x5 FILLER_261_1723 ();
 b15zdnd11an1n64x5 FILLER_261_1787 ();
 b15zdnd11an1n64x5 FILLER_261_1851 ();
 b15zdnd11an1n64x5 FILLER_261_1915 ();
 b15zdnd11an1n64x5 FILLER_261_1979 ();
 b15zdnd11an1n64x5 FILLER_261_2043 ();
 b15zdnd11an1n64x5 FILLER_261_2107 ();
 b15zdnd11an1n32x5 FILLER_261_2171 ();
 b15zdnd11an1n08x5 FILLER_261_2203 ();
 b15zdnd00an1n02x5 FILLER_261_2211 ();
 b15zdnd11an1n64x5 FILLER_261_2217 ();
 b15zdnd00an1n02x5 FILLER_261_2281 ();
 b15zdnd00an1n01x5 FILLER_261_2283 ();
 b15zdnd11an1n16x5 FILLER_262_8 ();
 b15zdnd11an1n04x5 FILLER_262_24 ();
 b15zdnd00an1n01x5 FILLER_262_28 ();
 b15zdnd11an1n64x5 FILLER_262_49 ();
 b15zdnd11an1n32x5 FILLER_262_113 ();
 b15zdnd11an1n08x5 FILLER_262_145 ();
 b15zdnd11an1n04x5 FILLER_262_153 ();
 b15zdnd11an1n04x5 FILLER_262_160 ();
 b15zdnd11an1n64x5 FILLER_262_167 ();
 b15zdnd11an1n64x5 FILLER_262_231 ();
 b15zdnd11an1n64x5 FILLER_262_295 ();
 b15zdnd11an1n64x5 FILLER_262_359 ();
 b15zdnd11an1n64x5 FILLER_262_423 ();
 b15zdnd11an1n32x5 FILLER_262_487 ();
 b15zdnd11an1n08x5 FILLER_262_519 ();
 b15zdnd00an1n01x5 FILLER_262_527 ();
 b15zdnd11an1n16x5 FILLER_262_538 ();
 b15zdnd00an1n01x5 FILLER_262_554 ();
 b15zdnd11an1n16x5 FILLER_262_565 ();
 b15zdnd11an1n08x5 FILLER_262_581 ();
 b15zdnd11an1n04x5 FILLER_262_589 ();
 b15zdnd00an1n01x5 FILLER_262_593 ();
 b15zdnd11an1n04x5 FILLER_262_600 ();
 b15zdnd11an1n64x5 FILLER_262_646 ();
 b15zdnd11an1n08x5 FILLER_262_710 ();
 b15zdnd11an1n64x5 FILLER_262_726 ();
 b15zdnd11an1n64x5 FILLER_262_790 ();
 b15zdnd11an1n16x5 FILLER_262_854 ();
 b15zdnd11an1n08x5 FILLER_262_870 ();
 b15zdnd11an1n04x5 FILLER_262_878 ();
 b15zdnd00an1n02x5 FILLER_262_882 ();
 b15zdnd00an1n01x5 FILLER_262_884 ();
 b15zdnd11an1n64x5 FILLER_262_927 ();
 b15zdnd11an1n16x5 FILLER_262_991 ();
 b15zdnd11an1n08x5 FILLER_262_1007 ();
 b15zdnd11an1n64x5 FILLER_262_1024 ();
 b15zdnd11an1n64x5 FILLER_262_1088 ();
 b15zdnd11an1n64x5 FILLER_262_1152 ();
 b15zdnd11an1n64x5 FILLER_262_1216 ();
 b15zdnd11an1n64x5 FILLER_262_1280 ();
 b15zdnd11an1n64x5 FILLER_262_1344 ();
 b15zdnd11an1n64x5 FILLER_262_1408 ();
 b15zdnd11an1n64x5 FILLER_262_1472 ();
 b15zdnd11an1n64x5 FILLER_262_1536 ();
 b15zdnd11an1n64x5 FILLER_262_1600 ();
 b15zdnd11an1n64x5 FILLER_262_1664 ();
 b15zdnd11an1n64x5 FILLER_262_1728 ();
 b15zdnd11an1n64x5 FILLER_262_1792 ();
 b15zdnd11an1n64x5 FILLER_262_1856 ();
 b15zdnd11an1n64x5 FILLER_262_1920 ();
 b15zdnd11an1n64x5 FILLER_262_1984 ();
 b15zdnd11an1n64x5 FILLER_262_2048 ();
 b15zdnd11an1n32x5 FILLER_262_2112 ();
 b15zdnd11an1n08x5 FILLER_262_2144 ();
 b15zdnd00an1n02x5 FILLER_262_2152 ();
 b15zdnd11an1n64x5 FILLER_262_2162 ();
 b15zdnd11an1n32x5 FILLER_262_2226 ();
 b15zdnd11an1n16x5 FILLER_262_2258 ();
 b15zdnd00an1n02x5 FILLER_262_2274 ();
 b15zdnd11an1n32x5 FILLER_263_0 ();
 b15zdnd11an1n64x5 FILLER_263_52 ();
 b15zdnd11an1n64x5 FILLER_263_116 ();
 b15zdnd11an1n64x5 FILLER_263_180 ();
 b15zdnd11an1n64x5 FILLER_263_244 ();
 b15zdnd11an1n64x5 FILLER_263_308 ();
 b15zdnd11an1n64x5 FILLER_263_372 ();
 b15zdnd11an1n64x5 FILLER_263_436 ();
 b15zdnd11an1n16x5 FILLER_263_500 ();
 b15zdnd11an1n08x5 FILLER_263_516 ();
 b15zdnd11an1n04x5 FILLER_263_524 ();
 b15zdnd00an1n02x5 FILLER_263_528 ();
 b15zdnd11an1n08x5 FILLER_263_538 ();
 b15zdnd11an1n04x5 FILLER_263_546 ();
 b15zdnd00an1n02x5 FILLER_263_550 ();
 b15zdnd11an1n16x5 FILLER_263_558 ();
 b15zdnd11an1n04x5 FILLER_263_574 ();
 b15zdnd00an1n01x5 FILLER_263_578 ();
 b15zdnd11an1n64x5 FILLER_263_631 ();
 b15zdnd11an1n64x5 FILLER_263_695 ();
 b15zdnd11an1n64x5 FILLER_263_759 ();
 b15zdnd11an1n64x5 FILLER_263_823 ();
 b15zdnd11an1n64x5 FILLER_263_887 ();
 b15zdnd11an1n64x5 FILLER_263_951 ();
 b15zdnd11an1n32x5 FILLER_263_1015 ();
 b15zdnd11an1n08x5 FILLER_263_1047 ();
 b15zdnd00an1n02x5 FILLER_263_1055 ();
 b15zdnd00an1n01x5 FILLER_263_1057 ();
 b15zdnd11an1n32x5 FILLER_263_1064 ();
 b15zdnd11an1n04x5 FILLER_263_1096 ();
 b15zdnd00an1n02x5 FILLER_263_1100 ();
 b15zdnd11an1n64x5 FILLER_263_1105 ();
 b15zdnd11an1n64x5 FILLER_263_1169 ();
 b15zdnd11an1n64x5 FILLER_263_1233 ();
 b15zdnd11an1n64x5 FILLER_263_1297 ();
 b15zdnd11an1n64x5 FILLER_263_1361 ();
 b15zdnd11an1n64x5 FILLER_263_1425 ();
 b15zdnd11an1n64x5 FILLER_263_1489 ();
 b15zdnd11an1n64x5 FILLER_263_1553 ();
 b15zdnd11an1n64x5 FILLER_263_1617 ();
 b15zdnd11an1n64x5 FILLER_263_1681 ();
 b15zdnd11an1n64x5 FILLER_263_1745 ();
 b15zdnd11an1n04x5 FILLER_263_1809 ();
 b15zdnd00an1n02x5 FILLER_263_1813 ();
 b15zdnd00an1n01x5 FILLER_263_1815 ();
 b15zdnd11an1n64x5 FILLER_263_1858 ();
 b15zdnd11an1n64x5 FILLER_263_1922 ();
 b15zdnd11an1n64x5 FILLER_263_1986 ();
 b15zdnd11an1n64x5 FILLER_263_2050 ();
 b15zdnd11an1n64x5 FILLER_263_2114 ();
 b15zdnd11an1n64x5 FILLER_263_2178 ();
 b15zdnd11an1n32x5 FILLER_263_2242 ();
 b15zdnd11an1n08x5 FILLER_263_2274 ();
 b15zdnd00an1n02x5 FILLER_263_2282 ();
 b15zdnd11an1n64x5 FILLER_264_8 ();
 b15zdnd11an1n64x5 FILLER_264_72 ();
 b15zdnd11an1n64x5 FILLER_264_136 ();
 b15zdnd11an1n64x5 FILLER_264_200 ();
 b15zdnd11an1n64x5 FILLER_264_264 ();
 b15zdnd11an1n64x5 FILLER_264_328 ();
 b15zdnd11an1n16x5 FILLER_264_392 ();
 b15zdnd11an1n08x5 FILLER_264_408 ();
 b15zdnd00an1n02x5 FILLER_264_416 ();
 b15zdnd11an1n64x5 FILLER_264_441 ();
 b15zdnd11an1n08x5 FILLER_264_505 ();
 b15zdnd11an1n04x5 FILLER_264_513 ();
 b15zdnd00an1n02x5 FILLER_264_517 ();
 b15zdnd00an1n01x5 FILLER_264_519 ();
 b15zdnd11an1n32x5 FILLER_264_533 ();
 b15zdnd11an1n04x5 FILLER_264_565 ();
 b15zdnd11an1n64x5 FILLER_264_611 ();
 b15zdnd11an1n32x5 FILLER_264_675 ();
 b15zdnd11an1n08x5 FILLER_264_707 ();
 b15zdnd00an1n02x5 FILLER_264_715 ();
 b15zdnd00an1n01x5 FILLER_264_717 ();
 b15zdnd11an1n64x5 FILLER_264_726 ();
 b15zdnd11an1n64x5 FILLER_264_790 ();
 b15zdnd11an1n64x5 FILLER_264_854 ();
 b15zdnd11an1n64x5 FILLER_264_918 ();
 b15zdnd11an1n64x5 FILLER_264_982 ();
 b15zdnd11an1n16x5 FILLER_264_1046 ();
 b15zdnd11an1n16x5 FILLER_264_1068 ();
 b15zdnd11an1n04x5 FILLER_264_1084 ();
 b15zdnd00an1n02x5 FILLER_264_1088 ();
 b15zdnd00an1n01x5 FILLER_264_1090 ();
 b15zdnd11an1n64x5 FILLER_264_1101 ();
 b15zdnd11an1n64x5 FILLER_264_1165 ();
 b15zdnd11an1n64x5 FILLER_264_1229 ();
 b15zdnd11an1n64x5 FILLER_264_1293 ();
 b15zdnd11an1n64x5 FILLER_264_1357 ();
 b15zdnd11an1n64x5 FILLER_264_1421 ();
 b15zdnd11an1n64x5 FILLER_264_1485 ();
 b15zdnd11an1n64x5 FILLER_264_1549 ();
 b15zdnd11an1n64x5 FILLER_264_1613 ();
 b15zdnd11an1n64x5 FILLER_264_1677 ();
 b15zdnd11an1n64x5 FILLER_264_1741 ();
 b15zdnd11an1n64x5 FILLER_264_1805 ();
 b15zdnd11an1n64x5 FILLER_264_1869 ();
 b15zdnd11an1n64x5 FILLER_264_1933 ();
 b15zdnd11an1n64x5 FILLER_264_1997 ();
 b15zdnd11an1n04x5 FILLER_264_2061 ();
 b15zdnd00an1n02x5 FILLER_264_2065 ();
 b15zdnd00an1n01x5 FILLER_264_2067 ();
 b15zdnd11an1n32x5 FILLER_264_2110 ();
 b15zdnd11an1n08x5 FILLER_264_2142 ();
 b15zdnd11an1n04x5 FILLER_264_2150 ();
 b15zdnd11an1n64x5 FILLER_264_2162 ();
 b15zdnd11an1n32x5 FILLER_264_2226 ();
 b15zdnd11an1n16x5 FILLER_264_2258 ();
 b15zdnd00an1n02x5 FILLER_264_2274 ();
 b15zdnd11an1n64x5 FILLER_265_0 ();
 b15zdnd11an1n64x5 FILLER_265_64 ();
 b15zdnd11an1n64x5 FILLER_265_128 ();
 b15zdnd11an1n64x5 FILLER_265_192 ();
 b15zdnd11an1n64x5 FILLER_265_256 ();
 b15zdnd11an1n64x5 FILLER_265_320 ();
 b15zdnd11an1n32x5 FILLER_265_384 ();
 b15zdnd11an1n08x5 FILLER_265_416 ();
 b15zdnd00an1n02x5 FILLER_265_424 ();
 b15zdnd11an1n16x5 FILLER_265_429 ();
 b15zdnd00an1n02x5 FILLER_265_445 ();
 b15zdnd00an1n01x5 FILLER_265_447 ();
 b15zdnd11an1n64x5 FILLER_265_454 ();
 b15zdnd11an1n64x5 FILLER_265_518 ();
 b15zdnd11an1n16x5 FILLER_265_582 ();
 b15zdnd11an1n04x5 FILLER_265_598 ();
 b15zdnd00an1n02x5 FILLER_265_602 ();
 b15zdnd11an1n04x5 FILLER_265_607 ();
 b15zdnd11an1n64x5 FILLER_265_614 ();
 b15zdnd11an1n64x5 FILLER_265_678 ();
 b15zdnd11an1n32x5 FILLER_265_742 ();
 b15zdnd11an1n16x5 FILLER_265_774 ();
 b15zdnd11an1n08x5 FILLER_265_790 ();
 b15zdnd11an1n04x5 FILLER_265_801 ();
 b15zdnd11an1n64x5 FILLER_265_808 ();
 b15zdnd11an1n64x5 FILLER_265_872 ();
 b15zdnd11an1n64x5 FILLER_265_936 ();
 b15zdnd11an1n32x5 FILLER_265_1000 ();
 b15zdnd11an1n16x5 FILLER_265_1032 ();
 b15zdnd11an1n08x5 FILLER_265_1048 ();
 b15zdnd00an1n01x5 FILLER_265_1056 ();
 b15zdnd11an1n04x5 FILLER_265_1061 ();
 b15zdnd11an1n64x5 FILLER_265_1068 ();
 b15zdnd11an1n32x5 FILLER_265_1132 ();
 b15zdnd11an1n16x5 FILLER_265_1164 ();
 b15zdnd00an1n01x5 FILLER_265_1180 ();
 b15zdnd11an1n64x5 FILLER_265_1186 ();
 b15zdnd11an1n64x5 FILLER_265_1250 ();
 b15zdnd11an1n16x5 FILLER_265_1314 ();
 b15zdnd11an1n08x5 FILLER_265_1330 ();
 b15zdnd11an1n04x5 FILLER_265_1338 ();
 b15zdnd00an1n01x5 FILLER_265_1342 ();
 b15zdnd11an1n32x5 FILLER_265_1354 ();
 b15zdnd11an1n04x5 FILLER_265_1386 ();
 b15zdnd00an1n01x5 FILLER_265_1390 ();
 b15zdnd11an1n04x5 FILLER_265_1431 ();
 b15zdnd11an1n64x5 FILLER_265_1438 ();
 b15zdnd11an1n64x5 FILLER_265_1502 ();
 b15zdnd00an1n01x5 FILLER_265_1566 ();
 b15zdnd11an1n64x5 FILLER_265_1576 ();
 b15zdnd11an1n64x5 FILLER_265_1640 ();
 b15zdnd11an1n64x5 FILLER_265_1704 ();
 b15zdnd11an1n32x5 FILLER_265_1768 ();
 b15zdnd11an1n08x5 FILLER_265_1800 ();
 b15zdnd00an1n02x5 FILLER_265_1808 ();
 b15zdnd11an1n64x5 FILLER_265_1852 ();
 b15zdnd11an1n64x5 FILLER_265_1916 ();
 b15zdnd11an1n64x5 FILLER_265_1980 ();
 b15zdnd11an1n64x5 FILLER_265_2044 ();
 b15zdnd11an1n64x5 FILLER_265_2108 ();
 b15zdnd11an1n32x5 FILLER_265_2172 ();
 b15zdnd11an1n08x5 FILLER_265_2204 ();
 b15zdnd11an1n04x5 FILLER_265_2212 ();
 b15zdnd00an1n01x5 FILLER_265_2216 ();
 b15zdnd11an1n32x5 FILLER_265_2222 ();
 b15zdnd11an1n16x5 FILLER_265_2254 ();
 b15zdnd11an1n08x5 FILLER_265_2270 ();
 b15zdnd11an1n04x5 FILLER_265_2278 ();
 b15zdnd00an1n02x5 FILLER_265_2282 ();
 b15zdnd11an1n64x5 FILLER_266_8 ();
 b15zdnd11an1n64x5 FILLER_266_72 ();
 b15zdnd11an1n64x5 FILLER_266_136 ();
 b15zdnd11an1n64x5 FILLER_266_200 ();
 b15zdnd11an1n64x5 FILLER_266_264 ();
 b15zdnd11an1n64x5 FILLER_266_328 ();
 b15zdnd11an1n04x5 FILLER_266_392 ();
 b15zdnd00an1n02x5 FILLER_266_396 ();
 b15zdnd00an1n01x5 FILLER_266_398 ();
 b15zdnd11an1n04x5 FILLER_266_451 ();
 b15zdnd11an1n64x5 FILLER_266_497 ();
 b15zdnd11an1n64x5 FILLER_266_561 ();
 b15zdnd11an1n64x5 FILLER_266_625 ();
 b15zdnd11an1n16x5 FILLER_266_689 ();
 b15zdnd11an1n08x5 FILLER_266_705 ();
 b15zdnd11an1n04x5 FILLER_266_713 ();
 b15zdnd00an1n01x5 FILLER_266_717 ();
 b15zdnd11an1n32x5 FILLER_266_726 ();
 b15zdnd11an1n16x5 FILLER_266_758 ();
 b15zdnd11an1n04x5 FILLER_266_774 ();
 b15zdnd11an1n64x5 FILLER_266_830 ();
 b15zdnd11an1n64x5 FILLER_266_894 ();
 b15zdnd11an1n64x5 FILLER_266_958 ();
 b15zdnd11an1n64x5 FILLER_266_1022 ();
 b15zdnd11an1n64x5 FILLER_266_1086 ();
 b15zdnd11an1n64x5 FILLER_266_1150 ();
 b15zdnd11an1n64x5 FILLER_266_1214 ();
 b15zdnd11an1n32x5 FILLER_266_1278 ();
 b15zdnd11an1n16x5 FILLER_266_1310 ();
 b15zdnd11an1n04x5 FILLER_266_1326 ();
 b15zdnd11an1n64x5 FILLER_266_1340 ();
 b15zdnd11an1n16x5 FILLER_266_1404 ();
 b15zdnd11an1n08x5 FILLER_266_1420 ();
 b15zdnd11an1n64x5 FILLER_266_1431 ();
 b15zdnd11an1n64x5 FILLER_266_1495 ();
 b15zdnd11an1n64x5 FILLER_266_1559 ();
 b15zdnd11an1n64x5 FILLER_266_1623 ();
 b15zdnd11an1n64x5 FILLER_266_1687 ();
 b15zdnd11an1n32x5 FILLER_266_1751 ();
 b15zdnd11an1n16x5 FILLER_266_1783 ();
 b15zdnd11an1n04x5 FILLER_266_1799 ();
 b15zdnd11an1n64x5 FILLER_266_1845 ();
 b15zdnd11an1n64x5 FILLER_266_1909 ();
 b15zdnd11an1n64x5 FILLER_266_1973 ();
 b15zdnd11an1n64x5 FILLER_266_2037 ();
 b15zdnd11an1n32x5 FILLER_266_2101 ();
 b15zdnd11an1n16x5 FILLER_266_2133 ();
 b15zdnd11an1n04x5 FILLER_266_2149 ();
 b15zdnd00an1n01x5 FILLER_266_2153 ();
 b15zdnd11an1n64x5 FILLER_266_2162 ();
 b15zdnd11an1n32x5 FILLER_266_2226 ();
 b15zdnd11an1n16x5 FILLER_266_2258 ();
 b15zdnd00an1n02x5 FILLER_266_2274 ();
 b15zdnd11an1n16x5 FILLER_267_0 ();
 b15zdnd11an1n08x5 FILLER_267_16 ();
 b15zdnd00an1n02x5 FILLER_267_24 ();
 b15zdnd11an1n64x5 FILLER_267_30 ();
 b15zdnd11an1n64x5 FILLER_267_94 ();
 b15zdnd11an1n64x5 FILLER_267_158 ();
 b15zdnd11an1n64x5 FILLER_267_222 ();
 b15zdnd11an1n64x5 FILLER_267_286 ();
 b15zdnd11an1n32x5 FILLER_267_350 ();
 b15zdnd11an1n16x5 FILLER_267_382 ();
 b15zdnd00an1n02x5 FILLER_267_398 ();
 b15zdnd11an1n04x5 FILLER_267_417 ();
 b15zdnd00an1n01x5 FILLER_267_421 ();
 b15zdnd11an1n04x5 FILLER_267_425 ();
 b15zdnd00an1n01x5 FILLER_267_429 ();
 b15zdnd11an1n64x5 FILLER_267_433 ();
 b15zdnd11an1n64x5 FILLER_267_497 ();
 b15zdnd11an1n64x5 FILLER_267_561 ();
 b15zdnd11an1n64x5 FILLER_267_625 ();
 b15zdnd11an1n64x5 FILLER_267_689 ();
 b15zdnd11an1n32x5 FILLER_267_753 ();
 b15zdnd11an1n08x5 FILLER_267_785 ();
 b15zdnd00an1n01x5 FILLER_267_793 ();
 b15zdnd11an1n04x5 FILLER_267_797 ();
 b15zdnd11an1n04x5 FILLER_267_804 ();
 b15zdnd11an1n64x5 FILLER_267_811 ();
 b15zdnd11an1n64x5 FILLER_267_875 ();
 b15zdnd11an1n64x5 FILLER_267_939 ();
 b15zdnd11an1n64x5 FILLER_267_1003 ();
 b15zdnd11an1n64x5 FILLER_267_1067 ();
 b15zdnd11an1n32x5 FILLER_267_1131 ();
 b15zdnd11an1n16x5 FILLER_267_1163 ();
 b15zdnd11an1n04x5 FILLER_267_1179 ();
 b15zdnd11an1n64x5 FILLER_267_1187 ();
 b15zdnd11an1n64x5 FILLER_267_1251 ();
 b15zdnd11an1n16x5 FILLER_267_1315 ();
 b15zdnd11an1n04x5 FILLER_267_1331 ();
 b15zdnd00an1n02x5 FILLER_267_1335 ();
 b15zdnd00an1n01x5 FILLER_267_1337 ();
 b15zdnd11an1n64x5 FILLER_267_1342 ();
 b15zdnd11an1n64x5 FILLER_267_1406 ();
 b15zdnd11an1n64x5 FILLER_267_1470 ();
 b15zdnd11an1n64x5 FILLER_267_1534 ();
 b15zdnd11an1n64x5 FILLER_267_1598 ();
 b15zdnd11an1n64x5 FILLER_267_1662 ();
 b15zdnd11an1n64x5 FILLER_267_1726 ();
 b15zdnd11an1n16x5 FILLER_267_1790 ();
 b15zdnd11an1n08x5 FILLER_267_1806 ();
 b15zdnd11an1n64x5 FILLER_267_1820 ();
 b15zdnd11an1n64x5 FILLER_267_1884 ();
 b15zdnd00an1n02x5 FILLER_267_1948 ();
 b15zdnd00an1n01x5 FILLER_267_1950 ();
 b15zdnd11an1n64x5 FILLER_267_1955 ();
 b15zdnd11an1n32x5 FILLER_267_2019 ();
 b15zdnd11an1n16x5 FILLER_267_2051 ();
 b15zdnd11an1n08x5 FILLER_267_2067 ();
 b15zdnd11an1n04x5 FILLER_267_2075 ();
 b15zdnd11an1n64x5 FILLER_267_2121 ();
 b15zdnd11an1n16x5 FILLER_267_2185 ();
 b15zdnd11an1n04x5 FILLER_267_2201 ();
 b15zdnd00an1n02x5 FILLER_267_2205 ();
 b15zdnd00an1n01x5 FILLER_267_2207 ();
 b15zdnd11an1n64x5 FILLER_267_2214 ();
 b15zdnd11an1n04x5 FILLER_267_2278 ();
 b15zdnd00an1n02x5 FILLER_267_2282 ();
 b15zdnd11an1n64x5 FILLER_268_8 ();
 b15zdnd11an1n64x5 FILLER_268_72 ();
 b15zdnd11an1n64x5 FILLER_268_136 ();
 b15zdnd11an1n64x5 FILLER_268_200 ();
 b15zdnd11an1n64x5 FILLER_268_264 ();
 b15zdnd00an1n01x5 FILLER_268_328 ();
 b15zdnd11an1n04x5 FILLER_268_332 ();
 b15zdnd11an1n32x5 FILLER_268_339 ();
 b15zdnd11an1n08x5 FILLER_268_371 ();
 b15zdnd11an1n04x5 FILLER_268_379 ();
 b15zdnd11an1n04x5 FILLER_268_387 ();
 b15zdnd11an1n04x5 FILLER_268_396 ();
 b15zdnd00an1n01x5 FILLER_268_400 ();
 b15zdnd11an1n04x5 FILLER_268_417 ();
 b15zdnd00an1n02x5 FILLER_268_421 ();
 b15zdnd00an1n01x5 FILLER_268_423 ();
 b15zdnd11an1n64x5 FILLER_268_429 ();
 b15zdnd11an1n64x5 FILLER_268_493 ();
 b15zdnd11an1n64x5 FILLER_268_557 ();
 b15zdnd11an1n64x5 FILLER_268_621 ();
 b15zdnd11an1n32x5 FILLER_268_685 ();
 b15zdnd00an1n01x5 FILLER_268_717 ();
 b15zdnd11an1n64x5 FILLER_268_726 ();
 b15zdnd11an1n64x5 FILLER_268_790 ();
 b15zdnd11an1n64x5 FILLER_268_854 ();
 b15zdnd11an1n64x5 FILLER_268_918 ();
 b15zdnd11an1n64x5 FILLER_268_982 ();
 b15zdnd11an1n64x5 FILLER_268_1046 ();
 b15zdnd11an1n64x5 FILLER_268_1110 ();
 b15zdnd11an1n64x5 FILLER_268_1216 ();
 b15zdnd11an1n64x5 FILLER_268_1280 ();
 b15zdnd11an1n64x5 FILLER_268_1344 ();
 b15zdnd11an1n64x5 FILLER_268_1408 ();
 b15zdnd11an1n64x5 FILLER_268_1472 ();
 b15zdnd11an1n64x5 FILLER_268_1536 ();
 b15zdnd11an1n64x5 FILLER_268_1600 ();
 b15zdnd11an1n64x5 FILLER_268_1664 ();
 b15zdnd11an1n64x5 FILLER_268_1728 ();
 b15zdnd11an1n64x5 FILLER_268_1792 ();
 b15zdnd11an1n64x5 FILLER_268_1856 ();
 b15zdnd11an1n16x5 FILLER_268_1920 ();
 b15zdnd11an1n08x5 FILLER_268_1936 ();
 b15zdnd11an1n04x5 FILLER_268_1944 ();
 b15zdnd00an1n02x5 FILLER_268_1948 ();
 b15zdnd00an1n01x5 FILLER_268_1950 ();
 b15zdnd11an1n64x5 FILLER_268_1958 ();
 b15zdnd11an1n64x5 FILLER_268_2022 ();
 b15zdnd11an1n64x5 FILLER_268_2086 ();
 b15zdnd11an1n04x5 FILLER_268_2150 ();
 b15zdnd11an1n64x5 FILLER_268_2162 ();
 b15zdnd11an1n32x5 FILLER_268_2226 ();
 b15zdnd11an1n16x5 FILLER_268_2258 ();
 b15zdnd00an1n02x5 FILLER_268_2274 ();
 b15zdnd11an1n64x5 FILLER_269_0 ();
 b15zdnd11an1n64x5 FILLER_269_64 ();
 b15zdnd11an1n64x5 FILLER_269_128 ();
 b15zdnd11an1n64x5 FILLER_269_192 ();
 b15zdnd11an1n32x5 FILLER_269_256 ();
 b15zdnd11an1n16x5 FILLER_269_288 ();
 b15zdnd00an1n02x5 FILLER_269_304 ();
 b15zdnd00an1n01x5 FILLER_269_306 ();
 b15zdnd11an1n04x5 FILLER_269_359 ();
 b15zdnd11an1n08x5 FILLER_269_405 ();
 b15zdnd11an1n04x5 FILLER_269_413 ();
 b15zdnd11an1n64x5 FILLER_269_424 ();
 b15zdnd11an1n64x5 FILLER_269_488 ();
 b15zdnd11an1n64x5 FILLER_269_552 ();
 b15zdnd11an1n64x5 FILLER_269_616 ();
 b15zdnd11an1n64x5 FILLER_269_680 ();
 b15zdnd11an1n64x5 FILLER_269_744 ();
 b15zdnd11an1n32x5 FILLER_269_808 ();
 b15zdnd11an1n08x5 FILLER_269_840 ();
 b15zdnd00an1n01x5 FILLER_269_848 ();
 b15zdnd11an1n64x5 FILLER_269_852 ();
 b15zdnd11an1n32x5 FILLER_269_916 ();
 b15zdnd00an1n01x5 FILLER_269_948 ();
 b15zdnd11an1n64x5 FILLER_269_991 ();
 b15zdnd11an1n64x5 FILLER_269_1055 ();
 b15zdnd11an1n64x5 FILLER_269_1119 ();
 b15zdnd11an1n64x5 FILLER_269_1183 ();
 b15zdnd11an1n64x5 FILLER_269_1247 ();
 b15zdnd11an1n64x5 FILLER_269_1311 ();
 b15zdnd11an1n64x5 FILLER_269_1375 ();
 b15zdnd11an1n64x5 FILLER_269_1439 ();
 b15zdnd11an1n32x5 FILLER_269_1503 ();
 b15zdnd11an1n16x5 FILLER_269_1535 ();
 b15zdnd11an1n08x5 FILLER_269_1551 ();
 b15zdnd11an1n04x5 FILLER_269_1559 ();
 b15zdnd11an1n64x5 FILLER_269_1568 ();
 b15zdnd11an1n64x5 FILLER_269_1632 ();
 b15zdnd11an1n64x5 FILLER_269_1696 ();
 b15zdnd11an1n64x5 FILLER_269_1760 ();
 b15zdnd11an1n64x5 FILLER_269_1824 ();
 b15zdnd11an1n64x5 FILLER_269_1888 ();
 b15zdnd11an1n64x5 FILLER_269_1952 ();
 b15zdnd11an1n64x5 FILLER_269_2016 ();
 b15zdnd11an1n64x5 FILLER_269_2080 ();
 b15zdnd11an1n64x5 FILLER_269_2144 ();
 b15zdnd11an1n16x5 FILLER_269_2208 ();
 b15zdnd11an1n08x5 FILLER_269_2224 ();
 b15zdnd00an1n02x5 FILLER_269_2232 ();
 b15zdnd11an1n08x5 FILLER_269_2276 ();
 b15zdnd11an1n64x5 FILLER_270_8 ();
 b15zdnd11an1n64x5 FILLER_270_72 ();
 b15zdnd11an1n64x5 FILLER_270_136 ();
 b15zdnd11an1n64x5 FILLER_270_200 ();
 b15zdnd11an1n64x5 FILLER_270_264 ();
 b15zdnd11an1n32x5 FILLER_270_331 ();
 b15zdnd11an1n16x5 FILLER_270_363 ();
 b15zdnd11an1n08x5 FILLER_270_379 ();
 b15zdnd00an1n01x5 FILLER_270_387 ();
 b15zdnd11an1n04x5 FILLER_270_393 ();
 b15zdnd11an1n04x5 FILLER_270_413 ();
 b15zdnd00an1n02x5 FILLER_270_417 ();
 b15zdnd11an1n64x5 FILLER_270_422 ();
 b15zdnd11an1n64x5 FILLER_270_486 ();
 b15zdnd11an1n64x5 FILLER_270_550 ();
 b15zdnd11an1n64x5 FILLER_270_614 ();
 b15zdnd11an1n32x5 FILLER_270_678 ();
 b15zdnd11an1n08x5 FILLER_270_710 ();
 b15zdnd11an1n64x5 FILLER_270_726 ();
 b15zdnd11an1n16x5 FILLER_270_790 ();
 b15zdnd11an1n04x5 FILLER_270_806 ();
 b15zdnd00an1n02x5 FILLER_270_810 ();
 b15zdnd00an1n01x5 FILLER_270_812 ();
 b15zdnd11an1n64x5 FILLER_270_853 ();
 b15zdnd11an1n64x5 FILLER_270_917 ();
 b15zdnd11an1n64x5 FILLER_270_981 ();
 b15zdnd11an1n64x5 FILLER_270_1045 ();
 b15zdnd11an1n64x5 FILLER_270_1109 ();
 b15zdnd11an1n64x5 FILLER_270_1173 ();
 b15zdnd11an1n64x5 FILLER_270_1237 ();
 b15zdnd11an1n64x5 FILLER_270_1301 ();
 b15zdnd11an1n64x5 FILLER_270_1365 ();
 b15zdnd11an1n64x5 FILLER_270_1429 ();
 b15zdnd11an1n32x5 FILLER_270_1493 ();
 b15zdnd11an1n16x5 FILLER_270_1525 ();
 b15zdnd11an1n08x5 FILLER_270_1541 ();
 b15zdnd00an1n01x5 FILLER_270_1549 ();
 b15zdnd11an1n08x5 FILLER_270_1555 ();
 b15zdnd00an1n01x5 FILLER_270_1563 ();
 b15zdnd11an1n04x5 FILLER_270_1571 ();
 b15zdnd11an1n64x5 FILLER_270_1578 ();
 b15zdnd11an1n64x5 FILLER_270_1642 ();
 b15zdnd11an1n64x5 FILLER_270_1706 ();
 b15zdnd11an1n32x5 FILLER_270_1770 ();
 b15zdnd11an1n08x5 FILLER_270_1802 ();
 b15zdnd11an1n04x5 FILLER_270_1810 ();
 b15zdnd00an1n01x5 FILLER_270_1814 ();
 b15zdnd11an1n64x5 FILLER_270_1818 ();
 b15zdnd11an1n64x5 FILLER_270_1882 ();
 b15zdnd11an1n64x5 FILLER_270_1946 ();
 b15zdnd11an1n64x5 FILLER_270_2010 ();
 b15zdnd11an1n64x5 FILLER_270_2074 ();
 b15zdnd11an1n16x5 FILLER_270_2138 ();
 b15zdnd11an1n32x5 FILLER_270_2162 ();
 b15zdnd11an1n16x5 FILLER_270_2194 ();
 b15zdnd11an1n08x5 FILLER_270_2210 ();
 b15zdnd11an1n04x5 FILLER_270_2218 ();
 b15zdnd00an1n02x5 FILLER_270_2222 ();
 b15zdnd00an1n01x5 FILLER_270_2224 ();
 b15zdnd11an1n08x5 FILLER_270_2267 ();
 b15zdnd00an1n01x5 FILLER_270_2275 ();
 b15zdnd11an1n64x5 FILLER_271_0 ();
 b15zdnd11an1n04x5 FILLER_271_64 ();
 b15zdnd00an1n02x5 FILLER_271_68 ();
 b15zdnd00an1n01x5 FILLER_271_70 ();
 b15zdnd11an1n64x5 FILLER_271_82 ();
 b15zdnd11an1n32x5 FILLER_271_146 ();
 b15zdnd00an1n02x5 FILLER_271_178 ();
 b15zdnd11an1n04x5 FILLER_271_183 ();
 b15zdnd11an1n08x5 FILLER_271_190 ();
 b15zdnd00an1n02x5 FILLER_271_198 ();
 b15zdnd11an1n64x5 FILLER_271_203 ();
 b15zdnd11an1n64x5 FILLER_271_267 ();
 b15zdnd11an1n32x5 FILLER_271_331 ();
 b15zdnd11an1n16x5 FILLER_271_363 ();
 b15zdnd11an1n08x5 FILLER_271_379 ();
 b15zdnd00an1n01x5 FILLER_271_387 ();
 b15zdnd11an1n64x5 FILLER_271_399 ();
 b15zdnd11an1n64x5 FILLER_271_463 ();
 b15zdnd11an1n64x5 FILLER_271_527 ();
 b15zdnd11an1n64x5 FILLER_271_591 ();
 b15zdnd11an1n64x5 FILLER_271_655 ();
 b15zdnd11an1n64x5 FILLER_271_719 ();
 b15zdnd11an1n64x5 FILLER_271_783 ();
 b15zdnd00an1n02x5 FILLER_271_847 ();
 b15zdnd00an1n01x5 FILLER_271_849 ();
 b15zdnd11an1n64x5 FILLER_271_853 ();
 b15zdnd11an1n08x5 FILLER_271_917 ();
 b15zdnd00an1n02x5 FILLER_271_925 ();
 b15zdnd00an1n01x5 FILLER_271_927 ();
 b15zdnd11an1n64x5 FILLER_271_931 ();
 b15zdnd11an1n64x5 FILLER_271_995 ();
 b15zdnd11an1n64x5 FILLER_271_1059 ();
 b15zdnd11an1n64x5 FILLER_271_1123 ();
 b15zdnd11an1n64x5 FILLER_271_1187 ();
 b15zdnd11an1n64x5 FILLER_271_1251 ();
 b15zdnd11an1n64x5 FILLER_271_1315 ();
 b15zdnd11an1n64x5 FILLER_271_1379 ();
 b15zdnd11an1n64x5 FILLER_271_1443 ();
 b15zdnd11an1n32x5 FILLER_271_1507 ();
 b15zdnd11an1n08x5 FILLER_271_1539 ();
 b15zdnd11an1n04x5 FILLER_271_1560 ();
 b15zdnd11an1n04x5 FILLER_271_1574 ();
 b15zdnd00an1n02x5 FILLER_271_1578 ();
 b15zdnd00an1n01x5 FILLER_271_1580 ();
 b15zdnd11an1n64x5 FILLER_271_1623 ();
 b15zdnd11an1n64x5 FILLER_271_1687 ();
 b15zdnd11an1n64x5 FILLER_271_1751 ();
 b15zdnd11an1n64x5 FILLER_271_1815 ();
 b15zdnd11an1n64x5 FILLER_271_1879 ();
 b15zdnd11an1n64x5 FILLER_271_1943 ();
 b15zdnd11an1n64x5 FILLER_271_2007 ();
 b15zdnd11an1n64x5 FILLER_271_2071 ();
 b15zdnd11an1n32x5 FILLER_271_2135 ();
 b15zdnd11an1n16x5 FILLER_271_2167 ();
 b15zdnd11an1n08x5 FILLER_271_2183 ();
 b15zdnd00an1n02x5 FILLER_271_2191 ();
 b15zdnd00an1n01x5 FILLER_271_2193 ();
 b15zdnd11an1n32x5 FILLER_271_2236 ();
 b15zdnd11an1n16x5 FILLER_271_2268 ();
 b15zdnd11an1n64x5 FILLER_272_8 ();
 b15zdnd11an1n64x5 FILLER_272_72 ();
 b15zdnd11an1n16x5 FILLER_272_136 ();
 b15zdnd11an1n04x5 FILLER_272_152 ();
 b15zdnd00an1n01x5 FILLER_272_156 ();
 b15zdnd11an1n32x5 FILLER_272_209 ();
 b15zdnd11an1n16x5 FILLER_272_241 ();
 b15zdnd11an1n08x5 FILLER_272_257 ();
 b15zdnd11an1n04x5 FILLER_272_265 ();
 b15zdnd00an1n02x5 FILLER_272_269 ();
 b15zdnd00an1n01x5 FILLER_272_271 ();
 b15zdnd11an1n04x5 FILLER_272_275 ();
 b15zdnd11an1n64x5 FILLER_272_282 ();
 b15zdnd11an1n64x5 FILLER_272_346 ();
 b15zdnd11an1n64x5 FILLER_272_410 ();
 b15zdnd11an1n32x5 FILLER_272_474 ();
 b15zdnd11an1n16x5 FILLER_272_506 ();
 b15zdnd11an1n04x5 FILLER_272_522 ();
 b15zdnd00an1n02x5 FILLER_272_526 ();
 b15zdnd00an1n01x5 FILLER_272_528 ();
 b15zdnd11an1n64x5 FILLER_272_571 ();
 b15zdnd11an1n64x5 FILLER_272_635 ();
 b15zdnd11an1n16x5 FILLER_272_699 ();
 b15zdnd00an1n02x5 FILLER_272_715 ();
 b15zdnd00an1n01x5 FILLER_272_717 ();
 b15zdnd11an1n64x5 FILLER_272_726 ();
 b15zdnd11an1n64x5 FILLER_272_790 ();
 b15zdnd11an1n32x5 FILLER_272_854 ();
 b15zdnd11an1n04x5 FILLER_272_886 ();
 b15zdnd00an1n02x5 FILLER_272_890 ();
 b15zdnd11an1n04x5 FILLER_272_932 ();
 b15zdnd11an1n64x5 FILLER_272_939 ();
 b15zdnd11an1n64x5 FILLER_272_1003 ();
 b15zdnd11an1n64x5 FILLER_272_1067 ();
 b15zdnd11an1n64x5 FILLER_272_1131 ();
 b15zdnd11an1n64x5 FILLER_272_1195 ();
 b15zdnd11an1n16x5 FILLER_272_1259 ();
 b15zdnd11an1n08x5 FILLER_272_1275 ();
 b15zdnd11an1n04x5 FILLER_272_1283 ();
 b15zdnd00an1n02x5 FILLER_272_1287 ();
 b15zdnd11an1n32x5 FILLER_272_1292 ();
 b15zdnd11an1n04x5 FILLER_272_1324 ();
 b15zdnd00an1n02x5 FILLER_272_1328 ();
 b15zdnd00an1n01x5 FILLER_272_1330 ();
 b15zdnd11an1n64x5 FILLER_272_1334 ();
 b15zdnd11an1n64x5 FILLER_272_1398 ();
 b15zdnd11an1n64x5 FILLER_272_1462 ();
 b15zdnd11an1n04x5 FILLER_272_1526 ();
 b15zdnd11an1n04x5 FILLER_272_1534 ();
 b15zdnd11an1n04x5 FILLER_272_1551 ();
 b15zdnd11an1n04x5 FILLER_272_1597 ();
 b15zdnd00an1n02x5 FILLER_272_1601 ();
 b15zdnd00an1n01x5 FILLER_272_1603 ();
 b15zdnd11an1n64x5 FILLER_272_1608 ();
 b15zdnd11an1n32x5 FILLER_272_1672 ();
 b15zdnd11an1n16x5 FILLER_272_1704 ();
 b15zdnd11an1n08x5 FILLER_272_1720 ();
 b15zdnd11an1n04x5 FILLER_272_1728 ();
 b15zdnd00an1n01x5 FILLER_272_1732 ();
 b15zdnd11an1n04x5 FILLER_272_1736 ();
 b15zdnd11an1n04x5 FILLER_272_1743 ();
 b15zdnd11an1n64x5 FILLER_272_1750 ();
 b15zdnd11an1n64x5 FILLER_272_1814 ();
 b15zdnd11an1n64x5 FILLER_272_1878 ();
 b15zdnd11an1n04x5 FILLER_272_1942 ();
 b15zdnd11an1n16x5 FILLER_272_1949 ();
 b15zdnd11an1n08x5 FILLER_272_1965 ();
 b15zdnd00an1n01x5 FILLER_272_1973 ();
 b15zdnd11an1n64x5 FILLER_272_2016 ();
 b15zdnd11an1n64x5 FILLER_272_2080 ();
 b15zdnd11an1n08x5 FILLER_272_2144 ();
 b15zdnd00an1n02x5 FILLER_272_2152 ();
 b15zdnd11an1n32x5 FILLER_272_2162 ();
 b15zdnd11an1n04x5 FILLER_272_2194 ();
 b15zdnd11an1n32x5 FILLER_272_2229 ();
 b15zdnd11an1n08x5 FILLER_272_2261 ();
 b15zdnd11an1n04x5 FILLER_272_2269 ();
 b15zdnd00an1n02x5 FILLER_272_2273 ();
 b15zdnd00an1n01x5 FILLER_272_2275 ();
 b15zdnd11an1n64x5 FILLER_273_0 ();
 b15zdnd11an1n64x5 FILLER_273_64 ();
 b15zdnd11an1n64x5 FILLER_273_128 ();
 b15zdnd11an1n32x5 FILLER_273_192 ();
 b15zdnd11an1n16x5 FILLER_273_224 ();
 b15zdnd11an1n04x5 FILLER_273_240 ();
 b15zdnd11an1n64x5 FILLER_273_286 ();
 b15zdnd11an1n64x5 FILLER_273_350 ();
 b15zdnd11an1n64x5 FILLER_273_414 ();
 b15zdnd11an1n64x5 FILLER_273_478 ();
 b15zdnd11an1n64x5 FILLER_273_542 ();
 b15zdnd11an1n64x5 FILLER_273_606 ();
 b15zdnd11an1n64x5 FILLER_273_670 ();
 b15zdnd11an1n64x5 FILLER_273_734 ();
 b15zdnd11an1n64x5 FILLER_273_798 ();
 b15zdnd11an1n64x5 FILLER_273_862 ();
 b15zdnd11an1n64x5 FILLER_273_926 ();
 b15zdnd11an1n64x5 FILLER_273_990 ();
 b15zdnd11an1n64x5 FILLER_273_1054 ();
 b15zdnd11an1n64x5 FILLER_273_1118 ();
 b15zdnd11an1n64x5 FILLER_273_1182 ();
 b15zdnd11an1n16x5 FILLER_273_1246 ();
 b15zdnd11an1n08x5 FILLER_273_1262 ();
 b15zdnd00an1n01x5 FILLER_273_1270 ();
 b15zdnd11an1n08x5 FILLER_273_1278 ();
 b15zdnd11an1n04x5 FILLER_273_1289 ();
 b15zdnd11an1n64x5 FILLER_273_1296 ();
 b15zdnd11an1n64x5 FILLER_273_1360 ();
 b15zdnd11an1n64x5 FILLER_273_1424 ();
 b15zdnd11an1n16x5 FILLER_273_1488 ();
 b15zdnd00an1n02x5 FILLER_273_1504 ();
 b15zdnd11an1n08x5 FILLER_273_1509 ();
 b15zdnd00an1n02x5 FILLER_273_1517 ();
 b15zdnd00an1n01x5 FILLER_273_1519 ();
 b15zdnd11an1n04x5 FILLER_273_1562 ();
 b15zdnd11an1n04x5 FILLER_273_1571 ();
 b15zdnd00an1n01x5 FILLER_273_1575 ();
 b15zdnd11an1n64x5 FILLER_273_1628 ();
 b15zdnd11an1n16x5 FILLER_273_1692 ();
 b15zdnd11an1n04x5 FILLER_273_1708 ();
 b15zdnd11an1n64x5 FILLER_273_1764 ();
 b15zdnd11an1n64x5 FILLER_273_1828 ();
 b15zdnd11an1n32x5 FILLER_273_1892 ();
 b15zdnd11an1n04x5 FILLER_273_1924 ();
 b15zdnd00an1n01x5 FILLER_273_1928 ();
 b15zdnd11an1n04x5 FILLER_273_1932 ();
 b15zdnd11an1n04x5 FILLER_273_1939 ();
 b15zdnd11an1n08x5 FILLER_273_1949 ();
 b15zdnd11an1n04x5 FILLER_273_1957 ();
 b15zdnd11an1n64x5 FILLER_273_1965 ();
 b15zdnd11an1n32x5 FILLER_273_2029 ();
 b15zdnd11an1n04x5 FILLER_273_2061 ();
 b15zdnd00an1n01x5 FILLER_273_2065 ();
 b15zdnd11an1n64x5 FILLER_273_2084 ();
 b15zdnd11an1n64x5 FILLER_273_2148 ();
 b15zdnd11an1n04x5 FILLER_273_2212 ();
 b15zdnd00an1n01x5 FILLER_273_2216 ();
 b15zdnd11an1n04x5 FILLER_273_2220 ();
 b15zdnd11an1n32x5 FILLER_273_2227 ();
 b15zdnd11an1n16x5 FILLER_273_2259 ();
 b15zdnd11an1n08x5 FILLER_273_2275 ();
 b15zdnd00an1n01x5 FILLER_273_2283 ();
 b15zdnd11an1n64x5 FILLER_274_8 ();
 b15zdnd11an1n64x5 FILLER_274_72 ();
 b15zdnd11an1n64x5 FILLER_274_136 ();
 b15zdnd11an1n32x5 FILLER_274_200 ();
 b15zdnd11an1n16x5 FILLER_274_232 ();
 b15zdnd00an1n01x5 FILLER_274_248 ();
 b15zdnd11an1n64x5 FILLER_274_301 ();
 b15zdnd11an1n64x5 FILLER_274_365 ();
 b15zdnd11an1n64x5 FILLER_274_429 ();
 b15zdnd11an1n64x5 FILLER_274_493 ();
 b15zdnd11an1n64x5 FILLER_274_557 ();
 b15zdnd11an1n64x5 FILLER_274_621 ();
 b15zdnd11an1n32x5 FILLER_274_685 ();
 b15zdnd00an1n01x5 FILLER_274_717 ();
 b15zdnd11an1n64x5 FILLER_274_726 ();
 b15zdnd11an1n64x5 FILLER_274_790 ();
 b15zdnd11an1n64x5 FILLER_274_854 ();
 b15zdnd11an1n64x5 FILLER_274_918 ();
 b15zdnd11an1n64x5 FILLER_274_982 ();
 b15zdnd11an1n64x5 FILLER_274_1046 ();
 b15zdnd11an1n32x5 FILLER_274_1110 ();
 b15zdnd11an1n08x5 FILLER_274_1142 ();
 b15zdnd11an1n04x5 FILLER_274_1150 ();
 b15zdnd00an1n02x5 FILLER_274_1154 ();
 b15zdnd00an1n01x5 FILLER_274_1156 ();
 b15zdnd11an1n04x5 FILLER_274_1160 ();
 b15zdnd11an1n64x5 FILLER_274_1167 ();
 b15zdnd11an1n32x5 FILLER_274_1231 ();
 b15zdnd11an1n08x5 FILLER_274_1315 ();
 b15zdnd00an1n02x5 FILLER_274_1323 ();
 b15zdnd11an1n64x5 FILLER_274_1332 ();
 b15zdnd11an1n64x5 FILLER_274_1396 ();
 b15zdnd11an1n16x5 FILLER_274_1460 ();
 b15zdnd11an1n08x5 FILLER_274_1476 ();
 b15zdnd00an1n02x5 FILLER_274_1484 ();
 b15zdnd11an1n04x5 FILLER_274_1538 ();
 b15zdnd11an1n04x5 FILLER_274_1584 ();
 b15zdnd11an1n64x5 FILLER_274_1630 ();
 b15zdnd11an1n32x5 FILLER_274_1694 ();
 b15zdnd11an1n04x5 FILLER_274_1726 ();
 b15zdnd11an1n04x5 FILLER_274_1733 ();
 b15zdnd11an1n64x5 FILLER_274_1740 ();
 b15zdnd11an1n64x5 FILLER_274_1804 ();
 b15zdnd11an1n32x5 FILLER_274_1868 ();
 b15zdnd11an1n08x5 FILLER_274_1900 ();
 b15zdnd00an1n01x5 FILLER_274_1908 ();
 b15zdnd11an1n64x5 FILLER_274_1961 ();
 b15zdnd11an1n32x5 FILLER_274_2025 ();
 b15zdnd11an1n16x5 FILLER_274_2057 ();
 b15zdnd11an1n08x5 FILLER_274_2073 ();
 b15zdnd00an1n01x5 FILLER_274_2081 ();
 b15zdnd11an1n32x5 FILLER_274_2113 ();
 b15zdnd11an1n08x5 FILLER_274_2145 ();
 b15zdnd00an1n01x5 FILLER_274_2153 ();
 b15zdnd11an1n16x5 FILLER_274_2162 ();
 b15zdnd11an1n08x5 FILLER_274_2178 ();
 b15zdnd11an1n04x5 FILLER_274_2193 ();
 b15zdnd00an1n02x5 FILLER_274_2197 ();
 b15zdnd11an1n16x5 FILLER_274_2251 ();
 b15zdnd11an1n08x5 FILLER_274_2267 ();
 b15zdnd00an1n01x5 FILLER_274_2275 ();
 b15zdnd11an1n64x5 FILLER_275_0 ();
 b15zdnd11an1n64x5 FILLER_275_64 ();
 b15zdnd11an1n64x5 FILLER_275_128 ();
 b15zdnd11an1n64x5 FILLER_275_192 ();
 b15zdnd11an1n08x5 FILLER_275_256 ();
 b15zdnd11an1n04x5 FILLER_275_264 ();
 b15zdnd00an1n01x5 FILLER_275_268 ();
 b15zdnd11an1n04x5 FILLER_275_272 ();
 b15zdnd11an1n04x5 FILLER_275_279 ();
 b15zdnd11an1n64x5 FILLER_275_286 ();
 b15zdnd11an1n64x5 FILLER_275_350 ();
 b15zdnd11an1n64x5 FILLER_275_414 ();
 b15zdnd11an1n64x5 FILLER_275_478 ();
 b15zdnd11an1n64x5 FILLER_275_542 ();
 b15zdnd11an1n64x5 FILLER_275_606 ();
 b15zdnd11an1n64x5 FILLER_275_670 ();
 b15zdnd11an1n64x5 FILLER_275_734 ();
 b15zdnd11an1n64x5 FILLER_275_798 ();
 b15zdnd11an1n64x5 FILLER_275_862 ();
 b15zdnd11an1n64x5 FILLER_275_926 ();
 b15zdnd11an1n16x5 FILLER_275_990 ();
 b15zdnd11an1n08x5 FILLER_275_1006 ();
 b15zdnd11an1n04x5 FILLER_275_1014 ();
 b15zdnd11an1n32x5 FILLER_275_1070 ();
 b15zdnd11an1n16x5 FILLER_275_1102 ();
 b15zdnd11an1n08x5 FILLER_275_1118 ();
 b15zdnd11an1n04x5 FILLER_275_1126 ();
 b15zdnd00an1n02x5 FILLER_275_1130 ();
 b15zdnd11an1n64x5 FILLER_275_1184 ();
 b15zdnd11an1n16x5 FILLER_275_1248 ();
 b15zdnd11an1n08x5 FILLER_275_1264 ();
 b15zdnd11an1n04x5 FILLER_275_1285 ();
 b15zdnd11an1n64x5 FILLER_275_1331 ();
 b15zdnd11an1n08x5 FILLER_275_1395 ();
 b15zdnd11an1n04x5 FILLER_275_1403 ();
 b15zdnd00an1n01x5 FILLER_275_1407 ();
 b15zdnd11an1n64x5 FILLER_275_1411 ();
 b15zdnd11an1n32x5 FILLER_275_1475 ();
 b15zdnd00an1n01x5 FILLER_275_1507 ();
 b15zdnd11an1n04x5 FILLER_275_1511 ();
 b15zdnd00an1n01x5 FILLER_275_1515 ();
 b15zdnd11an1n16x5 FILLER_275_1519 ();
 b15zdnd11an1n04x5 FILLER_275_1535 ();
 b15zdnd00an1n02x5 FILLER_275_1539 ();
 b15zdnd00an1n01x5 FILLER_275_1541 ();
 b15zdnd11an1n16x5 FILLER_275_1584 ();
 b15zdnd00an1n02x5 FILLER_275_1600 ();
 b15zdnd00an1n01x5 FILLER_275_1602 ();
 b15zdnd11an1n04x5 FILLER_275_1606 ();
 b15zdnd00an1n01x5 FILLER_275_1610 ();
 b15zdnd11an1n64x5 FILLER_275_1614 ();
 b15zdnd11an1n64x5 FILLER_275_1678 ();
 b15zdnd11an1n64x5 FILLER_275_1742 ();
 b15zdnd11an1n64x5 FILLER_275_1806 ();
 b15zdnd11an1n32x5 FILLER_275_1870 ();
 b15zdnd11an1n16x5 FILLER_275_1902 ();
 b15zdnd11an1n08x5 FILLER_275_1918 ();
 b15zdnd00an1n01x5 FILLER_275_1926 ();
 b15zdnd11an1n04x5 FILLER_275_1930 ();
 b15zdnd11an1n04x5 FILLER_275_1937 ();
 b15zdnd11an1n64x5 FILLER_275_1944 ();
 b15zdnd11an1n64x5 FILLER_275_2008 ();
 b15zdnd00an1n02x5 FILLER_275_2072 ();
 b15zdnd11an1n08x5 FILLER_275_2077 ();
 b15zdnd11an1n04x5 FILLER_275_2085 ();
 b15zdnd11an1n32x5 FILLER_275_2131 ();
 b15zdnd11an1n08x5 FILLER_275_2163 ();
 b15zdnd11an1n04x5 FILLER_275_2171 ();
 b15zdnd00an1n01x5 FILLER_275_2175 ();
 b15zdnd11an1n04x5 FILLER_275_2228 ();
 b15zdnd11an1n32x5 FILLER_275_2235 ();
 b15zdnd11an1n16x5 FILLER_275_2267 ();
 b15zdnd00an1n01x5 FILLER_275_2283 ();
 b15zdnd11an1n64x5 FILLER_276_8 ();
 b15zdnd11an1n64x5 FILLER_276_72 ();
 b15zdnd11an1n08x5 FILLER_276_136 ();
 b15zdnd00an1n02x5 FILLER_276_144 ();
 b15zdnd11an1n64x5 FILLER_276_150 ();
 b15zdnd11an1n64x5 FILLER_276_214 ();
 b15zdnd11an1n64x5 FILLER_276_278 ();
 b15zdnd11an1n64x5 FILLER_276_342 ();
 b15zdnd11an1n64x5 FILLER_276_406 ();
 b15zdnd11an1n64x5 FILLER_276_470 ();
 b15zdnd11an1n64x5 FILLER_276_534 ();
 b15zdnd11an1n64x5 FILLER_276_598 ();
 b15zdnd11an1n32x5 FILLER_276_662 ();
 b15zdnd11an1n16x5 FILLER_276_694 ();
 b15zdnd11an1n08x5 FILLER_276_710 ();
 b15zdnd00an1n02x5 FILLER_276_726 ();
 b15zdnd11an1n64x5 FILLER_276_731 ();
 b15zdnd11an1n64x5 FILLER_276_795 ();
 b15zdnd11an1n64x5 FILLER_276_859 ();
 b15zdnd11an1n64x5 FILLER_276_923 ();
 b15zdnd11an1n32x5 FILLER_276_987 ();
 b15zdnd11an1n16x5 FILLER_276_1019 ();
 b15zdnd11an1n08x5 FILLER_276_1035 ();
 b15zdnd11an1n04x5 FILLER_276_1046 ();
 b15zdnd11an1n64x5 FILLER_276_1053 ();
 b15zdnd11an1n32x5 FILLER_276_1117 ();
 b15zdnd11an1n08x5 FILLER_276_1149 ();
 b15zdnd11an1n64x5 FILLER_276_1160 ();
 b15zdnd11an1n32x5 FILLER_276_1224 ();
 b15zdnd11an1n16x5 FILLER_276_1256 ();
 b15zdnd11an1n04x5 FILLER_276_1272 ();
 b15zdnd00an1n02x5 FILLER_276_1276 ();
 b15zdnd00an1n01x5 FILLER_276_1278 ();
 b15zdnd11an1n64x5 FILLER_276_1321 ();
 b15zdnd11an1n08x5 FILLER_276_1385 ();
 b15zdnd11an1n04x5 FILLER_276_1393 ();
 b15zdnd00an1n02x5 FILLER_276_1397 ();
 b15zdnd00an1n01x5 FILLER_276_1399 ();
 b15zdnd11an1n04x5 FILLER_276_1403 ();
 b15zdnd11an1n64x5 FILLER_276_1410 ();
 b15zdnd11an1n64x5 FILLER_276_1474 ();
 b15zdnd11an1n04x5 FILLER_276_1538 ();
 b15zdnd11an1n32x5 FILLER_276_1553 ();
 b15zdnd11an1n16x5 FILLER_276_1585 ();
 b15zdnd11an1n04x5 FILLER_276_1601 ();
 b15zdnd00an1n02x5 FILLER_276_1605 ();
 b15zdnd00an1n01x5 FILLER_276_1607 ();
 b15zdnd11an1n64x5 FILLER_276_1611 ();
 b15zdnd11an1n64x5 FILLER_276_1675 ();
 b15zdnd11an1n64x5 FILLER_276_1739 ();
 b15zdnd11an1n64x5 FILLER_276_1803 ();
 b15zdnd11an1n64x5 FILLER_276_1867 ();
 b15zdnd11an1n08x5 FILLER_276_1931 ();
 b15zdnd11an1n04x5 FILLER_276_1939 ();
 b15zdnd00an1n02x5 FILLER_276_1943 ();
 b15zdnd00an1n01x5 FILLER_276_1945 ();
 b15zdnd11an1n64x5 FILLER_276_1950 ();
 b15zdnd11an1n32x5 FILLER_276_2014 ();
 b15zdnd00an1n01x5 FILLER_276_2046 ();
 b15zdnd11an1n32x5 FILLER_276_2099 ();
 b15zdnd11an1n16x5 FILLER_276_2131 ();
 b15zdnd11an1n04x5 FILLER_276_2147 ();
 b15zdnd00an1n02x5 FILLER_276_2151 ();
 b15zdnd00an1n01x5 FILLER_276_2153 ();
 b15zdnd11an1n16x5 FILLER_276_2162 ();
 b15zdnd11an1n04x5 FILLER_276_2178 ();
 b15zdnd11an1n04x5 FILLER_276_2188 ();
 b15zdnd00an1n02x5 FILLER_276_2192 ();
 b15zdnd11an1n32x5 FILLER_276_2236 ();
 b15zdnd11an1n08x5 FILLER_276_2268 ();
 b15zdnd11an1n64x5 FILLER_277_0 ();
 b15zdnd11an1n64x5 FILLER_277_64 ();
 b15zdnd11an1n16x5 FILLER_277_128 ();
 b15zdnd11an1n04x5 FILLER_277_149 ();
 b15zdnd11an1n64x5 FILLER_277_195 ();
 b15zdnd11an1n64x5 FILLER_277_259 ();
 b15zdnd11an1n64x5 FILLER_277_323 ();
 b15zdnd11an1n64x5 FILLER_277_387 ();
 b15zdnd11an1n64x5 FILLER_277_451 ();
 b15zdnd11an1n64x5 FILLER_277_515 ();
 b15zdnd11an1n64x5 FILLER_277_579 ();
 b15zdnd11an1n32x5 FILLER_277_643 ();
 b15zdnd11an1n16x5 FILLER_277_675 ();
 b15zdnd11an1n08x5 FILLER_277_691 ();
 b15zdnd00an1n02x5 FILLER_277_699 ();
 b15zdnd11an1n04x5 FILLER_277_717 ();
 b15zdnd00an1n02x5 FILLER_277_721 ();
 b15zdnd11an1n04x5 FILLER_277_726 ();
 b15zdnd11an1n04x5 FILLER_277_734 ();
 b15zdnd11an1n64x5 FILLER_277_741 ();
 b15zdnd11an1n64x5 FILLER_277_805 ();
 b15zdnd11an1n64x5 FILLER_277_869 ();
 b15zdnd11an1n64x5 FILLER_277_933 ();
 b15zdnd11an1n32x5 FILLER_277_997 ();
 b15zdnd11an1n08x5 FILLER_277_1029 ();
 b15zdnd11an1n04x5 FILLER_277_1037 ();
 b15zdnd11an1n64x5 FILLER_277_1044 ();
 b15zdnd11an1n64x5 FILLER_277_1108 ();
 b15zdnd11an1n64x5 FILLER_277_1172 ();
 b15zdnd11an1n32x5 FILLER_277_1236 ();
 b15zdnd00an1n01x5 FILLER_277_1268 ();
 b15zdnd11an1n64x5 FILLER_277_1311 ();
 b15zdnd11an1n04x5 FILLER_277_1375 ();
 b15zdnd00an1n01x5 FILLER_277_1379 ();
 b15zdnd11an1n64x5 FILLER_277_1432 ();
 b15zdnd11an1n64x5 FILLER_277_1496 ();
 b15zdnd11an1n64x5 FILLER_277_1560 ();
 b15zdnd11an1n64x5 FILLER_277_1624 ();
 b15zdnd11an1n64x5 FILLER_277_1688 ();
 b15zdnd11an1n64x5 FILLER_277_1752 ();
 b15zdnd11an1n64x5 FILLER_277_1816 ();
 b15zdnd11an1n64x5 FILLER_277_1880 ();
 b15zdnd11an1n64x5 FILLER_277_1944 ();
 b15zdnd11an1n32x5 FILLER_277_2008 ();
 b15zdnd11an1n16x5 FILLER_277_2040 ();
 b15zdnd11an1n04x5 FILLER_277_2056 ();
 b15zdnd00an1n02x5 FILLER_277_2060 ();
 b15zdnd11an1n08x5 FILLER_277_2065 ();
 b15zdnd00an1n01x5 FILLER_277_2073 ();
 b15zdnd11an1n04x5 FILLER_277_2078 ();
 b15zdnd11an1n64x5 FILLER_277_2124 ();
 b15zdnd11an1n08x5 FILLER_277_2188 ();
 b15zdnd00an1n02x5 FILLER_277_2196 ();
 b15zdnd00an1n01x5 FILLER_277_2198 ();
 b15zdnd11an1n04x5 FILLER_277_2202 ();
 b15zdnd11an1n04x5 FILLER_277_2209 ();
 b15zdnd11an1n64x5 FILLER_277_2216 ();
 b15zdnd11an1n04x5 FILLER_277_2280 ();
 b15zdnd11an1n64x5 FILLER_278_8 ();
 b15zdnd11an1n64x5 FILLER_278_72 ();
 b15zdnd11an1n64x5 FILLER_278_136 ();
 b15zdnd11an1n64x5 FILLER_278_200 ();
 b15zdnd11an1n64x5 FILLER_278_264 ();
 b15zdnd11an1n64x5 FILLER_278_328 ();
 b15zdnd11an1n32x5 FILLER_278_392 ();
 b15zdnd11an1n16x5 FILLER_278_424 ();
 b15zdnd11an1n04x5 FILLER_278_440 ();
 b15zdnd00an1n02x5 FILLER_278_444 ();
 b15zdnd00an1n01x5 FILLER_278_446 ();
 b15zdnd11an1n16x5 FILLER_278_489 ();
 b15zdnd00an1n02x5 FILLER_278_505 ();
 b15zdnd11an1n64x5 FILLER_278_510 ();
 b15zdnd11an1n64x5 FILLER_278_574 ();
 b15zdnd11an1n64x5 FILLER_278_638 ();
 b15zdnd00an1n02x5 FILLER_278_702 ();
 b15zdnd00an1n01x5 FILLER_278_704 ();
 b15zdnd00an1n02x5 FILLER_278_716 ();
 b15zdnd00an1n02x5 FILLER_278_726 ();
 b15zdnd11an1n08x5 FILLER_278_734 ();
 b15zdnd11an1n64x5 FILLER_278_784 ();
 b15zdnd11an1n64x5 FILLER_278_848 ();
 b15zdnd11an1n64x5 FILLER_278_912 ();
 b15zdnd11an1n64x5 FILLER_278_976 ();
 b15zdnd11an1n64x5 FILLER_278_1040 ();
 b15zdnd11an1n64x5 FILLER_278_1104 ();
 b15zdnd11an1n64x5 FILLER_278_1168 ();
 b15zdnd11an1n16x5 FILLER_278_1232 ();
 b15zdnd11an1n08x5 FILLER_278_1248 ();
 b15zdnd11an1n04x5 FILLER_278_1256 ();
 b15zdnd00an1n02x5 FILLER_278_1260 ();
 b15zdnd00an1n01x5 FILLER_278_1262 ();
 b15zdnd11an1n04x5 FILLER_278_1270 ();
 b15zdnd11an1n64x5 FILLER_278_1316 ();
 b15zdnd11an1n16x5 FILLER_278_1380 ();
 b15zdnd11an1n08x5 FILLER_278_1396 ();
 b15zdnd00an1n01x5 FILLER_278_1404 ();
 b15zdnd11an1n04x5 FILLER_278_1408 ();
 b15zdnd11an1n08x5 FILLER_278_1415 ();
 b15zdnd00an1n02x5 FILLER_278_1423 ();
 b15zdnd00an1n01x5 FILLER_278_1425 ();
 b15zdnd11an1n64x5 FILLER_278_1433 ();
 b15zdnd11an1n64x5 FILLER_278_1497 ();
 b15zdnd11an1n64x5 FILLER_278_1561 ();
 b15zdnd11an1n64x5 FILLER_278_1625 ();
 b15zdnd11an1n64x5 FILLER_278_1689 ();
 b15zdnd11an1n32x5 FILLER_278_1753 ();
 b15zdnd11an1n16x5 FILLER_278_1785 ();
 b15zdnd11an1n04x5 FILLER_278_1801 ();
 b15zdnd11an1n64x5 FILLER_278_1809 ();
 b15zdnd11an1n64x5 FILLER_278_1873 ();
 b15zdnd11an1n64x5 FILLER_278_1937 ();
 b15zdnd11an1n64x5 FILLER_278_2001 ();
 b15zdnd00an1n02x5 FILLER_278_2065 ();
 b15zdnd11an1n04x5 FILLER_278_2070 ();
 b15zdnd11an1n16x5 FILLER_278_2094 ();
 b15zdnd11an1n08x5 FILLER_278_2110 ();
 b15zdnd11an1n04x5 FILLER_278_2118 ();
 b15zdnd00an1n02x5 FILLER_278_2122 ();
 b15zdnd00an1n01x5 FILLER_278_2124 ();
 b15zdnd11an1n16x5 FILLER_278_2128 ();
 b15zdnd11an1n08x5 FILLER_278_2144 ();
 b15zdnd00an1n02x5 FILLER_278_2152 ();
 b15zdnd11an1n64x5 FILLER_278_2162 ();
 b15zdnd11an1n32x5 FILLER_278_2226 ();
 b15zdnd11an1n16x5 FILLER_278_2258 ();
 b15zdnd00an1n02x5 FILLER_278_2274 ();
 b15zdnd11an1n64x5 FILLER_279_0 ();
 b15zdnd11an1n64x5 FILLER_279_64 ();
 b15zdnd11an1n08x5 FILLER_279_128 ();
 b15zdnd11an1n04x5 FILLER_279_136 ();
 b15zdnd00an1n01x5 FILLER_279_140 ();
 b15zdnd11an1n04x5 FILLER_279_157 ();
 b15zdnd11an1n64x5 FILLER_279_172 ();
 b15zdnd11an1n64x5 FILLER_279_236 ();
 b15zdnd11an1n64x5 FILLER_279_300 ();
 b15zdnd11an1n64x5 FILLER_279_364 ();
 b15zdnd11an1n32x5 FILLER_279_428 ();
 b15zdnd11an1n16x5 FILLER_279_460 ();
 b15zdnd11an1n04x5 FILLER_279_476 ();
 b15zdnd11an1n32x5 FILLER_279_532 ();
 b15zdnd11an1n16x5 FILLER_279_564 ();
 b15zdnd00an1n02x5 FILLER_279_580 ();
 b15zdnd11an1n64x5 FILLER_279_589 ();
 b15zdnd11an1n32x5 FILLER_279_653 ();
 b15zdnd11an1n04x5 FILLER_279_685 ();
 b15zdnd00an1n02x5 FILLER_279_689 ();
 b15zdnd00an1n01x5 FILLER_279_691 ();
 b15zdnd11an1n04x5 FILLER_279_699 ();
 b15zdnd11an1n64x5 FILLER_279_755 ();
 b15zdnd11an1n64x5 FILLER_279_819 ();
 b15zdnd11an1n64x5 FILLER_279_883 ();
 b15zdnd11an1n16x5 FILLER_279_947 ();
 b15zdnd11an1n08x5 FILLER_279_963 ();
 b15zdnd00an1n01x5 FILLER_279_971 ();
 b15zdnd11an1n32x5 FILLER_279_975 ();
 b15zdnd11an1n64x5 FILLER_279_1011 ();
 b15zdnd11an1n64x5 FILLER_279_1075 ();
 b15zdnd11an1n32x5 FILLER_279_1139 ();
 b15zdnd11an1n16x5 FILLER_279_1171 ();
 b15zdnd11an1n08x5 FILLER_279_1187 ();
 b15zdnd00an1n02x5 FILLER_279_1195 ();
 b15zdnd00an1n01x5 FILLER_279_1197 ();
 b15zdnd11an1n32x5 FILLER_279_1240 ();
 b15zdnd11an1n04x5 FILLER_279_1272 ();
 b15zdnd00an1n02x5 FILLER_279_1276 ();
 b15zdnd11an1n04x5 FILLER_279_1290 ();
 b15zdnd11an1n64x5 FILLER_279_1299 ();
 b15zdnd11an1n32x5 FILLER_279_1363 ();
 b15zdnd11an1n04x5 FILLER_279_1395 ();
 b15zdnd00an1n02x5 FILLER_279_1399 ();
 b15zdnd11an1n64x5 FILLER_279_1443 ();
 b15zdnd11an1n64x5 FILLER_279_1507 ();
 b15zdnd11an1n64x5 FILLER_279_1571 ();
 b15zdnd11an1n64x5 FILLER_279_1635 ();
 b15zdnd11an1n64x5 FILLER_279_1699 ();
 b15zdnd11an1n32x5 FILLER_279_1763 ();
 b15zdnd11an1n04x5 FILLER_279_1799 ();
 b15zdnd00an1n02x5 FILLER_279_1803 ();
 b15zdnd11an1n04x5 FILLER_279_1809 ();
 b15zdnd11an1n08x5 FILLER_279_1820 ();
 b15zdnd11an1n04x5 FILLER_279_1831 ();
 b15zdnd11an1n64x5 FILLER_279_1838 ();
 b15zdnd11an1n64x5 FILLER_279_1902 ();
 b15zdnd11an1n64x5 FILLER_279_1966 ();
 b15zdnd11an1n64x5 FILLER_279_2030 ();
 b15zdnd11an1n08x5 FILLER_279_2094 ();
 b15zdnd11an1n04x5 FILLER_279_2134 ();
 b15zdnd11an1n64x5 FILLER_279_2141 ();
 b15zdnd11an1n64x5 FILLER_279_2205 ();
 b15zdnd11an1n08x5 FILLER_279_2269 ();
 b15zdnd11an1n04x5 FILLER_279_2277 ();
 b15zdnd00an1n02x5 FILLER_279_2281 ();
 b15zdnd00an1n01x5 FILLER_279_2283 ();
 b15zdnd11an1n64x5 FILLER_280_8 ();
 b15zdnd11an1n64x5 FILLER_280_72 ();
 b15zdnd11an1n04x5 FILLER_280_136 ();
 b15zdnd00an1n01x5 FILLER_280_140 ();
 b15zdnd11an1n04x5 FILLER_280_157 ();
 b15zdnd11an1n04x5 FILLER_280_166 ();
 b15zdnd11an1n64x5 FILLER_280_176 ();
 b15zdnd11an1n64x5 FILLER_280_240 ();
 b15zdnd11an1n64x5 FILLER_280_304 ();
 b15zdnd11an1n64x5 FILLER_280_368 ();
 b15zdnd11an1n64x5 FILLER_280_432 ();
 b15zdnd00an1n02x5 FILLER_280_496 ();
 b15zdnd11an1n04x5 FILLER_280_501 ();
 b15zdnd11an1n32x5 FILLER_280_508 ();
 b15zdnd11an1n08x5 FILLER_280_540 ();
 b15zdnd11an1n04x5 FILLER_280_548 ();
 b15zdnd11an1n16x5 FILLER_280_559 ();
 b15zdnd11an1n08x5 FILLER_280_575 ();
 b15zdnd11an1n32x5 FILLER_280_622 ();
 b15zdnd11an1n16x5 FILLER_280_654 ();
 b15zdnd11an1n08x5 FILLER_280_670 ();
 b15zdnd00an1n02x5 FILLER_280_678 ();
 b15zdnd11an1n04x5 FILLER_280_695 ();
 b15zdnd11an1n04x5 FILLER_280_712 ();
 b15zdnd00an1n02x5 FILLER_280_716 ();
 b15zdnd00an1n02x5 FILLER_280_726 ();
 b15zdnd11an1n64x5 FILLER_280_770 ();
 b15zdnd11an1n32x5 FILLER_280_834 ();
 b15zdnd11an1n16x5 FILLER_280_866 ();
 b15zdnd11an1n08x5 FILLER_280_882 ();
 b15zdnd11an1n04x5 FILLER_280_893 ();
 b15zdnd11an1n32x5 FILLER_280_903 ();
 b15zdnd11an1n08x5 FILLER_280_935 ();
 b15zdnd00an1n02x5 FILLER_280_943 ();
 b15zdnd00an1n01x5 FILLER_280_945 ();
 b15zdnd11an1n64x5 FILLER_280_988 ();
 b15zdnd11an1n64x5 FILLER_280_1052 ();
 b15zdnd11an1n32x5 FILLER_280_1116 ();
 b15zdnd11an1n16x5 FILLER_280_1148 ();
 b15zdnd11an1n64x5 FILLER_280_1189 ();
 b15zdnd11an1n08x5 FILLER_280_1253 ();
 b15zdnd11an1n04x5 FILLER_280_1264 ();
 b15zdnd00an1n01x5 FILLER_280_1268 ();
 b15zdnd11an1n04x5 FILLER_280_1273 ();
 b15zdnd11an1n64x5 FILLER_280_1287 ();
 b15zdnd11an1n64x5 FILLER_280_1351 ();
 b15zdnd11an1n64x5 FILLER_280_1457 ();
 b15zdnd11an1n64x5 FILLER_280_1521 ();
 b15zdnd11an1n64x5 FILLER_280_1585 ();
 b15zdnd11an1n64x5 FILLER_280_1649 ();
 b15zdnd11an1n64x5 FILLER_280_1713 ();
 b15zdnd11an1n16x5 FILLER_280_1777 ();
 b15zdnd00an1n02x5 FILLER_280_1793 ();
 b15zdnd11an1n04x5 FILLER_280_1800 ();
 b15zdnd00an1n02x5 FILLER_280_1804 ();
 b15zdnd00an1n01x5 FILLER_280_1806 ();
 b15zdnd11an1n04x5 FILLER_280_1812 ();
 b15zdnd11an1n64x5 FILLER_280_1858 ();
 b15zdnd11an1n64x5 FILLER_280_1922 ();
 b15zdnd11an1n64x5 FILLER_280_1986 ();
 b15zdnd11an1n16x5 FILLER_280_2050 ();
 b15zdnd11an1n08x5 FILLER_280_2066 ();
 b15zdnd00an1n02x5 FILLER_280_2074 ();
 b15zdnd11an1n04x5 FILLER_280_2084 ();
 b15zdnd11an1n32x5 FILLER_280_2092 ();
 b15zdnd11an1n16x5 FILLER_280_2124 ();
 b15zdnd11an1n08x5 FILLER_280_2140 ();
 b15zdnd11an1n04x5 FILLER_280_2148 ();
 b15zdnd00an1n02x5 FILLER_280_2152 ();
 b15zdnd11an1n64x5 FILLER_280_2162 ();
 b15zdnd11an1n32x5 FILLER_280_2226 ();
 b15zdnd11an1n16x5 FILLER_280_2258 ();
 b15zdnd00an1n02x5 FILLER_280_2274 ();
 b15zdnd11an1n64x5 FILLER_281_0 ();
 b15zdnd11an1n64x5 FILLER_281_64 ();
 b15zdnd11an1n64x5 FILLER_281_128 ();
 b15zdnd11an1n64x5 FILLER_281_192 ();
 b15zdnd11an1n64x5 FILLER_281_256 ();
 b15zdnd11an1n64x5 FILLER_281_320 ();
 b15zdnd11an1n32x5 FILLER_281_384 ();
 b15zdnd11an1n16x5 FILLER_281_416 ();
 b15zdnd00an1n02x5 FILLER_281_432 ();
 b15zdnd11an1n64x5 FILLER_281_448 ();
 b15zdnd11an1n32x5 FILLER_281_512 ();
 b15zdnd11an1n16x5 FILLER_281_544 ();
 b15zdnd11an1n04x5 FILLER_281_560 ();
 b15zdnd00an1n01x5 FILLER_281_564 ();
 b15zdnd11an1n04x5 FILLER_281_607 ();
 b15zdnd11an1n64x5 FILLER_281_614 ();
 b15zdnd00an1n02x5 FILLER_281_678 ();
 b15zdnd00an1n01x5 FILLER_281_680 ();
 b15zdnd11an1n08x5 FILLER_281_687 ();
 b15zdnd00an1n01x5 FILLER_281_695 ();
 b15zdnd11an1n04x5 FILLER_281_705 ();
 b15zdnd11an1n04x5 FILLER_281_713 ();
 b15zdnd11an1n64x5 FILLER_281_759 ();
 b15zdnd11an1n32x5 FILLER_281_823 ();
 b15zdnd11an1n08x5 FILLER_281_855 ();
 b15zdnd11an1n04x5 FILLER_281_863 ();
 b15zdnd11an1n16x5 FILLER_281_919 ();
 b15zdnd11an1n08x5 FILLER_281_935 ();
 b15zdnd00an1n02x5 FILLER_281_943 ();
 b15zdnd11an1n04x5 FILLER_281_997 ();
 b15zdnd00an1n01x5 FILLER_281_1001 ();
 b15zdnd11an1n64x5 FILLER_281_1054 ();
 b15zdnd11an1n32x5 FILLER_281_1118 ();
 b15zdnd11an1n64x5 FILLER_281_1153 ();
 b15zdnd11an1n32x5 FILLER_281_1217 ();
 b15zdnd11an1n16x5 FILLER_281_1249 ();
 b15zdnd00an1n02x5 FILLER_281_1265 ();
 b15zdnd00an1n01x5 FILLER_281_1267 ();
 b15zdnd11an1n08x5 FILLER_281_1271 ();
 b15zdnd00an1n01x5 FILLER_281_1279 ();
 b15zdnd11an1n64x5 FILLER_281_1285 ();
 b15zdnd11an1n32x5 FILLER_281_1349 ();
 b15zdnd11an1n16x5 FILLER_281_1381 ();
 b15zdnd00an1n02x5 FILLER_281_1397 ();
 b15zdnd00an1n01x5 FILLER_281_1399 ();
 b15zdnd11an1n64x5 FILLER_281_1452 ();
 b15zdnd11an1n64x5 FILLER_281_1516 ();
 b15zdnd11an1n64x5 FILLER_281_1580 ();
 b15zdnd11an1n32x5 FILLER_281_1644 ();
 b15zdnd11an1n16x5 FILLER_281_1676 ();
 b15zdnd11an1n08x5 FILLER_281_1692 ();
 b15zdnd11an1n04x5 FILLER_281_1700 ();
 b15zdnd00an1n02x5 FILLER_281_1704 ();
 b15zdnd00an1n01x5 FILLER_281_1706 ();
 b15zdnd11an1n64x5 FILLER_281_1710 ();
 b15zdnd11an1n16x5 FILLER_281_1774 ();
 b15zdnd00an1n02x5 FILLER_281_1790 ();
 b15zdnd00an1n01x5 FILLER_281_1792 ();
 b15zdnd11an1n04x5 FILLER_281_1803 ();
 b15zdnd11an1n04x5 FILLER_281_1813 ();
 b15zdnd00an1n01x5 FILLER_281_1817 ();
 b15zdnd11an1n64x5 FILLER_281_1860 ();
 b15zdnd11an1n64x5 FILLER_281_1924 ();
 b15zdnd11an1n64x5 FILLER_281_1988 ();
 b15zdnd11an1n08x5 FILLER_281_2052 ();
 b15zdnd11an1n04x5 FILLER_281_2060 ();
 b15zdnd00an1n02x5 FILLER_281_2064 ();
 b15zdnd00an1n01x5 FILLER_281_2066 ();
 b15zdnd11an1n64x5 FILLER_281_2078 ();
 b15zdnd11an1n64x5 FILLER_281_2142 ();
 b15zdnd11an1n64x5 FILLER_281_2206 ();
 b15zdnd11an1n08x5 FILLER_281_2270 ();
 b15zdnd11an1n04x5 FILLER_281_2278 ();
 b15zdnd00an1n02x5 FILLER_281_2282 ();
 b15zdnd11an1n64x5 FILLER_282_8 ();
 b15zdnd11an1n64x5 FILLER_282_72 ();
 b15zdnd11an1n64x5 FILLER_282_136 ();
 b15zdnd11an1n64x5 FILLER_282_200 ();
 b15zdnd11an1n64x5 FILLER_282_264 ();
 b15zdnd11an1n64x5 FILLER_282_328 ();
 b15zdnd11an1n16x5 FILLER_282_392 ();
 b15zdnd11an1n08x5 FILLER_282_408 ();
 b15zdnd11an1n64x5 FILLER_282_424 ();
 b15zdnd11an1n64x5 FILLER_282_488 ();
 b15zdnd11an1n16x5 FILLER_282_552 ();
 b15zdnd11an1n04x5 FILLER_282_568 ();
 b15zdnd00an1n02x5 FILLER_282_572 ();
 b15zdnd00an1n01x5 FILLER_282_574 ();
 b15zdnd11an1n16x5 FILLER_282_627 ();
 b15zdnd11an1n08x5 FILLER_282_643 ();
 b15zdnd00an1n02x5 FILLER_282_651 ();
 b15zdnd00an1n01x5 FILLER_282_653 ();
 b15zdnd11an1n04x5 FILLER_282_696 ();
 b15zdnd11an1n04x5 FILLER_282_711 ();
 b15zdnd00an1n02x5 FILLER_282_715 ();
 b15zdnd00an1n01x5 FILLER_282_717 ();
 b15zdnd00an1n02x5 FILLER_282_726 ();
 b15zdnd11an1n64x5 FILLER_282_731 ();
 b15zdnd11an1n64x5 FILLER_282_795 ();
 b15zdnd11an1n16x5 FILLER_282_859 ();
 b15zdnd11an1n08x5 FILLER_282_875 ();
 b15zdnd11an1n04x5 FILLER_282_883 ();
 b15zdnd11an1n08x5 FILLER_282_890 ();
 b15zdnd11an1n32x5 FILLER_282_901 ();
 b15zdnd11an1n16x5 FILLER_282_933 ();
 b15zdnd11an1n08x5 FILLER_282_949 ();
 b15zdnd11an1n04x5 FILLER_282_957 ();
 b15zdnd00an1n02x5 FILLER_282_961 ();
 b15zdnd11an1n04x5 FILLER_282_966 ();
 b15zdnd11an1n32x5 FILLER_282_973 ();
 b15zdnd11an1n08x5 FILLER_282_1005 ();
 b15zdnd00an1n01x5 FILLER_282_1013 ();
 b15zdnd11an1n64x5 FILLER_282_1056 ();
 b15zdnd00an1n02x5 FILLER_282_1120 ();
 b15zdnd00an1n01x5 FILLER_282_1122 ();
 b15zdnd11an1n16x5 FILLER_282_1175 ();
 b15zdnd11an1n08x5 FILLER_282_1191 ();
 b15zdnd11an1n04x5 FILLER_282_1199 ();
 b15zdnd00an1n02x5 FILLER_282_1203 ();
 b15zdnd11an1n08x5 FILLER_282_1247 ();
 b15zdnd11an1n04x5 FILLER_282_1255 ();
 b15zdnd00an1n01x5 FILLER_282_1259 ();
 b15zdnd11an1n04x5 FILLER_282_1269 ();
 b15zdnd11an1n64x5 FILLER_282_1315 ();
 b15zdnd11an1n32x5 FILLER_282_1379 ();
 b15zdnd11an1n08x5 FILLER_282_1411 ();
 b15zdnd11an1n04x5 FILLER_282_1419 ();
 b15zdnd00an1n02x5 FILLER_282_1423 ();
 b15zdnd11an1n04x5 FILLER_282_1428 ();
 b15zdnd11an1n64x5 FILLER_282_1435 ();
 b15zdnd11an1n64x5 FILLER_282_1499 ();
 b15zdnd11an1n64x5 FILLER_282_1563 ();
 b15zdnd11an1n64x5 FILLER_282_1627 ();
 b15zdnd11an1n16x5 FILLER_282_1691 ();
 b15zdnd11an1n64x5 FILLER_282_1710 ();
 b15zdnd11an1n08x5 FILLER_282_1774 ();
 b15zdnd11an1n04x5 FILLER_282_1789 ();
 b15zdnd11an1n04x5 FILLER_282_1801 ();
 b15zdnd11an1n04x5 FILLER_282_1847 ();
 b15zdnd11an1n32x5 FILLER_282_1893 ();
 b15zdnd11an1n16x5 FILLER_282_1925 ();
 b15zdnd11an1n08x5 FILLER_282_1941 ();
 b15zdnd11an1n04x5 FILLER_282_1949 ();
 b15zdnd00an1n02x5 FILLER_282_1953 ();
 b15zdnd00an1n01x5 FILLER_282_1955 ();
 b15zdnd11an1n64x5 FILLER_282_2008 ();
 b15zdnd11an1n64x5 FILLER_282_2072 ();
 b15zdnd11an1n16x5 FILLER_282_2136 ();
 b15zdnd00an1n02x5 FILLER_282_2152 ();
 b15zdnd11an1n64x5 FILLER_282_2162 ();
 b15zdnd11an1n32x5 FILLER_282_2226 ();
 b15zdnd11an1n16x5 FILLER_282_2258 ();
 b15zdnd00an1n02x5 FILLER_282_2274 ();
 b15zdnd11an1n64x5 FILLER_283_0 ();
 b15zdnd11an1n64x5 FILLER_283_64 ();
 b15zdnd11an1n64x5 FILLER_283_128 ();
 b15zdnd11an1n64x5 FILLER_283_192 ();
 b15zdnd11an1n64x5 FILLER_283_256 ();
 b15zdnd11an1n64x5 FILLER_283_320 ();
 b15zdnd11an1n64x5 FILLER_283_384 ();
 b15zdnd11an1n32x5 FILLER_283_448 ();
 b15zdnd11an1n16x5 FILLER_283_480 ();
 b15zdnd11an1n08x5 FILLER_283_496 ();
 b15zdnd00an1n01x5 FILLER_283_504 ();
 b15zdnd11an1n32x5 FILLER_283_509 ();
 b15zdnd11an1n04x5 FILLER_283_541 ();
 b15zdnd11an1n04x5 FILLER_283_597 ();
 b15zdnd11an1n04x5 FILLER_283_604 ();
 b15zdnd11an1n64x5 FILLER_283_616 ();
 b15zdnd11an1n32x5 FILLER_283_680 ();
 b15zdnd11an1n04x5 FILLER_283_712 ();
 b15zdnd00an1n01x5 FILLER_283_716 ();
 b15zdnd11an1n64x5 FILLER_283_720 ();
 b15zdnd11an1n64x5 FILLER_283_784 ();
 b15zdnd11an1n64x5 FILLER_283_848 ();
 b15zdnd11an1n64x5 FILLER_283_912 ();
 b15zdnd11an1n32x5 FILLER_283_976 ();
 b15zdnd11an1n08x5 FILLER_283_1008 ();
 b15zdnd00an1n02x5 FILLER_283_1016 ();
 b15zdnd11an1n04x5 FILLER_283_1021 ();
 b15zdnd11an1n04x5 FILLER_283_1028 ();
 b15zdnd11an1n04x5 FILLER_283_1035 ();
 b15zdnd11an1n64x5 FILLER_283_1042 ();
 b15zdnd11an1n32x5 FILLER_283_1106 ();
 b15zdnd00an1n02x5 FILLER_283_1138 ();
 b15zdnd00an1n01x5 FILLER_283_1140 ();
 b15zdnd11an1n04x5 FILLER_283_1144 ();
 b15zdnd11an1n64x5 FILLER_283_1151 ();
 b15zdnd11an1n64x5 FILLER_283_1215 ();
 b15zdnd00an1n01x5 FILLER_283_1279 ();
 b15zdnd11an1n64x5 FILLER_283_1286 ();
 b15zdnd11an1n64x5 FILLER_283_1350 ();
 b15zdnd11an1n08x5 FILLER_283_1414 ();
 b15zdnd00an1n02x5 FILLER_283_1422 ();
 b15zdnd00an1n01x5 FILLER_283_1424 ();
 b15zdnd11an1n64x5 FILLER_283_1428 ();
 b15zdnd11an1n64x5 FILLER_283_1492 ();
 b15zdnd11an1n64x5 FILLER_283_1556 ();
 b15zdnd11an1n32x5 FILLER_283_1620 ();
 b15zdnd11an1n16x5 FILLER_283_1652 ();
 b15zdnd11an1n08x5 FILLER_283_1668 ();
 b15zdnd11an1n04x5 FILLER_283_1676 ();
 b15zdnd00an1n02x5 FILLER_283_1680 ();
 b15zdnd11an1n16x5 FILLER_283_1734 ();
 b15zdnd00an1n02x5 FILLER_283_1750 ();
 b15zdnd11an1n16x5 FILLER_283_1794 ();
 b15zdnd11an1n64x5 FILLER_283_1862 ();
 b15zdnd11an1n32x5 FILLER_283_1926 ();
 b15zdnd11an1n16x5 FILLER_283_1958 ();
 b15zdnd11an1n04x5 FILLER_283_1974 ();
 b15zdnd00an1n01x5 FILLER_283_1978 ();
 b15zdnd11an1n04x5 FILLER_283_1982 ();
 b15zdnd11an1n64x5 FILLER_283_1989 ();
 b15zdnd11an1n64x5 FILLER_283_2053 ();
 b15zdnd11an1n64x5 FILLER_283_2117 ();
 b15zdnd11an1n64x5 FILLER_283_2181 ();
 b15zdnd11an1n32x5 FILLER_283_2245 ();
 b15zdnd11an1n04x5 FILLER_283_2277 ();
 b15zdnd00an1n02x5 FILLER_283_2281 ();
 b15zdnd00an1n01x5 FILLER_283_2283 ();
 b15zdnd11an1n64x5 FILLER_284_8 ();
 b15zdnd11an1n64x5 FILLER_284_72 ();
 b15zdnd11an1n32x5 FILLER_284_136 ();
 b15zdnd00an1n02x5 FILLER_284_168 ();
 b15zdnd11an1n64x5 FILLER_284_212 ();
 b15zdnd11an1n64x5 FILLER_284_276 ();
 b15zdnd11an1n64x5 FILLER_284_340 ();
 b15zdnd11an1n64x5 FILLER_284_404 ();
 b15zdnd11an1n64x5 FILLER_284_468 ();
 b15zdnd11an1n32x5 FILLER_284_532 ();
 b15zdnd00an1n01x5 FILLER_284_564 ();
 b15zdnd11an1n04x5 FILLER_284_568 ();
 b15zdnd11an1n08x5 FILLER_284_575 ();
 b15zdnd11an1n04x5 FILLER_284_583 ();
 b15zdnd00an1n02x5 FILLER_284_587 ();
 b15zdnd00an1n01x5 FILLER_284_589 ();
 b15zdnd11an1n64x5 FILLER_284_593 ();
 b15zdnd11an1n32x5 FILLER_284_657 ();
 b15zdnd11an1n16x5 FILLER_284_689 ();
 b15zdnd11an1n08x5 FILLER_284_705 ();
 b15zdnd11an1n04x5 FILLER_284_713 ();
 b15zdnd00an1n01x5 FILLER_284_717 ();
 b15zdnd11an1n64x5 FILLER_284_726 ();
 b15zdnd11an1n64x5 FILLER_284_790 ();
 b15zdnd11an1n64x5 FILLER_284_854 ();
 b15zdnd11an1n64x5 FILLER_284_918 ();
 b15zdnd11an1n32x5 FILLER_284_982 ();
 b15zdnd11an1n08x5 FILLER_284_1014 ();
 b15zdnd11an1n04x5 FILLER_284_1022 ();
 b15zdnd00an1n01x5 FILLER_284_1026 ();
 b15zdnd11an1n64x5 FILLER_284_1030 ();
 b15zdnd11an1n64x5 FILLER_284_1094 ();
 b15zdnd11an1n64x5 FILLER_284_1158 ();
 b15zdnd11an1n64x5 FILLER_284_1222 ();
 b15zdnd11an1n64x5 FILLER_284_1286 ();
 b15zdnd11an1n64x5 FILLER_284_1350 ();
 b15zdnd11an1n64x5 FILLER_284_1414 ();
 b15zdnd11an1n64x5 FILLER_284_1478 ();
 b15zdnd11an1n64x5 FILLER_284_1542 ();
 b15zdnd11an1n64x5 FILLER_284_1606 ();
 b15zdnd11an1n32x5 FILLER_284_1670 ();
 b15zdnd11an1n04x5 FILLER_284_1702 ();
 b15zdnd00an1n02x5 FILLER_284_1706 ();
 b15zdnd11an1n64x5 FILLER_284_1711 ();
 b15zdnd11an1n32x5 FILLER_284_1775 ();
 b15zdnd11an1n16x5 FILLER_284_1807 ();
 b15zdnd11an1n04x5 FILLER_284_1823 ();
 b15zdnd11an1n64x5 FILLER_284_1869 ();
 b15zdnd11an1n32x5 FILLER_284_1933 ();
 b15zdnd11an1n16x5 FILLER_284_1965 ();
 b15zdnd11an1n64x5 FILLER_284_1984 ();
 b15zdnd11an1n64x5 FILLER_284_2048 ();
 b15zdnd11an1n32x5 FILLER_284_2112 ();
 b15zdnd11an1n08x5 FILLER_284_2144 ();
 b15zdnd00an1n02x5 FILLER_284_2152 ();
 b15zdnd11an1n64x5 FILLER_284_2162 ();
 b15zdnd11an1n32x5 FILLER_284_2226 ();
 b15zdnd11an1n16x5 FILLER_284_2258 ();
 b15zdnd00an1n02x5 FILLER_284_2274 ();
 b15zdnd11an1n64x5 FILLER_285_0 ();
 b15zdnd11an1n64x5 FILLER_285_64 ();
 b15zdnd11an1n32x5 FILLER_285_128 ();
 b15zdnd00an1n02x5 FILLER_285_160 ();
 b15zdnd00an1n01x5 FILLER_285_162 ();
 b15zdnd11an1n04x5 FILLER_285_166 ();
 b15zdnd11an1n04x5 FILLER_285_181 ();
 b15zdnd00an1n02x5 FILLER_285_185 ();
 b15zdnd11an1n04x5 FILLER_285_190 ();
 b15zdnd11an1n08x5 FILLER_285_197 ();
 b15zdnd11an1n04x5 FILLER_285_205 ();
 b15zdnd00an1n02x5 FILLER_285_209 ();
 b15zdnd11an1n64x5 FILLER_285_215 ();
 b15zdnd11an1n64x5 FILLER_285_279 ();
 b15zdnd11an1n64x5 FILLER_285_343 ();
 b15zdnd11an1n64x5 FILLER_285_407 ();
 b15zdnd11an1n64x5 FILLER_285_471 ();
 b15zdnd11an1n32x5 FILLER_285_535 ();
 b15zdnd11an1n04x5 FILLER_285_567 ();
 b15zdnd11an1n64x5 FILLER_285_574 ();
 b15zdnd11an1n64x5 FILLER_285_638 ();
 b15zdnd11an1n64x5 FILLER_285_702 ();
 b15zdnd11an1n64x5 FILLER_285_766 ();
 b15zdnd11an1n64x5 FILLER_285_830 ();
 b15zdnd11an1n64x5 FILLER_285_894 ();
 b15zdnd11an1n64x5 FILLER_285_958 ();
 b15zdnd11an1n64x5 FILLER_285_1022 ();
 b15zdnd11an1n64x5 FILLER_285_1086 ();
 b15zdnd11an1n64x5 FILLER_285_1150 ();
 b15zdnd11an1n64x5 FILLER_285_1214 ();
 b15zdnd11an1n64x5 FILLER_285_1278 ();
 b15zdnd11an1n64x5 FILLER_285_1342 ();
 b15zdnd11an1n64x5 FILLER_285_1406 ();
 b15zdnd11an1n64x5 FILLER_285_1470 ();
 b15zdnd11an1n64x5 FILLER_285_1534 ();
 b15zdnd11an1n64x5 FILLER_285_1598 ();
 b15zdnd11an1n64x5 FILLER_285_1662 ();
 b15zdnd11an1n64x5 FILLER_285_1726 ();
 b15zdnd11an1n32x5 FILLER_285_1790 ();
 b15zdnd11an1n08x5 FILLER_285_1822 ();
 b15zdnd11an1n04x5 FILLER_285_1830 ();
 b15zdnd00an1n01x5 FILLER_285_1834 ();
 b15zdnd11an1n64x5 FILLER_285_1838 ();
 b15zdnd11an1n64x5 FILLER_285_1902 ();
 b15zdnd11an1n64x5 FILLER_285_1966 ();
 b15zdnd11an1n64x5 FILLER_285_2030 ();
 b15zdnd11an1n64x5 FILLER_285_2094 ();
 b15zdnd11an1n64x5 FILLER_285_2158 ();
 b15zdnd11an1n32x5 FILLER_285_2222 ();
 b15zdnd11an1n16x5 FILLER_285_2254 ();
 b15zdnd11an1n08x5 FILLER_285_2270 ();
 b15zdnd11an1n04x5 FILLER_285_2278 ();
 b15zdnd00an1n02x5 FILLER_285_2282 ();
 b15zdnd11an1n64x5 FILLER_286_8 ();
 b15zdnd11an1n64x5 FILLER_286_72 ();
 b15zdnd11an1n32x5 FILLER_286_136 ();
 b15zdnd00an1n02x5 FILLER_286_168 ();
 b15zdnd00an1n01x5 FILLER_286_170 ();
 b15zdnd11an1n08x5 FILLER_286_176 ();
 b15zdnd00an1n02x5 FILLER_286_184 ();
 b15zdnd11an1n64x5 FILLER_286_228 ();
 b15zdnd11an1n64x5 FILLER_286_292 ();
 b15zdnd11an1n08x5 FILLER_286_356 ();
 b15zdnd11an1n04x5 FILLER_286_364 ();
 b15zdnd00an1n02x5 FILLER_286_368 ();
 b15zdnd11an1n64x5 FILLER_286_395 ();
 b15zdnd11an1n16x5 FILLER_286_459 ();
 b15zdnd11an1n08x5 FILLER_286_475 ();
 b15zdnd11an1n04x5 FILLER_286_483 ();
 b15zdnd11an1n64x5 FILLER_286_529 ();
 b15zdnd11an1n64x5 FILLER_286_593 ();
 b15zdnd11an1n32x5 FILLER_286_657 ();
 b15zdnd11an1n16x5 FILLER_286_689 ();
 b15zdnd11an1n08x5 FILLER_286_705 ();
 b15zdnd11an1n04x5 FILLER_286_713 ();
 b15zdnd00an1n01x5 FILLER_286_717 ();
 b15zdnd11an1n64x5 FILLER_286_726 ();
 b15zdnd11an1n32x5 FILLER_286_790 ();
 b15zdnd11an1n08x5 FILLER_286_822 ();
 b15zdnd11an1n04x5 FILLER_286_830 ();
 b15zdnd11an1n64x5 FILLER_286_837 ();
 b15zdnd11an1n64x5 FILLER_286_901 ();
 b15zdnd11an1n64x5 FILLER_286_965 ();
 b15zdnd11an1n64x5 FILLER_286_1029 ();
 b15zdnd11an1n64x5 FILLER_286_1093 ();
 b15zdnd11an1n64x5 FILLER_286_1157 ();
 b15zdnd11an1n64x5 FILLER_286_1221 ();
 b15zdnd11an1n64x5 FILLER_286_1285 ();
 b15zdnd11an1n64x5 FILLER_286_1349 ();
 b15zdnd11an1n64x5 FILLER_286_1413 ();
 b15zdnd11an1n64x5 FILLER_286_1477 ();
 b15zdnd11an1n64x5 FILLER_286_1541 ();
 b15zdnd11an1n64x5 FILLER_286_1605 ();
 b15zdnd11an1n64x5 FILLER_286_1669 ();
 b15zdnd11an1n64x5 FILLER_286_1733 ();
 b15zdnd11an1n64x5 FILLER_286_1797 ();
 b15zdnd11an1n32x5 FILLER_286_1861 ();
 b15zdnd11an1n16x5 FILLER_286_1893 ();
 b15zdnd11an1n04x5 FILLER_286_1909 ();
 b15zdnd00an1n02x5 FILLER_286_1913 ();
 b15zdnd11an1n04x5 FILLER_286_1918 ();
 b15zdnd11an1n64x5 FILLER_286_1925 ();
 b15zdnd11an1n64x5 FILLER_286_1989 ();
 b15zdnd11an1n64x5 FILLER_286_2053 ();
 b15zdnd11an1n32x5 FILLER_286_2117 ();
 b15zdnd11an1n04x5 FILLER_286_2149 ();
 b15zdnd00an1n01x5 FILLER_286_2153 ();
 b15zdnd11an1n64x5 FILLER_286_2162 ();
 b15zdnd11an1n32x5 FILLER_286_2226 ();
 b15zdnd11an1n16x5 FILLER_286_2258 ();
 b15zdnd00an1n02x5 FILLER_286_2274 ();
 b15zdnd11an1n64x5 FILLER_287_0 ();
 b15zdnd11an1n64x5 FILLER_287_64 ();
 b15zdnd11an1n32x5 FILLER_287_128 ();
 b15zdnd11an1n04x5 FILLER_287_160 ();
 b15zdnd00an1n02x5 FILLER_287_164 ();
 b15zdnd00an1n01x5 FILLER_287_166 ();
 b15zdnd11an1n04x5 FILLER_287_219 ();
 b15zdnd11an1n64x5 FILLER_287_265 ();
 b15zdnd11an1n64x5 FILLER_287_329 ();
 b15zdnd11an1n64x5 FILLER_287_393 ();
 b15zdnd11an1n64x5 FILLER_287_457 ();
 b15zdnd11an1n64x5 FILLER_287_521 ();
 b15zdnd11an1n64x5 FILLER_287_585 ();
 b15zdnd11an1n64x5 FILLER_287_649 ();
 b15zdnd11an1n64x5 FILLER_287_713 ();
 b15zdnd11an1n16x5 FILLER_287_777 ();
 b15zdnd11an1n08x5 FILLER_287_793 ();
 b15zdnd11an1n04x5 FILLER_287_801 ();
 b15zdnd00an1n02x5 FILLER_287_805 ();
 b15zdnd11an1n04x5 FILLER_287_859 ();
 b15zdnd11an1n64x5 FILLER_287_881 ();
 b15zdnd11an1n64x5 FILLER_287_945 ();
 b15zdnd11an1n64x5 FILLER_287_1009 ();
 b15zdnd11an1n64x5 FILLER_287_1073 ();
 b15zdnd11an1n64x5 FILLER_287_1137 ();
 b15zdnd11an1n64x5 FILLER_287_1201 ();
 b15zdnd11an1n64x5 FILLER_287_1265 ();
 b15zdnd11an1n64x5 FILLER_287_1329 ();
 b15zdnd11an1n64x5 FILLER_287_1393 ();
 b15zdnd11an1n64x5 FILLER_287_1457 ();
 b15zdnd11an1n64x5 FILLER_287_1521 ();
 b15zdnd11an1n08x5 FILLER_287_1585 ();
 b15zdnd00an1n02x5 FILLER_287_1593 ();
 b15zdnd00an1n01x5 FILLER_287_1595 ();
 b15zdnd11an1n08x5 FILLER_287_1636 ();
 b15zdnd00an1n02x5 FILLER_287_1644 ();
 b15zdnd11an1n04x5 FILLER_287_1649 ();
 b15zdnd11an1n64x5 FILLER_287_1656 ();
 b15zdnd11an1n64x5 FILLER_287_1720 ();
 b15zdnd11an1n64x5 FILLER_287_1784 ();
 b15zdnd11an1n32x5 FILLER_287_1848 ();
 b15zdnd11an1n16x5 FILLER_287_1880 ();
 b15zdnd00an1n01x5 FILLER_287_1896 ();
 b15zdnd11an1n64x5 FILLER_287_1949 ();
 b15zdnd11an1n64x5 FILLER_287_2013 ();
 b15zdnd11an1n64x5 FILLER_287_2077 ();
 b15zdnd11an1n64x5 FILLER_287_2141 ();
 b15zdnd11an1n64x5 FILLER_287_2205 ();
 b15zdnd11an1n08x5 FILLER_287_2269 ();
 b15zdnd11an1n04x5 FILLER_287_2277 ();
 b15zdnd00an1n02x5 FILLER_287_2281 ();
 b15zdnd00an1n01x5 FILLER_287_2283 ();
 b15zdnd11an1n64x5 FILLER_288_8 ();
 b15zdnd11an1n64x5 FILLER_288_72 ();
 b15zdnd11an1n32x5 FILLER_288_136 ();
 b15zdnd11an1n16x5 FILLER_288_168 ();
 b15zdnd11an1n08x5 FILLER_288_184 ();
 b15zdnd00an1n02x5 FILLER_288_192 ();
 b15zdnd00an1n01x5 FILLER_288_194 ();
 b15zdnd11an1n08x5 FILLER_288_198 ();
 b15zdnd11an1n04x5 FILLER_288_206 ();
 b15zdnd11an1n32x5 FILLER_288_214 ();
 b15zdnd11an1n16x5 FILLER_288_246 ();
 b15zdnd11an1n04x5 FILLER_288_262 ();
 b15zdnd00an1n02x5 FILLER_288_266 ();
 b15zdnd11an1n04x5 FILLER_288_308 ();
 b15zdnd11an1n64x5 FILLER_288_315 ();
 b15zdnd11an1n64x5 FILLER_288_421 ();
 b15zdnd11an1n64x5 FILLER_288_485 ();
 b15zdnd11an1n64x5 FILLER_288_549 ();
 b15zdnd11an1n64x5 FILLER_288_613 ();
 b15zdnd11an1n32x5 FILLER_288_677 ();
 b15zdnd11an1n08x5 FILLER_288_709 ();
 b15zdnd00an1n01x5 FILLER_288_717 ();
 b15zdnd11an1n64x5 FILLER_288_726 ();
 b15zdnd11an1n32x5 FILLER_288_790 ();
 b15zdnd00an1n02x5 FILLER_288_822 ();
 b15zdnd00an1n01x5 FILLER_288_824 ();
 b15zdnd11an1n04x5 FILLER_288_828 ();
 b15zdnd11an1n16x5 FILLER_288_835 ();
 b15zdnd11an1n08x5 FILLER_288_851 ();
 b15zdnd00an1n02x5 FILLER_288_859 ();
 b15zdnd11an1n64x5 FILLER_288_903 ();
 b15zdnd11an1n64x5 FILLER_288_967 ();
 b15zdnd11an1n64x5 FILLER_288_1031 ();
 b15zdnd11an1n64x5 FILLER_288_1095 ();
 b15zdnd11an1n64x5 FILLER_288_1159 ();
 b15zdnd11an1n64x5 FILLER_288_1223 ();
 b15zdnd11an1n08x5 FILLER_288_1287 ();
 b15zdnd11an1n04x5 FILLER_288_1295 ();
 b15zdnd00an1n01x5 FILLER_288_1299 ();
 b15zdnd11an1n64x5 FILLER_288_1342 ();
 b15zdnd11an1n64x5 FILLER_288_1406 ();
 b15zdnd11an1n08x5 FILLER_288_1470 ();
 b15zdnd11an1n64x5 FILLER_288_1520 ();
 b15zdnd11an1n16x5 FILLER_288_1584 ();
 b15zdnd11an1n08x5 FILLER_288_1600 ();
 b15zdnd11an1n04x5 FILLER_288_1608 ();
 b15zdnd00an1n02x5 FILLER_288_1612 ();
 b15zdnd00an1n01x5 FILLER_288_1614 ();
 b15zdnd11an1n64x5 FILLER_288_1655 ();
 b15zdnd11an1n64x5 FILLER_288_1719 ();
 b15zdnd11an1n64x5 FILLER_288_1783 ();
 b15zdnd11an1n32x5 FILLER_288_1847 ();
 b15zdnd11an1n16x5 FILLER_288_1879 ();
 b15zdnd11an1n08x5 FILLER_288_1895 ();
 b15zdnd00an1n02x5 FILLER_288_1903 ();
 b15zdnd00an1n01x5 FILLER_288_1905 ();
 b15zdnd11an1n64x5 FILLER_288_1948 ();
 b15zdnd11an1n64x5 FILLER_288_2012 ();
 b15zdnd11an1n64x5 FILLER_288_2076 ();
 b15zdnd11an1n08x5 FILLER_288_2140 ();
 b15zdnd11an1n04x5 FILLER_288_2148 ();
 b15zdnd00an1n02x5 FILLER_288_2152 ();
 b15zdnd11an1n64x5 FILLER_288_2162 ();
 b15zdnd11an1n32x5 FILLER_288_2226 ();
 b15zdnd11an1n16x5 FILLER_288_2258 ();
 b15zdnd00an1n02x5 FILLER_288_2274 ();
 b15zdnd11an1n64x5 FILLER_289_0 ();
 b15zdnd11an1n64x5 FILLER_289_64 ();
 b15zdnd11an1n64x5 FILLER_289_128 ();
 b15zdnd11an1n64x5 FILLER_289_192 ();
 b15zdnd11an1n32x5 FILLER_289_256 ();
 b15zdnd11an1n08x5 FILLER_289_288 ();
 b15zdnd11an1n04x5 FILLER_289_296 ();
 b15zdnd11an1n64x5 FILLER_289_303 ();
 b15zdnd11an1n32x5 FILLER_289_367 ();
 b15zdnd11an1n08x5 FILLER_289_399 ();
 b15zdnd11an1n64x5 FILLER_289_459 ();
 b15zdnd11an1n64x5 FILLER_289_523 ();
 b15zdnd11an1n64x5 FILLER_289_587 ();
 b15zdnd11an1n64x5 FILLER_289_651 ();
 b15zdnd11an1n64x5 FILLER_289_715 ();
 b15zdnd11an1n64x5 FILLER_289_779 ();
 b15zdnd11an1n64x5 FILLER_289_843 ();
 b15zdnd11an1n64x5 FILLER_289_907 ();
 b15zdnd11an1n64x5 FILLER_289_971 ();
 b15zdnd11an1n64x5 FILLER_289_1035 ();
 b15zdnd11an1n64x5 FILLER_289_1099 ();
 b15zdnd11an1n64x5 FILLER_289_1163 ();
 b15zdnd11an1n64x5 FILLER_289_1227 ();
 b15zdnd11an1n08x5 FILLER_289_1291 ();
 b15zdnd00an1n01x5 FILLER_289_1299 ();
 b15zdnd11an1n64x5 FILLER_289_1342 ();
 b15zdnd11an1n64x5 FILLER_289_1406 ();
 b15zdnd11an1n64x5 FILLER_289_1470 ();
 b15zdnd11an1n64x5 FILLER_289_1534 ();
 b15zdnd11an1n32x5 FILLER_289_1598 ();
 b15zdnd00an1n02x5 FILLER_289_1630 ();
 b15zdnd11an1n04x5 FILLER_289_1635 ();
 b15zdnd11an1n64x5 FILLER_289_1642 ();
 b15zdnd11an1n64x5 FILLER_289_1706 ();
 b15zdnd11an1n64x5 FILLER_289_1770 ();
 b15zdnd11an1n64x5 FILLER_289_1834 ();
 b15zdnd11an1n08x5 FILLER_289_1898 ();
 b15zdnd11an1n04x5 FILLER_289_1906 ();
 b15zdnd00an1n01x5 FILLER_289_1910 ();
 b15zdnd11an1n04x5 FILLER_289_1917 ();
 b15zdnd00an1n02x5 FILLER_289_1921 ();
 b15zdnd11an1n64x5 FILLER_289_1926 ();
 b15zdnd11an1n64x5 FILLER_289_1990 ();
 b15zdnd11an1n64x5 FILLER_289_2054 ();
 b15zdnd11an1n64x5 FILLER_289_2118 ();
 b15zdnd11an1n64x5 FILLER_289_2182 ();
 b15zdnd11an1n32x5 FILLER_289_2246 ();
 b15zdnd11an1n04x5 FILLER_289_2278 ();
 b15zdnd00an1n02x5 FILLER_289_2282 ();
 b15zdnd11an1n64x5 FILLER_290_8 ();
 b15zdnd11an1n64x5 FILLER_290_72 ();
 b15zdnd11an1n64x5 FILLER_290_136 ();
 b15zdnd11an1n64x5 FILLER_290_200 ();
 b15zdnd11an1n64x5 FILLER_290_264 ();
 b15zdnd11an1n64x5 FILLER_290_328 ();
 b15zdnd11an1n16x5 FILLER_290_392 ();
 b15zdnd00an1n01x5 FILLER_290_408 ();
 b15zdnd11an1n04x5 FILLER_290_412 ();
 b15zdnd11an1n04x5 FILLER_290_419 ();
 b15zdnd11an1n04x5 FILLER_290_426 ();
 b15zdnd11an1n04x5 FILLER_290_433 ();
 b15zdnd11an1n04x5 FILLER_290_440 ();
 b15zdnd11an1n64x5 FILLER_290_447 ();
 b15zdnd11an1n64x5 FILLER_290_511 ();
 b15zdnd11an1n64x5 FILLER_290_575 ();
 b15zdnd11an1n64x5 FILLER_290_639 ();
 b15zdnd11an1n08x5 FILLER_290_703 ();
 b15zdnd11an1n04x5 FILLER_290_711 ();
 b15zdnd00an1n02x5 FILLER_290_715 ();
 b15zdnd00an1n01x5 FILLER_290_717 ();
 b15zdnd11an1n64x5 FILLER_290_726 ();
 b15zdnd11an1n64x5 FILLER_290_790 ();
 b15zdnd11an1n64x5 FILLER_290_854 ();
 b15zdnd11an1n64x5 FILLER_290_918 ();
 b15zdnd11an1n64x5 FILLER_290_982 ();
 b15zdnd11an1n64x5 FILLER_290_1046 ();
 b15zdnd11an1n64x5 FILLER_290_1110 ();
 b15zdnd11an1n64x5 FILLER_290_1174 ();
 b15zdnd11an1n64x5 FILLER_290_1238 ();
 b15zdnd11an1n64x5 FILLER_290_1302 ();
 b15zdnd11an1n64x5 FILLER_290_1366 ();
 b15zdnd11an1n64x5 FILLER_290_1430 ();
 b15zdnd11an1n64x5 FILLER_290_1494 ();
 b15zdnd11an1n64x5 FILLER_290_1558 ();
 b15zdnd11an1n64x5 FILLER_290_1622 ();
 b15zdnd11an1n64x5 FILLER_290_1686 ();
 b15zdnd11an1n64x5 FILLER_290_1750 ();
 b15zdnd11an1n64x5 FILLER_290_1814 ();
 b15zdnd11an1n64x5 FILLER_290_1878 ();
 b15zdnd11an1n64x5 FILLER_290_1942 ();
 b15zdnd11an1n64x5 FILLER_290_2006 ();
 b15zdnd11an1n64x5 FILLER_290_2070 ();
 b15zdnd11an1n16x5 FILLER_290_2134 ();
 b15zdnd11an1n04x5 FILLER_290_2150 ();
 b15zdnd11an1n32x5 FILLER_290_2162 ();
 b15zdnd11an1n08x5 FILLER_290_2194 ();
 b15zdnd11an1n04x5 FILLER_290_2202 ();
 b15zdnd00an1n02x5 FILLER_290_2206 ();
 b15zdnd00an1n01x5 FILLER_290_2208 ();
 b15zdnd11an1n64x5 FILLER_290_2212 ();
 b15zdnd11an1n64x5 FILLER_291_0 ();
 b15zdnd11an1n64x5 FILLER_291_64 ();
 b15zdnd11an1n64x5 FILLER_291_128 ();
 b15zdnd11an1n64x5 FILLER_291_192 ();
 b15zdnd11an1n64x5 FILLER_291_256 ();
 b15zdnd11an1n64x5 FILLER_291_320 ();
 b15zdnd11an1n04x5 FILLER_291_436 ();
 b15zdnd11an1n64x5 FILLER_291_482 ();
 b15zdnd11an1n64x5 FILLER_291_546 ();
 b15zdnd11an1n64x5 FILLER_291_610 ();
 b15zdnd11an1n64x5 FILLER_291_674 ();
 b15zdnd11an1n64x5 FILLER_291_738 ();
 b15zdnd11an1n64x5 FILLER_291_802 ();
 b15zdnd11an1n32x5 FILLER_291_866 ();
 b15zdnd11an1n08x5 FILLER_291_898 ();
 b15zdnd11an1n64x5 FILLER_291_948 ();
 b15zdnd11an1n64x5 FILLER_291_1012 ();
 b15zdnd11an1n64x5 FILLER_291_1076 ();
 b15zdnd11an1n64x5 FILLER_291_1140 ();
 b15zdnd11an1n64x5 FILLER_291_1204 ();
 b15zdnd11an1n64x5 FILLER_291_1268 ();
 b15zdnd11an1n64x5 FILLER_291_1332 ();
 b15zdnd11an1n64x5 FILLER_291_1396 ();
 b15zdnd11an1n64x5 FILLER_291_1460 ();
 b15zdnd11an1n64x5 FILLER_291_1524 ();
 b15zdnd11an1n64x5 FILLER_291_1588 ();
 b15zdnd11an1n64x5 FILLER_291_1652 ();
 b15zdnd11an1n64x5 FILLER_291_1716 ();
 b15zdnd11an1n64x5 FILLER_291_1780 ();
 b15zdnd11an1n64x5 FILLER_291_1844 ();
 b15zdnd11an1n64x5 FILLER_291_1908 ();
 b15zdnd11an1n64x5 FILLER_291_1972 ();
 b15zdnd11an1n64x5 FILLER_291_2036 ();
 b15zdnd11an1n64x5 FILLER_291_2100 ();
 b15zdnd11an1n32x5 FILLER_291_2164 ();
 b15zdnd11an1n04x5 FILLER_291_2196 ();
 b15zdnd00an1n02x5 FILLER_291_2200 ();
 b15zdnd11an1n08x5 FILLER_291_2205 ();
 b15zdnd00an1n02x5 FILLER_291_2213 ();
 b15zdnd11an1n32x5 FILLER_291_2240 ();
 b15zdnd11an1n08x5 FILLER_291_2272 ();
 b15zdnd11an1n04x5 FILLER_291_2280 ();
 b15zdnd11an1n16x5 FILLER_292_8 ();
 b15zdnd11an1n04x5 FILLER_292_24 ();
 b15zdnd00an1n02x5 FILLER_292_28 ();
 b15zdnd00an1n01x5 FILLER_292_30 ();
 b15zdnd11an1n64x5 FILLER_292_36 ();
 b15zdnd11an1n64x5 FILLER_292_100 ();
 b15zdnd11an1n64x5 FILLER_292_164 ();
 b15zdnd11an1n64x5 FILLER_292_228 ();
 b15zdnd11an1n16x5 FILLER_292_292 ();
 b15zdnd00an1n01x5 FILLER_292_308 ();
 b15zdnd11an1n04x5 FILLER_292_312 ();
 b15zdnd11an1n64x5 FILLER_292_319 ();
 b15zdnd11an1n16x5 FILLER_292_383 ();
 b15zdnd11an1n04x5 FILLER_292_399 ();
 b15zdnd00an1n01x5 FILLER_292_403 ();
 b15zdnd11an1n04x5 FILLER_292_407 ();
 b15zdnd11an1n64x5 FILLER_292_414 ();
 b15zdnd11an1n64x5 FILLER_292_478 ();
 b15zdnd11an1n64x5 FILLER_292_542 ();
 b15zdnd11an1n64x5 FILLER_292_606 ();
 b15zdnd11an1n32x5 FILLER_292_670 ();
 b15zdnd11an1n16x5 FILLER_292_702 ();
 b15zdnd11an1n64x5 FILLER_292_726 ();
 b15zdnd11an1n64x5 FILLER_292_790 ();
 b15zdnd11an1n64x5 FILLER_292_854 ();
 b15zdnd11an1n64x5 FILLER_292_918 ();
 b15zdnd11an1n64x5 FILLER_292_982 ();
 b15zdnd11an1n64x5 FILLER_292_1046 ();
 b15zdnd11an1n64x5 FILLER_292_1110 ();
 b15zdnd11an1n64x5 FILLER_292_1174 ();
 b15zdnd11an1n64x5 FILLER_292_1238 ();
 b15zdnd11an1n64x5 FILLER_292_1302 ();
 b15zdnd11an1n64x5 FILLER_292_1366 ();
 b15zdnd11an1n64x5 FILLER_292_1430 ();
 b15zdnd11an1n64x5 FILLER_292_1494 ();
 b15zdnd11an1n64x5 FILLER_292_1558 ();
 b15zdnd11an1n64x5 FILLER_292_1622 ();
 b15zdnd11an1n64x5 FILLER_292_1686 ();
 b15zdnd11an1n64x5 FILLER_292_1750 ();
 b15zdnd11an1n64x5 FILLER_292_1814 ();
 b15zdnd11an1n64x5 FILLER_292_1878 ();
 b15zdnd11an1n64x5 FILLER_292_1942 ();
 b15zdnd11an1n64x5 FILLER_292_2006 ();
 b15zdnd11an1n64x5 FILLER_292_2070 ();
 b15zdnd11an1n16x5 FILLER_292_2134 ();
 b15zdnd11an1n04x5 FILLER_292_2150 ();
 b15zdnd11an1n08x5 FILLER_292_2162 ();
 b15zdnd11an1n04x5 FILLER_292_2170 ();
 b15zdnd00an1n02x5 FILLER_292_2174 ();
 b15zdnd00an1n01x5 FILLER_292_2176 ();
 b15zdnd11an1n32x5 FILLER_292_2229 ();
 b15zdnd11an1n08x5 FILLER_292_2261 ();
 b15zdnd11an1n04x5 FILLER_292_2269 ();
 b15zdnd00an1n02x5 FILLER_292_2273 ();
 b15zdnd00an1n01x5 FILLER_292_2275 ();
 b15zdnd11an1n16x5 FILLER_293_0 ();
 b15zdnd00an1n02x5 FILLER_293_16 ();
 b15zdnd11an1n64x5 FILLER_293_23 ();
 b15zdnd11an1n64x5 FILLER_293_87 ();
 b15zdnd11an1n64x5 FILLER_293_151 ();
 b15zdnd11an1n64x5 FILLER_293_215 ();
 b15zdnd11an1n04x5 FILLER_293_279 ();
 b15zdnd00an1n02x5 FILLER_293_283 ();
 b15zdnd00an1n01x5 FILLER_293_285 ();
 b15zdnd11an1n64x5 FILLER_293_338 ();
 b15zdnd11an1n64x5 FILLER_293_402 ();
 b15zdnd11an1n64x5 FILLER_293_466 ();
 b15zdnd11an1n64x5 FILLER_293_530 ();
 b15zdnd11an1n64x5 FILLER_293_594 ();
 b15zdnd11an1n64x5 FILLER_293_658 ();
 b15zdnd11an1n64x5 FILLER_293_722 ();
 b15zdnd11an1n64x5 FILLER_293_786 ();
 b15zdnd11an1n32x5 FILLER_293_850 ();
 b15zdnd11an1n16x5 FILLER_293_882 ();
 b15zdnd11an1n08x5 FILLER_293_898 ();
 b15zdnd00an1n02x5 FILLER_293_906 ();
 b15zdnd11an1n64x5 FILLER_293_950 ();
 b15zdnd11an1n64x5 FILLER_293_1014 ();
 b15zdnd11an1n64x5 FILLER_293_1078 ();
 b15zdnd11an1n64x5 FILLER_293_1142 ();
 b15zdnd11an1n64x5 FILLER_293_1206 ();
 b15zdnd11an1n32x5 FILLER_293_1270 ();
 b15zdnd11an1n16x5 FILLER_293_1302 ();
 b15zdnd00an1n02x5 FILLER_293_1318 ();
 b15zdnd00an1n01x5 FILLER_293_1320 ();
 b15zdnd11an1n64x5 FILLER_293_1332 ();
 b15zdnd11an1n64x5 FILLER_293_1396 ();
 b15zdnd11an1n64x5 FILLER_293_1460 ();
 b15zdnd11an1n64x5 FILLER_293_1524 ();
 b15zdnd11an1n64x5 FILLER_293_1588 ();
 b15zdnd11an1n32x5 FILLER_293_1652 ();
 b15zdnd11an1n64x5 FILLER_293_1726 ();
 b15zdnd11an1n64x5 FILLER_293_1790 ();
 b15zdnd11an1n64x5 FILLER_293_1854 ();
 b15zdnd11an1n64x5 FILLER_293_1918 ();
 b15zdnd11an1n64x5 FILLER_293_1982 ();
 b15zdnd11an1n16x5 FILLER_293_2046 ();
 b15zdnd11an1n08x5 FILLER_293_2062 ();
 b15zdnd00an1n02x5 FILLER_293_2070 ();
 b15zdnd00an1n01x5 FILLER_293_2072 ();
 b15zdnd11an1n64x5 FILLER_293_2115 ();
 b15zdnd11an1n16x5 FILLER_293_2179 ();
 b15zdnd11an1n04x5 FILLER_293_2195 ();
 b15zdnd00an1n02x5 FILLER_293_2199 ();
 b15zdnd00an1n01x5 FILLER_293_2201 ();
 b15zdnd11an1n04x5 FILLER_293_2207 ();
 b15zdnd11an1n08x5 FILLER_293_2214 ();
 b15zdnd11an1n16x5 FILLER_293_2264 ();
 b15zdnd11an1n04x5 FILLER_293_2280 ();
 b15zdnd11an1n16x5 FILLER_294_8 ();
 b15zdnd11an1n08x5 FILLER_294_24 ();
 b15zdnd11an1n04x5 FILLER_294_32 ();
 b15zdnd00an1n02x5 FILLER_294_36 ();
 b15zdnd11an1n64x5 FILLER_294_43 ();
 b15zdnd11an1n64x5 FILLER_294_107 ();
 b15zdnd11an1n64x5 FILLER_294_171 ();
 b15zdnd11an1n64x5 FILLER_294_235 ();
 b15zdnd11an1n04x5 FILLER_294_299 ();
 b15zdnd00an1n02x5 FILLER_294_303 ();
 b15zdnd00an1n01x5 FILLER_294_305 ();
 b15zdnd11an1n04x5 FILLER_294_309 ();
 b15zdnd11an1n64x5 FILLER_294_316 ();
 b15zdnd11an1n64x5 FILLER_294_380 ();
 b15zdnd11an1n64x5 FILLER_294_444 ();
 b15zdnd11an1n64x5 FILLER_294_508 ();
 b15zdnd11an1n64x5 FILLER_294_572 ();
 b15zdnd11an1n64x5 FILLER_294_636 ();
 b15zdnd11an1n16x5 FILLER_294_700 ();
 b15zdnd00an1n02x5 FILLER_294_716 ();
 b15zdnd11an1n64x5 FILLER_294_726 ();
 b15zdnd11an1n64x5 FILLER_294_790 ();
 b15zdnd11an1n64x5 FILLER_294_854 ();
 b15zdnd11an1n64x5 FILLER_294_918 ();
 b15zdnd11an1n64x5 FILLER_294_982 ();
 b15zdnd11an1n64x5 FILLER_294_1046 ();
 b15zdnd11an1n64x5 FILLER_294_1110 ();
 b15zdnd11an1n64x5 FILLER_294_1174 ();
 b15zdnd11an1n32x5 FILLER_294_1238 ();
 b15zdnd11an1n16x5 FILLER_294_1270 ();
 b15zdnd11an1n04x5 FILLER_294_1286 ();
 b15zdnd11an1n16x5 FILLER_294_1293 ();
 b15zdnd00an1n01x5 FILLER_294_1309 ();
 b15zdnd11an1n64x5 FILLER_294_1320 ();
 b15zdnd11an1n64x5 FILLER_294_1384 ();
 b15zdnd11an1n32x5 FILLER_294_1448 ();
 b15zdnd11an1n16x5 FILLER_294_1480 ();
 b15zdnd11an1n04x5 FILLER_294_1496 ();
 b15zdnd00an1n02x5 FILLER_294_1500 ();
 b15zdnd11an1n04x5 FILLER_294_1509 ();
 b15zdnd11an1n04x5 FILLER_294_1518 ();
 b15zdnd11an1n64x5 FILLER_294_1526 ();
 b15zdnd11an1n64x5 FILLER_294_1590 ();
 b15zdnd11an1n64x5 FILLER_294_1654 ();
 b15zdnd11an1n64x5 FILLER_294_1718 ();
 b15zdnd11an1n64x5 FILLER_294_1782 ();
 b15zdnd11an1n64x5 FILLER_294_1846 ();
 b15zdnd11an1n64x5 FILLER_294_1910 ();
 b15zdnd11an1n64x5 FILLER_294_1974 ();
 b15zdnd11an1n64x5 FILLER_294_2038 ();
 b15zdnd11an1n32x5 FILLER_294_2102 ();
 b15zdnd11an1n16x5 FILLER_294_2134 ();
 b15zdnd11an1n04x5 FILLER_294_2150 ();
 b15zdnd11an1n16x5 FILLER_294_2162 ();
 b15zdnd11an1n08x5 FILLER_294_2178 ();
 b15zdnd11an1n04x5 FILLER_294_2186 ();
 b15zdnd00an1n01x5 FILLER_294_2190 ();
 b15zdnd11an1n32x5 FILLER_294_2233 ();
 b15zdnd11an1n08x5 FILLER_294_2265 ();
 b15zdnd00an1n02x5 FILLER_294_2273 ();
 b15zdnd00an1n01x5 FILLER_294_2275 ();
 b15zdnd11an1n64x5 FILLER_295_0 ();
 b15zdnd11an1n64x5 FILLER_295_64 ();
 b15zdnd11an1n64x5 FILLER_295_128 ();
 b15zdnd11an1n64x5 FILLER_295_192 ();
 b15zdnd11an1n32x5 FILLER_295_256 ();
 b15zdnd11an1n16x5 FILLER_295_288 ();
 b15zdnd11an1n08x5 FILLER_295_304 ();
 b15zdnd11an1n64x5 FILLER_295_315 ();
 b15zdnd11an1n64x5 FILLER_295_379 ();
 b15zdnd11an1n64x5 FILLER_295_443 ();
 b15zdnd11an1n64x5 FILLER_295_507 ();
 b15zdnd11an1n64x5 FILLER_295_571 ();
 b15zdnd11an1n64x5 FILLER_295_635 ();
 b15zdnd11an1n64x5 FILLER_295_699 ();
 b15zdnd11an1n64x5 FILLER_295_763 ();
 b15zdnd00an1n02x5 FILLER_295_827 ();
 b15zdnd00an1n01x5 FILLER_295_829 ();
 b15zdnd11an1n64x5 FILLER_295_872 ();
 b15zdnd11an1n64x5 FILLER_295_936 ();
 b15zdnd11an1n64x5 FILLER_295_1000 ();
 b15zdnd11an1n64x5 FILLER_295_1064 ();
 b15zdnd11an1n32x5 FILLER_295_1128 ();
 b15zdnd11an1n04x5 FILLER_295_1160 ();
 b15zdnd11an1n04x5 FILLER_295_1167 ();
 b15zdnd11an1n64x5 FILLER_295_1174 ();
 b15zdnd11an1n32x5 FILLER_295_1238 ();
 b15zdnd11an1n16x5 FILLER_295_1270 ();
 b15zdnd11an1n04x5 FILLER_295_1286 ();
 b15zdnd11an1n08x5 FILLER_295_1293 ();
 b15zdnd11an1n04x5 FILLER_295_1301 ();
 b15zdnd00an1n02x5 FILLER_295_1305 ();
 b15zdnd11an1n04x5 FILLER_295_1310 ();
 b15zdnd11an1n64x5 FILLER_295_1318 ();
 b15zdnd11an1n64x5 FILLER_295_1382 ();
 b15zdnd11an1n32x5 FILLER_295_1446 ();
 b15zdnd11an1n16x5 FILLER_295_1478 ();
 b15zdnd11an1n04x5 FILLER_295_1494 ();
 b15zdnd00an1n01x5 FILLER_295_1498 ();
 b15zdnd11an1n08x5 FILLER_295_1509 ();
 b15zdnd00an1n02x5 FILLER_295_1517 ();
 b15zdnd11an1n04x5 FILLER_295_1529 ();
 b15zdnd11an1n64x5 FILLER_295_1536 ();
 b15zdnd11an1n64x5 FILLER_295_1600 ();
 b15zdnd11an1n64x5 FILLER_295_1664 ();
 b15zdnd11an1n64x5 FILLER_295_1728 ();
 b15zdnd11an1n64x5 FILLER_295_1792 ();
 b15zdnd11an1n64x5 FILLER_295_1856 ();
 b15zdnd11an1n64x5 FILLER_295_1920 ();
 b15zdnd11an1n64x5 FILLER_295_1984 ();
 b15zdnd11an1n64x5 FILLER_295_2048 ();
 b15zdnd11an1n64x5 FILLER_295_2112 ();
 b15zdnd11an1n64x5 FILLER_295_2176 ();
 b15zdnd11an1n32x5 FILLER_295_2240 ();
 b15zdnd11an1n08x5 FILLER_295_2272 ();
 b15zdnd11an1n04x5 FILLER_295_2280 ();
 b15zdnd11an1n04x5 FILLER_296_8 ();
 b15zdnd00an1n01x5 FILLER_296_12 ();
 b15zdnd11an1n08x5 FILLER_296_19 ();
 b15zdnd11an1n04x5 FILLER_296_27 ();
 b15zdnd11an1n64x5 FILLER_296_39 ();
 b15zdnd11an1n64x5 FILLER_296_103 ();
 b15zdnd11an1n64x5 FILLER_296_167 ();
 b15zdnd11an1n64x5 FILLER_296_231 ();
 b15zdnd11an1n64x5 FILLER_296_295 ();
 b15zdnd11an1n64x5 FILLER_296_359 ();
 b15zdnd11an1n64x5 FILLER_296_423 ();
 b15zdnd11an1n64x5 FILLER_296_487 ();
 b15zdnd11an1n64x5 FILLER_296_551 ();
 b15zdnd11an1n64x5 FILLER_296_615 ();
 b15zdnd11an1n32x5 FILLER_296_679 ();
 b15zdnd11an1n04x5 FILLER_296_711 ();
 b15zdnd00an1n02x5 FILLER_296_715 ();
 b15zdnd00an1n01x5 FILLER_296_717 ();
 b15zdnd11an1n64x5 FILLER_296_726 ();
 b15zdnd11an1n64x5 FILLER_296_790 ();
 b15zdnd11an1n64x5 FILLER_296_854 ();
 b15zdnd11an1n64x5 FILLER_296_918 ();
 b15zdnd11an1n64x5 FILLER_296_982 ();
 b15zdnd11an1n64x5 FILLER_296_1046 ();
 b15zdnd11an1n16x5 FILLER_296_1110 ();
 b15zdnd11an1n08x5 FILLER_296_1126 ();
 b15zdnd11an1n04x5 FILLER_296_1134 ();
 b15zdnd00an1n01x5 FILLER_296_1138 ();
 b15zdnd11an1n08x5 FILLER_296_1191 ();
 b15zdnd11an1n04x5 FILLER_296_1199 ();
 b15zdnd11an1n32x5 FILLER_296_1206 ();
 b15zdnd11an1n16x5 FILLER_296_1238 ();
 b15zdnd11an1n08x5 FILLER_296_1254 ();
 b15zdnd00an1n02x5 FILLER_296_1262 ();
 b15zdnd00an1n01x5 FILLER_296_1264 ();
 b15zdnd11an1n64x5 FILLER_296_1317 ();
 b15zdnd11an1n64x5 FILLER_296_1381 ();
 b15zdnd11an1n32x5 FILLER_296_1445 ();
 b15zdnd11an1n16x5 FILLER_296_1477 ();
 b15zdnd11an1n04x5 FILLER_296_1493 ();
 b15zdnd00an1n01x5 FILLER_296_1497 ();
 b15zdnd11an1n04x5 FILLER_296_1506 ();
 b15zdnd11an1n64x5 FILLER_296_1552 ();
 b15zdnd11an1n64x5 FILLER_296_1616 ();
 b15zdnd11an1n64x5 FILLER_296_1680 ();
 b15zdnd11an1n64x5 FILLER_296_1744 ();
 b15zdnd11an1n64x5 FILLER_296_1808 ();
 b15zdnd11an1n64x5 FILLER_296_1872 ();
 b15zdnd11an1n64x5 FILLER_296_1936 ();
 b15zdnd11an1n64x5 FILLER_296_2000 ();
 b15zdnd11an1n32x5 FILLER_296_2064 ();
 b15zdnd11an1n16x5 FILLER_296_2096 ();
 b15zdnd11an1n08x5 FILLER_296_2112 ();
 b15zdnd00an1n02x5 FILLER_296_2152 ();
 b15zdnd11an1n64x5 FILLER_296_2162 ();
 b15zdnd11an1n32x5 FILLER_296_2226 ();
 b15zdnd11an1n16x5 FILLER_296_2258 ();
 b15zdnd00an1n02x5 FILLER_296_2274 ();
 b15zdnd11an1n64x5 FILLER_297_0 ();
 b15zdnd11an1n16x5 FILLER_297_64 ();
 b15zdnd11an1n04x5 FILLER_297_80 ();
 b15zdnd00an1n02x5 FILLER_297_84 ();
 b15zdnd11an1n64x5 FILLER_297_90 ();
 b15zdnd11an1n64x5 FILLER_297_154 ();
 b15zdnd11an1n64x5 FILLER_297_218 ();
 b15zdnd11an1n32x5 FILLER_297_282 ();
 b15zdnd11an1n16x5 FILLER_297_314 ();
 b15zdnd00an1n02x5 FILLER_297_330 ();
 b15zdnd00an1n01x5 FILLER_297_332 ();
 b15zdnd11an1n64x5 FILLER_297_337 ();
 b15zdnd11an1n64x5 FILLER_297_401 ();
 b15zdnd11an1n64x5 FILLER_297_465 ();
 b15zdnd11an1n64x5 FILLER_297_529 ();
 b15zdnd11an1n64x5 FILLER_297_593 ();
 b15zdnd11an1n64x5 FILLER_297_657 ();
 b15zdnd11an1n64x5 FILLER_297_721 ();
 b15zdnd11an1n64x5 FILLER_297_785 ();
 b15zdnd11an1n64x5 FILLER_297_849 ();
 b15zdnd11an1n64x5 FILLER_297_913 ();
 b15zdnd11an1n32x5 FILLER_297_977 ();
 b15zdnd11an1n16x5 FILLER_297_1009 ();
 b15zdnd11an1n04x5 FILLER_297_1025 ();
 b15zdnd11an1n04x5 FILLER_297_1060 ();
 b15zdnd11an1n64x5 FILLER_297_1067 ();
 b15zdnd11an1n32x5 FILLER_297_1131 ();
 b15zdnd00an1n01x5 FILLER_297_1163 ();
 b15zdnd11an1n04x5 FILLER_297_1167 ();
 b15zdnd11an1n04x5 FILLER_297_1211 ();
 b15zdnd11an1n64x5 FILLER_297_1218 ();
 b15zdnd11an1n08x5 FILLER_297_1282 ();
 b15zdnd00an1n01x5 FILLER_297_1290 ();
 b15zdnd11an1n64x5 FILLER_297_1294 ();
 b15zdnd11an1n08x5 FILLER_297_1358 ();
 b15zdnd11an1n04x5 FILLER_297_1366 ();
 b15zdnd00an1n02x5 FILLER_297_1370 ();
 b15zdnd00an1n01x5 FILLER_297_1372 ();
 b15zdnd11an1n04x5 FILLER_297_1379 ();
 b15zdnd11an1n04x5 FILLER_297_1393 ();
 b15zdnd00an1n01x5 FILLER_297_1397 ();
 b15zdnd11an1n64x5 FILLER_297_1401 ();
 b15zdnd11an1n16x5 FILLER_297_1465 ();
 b15zdnd11an1n08x5 FILLER_297_1481 ();
 b15zdnd00an1n02x5 FILLER_297_1489 ();
 b15zdnd00an1n01x5 FILLER_297_1491 ();
 b15zdnd11an1n64x5 FILLER_297_1544 ();
 b15zdnd11an1n64x5 FILLER_297_1608 ();
 b15zdnd11an1n64x5 FILLER_297_1672 ();
 b15zdnd11an1n64x5 FILLER_297_1736 ();
 b15zdnd11an1n64x5 FILLER_297_1800 ();
 b15zdnd11an1n64x5 FILLER_297_1864 ();
 b15zdnd11an1n64x5 FILLER_297_1928 ();
 b15zdnd11an1n64x5 FILLER_297_1992 ();
 b15zdnd11an1n64x5 FILLER_297_2056 ();
 b15zdnd11an1n16x5 FILLER_297_2120 ();
 b15zdnd11an1n08x5 FILLER_297_2136 ();
 b15zdnd00an1n01x5 FILLER_297_2144 ();
 b15zdnd11an1n04x5 FILLER_297_2148 ();
 b15zdnd00an1n02x5 FILLER_297_2152 ();
 b15zdnd00an1n01x5 FILLER_297_2154 ();
 b15zdnd11an1n64x5 FILLER_297_2158 ();
 b15zdnd11an1n32x5 FILLER_297_2227 ();
 b15zdnd11an1n16x5 FILLER_297_2259 ();
 b15zdnd11an1n08x5 FILLER_297_2275 ();
 b15zdnd00an1n01x5 FILLER_297_2283 ();
 b15zdnd11an1n64x5 FILLER_298_8 ();
 b15zdnd11an1n64x5 FILLER_298_72 ();
 b15zdnd11an1n64x5 FILLER_298_136 ();
 b15zdnd11an1n64x5 FILLER_298_200 ();
 b15zdnd11an1n64x5 FILLER_298_264 ();
 b15zdnd11an1n64x5 FILLER_298_328 ();
 b15zdnd11an1n32x5 FILLER_298_392 ();
 b15zdnd11an1n16x5 FILLER_298_424 ();
 b15zdnd11an1n08x5 FILLER_298_440 ();
 b15zdnd00an1n02x5 FILLER_298_448 ();
 b15zdnd11an1n64x5 FILLER_298_492 ();
 b15zdnd11an1n64x5 FILLER_298_556 ();
 b15zdnd11an1n64x5 FILLER_298_620 ();
 b15zdnd11an1n32x5 FILLER_298_684 ();
 b15zdnd00an1n02x5 FILLER_298_716 ();
 b15zdnd11an1n16x5 FILLER_298_726 ();
 b15zdnd11an1n08x5 FILLER_298_742 ();
 b15zdnd11an1n04x5 FILLER_298_750 ();
 b15zdnd11an1n64x5 FILLER_298_766 ();
 b15zdnd11an1n64x5 FILLER_298_830 ();
 b15zdnd11an1n64x5 FILLER_298_894 ();
 b15zdnd11an1n32x5 FILLER_298_958 ();
 b15zdnd11an1n16x5 FILLER_298_990 ();
 b15zdnd11an1n08x5 FILLER_298_1006 ();
 b15zdnd11an1n04x5 FILLER_298_1017 ();
 b15zdnd11an1n04x5 FILLER_298_1061 ();
 b15zdnd11an1n64x5 FILLER_298_1068 ();
 b15zdnd11an1n64x5 FILLER_298_1132 ();
 b15zdnd11an1n64x5 FILLER_298_1196 ();
 b15zdnd11an1n64x5 FILLER_298_1260 ();
 b15zdnd11an1n32x5 FILLER_298_1324 ();
 b15zdnd11an1n04x5 FILLER_298_1356 ();
 b15zdnd00an1n02x5 FILLER_298_1360 ();
 b15zdnd00an1n01x5 FILLER_298_1362 ();
 b15zdnd11an1n04x5 FILLER_298_1379 ();
 b15zdnd11an1n04x5 FILLER_298_1388 ();
 b15zdnd11an1n64x5 FILLER_298_1407 ();
 b15zdnd11an1n32x5 FILLER_298_1471 ();
 b15zdnd11an1n04x5 FILLER_298_1503 ();
 b15zdnd00an1n02x5 FILLER_298_1507 ();
 b15zdnd11an1n04x5 FILLER_298_1512 ();
 b15zdnd11an1n08x5 FILLER_298_1522 ();
 b15zdnd00an1n02x5 FILLER_298_1530 ();
 b15zdnd11an1n64x5 FILLER_298_1574 ();
 b15zdnd11an1n64x5 FILLER_298_1638 ();
 b15zdnd11an1n64x5 FILLER_298_1702 ();
 b15zdnd11an1n64x5 FILLER_298_1766 ();
 b15zdnd11an1n64x5 FILLER_298_1830 ();
 b15zdnd11an1n64x5 FILLER_298_1894 ();
 b15zdnd11an1n32x5 FILLER_298_1958 ();
 b15zdnd11an1n16x5 FILLER_298_1990 ();
 b15zdnd11an1n08x5 FILLER_298_2006 ();
 b15zdnd11an1n04x5 FILLER_298_2014 ();
 b15zdnd11an1n64x5 FILLER_298_2070 ();
 b15zdnd11an1n16x5 FILLER_298_2134 ();
 b15zdnd11an1n04x5 FILLER_298_2150 ();
 b15zdnd11an1n64x5 FILLER_298_2162 ();
 b15zdnd11an1n32x5 FILLER_298_2226 ();
 b15zdnd11an1n16x5 FILLER_298_2258 ();
 b15zdnd00an1n02x5 FILLER_298_2274 ();
 b15zdnd11an1n64x5 FILLER_299_0 ();
 b15zdnd11an1n64x5 FILLER_299_64 ();
 b15zdnd11an1n64x5 FILLER_299_128 ();
 b15zdnd11an1n64x5 FILLER_299_192 ();
 b15zdnd11an1n64x5 FILLER_299_256 ();
 b15zdnd11an1n64x5 FILLER_299_320 ();
 b15zdnd11an1n64x5 FILLER_299_384 ();
 b15zdnd11an1n64x5 FILLER_299_448 ();
 b15zdnd11an1n64x5 FILLER_299_512 ();
 b15zdnd11an1n64x5 FILLER_299_576 ();
 b15zdnd11an1n08x5 FILLER_299_640 ();
 b15zdnd11an1n16x5 FILLER_299_652 ();
 b15zdnd11an1n04x5 FILLER_299_668 ();
 b15zdnd00an1n01x5 FILLER_299_672 ();
 b15zdnd11an1n64x5 FILLER_299_679 ();
 b15zdnd11an1n08x5 FILLER_299_748 ();
 b15zdnd00an1n02x5 FILLER_299_756 ();
 b15zdnd11an1n04x5 FILLER_299_800 ();
 b15zdnd11an1n64x5 FILLER_299_819 ();
 b15zdnd11an1n04x5 FILLER_299_883 ();
 b15zdnd00an1n02x5 FILLER_299_887 ();
 b15zdnd00an1n01x5 FILLER_299_889 ();
 b15zdnd11an1n64x5 FILLER_299_899 ();
 b15zdnd11an1n32x5 FILLER_299_963 ();
 b15zdnd11an1n16x5 FILLER_299_995 ();
 b15zdnd00an1n02x5 FILLER_299_1011 ();
 b15zdnd11an1n64x5 FILLER_299_1055 ();
 b15zdnd11an1n64x5 FILLER_299_1119 ();
 b15zdnd11an1n08x5 FILLER_299_1183 ();
 b15zdnd00an1n02x5 FILLER_299_1191 ();
 b15zdnd00an1n01x5 FILLER_299_1193 ();
 b15zdnd11an1n64x5 FILLER_299_1236 ();
 b15zdnd11an1n64x5 FILLER_299_1300 ();
 b15zdnd11an1n08x5 FILLER_299_1364 ();
 b15zdnd11an1n04x5 FILLER_299_1372 ();
 b15zdnd11an1n04x5 FILLER_299_1387 ();
 b15zdnd11an1n08x5 FILLER_299_1404 ();
 b15zdnd00an1n01x5 FILLER_299_1412 ();
 b15zdnd11an1n64x5 FILLER_299_1428 ();
 b15zdnd11an1n16x5 FILLER_299_1492 ();
 b15zdnd11an1n04x5 FILLER_299_1508 ();
 b15zdnd11an1n08x5 FILLER_299_1515 ();
 b15zdnd11an1n64x5 FILLER_299_1565 ();
 b15zdnd11an1n64x5 FILLER_299_1629 ();
 b15zdnd11an1n64x5 FILLER_299_1693 ();
 b15zdnd11an1n64x5 FILLER_299_1757 ();
 b15zdnd11an1n64x5 FILLER_299_1821 ();
 b15zdnd11an1n64x5 FILLER_299_1885 ();
 b15zdnd11an1n64x5 FILLER_299_1949 ();
 b15zdnd11an1n16x5 FILLER_299_2013 ();
 b15zdnd11an1n04x5 FILLER_299_2029 ();
 b15zdnd00an1n02x5 FILLER_299_2033 ();
 b15zdnd00an1n01x5 FILLER_299_2035 ();
 b15zdnd11an1n04x5 FILLER_299_2039 ();
 b15zdnd11an1n64x5 FILLER_299_2046 ();
 b15zdnd11an1n64x5 FILLER_299_2110 ();
 b15zdnd11an1n64x5 FILLER_299_2174 ();
 b15zdnd11an1n32x5 FILLER_299_2238 ();
 b15zdnd11an1n08x5 FILLER_299_2270 ();
 b15zdnd11an1n04x5 FILLER_299_2278 ();
 b15zdnd00an1n02x5 FILLER_299_2282 ();
 b15zdnd11an1n16x5 FILLER_300_8 ();
 b15zdnd11an1n08x5 FILLER_300_24 ();
 b15zdnd11an1n04x5 FILLER_300_32 ();
 b15zdnd00an1n02x5 FILLER_300_36 ();
 b15zdnd11an1n64x5 FILLER_300_43 ();
 b15zdnd11an1n64x5 FILLER_300_107 ();
 b15zdnd11an1n64x5 FILLER_300_171 ();
 b15zdnd11an1n64x5 FILLER_300_235 ();
 b15zdnd11an1n64x5 FILLER_300_299 ();
 b15zdnd11an1n64x5 FILLER_300_363 ();
 b15zdnd11an1n64x5 FILLER_300_427 ();
 b15zdnd11an1n64x5 FILLER_300_491 ();
 b15zdnd11an1n64x5 FILLER_300_555 ();
 b15zdnd11an1n16x5 FILLER_300_619 ();
 b15zdnd11an1n08x5 FILLER_300_635 ();
 b15zdnd00an1n02x5 FILLER_300_643 ();
 b15zdnd00an1n01x5 FILLER_300_645 ();
 b15zdnd11an1n04x5 FILLER_300_651 ();
 b15zdnd00an1n01x5 FILLER_300_655 ();
 b15zdnd11an1n04x5 FILLER_300_661 ();
 b15zdnd11an1n04x5 FILLER_300_669 ();
 b15zdnd11an1n04x5 FILLER_300_683 ();
 b15zdnd11an1n16x5 FILLER_300_691 ();
 b15zdnd11an1n08x5 FILLER_300_707 ();
 b15zdnd00an1n02x5 FILLER_300_715 ();
 b15zdnd00an1n01x5 FILLER_300_717 ();
 b15zdnd11an1n16x5 FILLER_300_726 ();
 b15zdnd00an1n01x5 FILLER_300_742 ();
 b15zdnd11an1n04x5 FILLER_300_746 ();
 b15zdnd11an1n04x5 FILLER_300_802 ();
 b15zdnd11an1n32x5 FILLER_300_848 ();
 b15zdnd11an1n16x5 FILLER_300_880 ();
 b15zdnd11an1n04x5 FILLER_300_896 ();
 b15zdnd11an1n04x5 FILLER_300_906 ();
 b15zdnd11an1n08x5 FILLER_300_914 ();
 b15zdnd00an1n01x5 FILLER_300_922 ();
 b15zdnd11an1n64x5 FILLER_300_926 ();
 b15zdnd00an1n01x5 FILLER_300_990 ();
 b15zdnd11an1n32x5 FILLER_300_1043 ();
 b15zdnd00an1n01x5 FILLER_300_1075 ();
 b15zdnd11an1n04x5 FILLER_300_1079 ();
 b15zdnd11an1n64x5 FILLER_300_1086 ();
 b15zdnd11an1n64x5 FILLER_300_1150 ();
 b15zdnd11an1n64x5 FILLER_300_1214 ();
 b15zdnd11an1n64x5 FILLER_300_1278 ();
 b15zdnd11an1n32x5 FILLER_300_1342 ();
 b15zdnd00an1n02x5 FILLER_300_1374 ();
 b15zdnd00an1n01x5 FILLER_300_1376 ();
 b15zdnd11an1n08x5 FILLER_300_1381 ();
 b15zdnd00an1n01x5 FILLER_300_1389 ();
 b15zdnd11an1n64x5 FILLER_300_1395 ();
 b15zdnd11an1n32x5 FILLER_300_1459 ();
 b15zdnd11an1n08x5 FILLER_300_1491 ();
 b15zdnd00an1n01x5 FILLER_300_1499 ();
 b15zdnd11an1n08x5 FILLER_300_1504 ();
 b15zdnd00an1n02x5 FILLER_300_1512 ();
 b15zdnd11an1n04x5 FILLER_300_1518 ();
 b15zdnd11an1n64x5 FILLER_300_1564 ();
 b15zdnd11an1n64x5 FILLER_300_1628 ();
 b15zdnd11an1n64x5 FILLER_300_1692 ();
 b15zdnd11an1n32x5 FILLER_300_1756 ();
 b15zdnd11an1n08x5 FILLER_300_1788 ();
 b15zdnd11an1n04x5 FILLER_300_1796 ();
 b15zdnd11an1n64x5 FILLER_300_1803 ();
 b15zdnd11an1n64x5 FILLER_300_1867 ();
 b15zdnd11an1n64x5 FILLER_300_1931 ();
 b15zdnd11an1n32x5 FILLER_300_1995 ();
 b15zdnd11an1n16x5 FILLER_300_2027 ();
 b15zdnd00an1n01x5 FILLER_300_2043 ();
 b15zdnd11an1n64x5 FILLER_300_2047 ();
 b15zdnd11an1n32x5 FILLER_300_2111 ();
 b15zdnd11an1n08x5 FILLER_300_2143 ();
 b15zdnd00an1n02x5 FILLER_300_2151 ();
 b15zdnd00an1n01x5 FILLER_300_2153 ();
 b15zdnd11an1n64x5 FILLER_300_2162 ();
 b15zdnd11an1n32x5 FILLER_300_2226 ();
 b15zdnd11an1n16x5 FILLER_300_2258 ();
 b15zdnd00an1n02x5 FILLER_300_2274 ();
 b15zdnd11an1n64x5 FILLER_301_0 ();
 b15zdnd11an1n64x5 FILLER_301_64 ();
 b15zdnd11an1n64x5 FILLER_301_128 ();
 b15zdnd11an1n64x5 FILLER_301_192 ();
 b15zdnd11an1n64x5 FILLER_301_256 ();
 b15zdnd11an1n64x5 FILLER_301_320 ();
 b15zdnd11an1n64x5 FILLER_301_384 ();
 b15zdnd11an1n64x5 FILLER_301_448 ();
 b15zdnd11an1n64x5 FILLER_301_512 ();
 b15zdnd11an1n32x5 FILLER_301_576 ();
 b15zdnd11an1n04x5 FILLER_301_608 ();
 b15zdnd11an1n04x5 FILLER_301_654 ();
 b15zdnd11an1n04x5 FILLER_301_664 ();
 b15zdnd00an1n02x5 FILLER_301_668 ();
 b15zdnd11an1n04x5 FILLER_301_680 ();
 b15zdnd11an1n32x5 FILLER_301_726 ();
 b15zdnd11an1n08x5 FILLER_301_758 ();
 b15zdnd11an1n04x5 FILLER_301_766 ();
 b15zdnd11an1n04x5 FILLER_301_773 ();
 b15zdnd11an1n04x5 FILLER_301_780 ();
 b15zdnd11an1n64x5 FILLER_301_787 ();
 b15zdnd11an1n16x5 FILLER_301_851 ();
 b15zdnd11an1n04x5 FILLER_301_867 ();
 b15zdnd00an1n01x5 FILLER_301_871 ();
 b15zdnd11an1n08x5 FILLER_301_876 ();
 b15zdnd11an1n04x5 FILLER_301_884 ();
 b15zdnd00an1n01x5 FILLER_301_888 ();
 b15zdnd11an1n04x5 FILLER_301_892 ();
 b15zdnd11an1n04x5 FILLER_301_902 ();
 b15zdnd11an1n32x5 FILLER_301_948 ();
 b15zdnd11an1n16x5 FILLER_301_980 ();
 b15zdnd11an1n08x5 FILLER_301_996 ();
 b15zdnd11an1n04x5 FILLER_301_1004 ();
 b15zdnd00an1n01x5 FILLER_301_1008 ();
 b15zdnd11an1n04x5 FILLER_301_1012 ();
 b15zdnd11an1n32x5 FILLER_301_1019 ();
 b15zdnd00an1n02x5 FILLER_301_1051 ();
 b15zdnd11an1n64x5 FILLER_301_1105 ();
 b15zdnd11an1n64x5 FILLER_301_1169 ();
 b15zdnd11an1n64x5 FILLER_301_1233 ();
 b15zdnd11an1n64x5 FILLER_301_1297 ();
 b15zdnd11an1n64x5 FILLER_301_1361 ();
 b15zdnd11an1n64x5 FILLER_301_1425 ();
 b15zdnd11an1n32x5 FILLER_301_1489 ();
 b15zdnd11an1n64x5 FILLER_301_1528 ();
 b15zdnd11an1n64x5 FILLER_301_1592 ();
 b15zdnd11an1n16x5 FILLER_301_1656 ();
 b15zdnd11an1n08x5 FILLER_301_1672 ();
 b15zdnd00an1n02x5 FILLER_301_1680 ();
 b15zdnd00an1n01x5 FILLER_301_1682 ();
 b15zdnd11an1n64x5 FILLER_301_1686 ();
 b15zdnd11an1n32x5 FILLER_301_1750 ();
 b15zdnd11an1n16x5 FILLER_301_1782 ();
 b15zdnd00an1n01x5 FILLER_301_1798 ();
 b15zdnd11an1n64x5 FILLER_301_1802 ();
 b15zdnd11an1n64x5 FILLER_301_1866 ();
 b15zdnd11an1n64x5 FILLER_301_1930 ();
 b15zdnd11an1n32x5 FILLER_301_1994 ();
 b15zdnd11an1n08x5 FILLER_301_2026 ();
 b15zdnd00an1n02x5 FILLER_301_2034 ();
 b15zdnd11an1n04x5 FILLER_301_2039 ();
 b15zdnd00an1n01x5 FILLER_301_2043 ();
 b15zdnd11an1n64x5 FILLER_301_2047 ();
 b15zdnd11an1n16x5 FILLER_301_2111 ();
 b15zdnd11an1n04x5 FILLER_301_2127 ();
 b15zdnd00an1n02x5 FILLER_301_2131 ();
 b15zdnd00an1n01x5 FILLER_301_2133 ();
 b15zdnd11an1n64x5 FILLER_301_2176 ();
 b15zdnd11an1n32x5 FILLER_301_2240 ();
 b15zdnd11an1n08x5 FILLER_301_2272 ();
 b15zdnd11an1n04x5 FILLER_301_2280 ();
 b15zdnd11an1n64x5 FILLER_302_8 ();
 b15zdnd11an1n64x5 FILLER_302_72 ();
 b15zdnd11an1n64x5 FILLER_302_136 ();
 b15zdnd11an1n64x5 FILLER_302_200 ();
 b15zdnd11an1n64x5 FILLER_302_264 ();
 b15zdnd11an1n64x5 FILLER_302_328 ();
 b15zdnd11an1n64x5 FILLER_302_392 ();
 b15zdnd11an1n32x5 FILLER_302_456 ();
 b15zdnd11an1n16x5 FILLER_302_488 ();
 b15zdnd11an1n08x5 FILLER_302_504 ();
 b15zdnd00an1n02x5 FILLER_302_512 ();
 b15zdnd11an1n04x5 FILLER_302_517 ();
 b15zdnd11an1n08x5 FILLER_302_524 ();
 b15zdnd11an1n04x5 FILLER_302_532 ();
 b15zdnd00an1n02x5 FILLER_302_536 ();
 b15zdnd11an1n32x5 FILLER_302_580 ();
 b15zdnd11an1n08x5 FILLER_302_612 ();
 b15zdnd00an1n02x5 FILLER_302_620 ();
 b15zdnd11an1n04x5 FILLER_302_664 ();
 b15zdnd00an1n02x5 FILLER_302_668 ();
 b15zdnd00an1n01x5 FILLER_302_670 ();
 b15zdnd11an1n04x5 FILLER_302_713 ();
 b15zdnd00an1n01x5 FILLER_302_717 ();
 b15zdnd11an1n64x5 FILLER_302_726 ();
 b15zdnd11an1n64x5 FILLER_302_790 ();
 b15zdnd11an1n08x5 FILLER_302_854 ();
 b15zdnd00an1n01x5 FILLER_302_862 ();
 b15zdnd11an1n16x5 FILLER_302_866 ();
 b15zdnd00an1n02x5 FILLER_302_882 ();
 b15zdnd00an1n01x5 FILLER_302_884 ();
 b15zdnd11an1n04x5 FILLER_302_892 ();
 b15zdnd11an1n64x5 FILLER_302_948 ();
 b15zdnd11an1n16x5 FILLER_302_1012 ();
 b15zdnd11an1n08x5 FILLER_302_1028 ();
 b15zdnd00an1n02x5 FILLER_302_1036 ();
 b15zdnd11an1n04x5 FILLER_302_1080 ();
 b15zdnd00an1n02x5 FILLER_302_1084 ();
 b15zdnd00an1n01x5 FILLER_302_1086 ();
 b15zdnd11an1n64x5 FILLER_302_1090 ();
 b15zdnd11an1n64x5 FILLER_302_1154 ();
 b15zdnd11an1n64x5 FILLER_302_1218 ();
 b15zdnd11an1n64x5 FILLER_302_1282 ();
 b15zdnd11an1n64x5 FILLER_302_1346 ();
 b15zdnd11an1n64x5 FILLER_302_1410 ();
 b15zdnd11an1n64x5 FILLER_302_1474 ();
 b15zdnd11an1n64x5 FILLER_302_1538 ();
 b15zdnd11an1n64x5 FILLER_302_1602 ();
 b15zdnd11an1n08x5 FILLER_302_1666 ();
 b15zdnd00an1n02x5 FILLER_302_1674 ();
 b15zdnd00an1n01x5 FILLER_302_1676 ();
 b15zdnd11an1n04x5 FILLER_302_1680 ();
 b15zdnd11an1n04x5 FILLER_302_1687 ();
 b15zdnd11an1n64x5 FILLER_302_1694 ();
 b15zdnd11an1n16x5 FILLER_302_1758 ();
 b15zdnd11an1n64x5 FILLER_302_1826 ();
 b15zdnd11an1n08x5 FILLER_302_1890 ();
 b15zdnd00an1n02x5 FILLER_302_1898 ();
 b15zdnd11an1n64x5 FILLER_302_1904 ();
 b15zdnd11an1n32x5 FILLER_302_1968 ();
 b15zdnd11an1n04x5 FILLER_302_2000 ();
 b15zdnd00an1n01x5 FILLER_302_2004 ();
 b15zdnd11an1n16x5 FILLER_302_2045 ();
 b15zdnd11an1n04x5 FILLER_302_2061 ();
 b15zdnd00an1n02x5 FILLER_302_2065 ();
 b15zdnd00an1n01x5 FILLER_302_2067 ();
 b15zdnd11an1n04x5 FILLER_302_2071 ();
 b15zdnd11an1n64x5 FILLER_302_2078 ();
 b15zdnd11an1n08x5 FILLER_302_2142 ();
 b15zdnd11an1n04x5 FILLER_302_2150 ();
 b15zdnd11an1n64x5 FILLER_302_2162 ();
 b15zdnd11an1n32x5 FILLER_302_2226 ();
 b15zdnd11an1n16x5 FILLER_302_2258 ();
 b15zdnd00an1n02x5 FILLER_302_2274 ();
 b15zdnd11an1n32x5 FILLER_303_0 ();
 b15zdnd11an1n16x5 FILLER_303_32 ();
 b15zdnd11an1n08x5 FILLER_303_48 ();
 b15zdnd11an1n04x5 FILLER_303_56 ();
 b15zdnd00an1n01x5 FILLER_303_60 ();
 b15zdnd11an1n64x5 FILLER_303_73 ();
 b15zdnd11an1n64x5 FILLER_303_137 ();
 b15zdnd11an1n64x5 FILLER_303_201 ();
 b15zdnd11an1n04x5 FILLER_303_265 ();
 b15zdnd00an1n01x5 FILLER_303_269 ();
 b15zdnd11an1n64x5 FILLER_303_273 ();
 b15zdnd11an1n64x5 FILLER_303_337 ();
 b15zdnd11an1n64x5 FILLER_303_401 ();
 b15zdnd11an1n16x5 FILLER_303_465 ();
 b15zdnd11an1n04x5 FILLER_303_521 ();
 b15zdnd00an1n02x5 FILLER_303_525 ();
 b15zdnd00an1n01x5 FILLER_303_527 ();
 b15zdnd11an1n08x5 FILLER_303_534 ();
 b15zdnd00an1n02x5 FILLER_303_542 ();
 b15zdnd11an1n32x5 FILLER_303_596 ();
 b15zdnd11an1n08x5 FILLER_303_628 ();
 b15zdnd11an1n04x5 FILLER_303_636 ();
 b15zdnd00an1n01x5 FILLER_303_640 ();
 b15zdnd11an1n64x5 FILLER_303_693 ();
 b15zdnd11an1n64x5 FILLER_303_757 ();
 b15zdnd11an1n16x5 FILLER_303_821 ();
 b15zdnd11an1n08x5 FILLER_303_837 ();
 b15zdnd11an1n04x5 FILLER_303_845 ();
 b15zdnd00an1n01x5 FILLER_303_849 ();
 b15zdnd11an1n32x5 FILLER_303_856 ();
 b15zdnd11an1n04x5 FILLER_303_888 ();
 b15zdnd00an1n01x5 FILLER_303_892 ();
 b15zdnd11an1n04x5 FILLER_303_899 ();
 b15zdnd11an1n04x5 FILLER_303_908 ();
 b15zdnd00an1n02x5 FILLER_303_912 ();
 b15zdnd11an1n04x5 FILLER_303_917 ();
 b15zdnd11an1n64x5 FILLER_303_924 ();
 b15zdnd11an1n64x5 FILLER_303_988 ();
 b15zdnd11an1n16x5 FILLER_303_1052 ();
 b15zdnd11an1n04x5 FILLER_303_1068 ();
 b15zdnd00an1n01x5 FILLER_303_1072 ();
 b15zdnd11an1n04x5 FILLER_303_1076 ();
 b15zdnd11an1n64x5 FILLER_303_1083 ();
 b15zdnd11an1n64x5 FILLER_303_1147 ();
 b15zdnd11an1n64x5 FILLER_303_1211 ();
 b15zdnd11an1n64x5 FILLER_303_1275 ();
 b15zdnd11an1n64x5 FILLER_303_1339 ();
 b15zdnd11an1n64x5 FILLER_303_1403 ();
 b15zdnd11an1n64x5 FILLER_303_1467 ();
 b15zdnd11an1n64x5 FILLER_303_1531 ();
 b15zdnd11an1n64x5 FILLER_303_1595 ();
 b15zdnd11an1n04x5 FILLER_303_1659 ();
 b15zdnd11an1n64x5 FILLER_303_1715 ();
 b15zdnd11an1n08x5 FILLER_303_1779 ();
 b15zdnd11an1n04x5 FILLER_303_1787 ();
 b15zdnd00an1n01x5 FILLER_303_1791 ();
 b15zdnd11an1n04x5 FILLER_303_1795 ();
 b15zdnd11an1n04x5 FILLER_303_1802 ();
 b15zdnd11an1n64x5 FILLER_303_1813 ();
 b15zdnd11an1n08x5 FILLER_303_1877 ();
 b15zdnd11an1n04x5 FILLER_303_1896 ();
 b15zdnd11an1n16x5 FILLER_303_1905 ();
 b15zdnd11an1n04x5 FILLER_303_1921 ();
 b15zdnd00an1n02x5 FILLER_303_1925 ();
 b15zdnd00an1n01x5 FILLER_303_1927 ();
 b15zdnd11an1n04x5 FILLER_303_1931 ();
 b15zdnd11an1n64x5 FILLER_303_1938 ();
 b15zdnd11an1n16x5 FILLER_303_2002 ();
 b15zdnd11an1n04x5 FILLER_303_2018 ();
 b15zdnd00an1n02x5 FILLER_303_2022 ();
 b15zdnd00an1n01x5 FILLER_303_2024 ();
 b15zdnd11an1n32x5 FILLER_303_2034 ();
 b15zdnd00an1n02x5 FILLER_303_2066 ();
 b15zdnd11an1n64x5 FILLER_303_2110 ();
 b15zdnd11an1n32x5 FILLER_303_2174 ();
 b15zdnd11an1n16x5 FILLER_303_2206 ();
 b15zdnd11an1n04x5 FILLER_303_2222 ();
 b15zdnd11an1n32x5 FILLER_303_2242 ();
 b15zdnd11an1n08x5 FILLER_303_2274 ();
 b15zdnd00an1n02x5 FILLER_303_2282 ();
 b15zdnd11an1n32x5 FILLER_304_8 ();
 b15zdnd11an1n16x5 FILLER_304_40 ();
 b15zdnd11an1n04x5 FILLER_304_56 ();
 b15zdnd00an1n02x5 FILLER_304_60 ();
 b15zdnd00an1n01x5 FILLER_304_62 ();
 b15zdnd11an1n64x5 FILLER_304_70 ();
 b15zdnd11an1n64x5 FILLER_304_134 ();
 b15zdnd11an1n16x5 FILLER_304_198 ();
 b15zdnd11an1n04x5 FILLER_304_214 ();
 b15zdnd00an1n01x5 FILLER_304_218 ();
 b15zdnd11an1n08x5 FILLER_304_222 ();
 b15zdnd11an1n04x5 FILLER_304_230 ();
 b15zdnd00an1n02x5 FILLER_304_234 ();
 b15zdnd00an1n01x5 FILLER_304_236 ();
 b15zdnd11an1n64x5 FILLER_304_277 ();
 b15zdnd11an1n64x5 FILLER_304_341 ();
 b15zdnd11an1n64x5 FILLER_304_405 ();
 b15zdnd11an1n64x5 FILLER_304_469 ();
 b15zdnd11an1n16x5 FILLER_304_533 ();
 b15zdnd11an1n08x5 FILLER_304_549 ();
 b15zdnd11an1n04x5 FILLER_304_557 ();
 b15zdnd00an1n02x5 FILLER_304_561 ();
 b15zdnd00an1n01x5 FILLER_304_563 ();
 b15zdnd11an1n04x5 FILLER_304_567 ();
 b15zdnd11an1n32x5 FILLER_304_574 ();
 b15zdnd11an1n08x5 FILLER_304_606 ();
 b15zdnd11an1n04x5 FILLER_304_614 ();
 b15zdnd00an1n02x5 FILLER_304_618 ();
 b15zdnd00an1n01x5 FILLER_304_620 ();
 b15zdnd11an1n04x5 FILLER_304_663 ();
 b15zdnd00an1n01x5 FILLER_304_667 ();
 b15zdnd11an1n04x5 FILLER_304_671 ();
 b15zdnd11an1n32x5 FILLER_304_678 ();
 b15zdnd11an1n08x5 FILLER_304_710 ();
 b15zdnd11an1n64x5 FILLER_304_726 ();
 b15zdnd11an1n64x5 FILLER_304_790 ();
 b15zdnd11an1n32x5 FILLER_304_854 ();
 b15zdnd11an1n08x5 FILLER_304_886 ();
 b15zdnd00an1n02x5 FILLER_304_894 ();
 b15zdnd00an1n01x5 FILLER_304_896 ();
 b15zdnd11an1n64x5 FILLER_304_901 ();
 b15zdnd11an1n64x5 FILLER_304_965 ();
 b15zdnd11an1n64x5 FILLER_304_1029 ();
 b15zdnd11an1n64x5 FILLER_304_1093 ();
 b15zdnd11an1n64x5 FILLER_304_1157 ();
 b15zdnd11an1n64x5 FILLER_304_1221 ();
 b15zdnd11an1n64x5 FILLER_304_1285 ();
 b15zdnd11an1n32x5 FILLER_304_1349 ();
 b15zdnd11an1n16x5 FILLER_304_1381 ();
 b15zdnd11an1n04x5 FILLER_304_1397 ();
 b15zdnd11an1n08x5 FILLER_304_1404 ();
 b15zdnd00an1n01x5 FILLER_304_1412 ();
 b15zdnd11an1n64x5 FILLER_304_1416 ();
 b15zdnd11an1n64x5 FILLER_304_1480 ();
 b15zdnd11an1n64x5 FILLER_304_1544 ();
 b15zdnd11an1n32x5 FILLER_304_1608 ();
 b15zdnd11an1n16x5 FILLER_304_1640 ();
 b15zdnd00an1n02x5 FILLER_304_1656 ();
 b15zdnd00an1n01x5 FILLER_304_1658 ();
 b15zdnd11an1n32x5 FILLER_304_1711 ();
 b15zdnd11an1n08x5 FILLER_304_1743 ();
 b15zdnd11an1n04x5 FILLER_304_1751 ();
 b15zdnd00an1n02x5 FILLER_304_1755 ();
 b15zdnd00an1n01x5 FILLER_304_1757 ();
 b15zdnd11an1n04x5 FILLER_304_1798 ();
 b15zdnd11an1n04x5 FILLER_304_1805 ();
 b15zdnd11an1n32x5 FILLER_304_1815 ();
 b15zdnd11an1n16x5 FILLER_304_1847 ();
 b15zdnd11an1n08x5 FILLER_304_1863 ();
 b15zdnd11an1n04x5 FILLER_304_1877 ();
 b15zdnd11an1n04x5 FILLER_304_1890 ();
 b15zdnd11an1n08x5 FILLER_304_1899 ();
 b15zdnd00an1n02x5 FILLER_304_1907 ();
 b15zdnd11an1n64x5 FILLER_304_1951 ();
 b15zdnd11an1n32x5 FILLER_304_2015 ();
 b15zdnd00an1n02x5 FILLER_304_2047 ();
 b15zdnd00an1n01x5 FILLER_304_2049 ();
 b15zdnd11an1n32x5 FILLER_304_2102 ();
 b15zdnd11an1n16x5 FILLER_304_2134 ();
 b15zdnd11an1n04x5 FILLER_304_2150 ();
 b15zdnd11an1n32x5 FILLER_304_2162 ();
 b15zdnd11an1n16x5 FILLER_304_2194 ();
 b15zdnd11an1n32x5 FILLER_304_2219 ();
 b15zdnd11an1n16x5 FILLER_304_2251 ();
 b15zdnd11an1n08x5 FILLER_304_2267 ();
 b15zdnd00an1n01x5 FILLER_304_2275 ();
 b15zdnd11an1n32x5 FILLER_305_0 ();
 b15zdnd11an1n16x5 FILLER_305_32 ();
 b15zdnd11an1n08x5 FILLER_305_48 ();
 b15zdnd11an1n04x5 FILLER_305_56 ();
 b15zdnd00an1n02x5 FILLER_305_60 ();
 b15zdnd11an1n64x5 FILLER_305_68 ();
 b15zdnd11an1n32x5 FILLER_305_132 ();
 b15zdnd11an1n16x5 FILLER_305_164 ();
 b15zdnd11an1n04x5 FILLER_305_180 ();
 b15zdnd00an1n01x5 FILLER_305_184 ();
 b15zdnd11an1n04x5 FILLER_305_225 ();
 b15zdnd11an1n32x5 FILLER_305_232 ();
 b15zdnd11an1n08x5 FILLER_305_264 ();
 b15zdnd00an1n02x5 FILLER_305_272 ();
 b15zdnd00an1n01x5 FILLER_305_274 ();
 b15zdnd11an1n64x5 FILLER_305_278 ();
 b15zdnd11an1n64x5 FILLER_305_342 ();
 b15zdnd11an1n64x5 FILLER_305_406 ();
 b15zdnd11an1n64x5 FILLER_305_470 ();
 b15zdnd11an1n16x5 FILLER_305_534 ();
 b15zdnd00an1n01x5 FILLER_305_550 ();
 b15zdnd11an1n04x5 FILLER_305_554 ();
 b15zdnd11an1n04x5 FILLER_305_561 ();
 b15zdnd11an1n64x5 FILLER_305_568 ();
 b15zdnd11an1n32x5 FILLER_305_632 ();
 b15zdnd00an1n02x5 FILLER_305_664 ();
 b15zdnd00an1n01x5 FILLER_305_666 ();
 b15zdnd11an1n64x5 FILLER_305_670 ();
 b15zdnd11an1n64x5 FILLER_305_734 ();
 b15zdnd11an1n64x5 FILLER_305_798 ();
 b15zdnd11an1n64x5 FILLER_305_862 ();
 b15zdnd11an1n64x5 FILLER_305_926 ();
 b15zdnd11an1n64x5 FILLER_305_990 ();
 b15zdnd11an1n64x5 FILLER_305_1054 ();
 b15zdnd11an1n64x5 FILLER_305_1118 ();
 b15zdnd11an1n64x5 FILLER_305_1182 ();
 b15zdnd11an1n64x5 FILLER_305_1246 ();
 b15zdnd11an1n64x5 FILLER_305_1310 ();
 b15zdnd11an1n04x5 FILLER_305_1374 ();
 b15zdnd11an1n64x5 FILLER_305_1430 ();
 b15zdnd11an1n16x5 FILLER_305_1494 ();
 b15zdnd11an1n04x5 FILLER_305_1510 ();
 b15zdnd00an1n02x5 FILLER_305_1514 ();
 b15zdnd11an1n64x5 FILLER_305_1520 ();
 b15zdnd11an1n32x5 FILLER_305_1584 ();
 b15zdnd11an1n08x5 FILLER_305_1616 ();
 b15zdnd00an1n02x5 FILLER_305_1624 ();
 b15zdnd00an1n01x5 FILLER_305_1626 ();
 b15zdnd11an1n04x5 FILLER_305_1630 ();
 b15zdnd11an1n16x5 FILLER_305_1637 ();
 b15zdnd11an1n04x5 FILLER_305_1653 ();
 b15zdnd00an1n02x5 FILLER_305_1657 ();
 b15zdnd11an1n04x5 FILLER_305_1701 ();
 b15zdnd11an1n64x5 FILLER_305_1747 ();
 b15zdnd11an1n64x5 FILLER_305_1811 ();
 b15zdnd11an1n04x5 FILLER_305_1878 ();
 b15zdnd11an1n16x5 FILLER_305_1893 ();
 b15zdnd00an1n01x5 FILLER_305_1909 ();
 b15zdnd11an1n64x5 FILLER_305_1962 ();
 b15zdnd11an1n32x5 FILLER_305_2026 ();
 b15zdnd11an1n16x5 FILLER_305_2058 ();
 b15zdnd00an1n01x5 FILLER_305_2074 ();
 b15zdnd11an1n64x5 FILLER_305_2078 ();
 b15zdnd11an1n64x5 FILLER_305_2142 ();
 b15zdnd11an1n64x5 FILLER_305_2206 ();
 b15zdnd11an1n08x5 FILLER_305_2270 ();
 b15zdnd11an1n04x5 FILLER_305_2278 ();
 b15zdnd00an1n02x5 FILLER_305_2282 ();
 b15zdnd11an1n32x5 FILLER_306_8 ();
 b15zdnd11an1n16x5 FILLER_306_40 ();
 b15zdnd11an1n04x5 FILLER_306_56 ();
 b15zdnd00an1n02x5 FILLER_306_60 ();
 b15zdnd11an1n64x5 FILLER_306_67 ();
 b15zdnd11an1n32x5 FILLER_306_131 ();
 b15zdnd11an1n16x5 FILLER_306_163 ();
 b15zdnd11an1n04x5 FILLER_306_179 ();
 b15zdnd00an1n02x5 FILLER_306_183 ();
 b15zdnd00an1n01x5 FILLER_306_185 ();
 b15zdnd11an1n64x5 FILLER_306_206 ();
 b15zdnd11an1n64x5 FILLER_306_270 ();
 b15zdnd11an1n64x5 FILLER_306_334 ();
 b15zdnd11an1n64x5 FILLER_306_398 ();
 b15zdnd11an1n32x5 FILLER_306_462 ();
 b15zdnd11an1n16x5 FILLER_306_494 ();
 b15zdnd11an1n08x5 FILLER_306_510 ();
 b15zdnd11an1n04x5 FILLER_306_518 ();
 b15zdnd11an1n64x5 FILLER_306_562 ();
 b15zdnd11an1n64x5 FILLER_306_626 ();
 b15zdnd11an1n16x5 FILLER_306_690 ();
 b15zdnd11an1n08x5 FILLER_306_706 ();
 b15zdnd11an1n04x5 FILLER_306_714 ();
 b15zdnd11an1n64x5 FILLER_306_726 ();
 b15zdnd11an1n64x5 FILLER_306_790 ();
 b15zdnd11an1n64x5 FILLER_306_854 ();
 b15zdnd11an1n64x5 FILLER_306_918 ();
 b15zdnd11an1n64x5 FILLER_306_982 ();
 b15zdnd11an1n64x5 FILLER_306_1046 ();
 b15zdnd11an1n64x5 FILLER_306_1110 ();
 b15zdnd11an1n64x5 FILLER_306_1174 ();
 b15zdnd11an1n64x5 FILLER_306_1238 ();
 b15zdnd11an1n64x5 FILLER_306_1302 ();
 b15zdnd11an1n32x5 FILLER_306_1366 ();
 b15zdnd11an1n04x5 FILLER_306_1398 ();
 b15zdnd11an1n64x5 FILLER_306_1405 ();
 b15zdnd11an1n64x5 FILLER_306_1469 ();
 b15zdnd11an1n32x5 FILLER_306_1533 ();
 b15zdnd11an1n16x5 FILLER_306_1565 ();
 b15zdnd11an1n08x5 FILLER_306_1581 ();
 b15zdnd11an1n04x5 FILLER_306_1589 ();
 b15zdnd00an1n02x5 FILLER_306_1593 ();
 b15zdnd11an1n16x5 FILLER_306_1635 ();
 b15zdnd11an1n04x5 FILLER_306_1651 ();
 b15zdnd11an1n04x5 FILLER_306_1680 ();
 b15zdnd11an1n04x5 FILLER_306_1687 ();
 b15zdnd11an1n04x5 FILLER_306_1694 ();
 b15zdnd11an1n64x5 FILLER_306_1701 ();
 b15zdnd11an1n64x5 FILLER_306_1765 ();
 b15zdnd11an1n64x5 FILLER_306_1829 ();
 b15zdnd11an1n32x5 FILLER_306_1893 ();
 b15zdnd11an1n08x5 FILLER_306_1925 ();
 b15zdnd00an1n02x5 FILLER_306_1933 ();
 b15zdnd11an1n64x5 FILLER_306_1938 ();
 b15zdnd11an1n64x5 FILLER_306_2002 ();
 b15zdnd11an1n64x5 FILLER_306_2066 ();
 b15zdnd11an1n08x5 FILLER_306_2130 ();
 b15zdnd00an1n01x5 FILLER_306_2138 ();
 b15zdnd11an1n04x5 FILLER_306_2142 ();
 b15zdnd11an1n04x5 FILLER_306_2149 ();
 b15zdnd00an1n01x5 FILLER_306_2153 ();
 b15zdnd11an1n32x5 FILLER_306_2162 ();
 b15zdnd11an1n16x5 FILLER_306_2194 ();
 b15zdnd00an1n02x5 FILLER_306_2210 ();
 b15zdnd00an1n01x5 FILLER_306_2212 ();
 b15zdnd11an1n32x5 FILLER_306_2223 ();
 b15zdnd11an1n16x5 FILLER_306_2255 ();
 b15zdnd11an1n04x5 FILLER_306_2271 ();
 b15zdnd00an1n01x5 FILLER_306_2275 ();
 b15zdnd11an1n16x5 FILLER_307_0 ();
 b15zdnd11an1n04x5 FILLER_307_16 ();
 b15zdnd00an1n02x5 FILLER_307_20 ();
 b15zdnd11an1n32x5 FILLER_307_28 ();
 b15zdnd11an1n04x5 FILLER_307_60 ();
 b15zdnd11an1n04x5 FILLER_307_67 ();
 b15zdnd11an1n64x5 FILLER_307_74 ();
 b15zdnd11an1n32x5 FILLER_307_138 ();
 b15zdnd11an1n08x5 FILLER_307_170 ();
 b15zdnd11an1n04x5 FILLER_307_178 ();
 b15zdnd00an1n02x5 FILLER_307_182 ();
 b15zdnd11an1n04x5 FILLER_307_224 ();
 b15zdnd11an1n64x5 FILLER_307_231 ();
 b15zdnd11an1n64x5 FILLER_307_295 ();
 b15zdnd11an1n32x5 FILLER_307_359 ();
 b15zdnd11an1n04x5 FILLER_307_391 ();
 b15zdnd11an1n04x5 FILLER_307_399 ();
 b15zdnd11an1n64x5 FILLER_307_443 ();
 b15zdnd11an1n64x5 FILLER_307_507 ();
 b15zdnd11an1n64x5 FILLER_307_571 ();
 b15zdnd11an1n64x5 FILLER_307_635 ();
 b15zdnd11an1n64x5 FILLER_307_699 ();
 b15zdnd11an1n64x5 FILLER_307_763 ();
 b15zdnd11an1n64x5 FILLER_307_827 ();
 b15zdnd11an1n64x5 FILLER_307_891 ();
 b15zdnd11an1n64x5 FILLER_307_955 ();
 b15zdnd11an1n64x5 FILLER_307_1019 ();
 b15zdnd11an1n64x5 FILLER_307_1083 ();
 b15zdnd11an1n64x5 FILLER_307_1147 ();
 b15zdnd11an1n64x5 FILLER_307_1211 ();
 b15zdnd11an1n64x5 FILLER_307_1275 ();
 b15zdnd11an1n64x5 FILLER_307_1339 ();
 b15zdnd11an1n64x5 FILLER_307_1403 ();
 b15zdnd11an1n64x5 FILLER_307_1467 ();
 b15zdnd11an1n64x5 FILLER_307_1531 ();
 b15zdnd11an1n64x5 FILLER_307_1595 ();
 b15zdnd11an1n32x5 FILLER_307_1659 ();
 b15zdnd11an1n64x5 FILLER_307_1694 ();
 b15zdnd11an1n64x5 FILLER_307_1758 ();
 b15zdnd11an1n32x5 FILLER_307_1822 ();
 b15zdnd11an1n16x5 FILLER_307_1854 ();
 b15zdnd11an1n08x5 FILLER_307_1870 ();
 b15zdnd00an1n01x5 FILLER_307_1878 ();
 b15zdnd11an1n64x5 FILLER_307_1892 ();
 b15zdnd11an1n64x5 FILLER_307_1956 ();
 b15zdnd11an1n32x5 FILLER_307_2020 ();
 b15zdnd11an1n04x5 FILLER_307_2052 ();
 b15zdnd00an1n01x5 FILLER_307_2056 ();
 b15zdnd11an1n32x5 FILLER_307_2075 ();
 b15zdnd11an1n08x5 FILLER_307_2107 ();
 b15zdnd11an1n04x5 FILLER_307_2115 ();
 b15zdnd00an1n02x5 FILLER_307_2119 ();
 b15zdnd11an1n04x5 FILLER_307_2153 ();
 b15zdnd11an1n64x5 FILLER_307_2160 ();
 b15zdnd11an1n32x5 FILLER_307_2224 ();
 b15zdnd11an1n16x5 FILLER_307_2256 ();
 b15zdnd11an1n08x5 FILLER_307_2272 ();
 b15zdnd11an1n04x5 FILLER_307_2280 ();
 b15zdnd11an1n32x5 FILLER_308_8 ();
 b15zdnd11an1n16x5 FILLER_308_40 ();
 b15zdnd00an1n01x5 FILLER_308_56 ();
 b15zdnd11an1n04x5 FILLER_308_63 ();
 b15zdnd11an1n64x5 FILLER_308_74 ();
 b15zdnd11an1n32x5 FILLER_308_138 ();
 b15zdnd11an1n16x5 FILLER_308_170 ();
 b15zdnd00an1n01x5 FILLER_308_186 ();
 b15zdnd11an1n64x5 FILLER_308_229 ();
 b15zdnd11an1n64x5 FILLER_308_293 ();
 b15zdnd11an1n16x5 FILLER_308_357 ();
 b15zdnd00an1n02x5 FILLER_308_373 ();
 b15zdnd00an1n01x5 FILLER_308_375 ();
 b15zdnd11an1n04x5 FILLER_308_392 ();
 b15zdnd11an1n32x5 FILLER_308_399 ();
 b15zdnd00an1n02x5 FILLER_308_431 ();
 b15zdnd00an1n01x5 FILLER_308_433 ();
 b15zdnd11an1n04x5 FILLER_308_437 ();
 b15zdnd11an1n64x5 FILLER_308_444 ();
 b15zdnd11an1n64x5 FILLER_308_508 ();
 b15zdnd11an1n64x5 FILLER_308_572 ();
 b15zdnd11an1n64x5 FILLER_308_636 ();
 b15zdnd11an1n16x5 FILLER_308_700 ();
 b15zdnd00an1n02x5 FILLER_308_716 ();
 b15zdnd11an1n64x5 FILLER_308_726 ();
 b15zdnd11an1n64x5 FILLER_308_790 ();
 b15zdnd11an1n64x5 FILLER_308_854 ();
 b15zdnd11an1n64x5 FILLER_308_918 ();
 b15zdnd11an1n64x5 FILLER_308_982 ();
 b15zdnd11an1n64x5 FILLER_308_1046 ();
 b15zdnd11an1n64x5 FILLER_308_1110 ();
 b15zdnd11an1n64x5 FILLER_308_1174 ();
 b15zdnd11an1n64x5 FILLER_308_1238 ();
 b15zdnd11an1n64x5 FILLER_308_1302 ();
 b15zdnd11an1n64x5 FILLER_308_1366 ();
 b15zdnd11an1n64x5 FILLER_308_1430 ();
 b15zdnd11an1n64x5 FILLER_308_1494 ();
 b15zdnd11an1n64x5 FILLER_308_1558 ();
 b15zdnd11an1n64x5 FILLER_308_1622 ();
 b15zdnd11an1n64x5 FILLER_308_1686 ();
 b15zdnd11an1n16x5 FILLER_308_1750 ();
 b15zdnd11an1n08x5 FILLER_308_1766 ();
 b15zdnd00an1n02x5 FILLER_308_1774 ();
 b15zdnd11an1n08x5 FILLER_308_1785 ();
 b15zdnd11an1n04x5 FILLER_308_1793 ();
 b15zdnd00an1n02x5 FILLER_308_1797 ();
 b15zdnd11an1n64x5 FILLER_308_1808 ();
 b15zdnd11an1n64x5 FILLER_308_1872 ();
 b15zdnd11an1n64x5 FILLER_308_1936 ();
 b15zdnd11an1n64x5 FILLER_308_2000 ();
 b15zdnd11an1n64x5 FILLER_308_2064 ();
 b15zdnd11an1n16x5 FILLER_308_2128 ();
 b15zdnd11an1n08x5 FILLER_308_2144 ();
 b15zdnd00an1n02x5 FILLER_308_2152 ();
 b15zdnd11an1n32x5 FILLER_308_2162 ();
 b15zdnd11an1n16x5 FILLER_308_2194 ();
 b15zdnd11an1n08x5 FILLER_308_2210 ();
 b15zdnd11an1n04x5 FILLER_308_2218 ();
 b15zdnd00an1n02x5 FILLER_308_2222 ();
 b15zdnd11an1n04x5 FILLER_308_2227 ();
 b15zdnd11an1n32x5 FILLER_308_2244 ();
 b15zdnd11an1n16x5 FILLER_309_0 ();
 b15zdnd00an1n02x5 FILLER_309_16 ();
 b15zdnd00an1n01x5 FILLER_309_18 ();
 b15zdnd11an1n08x5 FILLER_309_24 ();
 b15zdnd00an1n02x5 FILLER_309_32 ();
 b15zdnd11an1n16x5 FILLER_309_39 ();
 b15zdnd11an1n04x5 FILLER_309_55 ();
 b15zdnd00an1n01x5 FILLER_309_59 ();
 b15zdnd11an1n08x5 FILLER_309_66 ();
 b15zdnd00an1n02x5 FILLER_309_74 ();
 b15zdnd11an1n16x5 FILLER_309_88 ();
 b15zdnd00an1n02x5 FILLER_309_104 ();
 b15zdnd00an1n01x5 FILLER_309_106 ();
 b15zdnd11an1n08x5 FILLER_309_110 ();
 b15zdnd00an1n02x5 FILLER_309_118 ();
 b15zdnd00an1n01x5 FILLER_309_120 ();
 b15zdnd11an1n64x5 FILLER_309_124 ();
 b15zdnd11an1n32x5 FILLER_309_188 ();
 b15zdnd11an1n64x5 FILLER_309_223 ();
 b15zdnd11an1n32x5 FILLER_309_287 ();
 b15zdnd11an1n08x5 FILLER_309_319 ();
 b15zdnd11an1n04x5 FILLER_309_327 ();
 b15zdnd00an1n02x5 FILLER_309_331 ();
 b15zdnd00an1n01x5 FILLER_309_333 ();
 b15zdnd11an1n16x5 FILLER_309_342 ();
 b15zdnd00an1n02x5 FILLER_309_358 ();
 b15zdnd11an1n64x5 FILLER_309_400 ();
 b15zdnd11an1n32x5 FILLER_309_464 ();
 b15zdnd11an1n16x5 FILLER_309_496 ();
 b15zdnd11an1n08x5 FILLER_309_512 ();
 b15zdnd11an1n04x5 FILLER_309_520 ();
 b15zdnd00an1n02x5 FILLER_309_524 ();
 b15zdnd00an1n01x5 FILLER_309_526 ();
 b15zdnd11an1n64x5 FILLER_309_530 ();
 b15zdnd11an1n64x5 FILLER_309_594 ();
 b15zdnd11an1n64x5 FILLER_309_658 ();
 b15zdnd11an1n64x5 FILLER_309_722 ();
 b15zdnd11an1n64x5 FILLER_309_786 ();
 b15zdnd11an1n64x5 FILLER_309_850 ();
 b15zdnd11an1n64x5 FILLER_309_914 ();
 b15zdnd11an1n64x5 FILLER_309_978 ();
 b15zdnd11an1n64x5 FILLER_309_1042 ();
 b15zdnd11an1n64x5 FILLER_309_1106 ();
 b15zdnd11an1n64x5 FILLER_309_1170 ();
 b15zdnd11an1n64x5 FILLER_309_1234 ();
 b15zdnd11an1n64x5 FILLER_309_1298 ();
 b15zdnd11an1n64x5 FILLER_309_1362 ();
 b15zdnd11an1n64x5 FILLER_309_1426 ();
 b15zdnd11an1n64x5 FILLER_309_1490 ();
 b15zdnd11an1n64x5 FILLER_309_1554 ();
 b15zdnd11an1n64x5 FILLER_309_1618 ();
 b15zdnd11an1n64x5 FILLER_309_1682 ();
 b15zdnd11an1n64x5 FILLER_309_1746 ();
 b15zdnd11an1n64x5 FILLER_309_1810 ();
 b15zdnd11an1n64x5 FILLER_309_1874 ();
 b15zdnd11an1n64x5 FILLER_309_1938 ();
 b15zdnd11an1n64x5 FILLER_309_2002 ();
 b15zdnd11an1n64x5 FILLER_309_2066 ();
 b15zdnd11an1n64x5 FILLER_309_2130 ();
 b15zdnd11an1n16x5 FILLER_309_2194 ();
 b15zdnd11an1n08x5 FILLER_309_2210 ();
 b15zdnd11an1n04x5 FILLER_309_2218 ();
 b15zdnd11an1n32x5 FILLER_309_2229 ();
 b15zdnd11an1n16x5 FILLER_309_2261 ();
 b15zdnd11an1n04x5 FILLER_309_2277 ();
 b15zdnd00an1n02x5 FILLER_309_2281 ();
 b15zdnd00an1n01x5 FILLER_309_2283 ();
 b15zdnd00an1n02x5 FILLER_310_8 ();
 b15zdnd11an1n04x5 FILLER_310_15 ();
 b15zdnd11an1n08x5 FILLER_310_23 ();
 b15zdnd11an1n16x5 FILLER_310_38 ();
 b15zdnd11an1n08x5 FILLER_310_54 ();
 b15zdnd11an1n64x5 FILLER_310_69 ();
 b15zdnd11an1n64x5 FILLER_310_133 ();
 b15zdnd11an1n64x5 FILLER_310_197 ();
 b15zdnd11an1n64x5 FILLER_310_261 ();
 b15zdnd11an1n32x5 FILLER_310_325 ();
 b15zdnd11an1n04x5 FILLER_310_357 ();
 b15zdnd00an1n01x5 FILLER_310_361 ();
 b15zdnd11an1n16x5 FILLER_310_372 ();
 b15zdnd11an1n04x5 FILLER_310_388 ();
 b15zdnd00an1n02x5 FILLER_310_392 ();
 b15zdnd00an1n01x5 FILLER_310_394 ();
 b15zdnd11an1n64x5 FILLER_310_398 ();
 b15zdnd11an1n16x5 FILLER_310_462 ();
 b15zdnd11an1n08x5 FILLER_310_478 ();
 b15zdnd11an1n04x5 FILLER_310_486 ();
 b15zdnd00an1n01x5 FILLER_310_490 ();
 b15zdnd11an1n64x5 FILLER_310_531 ();
 b15zdnd11an1n64x5 FILLER_310_595 ();
 b15zdnd11an1n32x5 FILLER_310_659 ();
 b15zdnd11an1n16x5 FILLER_310_691 ();
 b15zdnd11an1n08x5 FILLER_310_707 ();
 b15zdnd00an1n02x5 FILLER_310_715 ();
 b15zdnd00an1n01x5 FILLER_310_717 ();
 b15zdnd11an1n64x5 FILLER_310_726 ();
 b15zdnd11an1n64x5 FILLER_310_790 ();
 b15zdnd11an1n64x5 FILLER_310_854 ();
 b15zdnd11an1n64x5 FILLER_310_918 ();
 b15zdnd11an1n64x5 FILLER_310_982 ();
 b15zdnd11an1n64x5 FILLER_310_1046 ();
 b15zdnd11an1n64x5 FILLER_310_1110 ();
 b15zdnd11an1n64x5 FILLER_310_1174 ();
 b15zdnd11an1n64x5 FILLER_310_1238 ();
 b15zdnd11an1n64x5 FILLER_310_1302 ();
 b15zdnd11an1n64x5 FILLER_310_1366 ();
 b15zdnd11an1n64x5 FILLER_310_1430 ();
 b15zdnd11an1n32x5 FILLER_310_1494 ();
 b15zdnd11an1n08x5 FILLER_310_1526 ();
 b15zdnd00an1n02x5 FILLER_310_1534 ();
 b15zdnd11an1n64x5 FILLER_310_1539 ();
 b15zdnd11an1n64x5 FILLER_310_1603 ();
 b15zdnd11an1n64x5 FILLER_310_1667 ();
 b15zdnd11an1n64x5 FILLER_310_1731 ();
 b15zdnd11an1n64x5 FILLER_310_1795 ();
 b15zdnd11an1n64x5 FILLER_310_1859 ();
 b15zdnd11an1n64x5 FILLER_310_1923 ();
 b15zdnd11an1n64x5 FILLER_310_1987 ();
 b15zdnd11an1n64x5 FILLER_310_2051 ();
 b15zdnd11an1n32x5 FILLER_310_2115 ();
 b15zdnd11an1n04x5 FILLER_310_2147 ();
 b15zdnd00an1n02x5 FILLER_310_2151 ();
 b15zdnd00an1n01x5 FILLER_310_2153 ();
 b15zdnd11an1n32x5 FILLER_310_2162 ();
 b15zdnd11an1n16x5 FILLER_310_2194 ();
 b15zdnd11an1n04x5 FILLER_310_2210 ();
 b15zdnd00an1n02x5 FILLER_310_2214 ();
 b15zdnd00an1n01x5 FILLER_310_2216 ();
 b15zdnd11an1n04x5 FILLER_310_2228 ();
 b15zdnd11an1n32x5 FILLER_310_2237 ();
 b15zdnd11an1n04x5 FILLER_310_2269 ();
 b15zdnd00an1n02x5 FILLER_310_2273 ();
 b15zdnd00an1n01x5 FILLER_310_2275 ();
 b15zdnd11an1n64x5 FILLER_311_0 ();
 b15zdnd11an1n64x5 FILLER_311_64 ();
 b15zdnd11an1n64x5 FILLER_311_128 ();
 b15zdnd11an1n32x5 FILLER_311_192 ();
 b15zdnd00an1n01x5 FILLER_311_224 ();
 b15zdnd11an1n64x5 FILLER_311_228 ();
 b15zdnd11an1n64x5 FILLER_311_292 ();
 b15zdnd11an1n64x5 FILLER_311_356 ();
 b15zdnd11an1n64x5 FILLER_311_420 ();
 b15zdnd11an1n32x5 FILLER_311_484 ();
 b15zdnd11an1n08x5 FILLER_311_516 ();
 b15zdnd00an1n02x5 FILLER_311_524 ();
 b15zdnd00an1n01x5 FILLER_311_526 ();
 b15zdnd11an1n64x5 FILLER_311_530 ();
 b15zdnd11an1n64x5 FILLER_311_594 ();
 b15zdnd11an1n64x5 FILLER_311_658 ();
 b15zdnd11an1n64x5 FILLER_311_722 ();
 b15zdnd11an1n64x5 FILLER_311_786 ();
 b15zdnd11an1n64x5 FILLER_311_850 ();
 b15zdnd11an1n64x5 FILLER_311_914 ();
 b15zdnd11an1n64x5 FILLER_311_978 ();
 b15zdnd11an1n64x5 FILLER_311_1042 ();
 b15zdnd11an1n64x5 FILLER_311_1106 ();
 b15zdnd11an1n64x5 FILLER_311_1170 ();
 b15zdnd11an1n64x5 FILLER_311_1234 ();
 b15zdnd11an1n64x5 FILLER_311_1298 ();
 b15zdnd11an1n64x5 FILLER_311_1362 ();
 b15zdnd11an1n64x5 FILLER_311_1426 ();
 b15zdnd11an1n32x5 FILLER_311_1490 ();
 b15zdnd11an1n16x5 FILLER_311_1522 ();
 b15zdnd11an1n08x5 FILLER_311_1538 ();
 b15zdnd11an1n04x5 FILLER_311_1546 ();
 b15zdnd00an1n02x5 FILLER_311_1550 ();
 b15zdnd00an1n01x5 FILLER_311_1552 ();
 b15zdnd11an1n64x5 FILLER_311_1559 ();
 b15zdnd11an1n64x5 FILLER_311_1623 ();
 b15zdnd11an1n64x5 FILLER_311_1687 ();
 b15zdnd11an1n64x5 FILLER_311_1751 ();
 b15zdnd11an1n64x5 FILLER_311_1815 ();
 b15zdnd11an1n04x5 FILLER_311_1879 ();
 b15zdnd00an1n02x5 FILLER_311_1883 ();
 b15zdnd11an1n64x5 FILLER_311_1927 ();
 b15zdnd11an1n64x5 FILLER_311_1991 ();
 b15zdnd11an1n64x5 FILLER_311_2055 ();
 b15zdnd11an1n64x5 FILLER_311_2119 ();
 b15zdnd11an1n32x5 FILLER_311_2183 ();
 b15zdnd11an1n04x5 FILLER_311_2215 ();
 b15zdnd00an1n02x5 FILLER_311_2219 ();
 b15zdnd00an1n01x5 FILLER_311_2221 ();
 b15zdnd11an1n04x5 FILLER_311_2227 ();
 b15zdnd00an1n01x5 FILLER_311_2231 ();
 b15zdnd11an1n32x5 FILLER_311_2236 ();
 b15zdnd11an1n16x5 FILLER_311_2268 ();
 b15zdnd11an1n32x5 FILLER_312_8 ();
 b15zdnd11an1n16x5 FILLER_312_40 ();
 b15zdnd00an1n02x5 FILLER_312_56 ();
 b15zdnd00an1n01x5 FILLER_312_58 ();
 b15zdnd11an1n64x5 FILLER_312_68 ();
 b15zdnd11an1n32x5 FILLER_312_132 ();
 b15zdnd11an1n16x5 FILLER_312_164 ();
 b15zdnd11an1n08x5 FILLER_312_180 ();
 b15zdnd00an1n01x5 FILLER_312_188 ();
 b15zdnd11an1n64x5 FILLER_312_229 ();
 b15zdnd11an1n64x5 FILLER_312_293 ();
 b15zdnd11an1n64x5 FILLER_312_357 ();
 b15zdnd11an1n64x5 FILLER_312_421 ();
 b15zdnd11an1n64x5 FILLER_312_485 ();
 b15zdnd11an1n64x5 FILLER_312_549 ();
 b15zdnd11an1n64x5 FILLER_312_613 ();
 b15zdnd11an1n32x5 FILLER_312_677 ();
 b15zdnd11an1n08x5 FILLER_312_709 ();
 b15zdnd00an1n01x5 FILLER_312_717 ();
 b15zdnd11an1n64x5 FILLER_312_726 ();
 b15zdnd11an1n64x5 FILLER_312_790 ();
 b15zdnd11an1n64x5 FILLER_312_854 ();
 b15zdnd11an1n64x5 FILLER_312_918 ();
 b15zdnd11an1n64x5 FILLER_312_982 ();
 b15zdnd11an1n64x5 FILLER_312_1046 ();
 b15zdnd11an1n64x5 FILLER_312_1110 ();
 b15zdnd11an1n64x5 FILLER_312_1174 ();
 b15zdnd11an1n64x5 FILLER_312_1238 ();
 b15zdnd11an1n64x5 FILLER_312_1302 ();
 b15zdnd11an1n64x5 FILLER_312_1366 ();
 b15zdnd11an1n64x5 FILLER_312_1430 ();
 b15zdnd11an1n64x5 FILLER_312_1494 ();
 b15zdnd11an1n08x5 FILLER_312_1558 ();
 b15zdnd11an1n04x5 FILLER_312_1566 ();
 b15zdnd11an1n64x5 FILLER_312_1612 ();
 b15zdnd11an1n64x5 FILLER_312_1676 ();
 b15zdnd11an1n64x5 FILLER_312_1740 ();
 b15zdnd11an1n32x5 FILLER_312_1804 ();
 b15zdnd11an1n16x5 FILLER_312_1836 ();
 b15zdnd11an1n08x5 FILLER_312_1852 ();
 b15zdnd00an1n02x5 FILLER_312_1860 ();
 b15zdnd11an1n64x5 FILLER_312_1865 ();
 b15zdnd11an1n64x5 FILLER_312_1929 ();
 b15zdnd11an1n64x5 FILLER_312_1993 ();
 b15zdnd11an1n64x5 FILLER_312_2057 ();
 b15zdnd11an1n32x5 FILLER_312_2121 ();
 b15zdnd00an1n01x5 FILLER_312_2153 ();
 b15zdnd11an1n64x5 FILLER_312_2162 ();
 b15zdnd11an1n32x5 FILLER_312_2226 ();
 b15zdnd11an1n16x5 FILLER_312_2258 ();
 b15zdnd00an1n02x5 FILLER_312_2274 ();
 b15zdnd11an1n64x5 FILLER_313_0 ();
 b15zdnd11an1n64x5 FILLER_313_64 ();
 b15zdnd11an1n64x5 FILLER_313_128 ();
 b15zdnd11an1n32x5 FILLER_313_192 ();
 b15zdnd00an1n02x5 FILLER_313_224 ();
 b15zdnd00an1n01x5 FILLER_313_226 ();
 b15zdnd11an1n64x5 FILLER_313_230 ();
 b15zdnd11an1n64x5 FILLER_313_294 ();
 b15zdnd11an1n64x5 FILLER_313_358 ();
 b15zdnd11an1n64x5 FILLER_313_422 ();
 b15zdnd11an1n64x5 FILLER_313_486 ();
 b15zdnd11an1n64x5 FILLER_313_550 ();
 b15zdnd11an1n64x5 FILLER_313_614 ();
 b15zdnd11an1n64x5 FILLER_313_678 ();
 b15zdnd11an1n64x5 FILLER_313_742 ();
 b15zdnd11an1n64x5 FILLER_313_806 ();
 b15zdnd11an1n64x5 FILLER_313_870 ();
 b15zdnd11an1n64x5 FILLER_313_934 ();
 b15zdnd11an1n64x5 FILLER_313_998 ();
 b15zdnd11an1n64x5 FILLER_313_1062 ();
 b15zdnd11an1n64x5 FILLER_313_1126 ();
 b15zdnd11an1n64x5 FILLER_313_1190 ();
 b15zdnd11an1n64x5 FILLER_313_1254 ();
 b15zdnd11an1n64x5 FILLER_313_1318 ();
 b15zdnd11an1n64x5 FILLER_313_1382 ();
 b15zdnd11an1n64x5 FILLER_313_1446 ();
 b15zdnd11an1n32x5 FILLER_313_1510 ();
 b15zdnd11an1n16x5 FILLER_313_1542 ();
 b15zdnd00an1n01x5 FILLER_313_1558 ();
 b15zdnd11an1n04x5 FILLER_313_1601 ();
 b15zdnd11an1n64x5 FILLER_313_1636 ();
 b15zdnd11an1n64x5 FILLER_313_1700 ();
 b15zdnd11an1n64x5 FILLER_313_1764 ();
 b15zdnd11an1n32x5 FILLER_313_1828 ();
 b15zdnd00an1n01x5 FILLER_313_1860 ();
 b15zdnd11an1n64x5 FILLER_313_1864 ();
 b15zdnd11an1n64x5 FILLER_313_1928 ();
 b15zdnd11an1n64x5 FILLER_313_1992 ();
 b15zdnd11an1n64x5 FILLER_313_2056 ();
 b15zdnd11an1n64x5 FILLER_313_2120 ();
 b15zdnd11an1n32x5 FILLER_313_2184 ();
 b15zdnd11an1n04x5 FILLER_313_2216 ();
 b15zdnd11an1n16x5 FILLER_313_2262 ();
 b15zdnd11an1n04x5 FILLER_313_2278 ();
 b15zdnd00an1n02x5 FILLER_313_2282 ();
 b15zdnd11an1n64x5 FILLER_314_8 ();
 b15zdnd11an1n64x5 FILLER_314_72 ();
 b15zdnd11an1n64x5 FILLER_314_136 ();
 b15zdnd11an1n64x5 FILLER_314_200 ();
 b15zdnd11an1n64x5 FILLER_314_264 ();
 b15zdnd11an1n64x5 FILLER_314_328 ();
 b15zdnd11an1n64x5 FILLER_314_392 ();
 b15zdnd11an1n32x5 FILLER_314_456 ();
 b15zdnd11an1n04x5 FILLER_314_488 ();
 b15zdnd11an1n64x5 FILLER_314_501 ();
 b15zdnd11an1n64x5 FILLER_314_565 ();
 b15zdnd11an1n64x5 FILLER_314_629 ();
 b15zdnd11an1n16x5 FILLER_314_693 ();
 b15zdnd11an1n08x5 FILLER_314_709 ();
 b15zdnd00an1n01x5 FILLER_314_717 ();
 b15zdnd11an1n64x5 FILLER_314_726 ();
 b15zdnd11an1n64x5 FILLER_314_790 ();
 b15zdnd11an1n64x5 FILLER_314_854 ();
 b15zdnd11an1n64x5 FILLER_314_918 ();
 b15zdnd11an1n64x5 FILLER_314_982 ();
 b15zdnd11an1n64x5 FILLER_314_1046 ();
 b15zdnd11an1n64x5 FILLER_314_1110 ();
 b15zdnd11an1n64x5 FILLER_314_1174 ();
 b15zdnd11an1n64x5 FILLER_314_1238 ();
 b15zdnd11an1n64x5 FILLER_314_1302 ();
 b15zdnd11an1n64x5 FILLER_314_1366 ();
 b15zdnd11an1n64x5 FILLER_314_1430 ();
 b15zdnd11an1n64x5 FILLER_314_1494 ();
 b15zdnd11an1n04x5 FILLER_314_1558 ();
 b15zdnd11an1n64x5 FILLER_314_1614 ();
 b15zdnd11an1n64x5 FILLER_314_1678 ();
 b15zdnd11an1n64x5 FILLER_314_1742 ();
 b15zdnd11an1n16x5 FILLER_314_1806 ();
 b15zdnd11an1n08x5 FILLER_314_1822 ();
 b15zdnd11an1n04x5 FILLER_314_1830 ();
 b15zdnd00an1n02x5 FILLER_314_1834 ();
 b15zdnd11an1n64x5 FILLER_314_1888 ();
 b15zdnd11an1n64x5 FILLER_314_1952 ();
 b15zdnd11an1n64x5 FILLER_314_2016 ();
 b15zdnd11an1n64x5 FILLER_314_2080 ();
 b15zdnd11an1n08x5 FILLER_314_2144 ();
 b15zdnd00an1n02x5 FILLER_314_2152 ();
 b15zdnd11an1n64x5 FILLER_314_2162 ();
 b15zdnd11an1n32x5 FILLER_314_2226 ();
 b15zdnd11an1n16x5 FILLER_314_2258 ();
 b15zdnd00an1n02x5 FILLER_314_2274 ();
 b15zdnd11an1n64x5 FILLER_315_0 ();
 b15zdnd11an1n64x5 FILLER_315_68 ();
 b15zdnd11an1n64x5 FILLER_315_132 ();
 b15zdnd11an1n64x5 FILLER_315_196 ();
 b15zdnd11an1n64x5 FILLER_315_260 ();
 b15zdnd11an1n04x5 FILLER_315_324 ();
 b15zdnd00an1n02x5 FILLER_315_328 ();
 b15zdnd11an1n64x5 FILLER_315_338 ();
 b15zdnd11an1n64x5 FILLER_315_402 ();
 b15zdnd11an1n64x5 FILLER_315_466 ();
 b15zdnd11an1n64x5 FILLER_315_530 ();
 b15zdnd11an1n64x5 FILLER_315_594 ();
 b15zdnd11an1n64x5 FILLER_315_658 ();
 b15zdnd11an1n64x5 FILLER_315_722 ();
 b15zdnd11an1n64x5 FILLER_315_786 ();
 b15zdnd11an1n64x5 FILLER_315_850 ();
 b15zdnd11an1n64x5 FILLER_315_914 ();
 b15zdnd11an1n64x5 FILLER_315_978 ();
 b15zdnd11an1n64x5 FILLER_315_1042 ();
 b15zdnd11an1n32x5 FILLER_315_1106 ();
 b15zdnd11an1n04x5 FILLER_315_1138 ();
 b15zdnd00an1n02x5 FILLER_315_1142 ();
 b15zdnd11an1n64x5 FILLER_315_1196 ();
 b15zdnd11an1n64x5 FILLER_315_1260 ();
 b15zdnd11an1n64x5 FILLER_315_1324 ();
 b15zdnd11an1n64x5 FILLER_315_1388 ();
 b15zdnd11an1n64x5 FILLER_315_1452 ();
 b15zdnd11an1n32x5 FILLER_315_1516 ();
 b15zdnd11an1n16x5 FILLER_315_1548 ();
 b15zdnd11an1n08x5 FILLER_315_1564 ();
 b15zdnd11an1n04x5 FILLER_315_1572 ();
 b15zdnd00an1n02x5 FILLER_315_1576 ();
 b15zdnd11an1n04x5 FILLER_315_1581 ();
 b15zdnd11an1n64x5 FILLER_315_1588 ();
 b15zdnd11an1n64x5 FILLER_315_1652 ();
 b15zdnd11an1n64x5 FILLER_315_1716 ();
 b15zdnd11an1n64x5 FILLER_315_1780 ();
 b15zdnd11an1n16x5 FILLER_315_1844 ();
 b15zdnd00an1n01x5 FILLER_315_1860 ();
 b15zdnd11an1n64x5 FILLER_315_1864 ();
 b15zdnd11an1n32x5 FILLER_315_1928 ();
 b15zdnd11an1n08x5 FILLER_315_1960 ();
 b15zdnd11an1n64x5 FILLER_315_1978 ();
 b15zdnd11an1n64x5 FILLER_315_2042 ();
 b15zdnd11an1n64x5 FILLER_315_2106 ();
 b15zdnd11an1n32x5 FILLER_315_2170 ();
 b15zdnd11an1n08x5 FILLER_315_2202 ();
 b15zdnd11an1n64x5 FILLER_315_2213 ();
 b15zdnd11an1n04x5 FILLER_315_2277 ();
 b15zdnd00an1n02x5 FILLER_315_2281 ();
 b15zdnd00an1n01x5 FILLER_315_2283 ();
 b15zdnd11an1n32x5 FILLER_316_8 ();
 b15zdnd11an1n16x5 FILLER_316_40 ();
 b15zdnd11an1n04x5 FILLER_316_56 ();
 b15zdnd00an1n02x5 FILLER_316_60 ();
 b15zdnd11an1n64x5 FILLER_316_70 ();
 b15zdnd11an1n64x5 FILLER_316_134 ();
 b15zdnd11an1n64x5 FILLER_316_198 ();
 b15zdnd11an1n64x5 FILLER_316_262 ();
 b15zdnd11an1n64x5 FILLER_316_326 ();
 b15zdnd11an1n64x5 FILLER_316_390 ();
 b15zdnd11an1n64x5 FILLER_316_454 ();
 b15zdnd11an1n64x5 FILLER_316_518 ();
 b15zdnd11an1n64x5 FILLER_316_582 ();
 b15zdnd11an1n64x5 FILLER_316_646 ();
 b15zdnd11an1n08x5 FILLER_316_710 ();
 b15zdnd11an1n64x5 FILLER_316_726 ();
 b15zdnd11an1n64x5 FILLER_316_790 ();
 b15zdnd11an1n64x5 FILLER_316_854 ();
 b15zdnd11an1n64x5 FILLER_316_918 ();
 b15zdnd11an1n64x5 FILLER_316_982 ();
 b15zdnd11an1n64x5 FILLER_316_1046 ();
 b15zdnd11an1n32x5 FILLER_316_1110 ();
 b15zdnd11an1n08x5 FILLER_316_1142 ();
 b15zdnd00an1n02x5 FILLER_316_1150 ();
 b15zdnd00an1n01x5 FILLER_316_1152 ();
 b15zdnd11an1n64x5 FILLER_316_1205 ();
 b15zdnd11an1n16x5 FILLER_316_1269 ();
 b15zdnd11an1n04x5 FILLER_316_1285 ();
 b15zdnd00an1n02x5 FILLER_316_1289 ();
 b15zdnd00an1n01x5 FILLER_316_1291 ();
 b15zdnd11an1n64x5 FILLER_316_1295 ();
 b15zdnd11an1n64x5 FILLER_316_1359 ();
 b15zdnd11an1n64x5 FILLER_316_1423 ();
 b15zdnd11an1n64x5 FILLER_316_1487 ();
 b15zdnd11an1n32x5 FILLER_316_1551 ();
 b15zdnd00an1n02x5 FILLER_316_1583 ();
 b15zdnd00an1n01x5 FILLER_316_1585 ();
 b15zdnd11an1n64x5 FILLER_316_1589 ();
 b15zdnd11an1n64x5 FILLER_316_1653 ();
 b15zdnd11an1n64x5 FILLER_316_1717 ();
 b15zdnd11an1n64x5 FILLER_316_1781 ();
 b15zdnd11an1n64x5 FILLER_316_1845 ();
 b15zdnd11an1n64x5 FILLER_316_1909 ();
 b15zdnd11an1n64x5 FILLER_316_1973 ();
 b15zdnd11an1n64x5 FILLER_316_2037 ();
 b15zdnd11an1n32x5 FILLER_316_2101 ();
 b15zdnd11an1n16x5 FILLER_316_2133 ();
 b15zdnd11an1n04x5 FILLER_316_2149 ();
 b15zdnd00an1n01x5 FILLER_316_2153 ();
 b15zdnd11an1n32x5 FILLER_316_2162 ();
 b15zdnd11an1n16x5 FILLER_316_2194 ();
 b15zdnd00an1n01x5 FILLER_316_2210 ();
 b15zdnd11an1n32x5 FILLER_316_2214 ();
 b15zdnd11an1n16x5 FILLER_316_2246 ();
 b15zdnd11an1n08x5 FILLER_316_2262 ();
 b15zdnd11an1n04x5 FILLER_316_2270 ();
 b15zdnd00an1n02x5 FILLER_316_2274 ();
 b15zdnd11an1n64x5 FILLER_317_0 ();
 b15zdnd11an1n08x5 FILLER_317_64 ();
 b15zdnd11an1n04x5 FILLER_317_72 ();
 b15zdnd11an1n64x5 FILLER_317_80 ();
 b15zdnd11an1n64x5 FILLER_317_144 ();
 b15zdnd11an1n64x5 FILLER_317_208 ();
 b15zdnd11an1n64x5 FILLER_317_272 ();
 b15zdnd11an1n64x5 FILLER_317_336 ();
 b15zdnd11an1n64x5 FILLER_317_400 ();
 b15zdnd11an1n64x5 FILLER_317_464 ();
 b15zdnd11an1n64x5 FILLER_317_528 ();
 b15zdnd11an1n64x5 FILLER_317_592 ();
 b15zdnd11an1n64x5 FILLER_317_656 ();
 b15zdnd11an1n64x5 FILLER_317_720 ();
 b15zdnd11an1n64x5 FILLER_317_784 ();
 b15zdnd11an1n64x5 FILLER_317_848 ();
 b15zdnd11an1n64x5 FILLER_317_912 ();
 b15zdnd11an1n64x5 FILLER_317_976 ();
 b15zdnd11an1n64x5 FILLER_317_1040 ();
 b15zdnd11an1n32x5 FILLER_317_1104 ();
 b15zdnd11an1n16x5 FILLER_317_1136 ();
 b15zdnd11an1n08x5 FILLER_317_1152 ();
 b15zdnd00an1n02x5 FILLER_317_1160 ();
 b15zdnd11an1n04x5 FILLER_317_1165 ();
 b15zdnd11an1n04x5 FILLER_317_1172 ();
 b15zdnd11an1n04x5 FILLER_317_1179 ();
 b15zdnd11an1n08x5 FILLER_317_1186 ();
 b15zdnd11an1n04x5 FILLER_317_1194 ();
 b15zdnd00an1n02x5 FILLER_317_1198 ();
 b15zdnd11an1n32x5 FILLER_317_1242 ();
 b15zdnd11an1n16x5 FILLER_317_1274 ();
 b15zdnd00an1n01x5 FILLER_317_1290 ();
 b15zdnd11an1n64x5 FILLER_317_1294 ();
 b15zdnd11an1n64x5 FILLER_317_1358 ();
 b15zdnd11an1n64x5 FILLER_317_1422 ();
 b15zdnd11an1n64x5 FILLER_317_1486 ();
 b15zdnd11an1n64x5 FILLER_317_1550 ();
 b15zdnd11an1n64x5 FILLER_317_1614 ();
 b15zdnd11an1n64x5 FILLER_317_1678 ();
 b15zdnd11an1n64x5 FILLER_317_1742 ();
 b15zdnd11an1n64x5 FILLER_317_1806 ();
 b15zdnd11an1n64x5 FILLER_317_1870 ();
 b15zdnd11an1n64x5 FILLER_317_1934 ();
 b15zdnd11an1n64x5 FILLER_317_1998 ();
 b15zdnd11an1n64x5 FILLER_317_2062 ();
 b15zdnd11an1n32x5 FILLER_317_2126 ();
 b15zdnd11an1n16x5 FILLER_317_2158 ();
 b15zdnd11an1n08x5 FILLER_317_2174 ();
 b15zdnd11an1n04x5 FILLER_317_2182 ();
 b15zdnd11an1n32x5 FILLER_317_2238 ();
 b15zdnd11an1n08x5 FILLER_317_2270 ();
 b15zdnd11an1n04x5 FILLER_317_2278 ();
 b15zdnd00an1n02x5 FILLER_317_2282 ();
 b15zdnd11an1n64x5 FILLER_318_8 ();
 b15zdnd11an1n64x5 FILLER_318_72 ();
 b15zdnd11an1n64x5 FILLER_318_136 ();
 b15zdnd11an1n64x5 FILLER_318_200 ();
 b15zdnd11an1n64x5 FILLER_318_264 ();
 b15zdnd11an1n64x5 FILLER_318_328 ();
 b15zdnd11an1n64x5 FILLER_318_392 ();
 b15zdnd11an1n64x5 FILLER_318_456 ();
 b15zdnd11an1n64x5 FILLER_318_520 ();
 b15zdnd11an1n64x5 FILLER_318_584 ();
 b15zdnd11an1n64x5 FILLER_318_648 ();
 b15zdnd11an1n04x5 FILLER_318_712 ();
 b15zdnd00an1n02x5 FILLER_318_716 ();
 b15zdnd11an1n64x5 FILLER_318_726 ();
 b15zdnd11an1n64x5 FILLER_318_790 ();
 b15zdnd11an1n64x5 FILLER_318_854 ();
 b15zdnd11an1n64x5 FILLER_318_918 ();
 b15zdnd11an1n64x5 FILLER_318_982 ();
 b15zdnd11an1n64x5 FILLER_318_1046 ();
 b15zdnd11an1n32x5 FILLER_318_1110 ();
 b15zdnd11an1n16x5 FILLER_318_1142 ();
 b15zdnd11an1n08x5 FILLER_318_1158 ();
 b15zdnd00an1n02x5 FILLER_318_1166 ();
 b15zdnd00an1n01x5 FILLER_318_1168 ();
 b15zdnd11an1n04x5 FILLER_318_1172 ();
 b15zdnd11an1n16x5 FILLER_318_1179 ();
 b15zdnd11an1n32x5 FILLER_318_1203 ();
 b15zdnd11an1n16x5 FILLER_318_1235 ();
 b15zdnd11an1n08x5 FILLER_318_1251 ();
 b15zdnd11an1n04x5 FILLER_318_1259 ();
 b15zdnd00an1n02x5 FILLER_318_1263 ();
 b15zdnd00an1n01x5 FILLER_318_1265 ();
 b15zdnd11an1n64x5 FILLER_318_1318 ();
 b15zdnd11an1n64x5 FILLER_318_1382 ();
 b15zdnd11an1n64x5 FILLER_318_1446 ();
 b15zdnd11an1n64x5 FILLER_318_1510 ();
 b15zdnd11an1n64x5 FILLER_318_1574 ();
 b15zdnd11an1n64x5 FILLER_318_1638 ();
 b15zdnd11an1n64x5 FILLER_318_1702 ();
 b15zdnd11an1n64x5 FILLER_318_1766 ();
 b15zdnd11an1n64x5 FILLER_318_1830 ();
 b15zdnd11an1n64x5 FILLER_318_1894 ();
 b15zdnd11an1n64x5 FILLER_318_1958 ();
 b15zdnd11an1n64x5 FILLER_318_2022 ();
 b15zdnd11an1n64x5 FILLER_318_2086 ();
 b15zdnd11an1n04x5 FILLER_318_2150 ();
 b15zdnd11an1n32x5 FILLER_318_2162 ();
 b15zdnd11an1n16x5 FILLER_318_2194 ();
 b15zdnd00an1n02x5 FILLER_318_2210 ();
 b15zdnd11an1n32x5 FILLER_318_2215 ();
 b15zdnd11an1n16x5 FILLER_318_2247 ();
 b15zdnd11an1n08x5 FILLER_318_2263 ();
 b15zdnd11an1n04x5 FILLER_318_2271 ();
 b15zdnd00an1n01x5 FILLER_318_2275 ();
 b15zdnd11an1n32x5 FILLER_319_0 ();
 b15zdnd11an1n04x5 FILLER_319_32 ();
 b15zdnd00an1n01x5 FILLER_319_36 ();
 b15zdnd11an1n64x5 FILLER_319_43 ();
 b15zdnd11an1n64x5 FILLER_319_107 ();
 b15zdnd11an1n64x5 FILLER_319_171 ();
 b15zdnd11an1n64x5 FILLER_319_235 ();
 b15zdnd11an1n64x5 FILLER_319_299 ();
 b15zdnd11an1n64x5 FILLER_319_363 ();
 b15zdnd11an1n64x5 FILLER_319_427 ();
 b15zdnd11an1n64x5 FILLER_319_491 ();
 b15zdnd11an1n64x5 FILLER_319_555 ();
 b15zdnd11an1n64x5 FILLER_319_619 ();
 b15zdnd11an1n64x5 FILLER_319_683 ();
 b15zdnd11an1n64x5 FILLER_319_747 ();
 b15zdnd11an1n64x5 FILLER_319_811 ();
 b15zdnd11an1n64x5 FILLER_319_875 ();
 b15zdnd11an1n64x5 FILLER_319_939 ();
 b15zdnd11an1n64x5 FILLER_319_1003 ();
 b15zdnd11an1n64x5 FILLER_319_1067 ();
 b15zdnd11an1n16x5 FILLER_319_1131 ();
 b15zdnd00an1n02x5 FILLER_319_1147 ();
 b15zdnd00an1n01x5 FILLER_319_1149 ();
 b15zdnd11an1n04x5 FILLER_319_1153 ();
 b15zdnd11an1n64x5 FILLER_319_1184 ();
 b15zdnd11an1n16x5 FILLER_319_1248 ();
 b15zdnd11an1n04x5 FILLER_319_1264 ();
 b15zdnd11an1n64x5 FILLER_319_1320 ();
 b15zdnd11an1n64x5 FILLER_319_1384 ();
 b15zdnd11an1n64x5 FILLER_319_1448 ();
 b15zdnd11an1n64x5 FILLER_319_1512 ();
 b15zdnd11an1n64x5 FILLER_319_1576 ();
 b15zdnd11an1n64x5 FILLER_319_1640 ();
 b15zdnd11an1n64x5 FILLER_319_1704 ();
 b15zdnd11an1n64x5 FILLER_319_1768 ();
 b15zdnd11an1n64x5 FILLER_319_1832 ();
 b15zdnd11an1n64x5 FILLER_319_1896 ();
 b15zdnd11an1n64x5 FILLER_319_1960 ();
 b15zdnd11an1n64x5 FILLER_319_2024 ();
 b15zdnd11an1n64x5 FILLER_319_2088 ();
 b15zdnd11an1n64x5 FILLER_319_2152 ();
 b15zdnd11an1n64x5 FILLER_319_2216 ();
 b15zdnd11an1n04x5 FILLER_319_2280 ();
 b15zdnd11an1n16x5 FILLER_320_8 ();
 b15zdnd11an1n04x5 FILLER_320_24 ();
 b15zdnd00an1n02x5 FILLER_320_28 ();
 b15zdnd00an1n01x5 FILLER_320_30 ();
 b15zdnd11an1n32x5 FILLER_320_36 ();
 b15zdnd11an1n04x5 FILLER_320_68 ();
 b15zdnd00an1n02x5 FILLER_320_72 ();
 b15zdnd11an1n64x5 FILLER_320_80 ();
 b15zdnd11an1n64x5 FILLER_320_144 ();
 b15zdnd11an1n64x5 FILLER_320_208 ();
 b15zdnd11an1n64x5 FILLER_320_272 ();
 b15zdnd11an1n64x5 FILLER_320_336 ();
 b15zdnd11an1n64x5 FILLER_320_400 ();
 b15zdnd11an1n64x5 FILLER_320_464 ();
 b15zdnd11an1n64x5 FILLER_320_528 ();
 b15zdnd11an1n64x5 FILLER_320_592 ();
 b15zdnd11an1n32x5 FILLER_320_656 ();
 b15zdnd11an1n16x5 FILLER_320_688 ();
 b15zdnd11an1n08x5 FILLER_320_704 ();
 b15zdnd11an1n04x5 FILLER_320_712 ();
 b15zdnd00an1n02x5 FILLER_320_716 ();
 b15zdnd11an1n64x5 FILLER_320_726 ();
 b15zdnd11an1n64x5 FILLER_320_790 ();
 b15zdnd11an1n64x5 FILLER_320_854 ();
 b15zdnd11an1n64x5 FILLER_320_918 ();
 b15zdnd11an1n64x5 FILLER_320_982 ();
 b15zdnd11an1n64x5 FILLER_320_1046 ();
 b15zdnd11an1n64x5 FILLER_320_1110 ();
 b15zdnd11an1n64x5 FILLER_320_1174 ();
 b15zdnd11an1n32x5 FILLER_320_1238 ();
 b15zdnd11an1n08x5 FILLER_320_1270 ();
 b15zdnd11an1n04x5 FILLER_320_1278 ();
 b15zdnd00an1n02x5 FILLER_320_1282 ();
 b15zdnd00an1n01x5 FILLER_320_1284 ();
 b15zdnd11an1n04x5 FILLER_320_1288 ();
 b15zdnd11an1n04x5 FILLER_320_1295 ();
 b15zdnd11an1n04x5 FILLER_320_1302 ();
 b15zdnd11an1n04x5 FILLER_320_1309 ();
 b15zdnd11an1n64x5 FILLER_320_1316 ();
 b15zdnd11an1n64x5 FILLER_320_1380 ();
 b15zdnd11an1n64x5 FILLER_320_1444 ();
 b15zdnd11an1n64x5 FILLER_320_1508 ();
 b15zdnd11an1n64x5 FILLER_320_1572 ();
 b15zdnd11an1n64x5 FILLER_320_1636 ();
 b15zdnd11an1n64x5 FILLER_320_1700 ();
 b15zdnd11an1n64x5 FILLER_320_1764 ();
 b15zdnd11an1n64x5 FILLER_320_1828 ();
 b15zdnd11an1n64x5 FILLER_320_1892 ();
 b15zdnd11an1n64x5 FILLER_320_1956 ();
 b15zdnd11an1n64x5 FILLER_320_2020 ();
 b15zdnd11an1n64x5 FILLER_320_2084 ();
 b15zdnd11an1n04x5 FILLER_320_2148 ();
 b15zdnd00an1n02x5 FILLER_320_2152 ();
 b15zdnd11an1n64x5 FILLER_320_2162 ();
 b15zdnd11an1n32x5 FILLER_320_2226 ();
 b15zdnd11an1n16x5 FILLER_320_2258 ();
 b15zdnd00an1n02x5 FILLER_320_2274 ();
 b15zdnd11an1n64x5 FILLER_321_0 ();
 b15zdnd11an1n64x5 FILLER_321_64 ();
 b15zdnd11an1n64x5 FILLER_321_128 ();
 b15zdnd11an1n64x5 FILLER_321_192 ();
 b15zdnd11an1n64x5 FILLER_321_256 ();
 b15zdnd11an1n64x5 FILLER_321_320 ();
 b15zdnd11an1n64x5 FILLER_321_384 ();
 b15zdnd11an1n64x5 FILLER_321_448 ();
 b15zdnd11an1n64x5 FILLER_321_512 ();
 b15zdnd11an1n64x5 FILLER_321_576 ();
 b15zdnd11an1n64x5 FILLER_321_640 ();
 b15zdnd11an1n32x5 FILLER_321_704 ();
 b15zdnd11an1n16x5 FILLER_321_736 ();
 b15zdnd11an1n08x5 FILLER_321_752 ();
 b15zdnd11an1n04x5 FILLER_321_760 ();
 b15zdnd00an1n02x5 FILLER_321_764 ();
 b15zdnd11an1n64x5 FILLER_321_775 ();
 b15zdnd11an1n64x5 FILLER_321_839 ();
 b15zdnd11an1n64x5 FILLER_321_903 ();
 b15zdnd11an1n64x5 FILLER_321_967 ();
 b15zdnd11an1n64x5 FILLER_321_1031 ();
 b15zdnd11an1n64x5 FILLER_321_1095 ();
 b15zdnd11an1n16x5 FILLER_321_1159 ();
 b15zdnd11an1n04x5 FILLER_321_1175 ();
 b15zdnd00an1n02x5 FILLER_321_1179 ();
 b15zdnd00an1n01x5 FILLER_321_1181 ();
 b15zdnd11an1n32x5 FILLER_321_1191 ();
 b15zdnd11an1n08x5 FILLER_321_1223 ();
 b15zdnd11an1n04x5 FILLER_321_1231 ();
 b15zdnd00an1n02x5 FILLER_321_1235 ();
 b15zdnd00an1n01x5 FILLER_321_1237 ();
 b15zdnd11an1n16x5 FILLER_321_1247 ();
 b15zdnd11an1n04x5 FILLER_321_1263 ();
 b15zdnd00an1n01x5 FILLER_321_1267 ();
 b15zdnd11an1n64x5 FILLER_321_1320 ();
 b15zdnd11an1n64x5 FILLER_321_1384 ();
 b15zdnd11an1n64x5 FILLER_321_1448 ();
 b15zdnd11an1n64x5 FILLER_321_1512 ();
 b15zdnd11an1n64x5 FILLER_321_1576 ();
 b15zdnd11an1n64x5 FILLER_321_1640 ();
 b15zdnd11an1n64x5 FILLER_321_1704 ();
 b15zdnd11an1n64x5 FILLER_321_1768 ();
 b15zdnd11an1n64x5 FILLER_321_1832 ();
 b15zdnd11an1n64x5 FILLER_321_1896 ();
 b15zdnd00an1n01x5 FILLER_321_1960 ();
 b15zdnd11an1n64x5 FILLER_321_1965 ();
 b15zdnd11an1n64x5 FILLER_321_2029 ();
 b15zdnd11an1n64x5 FILLER_321_2093 ();
 b15zdnd11an1n64x5 FILLER_321_2157 ();
 b15zdnd11an1n32x5 FILLER_321_2221 ();
 b15zdnd11an1n16x5 FILLER_321_2253 ();
 b15zdnd11an1n08x5 FILLER_321_2269 ();
 b15zdnd11an1n04x5 FILLER_321_2277 ();
 b15zdnd00an1n02x5 FILLER_321_2281 ();
 b15zdnd00an1n01x5 FILLER_321_2283 ();
 b15zdnd11an1n32x5 FILLER_322_8 ();
 b15zdnd11an1n16x5 FILLER_322_40 ();
 b15zdnd11an1n04x5 FILLER_322_56 ();
 b15zdnd00an1n02x5 FILLER_322_60 ();
 b15zdnd00an1n01x5 FILLER_322_62 ();
 b15zdnd11an1n64x5 FILLER_322_75 ();
 b15zdnd11an1n64x5 FILLER_322_139 ();
 b15zdnd11an1n64x5 FILLER_322_203 ();
 b15zdnd11an1n64x5 FILLER_322_267 ();
 b15zdnd11an1n64x5 FILLER_322_331 ();
 b15zdnd11an1n64x5 FILLER_322_395 ();
 b15zdnd11an1n64x5 FILLER_322_459 ();
 b15zdnd11an1n64x5 FILLER_322_523 ();
 b15zdnd11an1n64x5 FILLER_322_587 ();
 b15zdnd11an1n64x5 FILLER_322_651 ();
 b15zdnd00an1n02x5 FILLER_322_715 ();
 b15zdnd00an1n01x5 FILLER_322_717 ();
 b15zdnd11an1n64x5 FILLER_322_726 ();
 b15zdnd11an1n64x5 FILLER_322_790 ();
 b15zdnd11an1n64x5 FILLER_322_854 ();
 b15zdnd11an1n64x5 FILLER_322_918 ();
 b15zdnd11an1n64x5 FILLER_322_982 ();
 b15zdnd11an1n64x5 FILLER_322_1046 ();
 b15zdnd11an1n64x5 FILLER_322_1110 ();
 b15zdnd11an1n32x5 FILLER_322_1174 ();
 b15zdnd11an1n16x5 FILLER_322_1206 ();
 b15zdnd11an1n08x5 FILLER_322_1222 ();
 b15zdnd00an1n02x5 FILLER_322_1230 ();
 b15zdnd11an1n16x5 FILLER_322_1241 ();
 b15zdnd11an1n08x5 FILLER_322_1257 ();
 b15zdnd00an1n02x5 FILLER_322_1265 ();
 b15zdnd00an1n01x5 FILLER_322_1267 ();
 b15zdnd11an1n64x5 FILLER_322_1320 ();
 b15zdnd11an1n64x5 FILLER_322_1384 ();
 b15zdnd11an1n64x5 FILLER_322_1448 ();
 b15zdnd11an1n64x5 FILLER_322_1512 ();
 b15zdnd11an1n64x5 FILLER_322_1576 ();
 b15zdnd11an1n64x5 FILLER_322_1640 ();
 b15zdnd11an1n64x5 FILLER_322_1704 ();
 b15zdnd11an1n08x5 FILLER_322_1768 ();
 b15zdnd11an1n64x5 FILLER_322_1818 ();
 b15zdnd11an1n64x5 FILLER_322_1882 ();
 b15zdnd11an1n08x5 FILLER_322_1946 ();
 b15zdnd11an1n04x5 FILLER_322_1954 ();
 b15zdnd00an1n01x5 FILLER_322_1958 ();
 b15zdnd11an1n64x5 FILLER_322_1966 ();
 b15zdnd11an1n64x5 FILLER_322_2030 ();
 b15zdnd11an1n32x5 FILLER_322_2094 ();
 b15zdnd11an1n16x5 FILLER_322_2126 ();
 b15zdnd11an1n08x5 FILLER_322_2142 ();
 b15zdnd11an1n04x5 FILLER_322_2150 ();
 b15zdnd11an1n64x5 FILLER_322_2162 ();
 b15zdnd11an1n32x5 FILLER_322_2226 ();
 b15zdnd11an1n16x5 FILLER_322_2258 ();
 b15zdnd00an1n02x5 FILLER_322_2274 ();
 b15zdnd11an1n64x5 FILLER_323_0 ();
 b15zdnd11an1n64x5 FILLER_323_64 ();
 b15zdnd11an1n64x5 FILLER_323_128 ();
 b15zdnd11an1n64x5 FILLER_323_192 ();
 b15zdnd11an1n64x5 FILLER_323_256 ();
 b15zdnd11an1n64x5 FILLER_323_320 ();
 b15zdnd11an1n64x5 FILLER_323_384 ();
 b15zdnd11an1n64x5 FILLER_323_448 ();
 b15zdnd11an1n64x5 FILLER_323_512 ();
 b15zdnd11an1n64x5 FILLER_323_576 ();
 b15zdnd11an1n64x5 FILLER_323_640 ();
 b15zdnd11an1n64x5 FILLER_323_704 ();
 b15zdnd11an1n64x5 FILLER_323_768 ();
 b15zdnd11an1n64x5 FILLER_323_832 ();
 b15zdnd11an1n64x5 FILLER_323_896 ();
 b15zdnd11an1n64x5 FILLER_323_960 ();
 b15zdnd11an1n64x5 FILLER_323_1024 ();
 b15zdnd11an1n64x5 FILLER_323_1088 ();
 b15zdnd11an1n64x5 FILLER_323_1152 ();
 b15zdnd11an1n64x5 FILLER_323_1216 ();
 b15zdnd11an1n04x5 FILLER_323_1280 ();
 b15zdnd00an1n02x5 FILLER_323_1284 ();
 b15zdnd11an1n04x5 FILLER_323_1289 ();
 b15zdnd11an1n04x5 FILLER_323_1296 ();
 b15zdnd11an1n64x5 FILLER_323_1303 ();
 b15zdnd11an1n64x5 FILLER_323_1367 ();
 b15zdnd11an1n64x5 FILLER_323_1431 ();
 b15zdnd11an1n64x5 FILLER_323_1495 ();
 b15zdnd11an1n64x5 FILLER_323_1559 ();
 b15zdnd11an1n64x5 FILLER_323_1623 ();
 b15zdnd11an1n16x5 FILLER_323_1687 ();
 b15zdnd11an1n08x5 FILLER_323_1703 ();
 b15zdnd11an1n04x5 FILLER_323_1711 ();
 b15zdnd00an1n01x5 FILLER_323_1715 ();
 b15zdnd11an1n04x5 FILLER_323_1719 ();
 b15zdnd11an1n32x5 FILLER_323_1726 ();
 b15zdnd11an1n16x5 FILLER_323_1758 ();
 b15zdnd00an1n01x5 FILLER_323_1774 ();
 b15zdnd11an1n64x5 FILLER_323_1780 ();
 b15zdnd11an1n64x5 FILLER_323_1844 ();
 b15zdnd11an1n32x5 FILLER_323_1908 ();
 b15zdnd11an1n16x5 FILLER_323_1940 ();
 b15zdnd11an1n04x5 FILLER_323_1956 ();
 b15zdnd00an1n01x5 FILLER_323_1960 ();
 b15zdnd11an1n04x5 FILLER_323_1971 ();
 b15zdnd11an1n04x5 FILLER_323_1978 ();
 b15zdnd00an1n02x5 FILLER_323_1982 ();
 b15zdnd11an1n64x5 FILLER_323_1987 ();
 b15zdnd11an1n64x5 FILLER_323_2051 ();
 b15zdnd11an1n64x5 FILLER_323_2115 ();
 b15zdnd11an1n64x5 FILLER_323_2179 ();
 b15zdnd11an1n32x5 FILLER_323_2243 ();
 b15zdnd11an1n08x5 FILLER_323_2275 ();
 b15zdnd00an1n01x5 FILLER_323_2283 ();
 b15zdnd11an1n32x5 FILLER_324_8 ();
 b15zdnd11an1n16x5 FILLER_324_40 ();
 b15zdnd11an1n04x5 FILLER_324_56 ();
 b15zdnd00an1n01x5 FILLER_324_60 ();
 b15zdnd11an1n64x5 FILLER_324_64 ();
 b15zdnd11an1n64x5 FILLER_324_128 ();
 b15zdnd11an1n64x5 FILLER_324_192 ();
 b15zdnd11an1n64x5 FILLER_324_256 ();
 b15zdnd11an1n64x5 FILLER_324_320 ();
 b15zdnd11an1n64x5 FILLER_324_384 ();
 b15zdnd11an1n64x5 FILLER_324_448 ();
 b15zdnd11an1n64x5 FILLER_324_512 ();
 b15zdnd11an1n64x5 FILLER_324_576 ();
 b15zdnd11an1n64x5 FILLER_324_640 ();
 b15zdnd11an1n08x5 FILLER_324_704 ();
 b15zdnd11an1n04x5 FILLER_324_712 ();
 b15zdnd00an1n02x5 FILLER_324_716 ();
 b15zdnd11an1n64x5 FILLER_324_726 ();
 b15zdnd11an1n64x5 FILLER_324_790 ();
 b15zdnd11an1n64x5 FILLER_324_854 ();
 b15zdnd11an1n64x5 FILLER_324_918 ();
 b15zdnd11an1n64x5 FILLER_324_982 ();
 b15zdnd11an1n64x5 FILLER_324_1046 ();
 b15zdnd11an1n32x5 FILLER_324_1110 ();
 b15zdnd11an1n16x5 FILLER_324_1142 ();
 b15zdnd11an1n08x5 FILLER_324_1158 ();
 b15zdnd00an1n01x5 FILLER_324_1166 ();
 b15zdnd11an1n04x5 FILLER_324_1170 ();
 b15zdnd11an1n64x5 FILLER_324_1177 ();
 b15zdnd11an1n32x5 FILLER_324_1241 ();
 b15zdnd11an1n08x5 FILLER_324_1273 ();
 b15zdnd11an1n04x5 FILLER_324_1281 ();
 b15zdnd00an1n01x5 FILLER_324_1285 ();
 b15zdnd11an1n04x5 FILLER_324_1289 ();
 b15zdnd11an1n64x5 FILLER_324_1296 ();
 b15zdnd11an1n64x5 FILLER_324_1360 ();
 b15zdnd11an1n64x5 FILLER_324_1424 ();
 b15zdnd11an1n64x5 FILLER_324_1488 ();
 b15zdnd11an1n64x5 FILLER_324_1552 ();
 b15zdnd11an1n64x5 FILLER_324_1616 ();
 b15zdnd11an1n16x5 FILLER_324_1680 ();
 b15zdnd00an1n02x5 FILLER_324_1696 ();
 b15zdnd11an1n08x5 FILLER_324_1750 ();
 b15zdnd11an1n04x5 FILLER_324_1758 ();
 b15zdnd11an1n64x5 FILLER_324_1804 ();
 b15zdnd11an1n64x5 FILLER_324_1868 ();
 b15zdnd11an1n16x5 FILLER_324_1932 ();
 b15zdnd11an1n04x5 FILLER_324_1948 ();
 b15zdnd11an1n64x5 FILLER_324_2004 ();
 b15zdnd11an1n64x5 FILLER_324_2068 ();
 b15zdnd11an1n16x5 FILLER_324_2132 ();
 b15zdnd11an1n04x5 FILLER_324_2148 ();
 b15zdnd00an1n02x5 FILLER_324_2152 ();
 b15zdnd11an1n64x5 FILLER_324_2162 ();
 b15zdnd11an1n32x5 FILLER_324_2226 ();
 b15zdnd11an1n16x5 FILLER_324_2258 ();
 b15zdnd00an1n02x5 FILLER_324_2274 ();
 b15zdnd11an1n64x5 FILLER_325_0 ();
 b15zdnd11an1n04x5 FILLER_325_71 ();
 b15zdnd11an1n64x5 FILLER_325_80 ();
 b15zdnd11an1n64x5 FILLER_325_144 ();
 b15zdnd11an1n64x5 FILLER_325_208 ();
 b15zdnd11an1n64x5 FILLER_325_272 ();
 b15zdnd11an1n32x5 FILLER_325_336 ();
 b15zdnd11an1n64x5 FILLER_325_371 ();
 b15zdnd11an1n64x5 FILLER_325_435 ();
 b15zdnd11an1n64x5 FILLER_325_499 ();
 b15zdnd11an1n64x5 FILLER_325_563 ();
 b15zdnd11an1n64x5 FILLER_325_627 ();
 b15zdnd11an1n64x5 FILLER_325_691 ();
 b15zdnd11an1n64x5 FILLER_325_755 ();
 b15zdnd11an1n64x5 FILLER_325_819 ();
 b15zdnd11an1n64x5 FILLER_325_883 ();
 b15zdnd11an1n64x5 FILLER_325_947 ();
 b15zdnd11an1n64x5 FILLER_325_1011 ();
 b15zdnd11an1n64x5 FILLER_325_1075 ();
 b15zdnd11an1n08x5 FILLER_325_1139 ();
 b15zdnd00an1n02x5 FILLER_325_1147 ();
 b15zdnd11an1n64x5 FILLER_325_1201 ();
 b15zdnd11an1n64x5 FILLER_325_1265 ();
 b15zdnd11an1n64x5 FILLER_325_1329 ();
 b15zdnd11an1n64x5 FILLER_325_1393 ();
 b15zdnd11an1n64x5 FILLER_325_1457 ();
 b15zdnd11an1n64x5 FILLER_325_1521 ();
 b15zdnd11an1n64x5 FILLER_325_1585 ();
 b15zdnd11an1n64x5 FILLER_325_1649 ();
 b15zdnd11an1n08x5 FILLER_325_1713 ();
 b15zdnd00an1n02x5 FILLER_325_1721 ();
 b15zdnd00an1n01x5 FILLER_325_1723 ();
 b15zdnd11an1n64x5 FILLER_325_1727 ();
 b15zdnd11an1n64x5 FILLER_325_1791 ();
 b15zdnd11an1n64x5 FILLER_325_1855 ();
 b15zdnd11an1n32x5 FILLER_325_1919 ();
 b15zdnd11an1n16x5 FILLER_325_1956 ();
 b15zdnd00an1n02x5 FILLER_325_1972 ();
 b15zdnd11an1n64x5 FILLER_325_1977 ();
 b15zdnd11an1n64x5 FILLER_325_2041 ();
 b15zdnd11an1n64x5 FILLER_325_2105 ();
 b15zdnd11an1n64x5 FILLER_325_2169 ();
 b15zdnd11an1n32x5 FILLER_325_2233 ();
 b15zdnd11an1n16x5 FILLER_325_2265 ();
 b15zdnd00an1n02x5 FILLER_325_2281 ();
 b15zdnd00an1n01x5 FILLER_325_2283 ();
 b15zdnd11an1n64x5 FILLER_326_8 ();
 b15zdnd11an1n64x5 FILLER_326_72 ();
 b15zdnd11an1n64x5 FILLER_326_136 ();
 b15zdnd11an1n64x5 FILLER_326_200 ();
 b15zdnd11an1n64x5 FILLER_326_264 ();
 b15zdnd00an1n02x5 FILLER_326_328 ();
 b15zdnd00an1n01x5 FILLER_326_330 ();
 b15zdnd11an1n64x5 FILLER_326_371 ();
 b15zdnd11an1n32x5 FILLER_326_435 ();
 b15zdnd11an1n16x5 FILLER_326_467 ();
 b15zdnd11an1n08x5 FILLER_326_483 ();
 b15zdnd00an1n02x5 FILLER_326_491 ();
 b15zdnd00an1n01x5 FILLER_326_493 ();
 b15zdnd11an1n64x5 FILLER_326_497 ();
 b15zdnd11an1n32x5 FILLER_326_561 ();
 b15zdnd11an1n04x5 FILLER_326_593 ();
 b15zdnd00an1n02x5 FILLER_326_597 ();
 b15zdnd11an1n16x5 FILLER_326_608 ();
 b15zdnd11an1n04x5 FILLER_326_624 ();
 b15zdnd11an1n16x5 FILLER_326_631 ();
 b15zdnd11an1n08x5 FILLER_326_647 ();
 b15zdnd11an1n32x5 FILLER_326_664 ();
 b15zdnd11an1n16x5 FILLER_326_696 ();
 b15zdnd11an1n04x5 FILLER_326_712 ();
 b15zdnd00an1n02x5 FILLER_326_716 ();
 b15zdnd11an1n16x5 FILLER_326_726 ();
 b15zdnd11an1n08x5 FILLER_326_742 ();
 b15zdnd11an1n04x5 FILLER_326_750 ();
 b15zdnd00an1n02x5 FILLER_326_754 ();
 b15zdnd00an1n01x5 FILLER_326_756 ();
 b15zdnd11an1n64x5 FILLER_326_784 ();
 b15zdnd11an1n64x5 FILLER_326_848 ();
 b15zdnd11an1n64x5 FILLER_326_912 ();
 b15zdnd11an1n32x5 FILLER_326_976 ();
 b15zdnd11an1n04x5 FILLER_326_1008 ();
 b15zdnd11an1n64x5 FILLER_326_1015 ();
 b15zdnd11an1n64x5 FILLER_326_1079 ();
 b15zdnd11an1n32x5 FILLER_326_1143 ();
 b15zdnd11an1n16x5 FILLER_326_1178 ();
 b15zdnd11an1n08x5 FILLER_326_1194 ();
 b15zdnd11an1n04x5 FILLER_326_1202 ();
 b15zdnd00an1n01x5 FILLER_326_1206 ();
 b15zdnd11an1n64x5 FILLER_326_1227 ();
 b15zdnd11an1n64x5 FILLER_326_1291 ();
 b15zdnd11an1n64x5 FILLER_326_1355 ();
 b15zdnd11an1n08x5 FILLER_326_1419 ();
 b15zdnd11an1n04x5 FILLER_326_1427 ();
 b15zdnd00an1n02x5 FILLER_326_1431 ();
 b15zdnd11an1n04x5 FILLER_326_1460 ();
 b15zdnd11an1n64x5 FILLER_326_1473 ();
 b15zdnd11an1n64x5 FILLER_326_1537 ();
 b15zdnd11an1n64x5 FILLER_326_1601 ();
 b15zdnd11an1n64x5 FILLER_326_1665 ();
 b15zdnd11an1n64x5 FILLER_326_1729 ();
 b15zdnd11an1n64x5 FILLER_326_1793 ();
 b15zdnd11an1n64x5 FILLER_326_1857 ();
 b15zdnd11an1n16x5 FILLER_326_1921 ();
 b15zdnd11an1n08x5 FILLER_326_1937 ();
 b15zdnd11an1n04x5 FILLER_326_1945 ();
 b15zdnd00an1n02x5 FILLER_326_1949 ();
 b15zdnd11an1n64x5 FILLER_326_1958 ();
 b15zdnd11an1n64x5 FILLER_326_2022 ();
 b15zdnd11an1n16x5 FILLER_326_2086 ();
 b15zdnd11an1n08x5 FILLER_326_2102 ();
 b15zdnd00an1n02x5 FILLER_326_2110 ();
 b15zdnd00an1n01x5 FILLER_326_2112 ();
 b15zdnd11an1n16x5 FILLER_326_2116 ();
 b15zdnd11an1n08x5 FILLER_326_2132 ();
 b15zdnd00an1n02x5 FILLER_326_2140 ();
 b15zdnd00an1n01x5 FILLER_326_2142 ();
 b15zdnd11an1n08x5 FILLER_326_2146 ();
 b15zdnd11an1n64x5 FILLER_326_2162 ();
 b15zdnd11an1n32x5 FILLER_326_2226 ();
 b15zdnd11an1n16x5 FILLER_326_2258 ();
 b15zdnd00an1n02x5 FILLER_326_2274 ();
 b15zdnd11an1n64x5 FILLER_327_0 ();
 b15zdnd11an1n04x5 FILLER_327_64 ();
 b15zdnd00an1n02x5 FILLER_327_68 ();
 b15zdnd00an1n01x5 FILLER_327_70 ();
 b15zdnd11an1n64x5 FILLER_327_76 ();
 b15zdnd11an1n64x5 FILLER_327_140 ();
 b15zdnd11an1n16x5 FILLER_327_204 ();
 b15zdnd11an1n08x5 FILLER_327_220 ();
 b15zdnd00an1n02x5 FILLER_327_228 ();
 b15zdnd11an1n64x5 FILLER_327_233 ();
 b15zdnd11an1n64x5 FILLER_327_297 ();
 b15zdnd11an1n04x5 FILLER_327_361 ();
 b15zdnd00an1n02x5 FILLER_327_365 ();
 b15zdnd11an1n04x5 FILLER_327_370 ();
 b15zdnd11an1n64x5 FILLER_327_377 ();
 b15zdnd11an1n32x5 FILLER_327_441 ();
 b15zdnd11an1n16x5 FILLER_327_473 ();
 b15zdnd11an1n04x5 FILLER_327_492 ();
 b15zdnd11an1n04x5 FILLER_327_499 ();
 b15zdnd00an1n01x5 FILLER_327_503 ();
 b15zdnd11an1n64x5 FILLER_327_507 ();
 b15zdnd11an1n32x5 FILLER_327_571 ();
 b15zdnd11an1n16x5 FILLER_327_603 ();
 b15zdnd00an1n02x5 FILLER_327_619 ();
 b15zdnd11an1n04x5 FILLER_327_624 ();
 b15zdnd11an1n64x5 FILLER_327_631 ();
 b15zdnd11an1n32x5 FILLER_327_695 ();
 b15zdnd11an1n16x5 FILLER_327_727 ();
 b15zdnd00an1n02x5 FILLER_327_743 ();
 b15zdnd00an1n01x5 FILLER_327_745 ();
 b15zdnd11an1n64x5 FILLER_327_798 ();
 b15zdnd11an1n32x5 FILLER_327_862 ();
 b15zdnd11an1n04x5 FILLER_327_894 ();
 b15zdnd11an1n64x5 FILLER_327_901 ();
 b15zdnd11an1n32x5 FILLER_327_965 ();
 b15zdnd11an1n08x5 FILLER_327_997 ();
 b15zdnd00an1n01x5 FILLER_327_1005 ();
 b15zdnd11an1n04x5 FILLER_327_1009 ();
 b15zdnd11an1n04x5 FILLER_327_1016 ();
 b15zdnd11an1n64x5 FILLER_327_1023 ();
 b15zdnd11an1n64x5 FILLER_327_1087 ();
 b15zdnd11an1n32x5 FILLER_327_1151 ();
 b15zdnd00an1n01x5 FILLER_327_1183 ();
 b15zdnd11an1n64x5 FILLER_327_1187 ();
 b15zdnd11an1n64x5 FILLER_327_1251 ();
 b15zdnd11an1n64x5 FILLER_327_1315 ();
 b15zdnd11an1n32x5 FILLER_327_1379 ();
 b15zdnd11an1n16x5 FILLER_327_1411 ();
 b15zdnd11an1n04x5 FILLER_327_1427 ();
 b15zdnd00an1n02x5 FILLER_327_1431 ();
 b15zdnd11an1n04x5 FILLER_327_1436 ();
 b15zdnd11an1n64x5 FILLER_327_1468 ();
 b15zdnd11an1n64x5 FILLER_327_1532 ();
 b15zdnd00an1n02x5 FILLER_327_1596 ();
 b15zdnd00an1n01x5 FILLER_327_1598 ();
 b15zdnd11an1n64x5 FILLER_327_1602 ();
 b15zdnd11an1n32x5 FILLER_327_1666 ();
 b15zdnd11an1n16x5 FILLER_327_1698 ();
 b15zdnd11an1n04x5 FILLER_327_1714 ();
 b15zdnd00an1n02x5 FILLER_327_1718 ();
 b15zdnd00an1n01x5 FILLER_327_1720 ();
 b15zdnd11an1n04x5 FILLER_327_1724 ();
 b15zdnd00an1n02x5 FILLER_327_1728 ();
 b15zdnd00an1n01x5 FILLER_327_1730 ();
 b15zdnd11an1n64x5 FILLER_327_1773 ();
 b15zdnd11an1n64x5 FILLER_327_1837 ();
 b15zdnd11an1n32x5 FILLER_327_1901 ();
 b15zdnd11an1n08x5 FILLER_327_1933 ();
 b15zdnd11an1n04x5 FILLER_327_1941 ();
 b15zdnd00an1n02x5 FILLER_327_1945 ();
 b15zdnd11an1n64x5 FILLER_327_1958 ();
 b15zdnd11an1n64x5 FILLER_327_2022 ();
 b15zdnd11an1n32x5 FILLER_327_2086 ();
 b15zdnd11an1n64x5 FILLER_327_2170 ();
 b15zdnd11an1n32x5 FILLER_327_2234 ();
 b15zdnd11an1n16x5 FILLER_327_2266 ();
 b15zdnd00an1n02x5 FILLER_327_2282 ();
 b15zdnd11an1n64x5 FILLER_328_8 ();
 b15zdnd11an1n64x5 FILLER_328_72 ();
 b15zdnd11an1n32x5 FILLER_328_136 ();
 b15zdnd11an1n08x5 FILLER_328_168 ();
 b15zdnd00an1n01x5 FILLER_328_176 ();
 b15zdnd11an1n04x5 FILLER_328_191 ();
 b15zdnd11an1n04x5 FILLER_328_235 ();
 b15zdnd11an1n64x5 FILLER_328_242 ();
 b15zdnd11an1n32x5 FILLER_328_306 ();
 b15zdnd11an1n04x5 FILLER_328_338 ();
 b15zdnd11an1n04x5 FILLER_328_382 ();
 b15zdnd00an1n01x5 FILLER_328_386 ();
 b15zdnd11an1n64x5 FILLER_328_390 ();
 b15zdnd11an1n08x5 FILLER_328_454 ();
 b15zdnd11an1n04x5 FILLER_328_462 ();
 b15zdnd00an1n02x5 FILLER_328_466 ();
 b15zdnd00an1n01x5 FILLER_328_468 ();
 b15zdnd11an1n32x5 FILLER_328_521 ();
 b15zdnd11an1n16x5 FILLER_328_553 ();
 b15zdnd11an1n08x5 FILLER_328_569 ();
 b15zdnd11an1n04x5 FILLER_328_577 ();
 b15zdnd00an1n02x5 FILLER_328_581 ();
 b15zdnd11an1n08x5 FILLER_328_610 ();
 b15zdnd00an1n02x5 FILLER_328_618 ();
 b15zdnd00an1n01x5 FILLER_328_620 ();
 b15zdnd11an1n32x5 FILLER_328_673 ();
 b15zdnd11an1n08x5 FILLER_328_705 ();
 b15zdnd11an1n04x5 FILLER_328_713 ();
 b15zdnd00an1n01x5 FILLER_328_717 ();
 b15zdnd11an1n08x5 FILLER_328_726 ();
 b15zdnd11an1n04x5 FILLER_328_734 ();
 b15zdnd00an1n02x5 FILLER_328_738 ();
 b15zdnd11an1n04x5 FILLER_328_743 ();
 b15zdnd11an1n04x5 FILLER_328_799 ();
 b15zdnd11an1n64x5 FILLER_328_806 ();
 b15zdnd11an1n16x5 FILLER_328_870 ();
 b15zdnd11an1n08x5 FILLER_328_886 ();
 b15zdnd11an1n04x5 FILLER_328_894 ();
 b15zdnd11an1n32x5 FILLER_328_925 ();
 b15zdnd11an1n16x5 FILLER_328_957 ();
 b15zdnd11an1n08x5 FILLER_328_973 ();
 b15zdnd11an1n04x5 FILLER_328_981 ();
 b15zdnd00an1n01x5 FILLER_328_985 ();
 b15zdnd11an1n64x5 FILLER_328_1038 ();
 b15zdnd11an1n32x5 FILLER_328_1102 ();
 b15zdnd11an1n16x5 FILLER_328_1134 ();
 b15zdnd11an1n08x5 FILLER_328_1150 ();
 b15zdnd11an1n16x5 FILLER_328_1210 ();
 b15zdnd11an1n08x5 FILLER_328_1226 ();
 b15zdnd11an1n04x5 FILLER_328_1234 ();
 b15zdnd11an1n64x5 FILLER_328_1252 ();
 b15zdnd11an1n64x5 FILLER_328_1316 ();
 b15zdnd11an1n32x5 FILLER_328_1380 ();
 b15zdnd11an1n16x5 FILLER_328_1412 ();
 b15zdnd11an1n04x5 FILLER_328_1428 ();
 b15zdnd00an1n01x5 FILLER_328_1432 ();
 b15zdnd11an1n04x5 FILLER_328_1485 ();
 b15zdnd11an1n64x5 FILLER_328_1492 ();
 b15zdnd11an1n32x5 FILLER_328_1556 ();
 b15zdnd00an1n02x5 FILLER_328_1588 ();
 b15zdnd11an1n04x5 FILLER_328_1593 ();
 b15zdnd00an1n02x5 FILLER_328_1597 ();
 b15zdnd00an1n01x5 FILLER_328_1599 ();
 b15zdnd11an1n64x5 FILLER_328_1603 ();
 b15zdnd11an1n32x5 FILLER_328_1667 ();
 b15zdnd11an1n08x5 FILLER_328_1699 ();
 b15zdnd11an1n04x5 FILLER_328_1707 ();
 b15zdnd00an1n01x5 FILLER_328_1711 ();
 b15zdnd11an1n04x5 FILLER_328_1715 ();
 b15zdnd00an1n02x5 FILLER_328_1719 ();
 b15zdnd00an1n01x5 FILLER_328_1721 ();
 b15zdnd11an1n16x5 FILLER_328_1725 ();
 b15zdnd11an1n04x5 FILLER_328_1741 ();
 b15zdnd11an1n64x5 FILLER_328_1765 ();
 b15zdnd11an1n32x5 FILLER_328_1829 ();
 b15zdnd11an1n08x5 FILLER_328_1877 ();
 b15zdnd00an1n01x5 FILLER_328_1885 ();
 b15zdnd11an1n16x5 FILLER_328_1897 ();
 b15zdnd11an1n04x5 FILLER_328_1913 ();
 b15zdnd00an1n02x5 FILLER_328_1917 ();
 b15zdnd11an1n64x5 FILLER_328_1961 ();
 b15zdnd11an1n16x5 FILLER_328_2025 ();
 b15zdnd11an1n04x5 FILLER_328_2041 ();
 b15zdnd11an1n08x5 FILLER_328_2048 ();
 b15zdnd11an1n16x5 FILLER_328_2062 ();
 b15zdnd00an1n02x5 FILLER_328_2078 ();
 b15zdnd11an1n16x5 FILLER_328_2085 ();
 b15zdnd11an1n08x5 FILLER_328_2101 ();
 b15zdnd00an1n02x5 FILLER_328_2109 ();
 b15zdnd00an1n01x5 FILLER_328_2111 ();
 b15zdnd11an1n08x5 FILLER_328_2119 ();
 b15zdnd00an1n01x5 FILLER_328_2127 ();
 b15zdnd11an1n04x5 FILLER_328_2132 ();
 b15zdnd11an1n04x5 FILLER_328_2142 ();
 b15zdnd11an1n04x5 FILLER_328_2149 ();
 b15zdnd00an1n01x5 FILLER_328_2153 ();
 b15zdnd00an1n02x5 FILLER_328_2162 ();
 b15zdnd11an1n64x5 FILLER_328_2206 ();
 b15zdnd11an1n04x5 FILLER_328_2270 ();
 b15zdnd00an1n02x5 FILLER_328_2274 ();
 b15zdnd11an1n64x5 FILLER_329_0 ();
 b15zdnd11an1n64x5 FILLER_329_64 ();
 b15zdnd11an1n64x5 FILLER_329_128 ();
 b15zdnd00an1n02x5 FILLER_329_192 ();
 b15zdnd00an1n01x5 FILLER_329_194 ();
 b15zdnd11an1n04x5 FILLER_329_235 ();
 b15zdnd11an1n04x5 FILLER_329_242 ();
 b15zdnd11an1n64x5 FILLER_329_249 ();
 b15zdnd11an1n16x5 FILLER_329_313 ();
 b15zdnd11an1n04x5 FILLER_329_343 ();
 b15zdnd11an1n04x5 FILLER_329_387 ();
 b15zdnd11an1n64x5 FILLER_329_394 ();
 b15zdnd11an1n08x5 FILLER_329_458 ();
 b15zdnd11an1n04x5 FILLER_329_506 ();
 b15zdnd11an1n16x5 FILLER_329_552 ();
 b15zdnd11an1n08x5 FILLER_329_568 ();
 b15zdnd11an1n04x5 FILLER_329_576 ();
 b15zdnd00an1n01x5 FILLER_329_580 ();
 b15zdnd11an1n16x5 FILLER_329_584 ();
 b15zdnd00an1n02x5 FILLER_329_600 ();
 b15zdnd11an1n04x5 FILLER_329_654 ();
 b15zdnd11an1n64x5 FILLER_329_661 ();
 b15zdnd11an1n16x5 FILLER_329_725 ();
 b15zdnd11an1n04x5 FILLER_329_741 ();
 b15zdnd00an1n02x5 FILLER_329_745 ();
 b15zdnd11an1n04x5 FILLER_329_799 ();
 b15zdnd11an1n64x5 FILLER_329_806 ();
 b15zdnd11an1n08x5 FILLER_329_870 ();
 b15zdnd00an1n02x5 FILLER_329_878 ();
 b15zdnd11an1n04x5 FILLER_329_932 ();
 b15zdnd11an1n32x5 FILLER_329_939 ();
 b15zdnd11an1n16x5 FILLER_329_971 ();
 b15zdnd11an1n08x5 FILLER_329_987 ();
 b15zdnd11an1n04x5 FILLER_329_995 ();
 b15zdnd00an1n01x5 FILLER_329_999 ();
 b15zdnd11an1n64x5 FILLER_329_1052 ();
 b15zdnd11an1n32x5 FILLER_329_1116 ();
 b15zdnd11an1n16x5 FILLER_329_1148 ();
 b15zdnd11an1n08x5 FILLER_329_1164 ();
 b15zdnd11an1n04x5 FILLER_329_1172 ();
 b15zdnd00an1n02x5 FILLER_329_1176 ();
 b15zdnd00an1n01x5 FILLER_329_1178 ();
 b15zdnd11an1n04x5 FILLER_329_1182 ();
 b15zdnd11an1n64x5 FILLER_329_1189 ();
 b15zdnd11an1n64x5 FILLER_329_1253 ();
 b15zdnd11an1n64x5 FILLER_329_1317 ();
 b15zdnd11an1n32x5 FILLER_329_1381 ();
 b15zdnd11an1n08x5 FILLER_329_1413 ();
 b15zdnd11an1n04x5 FILLER_329_1473 ();
 b15zdnd11an1n04x5 FILLER_329_1480 ();
 b15zdnd11an1n64x5 FILLER_329_1487 ();
 b15zdnd11an1n16x5 FILLER_329_1551 ();
 b15zdnd11an1n08x5 FILLER_329_1567 ();
 b15zdnd00an1n02x5 FILLER_329_1575 ();
 b15zdnd11an1n64x5 FILLER_329_1629 ();
 b15zdnd11an1n64x5 FILLER_329_1745 ();
 b15zdnd11an1n32x5 FILLER_329_1809 ();
 b15zdnd11an1n08x5 FILLER_329_1841 ();
 b15zdnd00an1n02x5 FILLER_329_1849 ();
 b15zdnd11an1n04x5 FILLER_329_1854 ();
 b15zdnd11an1n32x5 FILLER_329_1861 ();
 b15zdnd00an1n02x5 FILLER_329_1893 ();
 b15zdnd00an1n01x5 FILLER_329_1895 ();
 b15zdnd11an1n64x5 FILLER_329_1904 ();
 b15zdnd11an1n64x5 FILLER_329_1968 ();
 b15zdnd11an1n04x5 FILLER_329_2032 ();
 b15zdnd00an1n02x5 FILLER_329_2036 ();
 b15zdnd11an1n04x5 FILLER_329_2041 ();
 b15zdnd11an1n16x5 FILLER_329_2048 ();
 b15zdnd11an1n08x5 FILLER_329_2064 ();
 b15zdnd11an1n04x5 FILLER_329_2072 ();
 b15zdnd00an1n02x5 FILLER_329_2076 ();
 b15zdnd00an1n01x5 FILLER_329_2078 ();
 b15zdnd11an1n04x5 FILLER_329_2089 ();
 b15zdnd11an1n08x5 FILLER_329_2103 ();
 b15zdnd11an1n04x5 FILLER_329_2111 ();
 b15zdnd00an1n02x5 FILLER_329_2115 ();
 b15zdnd11an1n04x5 FILLER_329_2159 ();
 b15zdnd11an1n64x5 FILLER_329_2205 ();
 b15zdnd11an1n08x5 FILLER_329_2269 ();
 b15zdnd11an1n04x5 FILLER_329_2277 ();
 b15zdnd00an1n02x5 FILLER_329_2281 ();
 b15zdnd00an1n01x5 FILLER_329_2283 ();
 b15zdnd11an1n64x5 FILLER_330_8 ();
 b15zdnd00an1n01x5 FILLER_330_72 ();
 b15zdnd11an1n08x5 FILLER_330_77 ();
 b15zdnd00an1n01x5 FILLER_330_85 ();
 b15zdnd11an1n04x5 FILLER_330_95 ();
 b15zdnd11an1n64x5 FILLER_330_106 ();
 b15zdnd11an1n16x5 FILLER_330_170 ();
 b15zdnd11an1n04x5 FILLER_330_186 ();
 b15zdnd00an1n02x5 FILLER_330_190 ();
 b15zdnd00an1n01x5 FILLER_330_192 ();
 b15zdnd11an1n04x5 FILLER_330_233 ();
 b15zdnd11an1n08x5 FILLER_330_240 ();
 b15zdnd11an1n04x5 FILLER_330_248 ();
 b15zdnd00an1n02x5 FILLER_330_252 ();
 b15zdnd00an1n01x5 FILLER_330_254 ();
 b15zdnd11an1n64x5 FILLER_330_271 ();
 b15zdnd11an1n16x5 FILLER_330_335 ();
 b15zdnd11an1n08x5 FILLER_330_351 ();
 b15zdnd11an1n04x5 FILLER_330_359 ();
 b15zdnd00an1n02x5 FILLER_330_363 ();
 b15zdnd11an1n32x5 FILLER_330_407 ();
 b15zdnd11an1n16x5 FILLER_330_439 ();
 b15zdnd11an1n08x5 FILLER_330_455 ();
 b15zdnd11an1n04x5 FILLER_330_463 ();
 b15zdnd00an1n01x5 FILLER_330_467 ();
 b15zdnd11an1n04x5 FILLER_330_508 ();
 b15zdnd00an1n01x5 FILLER_330_512 ();
 b15zdnd11an1n08x5 FILLER_330_516 ();
 b15zdnd00an1n01x5 FILLER_330_524 ();
 b15zdnd11an1n32x5 FILLER_330_567 ();
 b15zdnd00an1n02x5 FILLER_330_599 ();
 b15zdnd00an1n01x5 FILLER_330_601 ();
 b15zdnd11an1n04x5 FILLER_330_654 ();
 b15zdnd11an1n04x5 FILLER_330_661 ();
 b15zdnd11an1n32x5 FILLER_330_668 ();
 b15zdnd11an1n16x5 FILLER_330_700 ();
 b15zdnd00an1n02x5 FILLER_330_716 ();
 b15zdnd11an1n16x5 FILLER_330_726 ();
 b15zdnd11an1n04x5 FILLER_330_742 ();
 b15zdnd00an1n02x5 FILLER_330_746 ();
 b15zdnd00an1n01x5 FILLER_330_748 ();
 b15zdnd11an1n64x5 FILLER_330_801 ();
 b15zdnd11an1n08x5 FILLER_330_865 ();
 b15zdnd11an1n04x5 FILLER_330_873 ();
 b15zdnd00an1n02x5 FILLER_330_877 ();
 b15zdnd00an1n01x5 FILLER_330_879 ();
 b15zdnd11an1n04x5 FILLER_330_932 ();
 b15zdnd11an1n32x5 FILLER_330_945 ();
 b15zdnd11an1n08x5 FILLER_330_977 ();
 b15zdnd00an1n02x5 FILLER_330_985 ();
 b15zdnd00an1n01x5 FILLER_330_987 ();
 b15zdnd11an1n08x5 FILLER_330_997 ();
 b15zdnd11an1n04x5 FILLER_330_1005 ();
 b15zdnd11an1n64x5 FILLER_330_1061 ();
 b15zdnd11an1n64x5 FILLER_330_1125 ();
 b15zdnd11an1n16x5 FILLER_330_1189 ();
 b15zdnd11an1n08x5 FILLER_330_1205 ();
 b15zdnd00an1n02x5 FILLER_330_1213 ();
 b15zdnd11an1n64x5 FILLER_330_1241 ();
 b15zdnd11an1n64x5 FILLER_330_1305 ();
 b15zdnd11an1n32x5 FILLER_330_1369 ();
 b15zdnd11an1n16x5 FILLER_330_1401 ();
 b15zdnd11an1n04x5 FILLER_330_1417 ();
 b15zdnd11an1n04x5 FILLER_330_1473 ();
 b15zdnd11an1n04x5 FILLER_330_1480 ();
 b15zdnd11an1n64x5 FILLER_330_1487 ();
 b15zdnd11an1n64x5 FILLER_330_1551 ();
 b15zdnd11an1n64x5 FILLER_330_1621 ();
 b15zdnd11an1n16x5 FILLER_330_1685 ();
 b15zdnd11an1n08x5 FILLER_330_1701 ();
 b15zdnd11an1n04x5 FILLER_330_1709 ();
 b15zdnd11an1n04x5 FILLER_330_1716 ();
 b15zdnd11an1n16x5 FILLER_330_1723 ();
 b15zdnd11an1n04x5 FILLER_330_1739 ();
 b15zdnd11an1n04x5 FILLER_330_1746 ();
 b15zdnd11an1n64x5 FILLER_330_1753 ();
 b15zdnd11an1n08x5 FILLER_330_1817 ();
 b15zdnd11an1n04x5 FILLER_330_1825 ();
 b15zdnd11an1n64x5 FILLER_330_1881 ();
 b15zdnd11an1n32x5 FILLER_330_1945 ();
 b15zdnd11an1n16x5 FILLER_330_1977 ();
 b15zdnd11an1n04x5 FILLER_330_1993 ();
 b15zdnd00an1n01x5 FILLER_330_1997 ();
 b15zdnd11an1n04x5 FILLER_330_2018 ();
 b15zdnd11an1n04x5 FILLER_330_2074 ();
 b15zdnd11an1n04x5 FILLER_330_2120 ();
 b15zdnd11an1n04x5 FILLER_330_2134 ();
 b15zdnd11an1n04x5 FILLER_330_2143 ();
 b15zdnd00an1n02x5 FILLER_330_2152 ();
 b15zdnd11an1n64x5 FILLER_330_2162 ();
 b15zdnd11an1n32x5 FILLER_330_2226 ();
 b15zdnd11an1n16x5 FILLER_330_2258 ();
 b15zdnd00an1n02x5 FILLER_330_2274 ();
 b15zdnd11an1n64x5 FILLER_331_0 ();
 b15zdnd11an1n16x5 FILLER_331_64 ();
 b15zdnd11an1n04x5 FILLER_331_80 ();
 b15zdnd00an1n02x5 FILLER_331_84 ();
 b15zdnd11an1n64x5 FILLER_331_106 ();
 b15zdnd11an1n16x5 FILLER_331_170 ();
 b15zdnd11an1n08x5 FILLER_331_186 ();
 b15zdnd00an1n02x5 FILLER_331_194 ();
 b15zdnd11an1n64x5 FILLER_331_238 ();
 b15zdnd11an1n32x5 FILLER_331_302 ();
 b15zdnd00an1n01x5 FILLER_331_334 ();
 b15zdnd11an1n08x5 FILLER_331_375 ();
 b15zdnd00an1n02x5 FILLER_331_383 ();
 b15zdnd11an1n04x5 FILLER_331_393 ();
 b15zdnd11an1n64x5 FILLER_331_400 ();
 b15zdnd11an1n32x5 FILLER_331_464 ();
 b15zdnd11an1n08x5 FILLER_331_496 ();
 b15zdnd00an1n01x5 FILLER_331_504 ();
 b15zdnd11an1n04x5 FILLER_331_508 ();
 b15zdnd11an1n64x5 FILLER_331_515 ();
 b15zdnd11an1n32x5 FILLER_331_579 ();
 b15zdnd11an1n04x5 FILLER_331_611 ();
 b15zdnd00an1n02x5 FILLER_331_615 ();
 b15zdnd00an1n01x5 FILLER_331_617 ();
 b15zdnd11an1n04x5 FILLER_331_621 ();
 b15zdnd11an1n64x5 FILLER_331_677 ();
 b15zdnd11an1n08x5 FILLER_331_741 ();
 b15zdnd00an1n02x5 FILLER_331_749 ();
 b15zdnd00an1n01x5 FILLER_331_751 ();
 b15zdnd11an1n04x5 FILLER_331_755 ();
 b15zdnd11an1n04x5 FILLER_331_762 ();
 b15zdnd11an1n04x5 FILLER_331_775 ();
 b15zdnd00an1n01x5 FILLER_331_779 ();
 b15zdnd11an1n04x5 FILLER_331_789 ();
 b15zdnd11an1n64x5 FILLER_331_796 ();
 b15zdnd11an1n16x5 FILLER_331_860 ();
 b15zdnd11an1n04x5 FILLER_331_876 ();
 b15zdnd11an1n32x5 FILLER_331_932 ();
 b15zdnd11an1n04x5 FILLER_331_964 ();
 b15zdnd00an1n02x5 FILLER_331_968 ();
 b15zdnd00an1n01x5 FILLER_331_970 ();
 b15zdnd11an1n32x5 FILLER_331_980 ();
 b15zdnd00an1n02x5 FILLER_331_1012 ();
 b15zdnd00an1n01x5 FILLER_331_1014 ();
 b15zdnd11an1n04x5 FILLER_331_1018 ();
 b15zdnd11an1n04x5 FILLER_331_1025 ();
 b15zdnd11an1n04x5 FILLER_331_1032 ();
 b15zdnd11an1n04x5 FILLER_331_1039 ();
 b15zdnd11an1n04x5 FILLER_331_1046 ();
 b15zdnd11an1n64x5 FILLER_331_1053 ();
 b15zdnd11an1n64x5 FILLER_331_1117 ();
 b15zdnd11an1n64x5 FILLER_331_1181 ();
 b15zdnd11an1n32x5 FILLER_331_1245 ();
 b15zdnd11an1n16x5 FILLER_331_1277 ();
 b15zdnd11an1n08x5 FILLER_331_1293 ();
 b15zdnd00an1n02x5 FILLER_331_1301 ();
 b15zdnd00an1n01x5 FILLER_331_1303 ();
 b15zdnd11an1n32x5 FILLER_331_1346 ();
 b15zdnd11an1n16x5 FILLER_331_1378 ();
 b15zdnd11an1n08x5 FILLER_331_1394 ();
 b15zdnd11an1n04x5 FILLER_331_1454 ();
 b15zdnd11an1n04x5 FILLER_331_1467 ();
 b15zdnd11an1n64x5 FILLER_331_1474 ();
 b15zdnd11an1n32x5 FILLER_331_1538 ();
 b15zdnd11an1n16x5 FILLER_331_1570 ();
 b15zdnd11an1n08x5 FILLER_331_1586 ();
 b15zdnd11an1n04x5 FILLER_331_1594 ();
 b15zdnd11an1n32x5 FILLER_331_1640 ();
 b15zdnd11an1n16x5 FILLER_331_1672 ();
 b15zdnd11an1n08x5 FILLER_331_1688 ();
 b15zdnd11an1n04x5 FILLER_331_1696 ();
 b15zdnd00an1n01x5 FILLER_331_1700 ();
 b15zdnd11an1n04x5 FILLER_331_1721 ();
 b15zdnd11an1n64x5 FILLER_331_1777 ();
 b15zdnd11an1n08x5 FILLER_331_1841 ();
 b15zdnd11an1n04x5 FILLER_331_1852 ();
 b15zdnd00an1n02x5 FILLER_331_1856 ();
 b15zdnd11an1n04x5 FILLER_331_1883 ();
 b15zdnd11an1n04x5 FILLER_331_1893 ();
 b15zdnd11an1n64x5 FILLER_331_1900 ();
 b15zdnd11an1n64x5 FILLER_331_1964 ();
 b15zdnd11an1n32x5 FILLER_331_2028 ();
 b15zdnd11an1n04x5 FILLER_331_2102 ();
 b15zdnd11an1n04x5 FILLER_331_2148 ();
 b15zdnd11an1n64x5 FILLER_331_2155 ();
 b15zdnd11an1n64x5 FILLER_331_2219 ();
 b15zdnd00an1n01x5 FILLER_331_2283 ();
 b15zdnd11an1n64x5 FILLER_332_8 ();
 b15zdnd11an1n16x5 FILLER_332_72 ();
 b15zdnd11an1n08x5 FILLER_332_88 ();
 b15zdnd11an1n04x5 FILLER_332_100 ();
 b15zdnd11an1n64x5 FILLER_332_108 ();
 b15zdnd11an1n04x5 FILLER_332_172 ();
 b15zdnd00an1n02x5 FILLER_332_176 ();
 b15zdnd00an1n01x5 FILLER_332_178 ();
 b15zdnd11an1n04x5 FILLER_332_207 ();
 b15zdnd11an1n04x5 FILLER_332_231 ();
 b15zdnd11an1n64x5 FILLER_332_238 ();
 b15zdnd11an1n32x5 FILLER_332_302 ();
 b15zdnd11an1n16x5 FILLER_332_334 ();
 b15zdnd00an1n02x5 FILLER_332_350 ();
 b15zdnd00an1n01x5 FILLER_332_352 ();
 b15zdnd11an1n16x5 FILLER_332_356 ();
 b15zdnd11an1n04x5 FILLER_332_372 ();
 b15zdnd00an1n02x5 FILLER_332_376 ();
 b15zdnd00an1n01x5 FILLER_332_378 ();
 b15zdnd11an1n04x5 FILLER_332_382 ();
 b15zdnd11an1n16x5 FILLER_332_389 ();
 b15zdnd11an1n64x5 FILLER_332_447 ();
 b15zdnd11an1n64x5 FILLER_332_511 ();
 b15zdnd11an1n32x5 FILLER_332_575 ();
 b15zdnd11an1n08x5 FILLER_332_607 ();
 b15zdnd11an1n04x5 FILLER_332_615 ();
 b15zdnd11an1n08x5 FILLER_332_622 ();
 b15zdnd00an1n01x5 FILLER_332_630 ();
 b15zdnd11an1n04x5 FILLER_332_634 ();
 b15zdnd11an1n08x5 FILLER_332_647 ();
 b15zdnd11an1n32x5 FILLER_332_675 ();
 b15zdnd11an1n08x5 FILLER_332_707 ();
 b15zdnd00an1n02x5 FILLER_332_715 ();
 b15zdnd00an1n01x5 FILLER_332_717 ();
 b15zdnd11an1n32x5 FILLER_332_726 ();
 b15zdnd00an1n02x5 FILLER_332_758 ();
 b15zdnd11an1n04x5 FILLER_332_763 ();
 b15zdnd11an1n04x5 FILLER_332_770 ();
 b15zdnd11an1n04x5 FILLER_332_777 ();
 b15zdnd11an1n04x5 FILLER_332_784 ();
 b15zdnd11an1n64x5 FILLER_332_791 ();
 b15zdnd11an1n32x5 FILLER_332_855 ();
 b15zdnd11an1n04x5 FILLER_332_887 ();
 b15zdnd00an1n01x5 FILLER_332_891 ();
 b15zdnd11an1n04x5 FILLER_332_895 ();
 b15zdnd11an1n04x5 FILLER_332_902 ();
 b15zdnd11an1n04x5 FILLER_332_909 ();
 b15zdnd11an1n04x5 FILLER_332_916 ();
 b15zdnd11an1n64x5 FILLER_332_923 ();
 b15zdnd11an1n16x5 FILLER_332_987 ();
 b15zdnd11an1n04x5 FILLER_332_1003 ();
 b15zdnd00an1n02x5 FILLER_332_1007 ();
 b15zdnd00an1n01x5 FILLER_332_1009 ();
 b15zdnd11an1n64x5 FILLER_332_1062 ();
 b15zdnd11an1n64x5 FILLER_332_1126 ();
 b15zdnd11an1n64x5 FILLER_332_1190 ();
 b15zdnd11an1n64x5 FILLER_332_1254 ();
 b15zdnd11an1n64x5 FILLER_332_1318 ();
 b15zdnd11an1n32x5 FILLER_332_1382 ();
 b15zdnd11an1n08x5 FILLER_332_1414 ();
 b15zdnd00an1n02x5 FILLER_332_1422 ();
 b15zdnd00an1n01x5 FILLER_332_1424 ();
 b15zdnd11an1n04x5 FILLER_332_1428 ();
 b15zdnd11an1n04x5 FILLER_332_1441 ();
 b15zdnd11an1n04x5 FILLER_332_1448 ();
 b15zdnd11an1n04x5 FILLER_332_1455 ();
 b15zdnd11an1n08x5 FILLER_332_1462 ();
 b15zdnd00an1n01x5 FILLER_332_1470 ();
 b15zdnd11an1n64x5 FILLER_332_1491 ();
 b15zdnd11an1n32x5 FILLER_332_1555 ();
 b15zdnd11an1n08x5 FILLER_332_1587 ();
 b15zdnd00an1n02x5 FILLER_332_1595 ();
 b15zdnd00an1n01x5 FILLER_332_1597 ();
 b15zdnd11an1n04x5 FILLER_332_1603 ();
 b15zdnd11an1n64x5 FILLER_332_1649 ();
 b15zdnd11an1n08x5 FILLER_332_1713 ();
 b15zdnd11an1n04x5 FILLER_332_1721 ();
 b15zdnd00an1n02x5 FILLER_332_1725 ();
 b15zdnd11an1n64x5 FILLER_332_1769 ();
 b15zdnd11an1n32x5 FILLER_332_1833 ();
 b15zdnd11an1n04x5 FILLER_332_1865 ();
 b15zdnd11an1n64x5 FILLER_332_1911 ();
 b15zdnd11an1n64x5 FILLER_332_1975 ();
 b15zdnd11an1n32x5 FILLER_332_2039 ();
 b15zdnd11an1n16x5 FILLER_332_2113 ();
 b15zdnd00an1n01x5 FILLER_332_2129 ();
 b15zdnd11an1n16x5 FILLER_332_2133 ();
 b15zdnd11an1n04x5 FILLER_332_2149 ();
 b15zdnd00an1n01x5 FILLER_332_2153 ();
 b15zdnd11an1n64x5 FILLER_332_2162 ();
 b15zdnd11an1n32x5 FILLER_332_2226 ();
 b15zdnd11an1n16x5 FILLER_332_2258 ();
 b15zdnd00an1n02x5 FILLER_332_2274 ();
 b15zdnd11an1n16x5 FILLER_333_0 ();
 b15zdnd11an1n04x5 FILLER_333_16 ();
 b15zdnd00an1n02x5 FILLER_333_20 ();
 b15zdnd00an1n01x5 FILLER_333_22 ();
 b15zdnd11an1n04x5 FILLER_333_27 ();
 b15zdnd11an1n64x5 FILLER_333_38 ();
 b15zdnd11an1n64x5 FILLER_333_102 ();
 b15zdnd11an1n16x5 FILLER_333_166 ();
 b15zdnd00an1n02x5 FILLER_333_182 ();
 b15zdnd00an1n01x5 FILLER_333_184 ();
 b15zdnd11an1n04x5 FILLER_333_207 ();
 b15zdnd11an1n64x5 FILLER_333_214 ();
 b15zdnd11an1n64x5 FILLER_333_278 ();
 b15zdnd11an1n64x5 FILLER_333_342 ();
 b15zdnd11an1n64x5 FILLER_333_406 ();
 b15zdnd11an1n64x5 FILLER_333_470 ();
 b15zdnd11an1n64x5 FILLER_333_534 ();
 b15zdnd11an1n16x5 FILLER_333_598 ();
 b15zdnd11an1n08x5 FILLER_333_614 ();
 b15zdnd11an1n04x5 FILLER_333_642 ();
 b15zdnd11an1n04x5 FILLER_333_649 ();
 b15zdnd11an1n64x5 FILLER_333_673 ();
 b15zdnd11an1n32x5 FILLER_333_737 ();
 b15zdnd00an1n02x5 FILLER_333_769 ();
 b15zdnd00an1n01x5 FILLER_333_771 ();
 b15zdnd11an1n04x5 FILLER_333_775 ();
 b15zdnd11an1n64x5 FILLER_333_782 ();
 b15zdnd11an1n32x5 FILLER_333_846 ();
 b15zdnd11an1n16x5 FILLER_333_878 ();
 b15zdnd11an1n04x5 FILLER_333_894 ();
 b15zdnd00an1n02x5 FILLER_333_898 ();
 b15zdnd11an1n04x5 FILLER_333_903 ();
 b15zdnd11an1n16x5 FILLER_333_910 ();
 b15zdnd11an1n04x5 FILLER_333_926 ();
 b15zdnd00an1n02x5 FILLER_333_930 ();
 b15zdnd00an1n01x5 FILLER_333_932 ();
 b15zdnd11an1n64x5 FILLER_333_953 ();
 b15zdnd11an1n64x5 FILLER_333_1069 ();
 b15zdnd11an1n64x5 FILLER_333_1133 ();
 b15zdnd11an1n32x5 FILLER_333_1197 ();
 b15zdnd11an1n16x5 FILLER_333_1229 ();
 b15zdnd11an1n04x5 FILLER_333_1245 ();
 b15zdnd00an1n02x5 FILLER_333_1249 ();
 b15zdnd11an1n64x5 FILLER_333_1293 ();
 b15zdnd11an1n64x5 FILLER_333_1357 ();
 b15zdnd00an1n02x5 FILLER_333_1421 ();
 b15zdnd00an1n01x5 FILLER_333_1423 ();
 b15zdnd11an1n16x5 FILLER_333_1427 ();
 b15zdnd00an1n02x5 FILLER_333_1443 ();
 b15zdnd00an1n01x5 FILLER_333_1445 ();
 b15zdnd11an1n04x5 FILLER_333_1449 ();
 b15zdnd00an1n02x5 FILLER_333_1453 ();
 b15zdnd00an1n01x5 FILLER_333_1455 ();
 b15zdnd11an1n04x5 FILLER_333_1459 ();
 b15zdnd11an1n64x5 FILLER_333_1466 ();
 b15zdnd11an1n64x5 FILLER_333_1530 ();
 b15zdnd11an1n04x5 FILLER_333_1594 ();
 b15zdnd00an1n02x5 FILLER_333_1598 ();
 b15zdnd00an1n01x5 FILLER_333_1600 ();
 b15zdnd11an1n08x5 FILLER_333_1610 ();
 b15zdnd00an1n01x5 FILLER_333_1618 ();
 b15zdnd11an1n32x5 FILLER_333_1661 ();
 b15zdnd11an1n08x5 FILLER_333_1693 ();
 b15zdnd00an1n01x5 FILLER_333_1701 ();
 b15zdnd11an1n04x5 FILLER_333_1744 ();
 b15zdnd00an1n02x5 FILLER_333_1748 ();
 b15zdnd00an1n01x5 FILLER_333_1750 ();
 b15zdnd11an1n64x5 FILLER_333_1754 ();
 b15zdnd11an1n64x5 FILLER_333_1818 ();
 b15zdnd11an1n64x5 FILLER_333_1882 ();
 b15zdnd11an1n64x5 FILLER_333_1946 ();
 b15zdnd11an1n64x5 FILLER_333_2010 ();
 b15zdnd11an1n64x5 FILLER_333_2074 ();
 b15zdnd11an1n64x5 FILLER_333_2138 ();
 b15zdnd11an1n64x5 FILLER_333_2202 ();
 b15zdnd11an1n16x5 FILLER_333_2266 ();
 b15zdnd00an1n02x5 FILLER_333_2282 ();
 b15zdnd00an1n02x5 FILLER_334_8 ();
 b15zdnd11an1n64x5 FILLER_334_52 ();
 b15zdnd11an1n32x5 FILLER_334_116 ();
 b15zdnd11an1n16x5 FILLER_334_148 ();
 b15zdnd11an1n08x5 FILLER_334_164 ();
 b15zdnd11an1n04x5 FILLER_334_172 ();
 b15zdnd11an1n04x5 FILLER_334_196 ();
 b15zdnd11an1n64x5 FILLER_334_203 ();
 b15zdnd11an1n64x5 FILLER_334_267 ();
 b15zdnd11an1n64x5 FILLER_334_331 ();
 b15zdnd11an1n64x5 FILLER_334_395 ();
 b15zdnd11an1n64x5 FILLER_334_459 ();
 b15zdnd11an1n64x5 FILLER_334_523 ();
 b15zdnd11an1n32x5 FILLER_334_587 ();
 b15zdnd11an1n16x5 FILLER_334_619 ();
 b15zdnd11an1n04x5 FILLER_334_635 ();
 b15zdnd00an1n01x5 FILLER_334_639 ();
 b15zdnd11an1n04x5 FILLER_334_643 ();
 b15zdnd11an1n64x5 FILLER_334_650 ();
 b15zdnd11an1n04x5 FILLER_334_714 ();
 b15zdnd11an1n64x5 FILLER_334_726 ();
 b15zdnd11an1n64x5 FILLER_334_790 ();
 b15zdnd11an1n32x5 FILLER_334_854 ();
 b15zdnd11an1n16x5 FILLER_334_886 ();
 b15zdnd11an1n04x5 FILLER_334_902 ();
 b15zdnd11an1n64x5 FILLER_334_909 ();
 b15zdnd11an1n32x5 FILLER_334_973 ();
 b15zdnd11an1n16x5 FILLER_334_1005 ();
 b15zdnd11an1n08x5 FILLER_334_1021 ();
 b15zdnd00an1n01x5 FILLER_334_1029 ();
 b15zdnd11an1n04x5 FILLER_334_1033 ();
 b15zdnd11an1n04x5 FILLER_334_1040 ();
 b15zdnd11an1n04x5 FILLER_334_1047 ();
 b15zdnd11an1n64x5 FILLER_334_1054 ();
 b15zdnd11an1n32x5 FILLER_334_1118 ();
 b15zdnd11an1n08x5 FILLER_334_1150 ();
 b15zdnd11an1n32x5 FILLER_334_1200 ();
 b15zdnd11an1n16x5 FILLER_334_1232 ();
 b15zdnd11an1n04x5 FILLER_334_1248 ();
 b15zdnd11an1n64x5 FILLER_334_1294 ();
 b15zdnd11an1n64x5 FILLER_334_1358 ();
 b15zdnd11an1n64x5 FILLER_334_1422 ();
 b15zdnd11an1n64x5 FILLER_334_1486 ();
 b15zdnd11an1n32x5 FILLER_334_1550 ();
 b15zdnd11an1n16x5 FILLER_334_1582 ();
 b15zdnd11an1n08x5 FILLER_334_1598 ();
 b15zdnd00an1n01x5 FILLER_334_1606 ();
 b15zdnd11an1n04x5 FILLER_334_1612 ();
 b15zdnd11an1n04x5 FILLER_334_1629 ();
 b15zdnd11an1n64x5 FILLER_334_1639 ();
 b15zdnd11an1n64x5 FILLER_334_1703 ();
 b15zdnd11an1n64x5 FILLER_334_1767 ();
 b15zdnd11an1n64x5 FILLER_334_1831 ();
 b15zdnd11an1n64x5 FILLER_334_1895 ();
 b15zdnd11an1n64x5 FILLER_334_1959 ();
 b15zdnd11an1n64x5 FILLER_334_2023 ();
 b15zdnd11an1n64x5 FILLER_334_2087 ();
 b15zdnd00an1n02x5 FILLER_334_2151 ();
 b15zdnd00an1n01x5 FILLER_334_2153 ();
 b15zdnd11an1n64x5 FILLER_334_2162 ();
 b15zdnd11an1n32x5 FILLER_334_2226 ();
 b15zdnd11an1n16x5 FILLER_334_2258 ();
 b15zdnd00an1n02x5 FILLER_334_2274 ();
 b15zdnd11an1n64x5 FILLER_335_0 ();
 b15zdnd11an1n64x5 FILLER_335_64 ();
 b15zdnd11an1n64x5 FILLER_335_128 ();
 b15zdnd11an1n64x5 FILLER_335_192 ();
 b15zdnd11an1n64x5 FILLER_335_256 ();
 b15zdnd11an1n64x5 FILLER_335_320 ();
 b15zdnd11an1n64x5 FILLER_335_384 ();
 b15zdnd11an1n32x5 FILLER_335_448 ();
 b15zdnd00an1n01x5 FILLER_335_480 ();
 b15zdnd11an1n64x5 FILLER_335_523 ();
 b15zdnd11an1n64x5 FILLER_335_587 ();
 b15zdnd11an1n64x5 FILLER_335_651 ();
 b15zdnd11an1n64x5 FILLER_335_715 ();
 b15zdnd11an1n64x5 FILLER_335_779 ();
 b15zdnd11an1n64x5 FILLER_335_843 ();
 b15zdnd11an1n64x5 FILLER_335_907 ();
 b15zdnd11an1n64x5 FILLER_335_971 ();
 b15zdnd11an1n04x5 FILLER_335_1035 ();
 b15zdnd00an1n02x5 FILLER_335_1039 ();
 b15zdnd00an1n01x5 FILLER_335_1041 ();
 b15zdnd11an1n64x5 FILLER_335_1045 ();
 b15zdnd11an1n64x5 FILLER_335_1109 ();
 b15zdnd11an1n64x5 FILLER_335_1173 ();
 b15zdnd11an1n64x5 FILLER_335_1237 ();
 b15zdnd11an1n64x5 FILLER_335_1301 ();
 b15zdnd11an1n64x5 FILLER_335_1365 ();
 b15zdnd11an1n64x5 FILLER_335_1429 ();
 b15zdnd11an1n64x5 FILLER_335_1493 ();
 b15zdnd11an1n32x5 FILLER_335_1557 ();
 b15zdnd11an1n16x5 FILLER_335_1589 ();
 b15zdnd11an1n04x5 FILLER_335_1605 ();
 b15zdnd11an1n04x5 FILLER_335_1612 ();
 b15zdnd00an1n01x5 FILLER_335_1616 ();
 b15zdnd11an1n04x5 FILLER_335_1627 ();
 b15zdnd00an1n01x5 FILLER_335_1631 ();
 b15zdnd11an1n32x5 FILLER_335_1642 ();
 b15zdnd00an1n02x5 FILLER_335_1674 ();
 b15zdnd00an1n01x5 FILLER_335_1676 ();
 b15zdnd11an1n64x5 FILLER_335_1683 ();
 b15zdnd11an1n64x5 FILLER_335_1747 ();
 b15zdnd11an1n64x5 FILLER_335_1811 ();
 b15zdnd11an1n64x5 FILLER_335_1875 ();
 b15zdnd11an1n64x5 FILLER_335_1939 ();
 b15zdnd11an1n64x5 FILLER_335_2003 ();
 b15zdnd11an1n64x5 FILLER_335_2067 ();
 b15zdnd11an1n64x5 FILLER_335_2131 ();
 b15zdnd11an1n64x5 FILLER_335_2195 ();
 b15zdnd11an1n16x5 FILLER_335_2259 ();
 b15zdnd11an1n08x5 FILLER_335_2275 ();
 b15zdnd00an1n01x5 FILLER_335_2283 ();
 b15zdnd11an1n64x5 FILLER_336_8 ();
 b15zdnd11an1n64x5 FILLER_336_72 ();
 b15zdnd11an1n64x5 FILLER_336_136 ();
 b15zdnd11an1n64x5 FILLER_336_200 ();
 b15zdnd11an1n64x5 FILLER_336_264 ();
 b15zdnd11an1n04x5 FILLER_336_328 ();
 b15zdnd11an1n64x5 FILLER_336_374 ();
 b15zdnd11an1n32x5 FILLER_336_438 ();
 b15zdnd11an1n04x5 FILLER_336_470 ();
 b15zdnd00an1n01x5 FILLER_336_474 ();
 b15zdnd11an1n08x5 FILLER_336_517 ();
 b15zdnd11an1n04x5 FILLER_336_525 ();
 b15zdnd00an1n01x5 FILLER_336_529 ();
 b15zdnd11an1n64x5 FILLER_336_572 ();
 b15zdnd11an1n64x5 FILLER_336_636 ();
 b15zdnd11an1n16x5 FILLER_336_700 ();
 b15zdnd00an1n02x5 FILLER_336_716 ();
 b15zdnd11an1n64x5 FILLER_336_726 ();
 b15zdnd11an1n64x5 FILLER_336_790 ();
 b15zdnd11an1n64x5 FILLER_336_854 ();
 b15zdnd11an1n64x5 FILLER_336_918 ();
 b15zdnd11an1n64x5 FILLER_336_982 ();
 b15zdnd11an1n64x5 FILLER_336_1046 ();
 b15zdnd11an1n64x5 FILLER_336_1110 ();
 b15zdnd11an1n32x5 FILLER_336_1174 ();
 b15zdnd11an1n08x5 FILLER_336_1206 ();
 b15zdnd00an1n02x5 FILLER_336_1214 ();
 b15zdnd11an1n64x5 FILLER_336_1258 ();
 b15zdnd11an1n64x5 FILLER_336_1322 ();
 b15zdnd11an1n64x5 FILLER_336_1386 ();
 b15zdnd11an1n64x5 FILLER_336_1450 ();
 b15zdnd11an1n64x5 FILLER_336_1514 ();
 b15zdnd11an1n32x5 FILLER_336_1578 ();
 b15zdnd11an1n08x5 FILLER_336_1610 ();
 b15zdnd00an1n02x5 FILLER_336_1618 ();
 b15zdnd00an1n01x5 FILLER_336_1620 ();
 b15zdnd11an1n64x5 FILLER_336_1625 ();
 b15zdnd11an1n64x5 FILLER_336_1689 ();
 b15zdnd11an1n64x5 FILLER_336_1753 ();
 b15zdnd11an1n64x5 FILLER_336_1817 ();
 b15zdnd11an1n64x5 FILLER_336_1881 ();
 b15zdnd11an1n64x5 FILLER_336_1945 ();
 b15zdnd11an1n64x5 FILLER_336_2009 ();
 b15zdnd11an1n64x5 FILLER_336_2073 ();
 b15zdnd11an1n16x5 FILLER_336_2137 ();
 b15zdnd00an1n01x5 FILLER_336_2153 ();
 b15zdnd11an1n64x5 FILLER_336_2162 ();
 b15zdnd11an1n32x5 FILLER_336_2226 ();
 b15zdnd11an1n16x5 FILLER_336_2258 ();
 b15zdnd00an1n02x5 FILLER_336_2274 ();
 b15zdnd11an1n64x5 FILLER_337_0 ();
 b15zdnd11an1n64x5 FILLER_337_64 ();
 b15zdnd11an1n64x5 FILLER_337_128 ();
 b15zdnd11an1n64x5 FILLER_337_192 ();
 b15zdnd11an1n64x5 FILLER_337_256 ();
 b15zdnd11an1n64x5 FILLER_337_320 ();
 b15zdnd11an1n64x5 FILLER_337_384 ();
 b15zdnd11an1n64x5 FILLER_337_448 ();
 b15zdnd11an1n64x5 FILLER_337_512 ();
 b15zdnd11an1n64x5 FILLER_337_576 ();
 b15zdnd11an1n64x5 FILLER_337_640 ();
 b15zdnd11an1n64x5 FILLER_337_704 ();
 b15zdnd11an1n64x5 FILLER_337_768 ();
 b15zdnd11an1n64x5 FILLER_337_832 ();
 b15zdnd11an1n64x5 FILLER_337_896 ();
 b15zdnd11an1n64x5 FILLER_337_960 ();
 b15zdnd11an1n16x5 FILLER_337_1024 ();
 b15zdnd11an1n04x5 FILLER_337_1040 ();
 b15zdnd00an1n02x5 FILLER_337_1044 ();
 b15zdnd11an1n04x5 FILLER_337_1088 ();
 b15zdnd11an1n64x5 FILLER_337_1134 ();
 b15zdnd11an1n64x5 FILLER_337_1198 ();
 b15zdnd11an1n64x5 FILLER_337_1262 ();
 b15zdnd11an1n64x5 FILLER_337_1326 ();
 b15zdnd11an1n64x5 FILLER_337_1390 ();
 b15zdnd11an1n64x5 FILLER_337_1454 ();
 b15zdnd11an1n64x5 FILLER_337_1518 ();
 b15zdnd11an1n32x5 FILLER_337_1582 ();
 b15zdnd11an1n08x5 FILLER_337_1614 ();
 b15zdnd11an1n04x5 FILLER_337_1622 ();
 b15zdnd00an1n01x5 FILLER_337_1626 ();
 b15zdnd11an1n64x5 FILLER_337_1630 ();
 b15zdnd11an1n64x5 FILLER_337_1694 ();
 b15zdnd11an1n64x5 FILLER_337_1758 ();
 b15zdnd11an1n64x5 FILLER_337_1822 ();
 b15zdnd11an1n64x5 FILLER_337_1886 ();
 b15zdnd11an1n64x5 FILLER_337_1950 ();
 b15zdnd11an1n64x5 FILLER_337_2014 ();
 b15zdnd11an1n64x5 FILLER_337_2078 ();
 b15zdnd11an1n64x5 FILLER_337_2142 ();
 b15zdnd11an1n64x5 FILLER_337_2206 ();
 b15zdnd11an1n08x5 FILLER_337_2270 ();
 b15zdnd11an1n04x5 FILLER_337_2278 ();
 b15zdnd00an1n02x5 FILLER_337_2282 ();
 b15zdnd11an1n64x5 FILLER_338_8 ();
 b15zdnd11an1n64x5 FILLER_338_72 ();
 b15zdnd11an1n64x5 FILLER_338_136 ();
 b15zdnd11an1n64x5 FILLER_338_200 ();
 b15zdnd11an1n64x5 FILLER_338_264 ();
 b15zdnd11an1n64x5 FILLER_338_328 ();
 b15zdnd11an1n64x5 FILLER_338_392 ();
 b15zdnd11an1n08x5 FILLER_338_456 ();
 b15zdnd00an1n02x5 FILLER_338_464 ();
 b15zdnd00an1n01x5 FILLER_338_466 ();
 b15zdnd11an1n64x5 FILLER_338_509 ();
 b15zdnd11an1n64x5 FILLER_338_573 ();
 b15zdnd11an1n64x5 FILLER_338_637 ();
 b15zdnd11an1n16x5 FILLER_338_701 ();
 b15zdnd00an1n01x5 FILLER_338_717 ();
 b15zdnd11an1n64x5 FILLER_338_726 ();
 b15zdnd11an1n64x5 FILLER_338_790 ();
 b15zdnd11an1n64x5 FILLER_338_854 ();
 b15zdnd11an1n64x5 FILLER_338_918 ();
 b15zdnd11an1n64x5 FILLER_338_982 ();
 b15zdnd11an1n08x5 FILLER_338_1046 ();
 b15zdnd00an1n02x5 FILLER_338_1054 ();
 b15zdnd11an1n16x5 FILLER_338_1098 ();
 b15zdnd11an1n08x5 FILLER_338_1114 ();
 b15zdnd11an1n04x5 FILLER_338_1122 ();
 b15zdnd00an1n02x5 FILLER_338_1126 ();
 b15zdnd00an1n01x5 FILLER_338_1128 ();
 b15zdnd11an1n64x5 FILLER_338_1171 ();
 b15zdnd11an1n64x5 FILLER_338_1235 ();
 b15zdnd11an1n64x5 FILLER_338_1299 ();
 b15zdnd11an1n04x5 FILLER_338_1363 ();
 b15zdnd00an1n02x5 FILLER_338_1367 ();
 b15zdnd11an1n64x5 FILLER_338_1411 ();
 b15zdnd11an1n64x5 FILLER_338_1475 ();
 b15zdnd11an1n64x5 FILLER_338_1539 ();
 b15zdnd11an1n64x5 FILLER_338_1603 ();
 b15zdnd11an1n64x5 FILLER_338_1667 ();
 b15zdnd11an1n64x5 FILLER_338_1731 ();
 b15zdnd11an1n64x5 FILLER_338_1795 ();
 b15zdnd11an1n64x5 FILLER_338_1859 ();
 b15zdnd11an1n64x5 FILLER_338_1923 ();
 b15zdnd11an1n64x5 FILLER_338_1987 ();
 b15zdnd11an1n64x5 FILLER_338_2051 ();
 b15zdnd11an1n32x5 FILLER_338_2115 ();
 b15zdnd11an1n04x5 FILLER_338_2147 ();
 b15zdnd00an1n02x5 FILLER_338_2151 ();
 b15zdnd00an1n01x5 FILLER_338_2153 ();
 b15zdnd11an1n64x5 FILLER_338_2162 ();
 b15zdnd11an1n32x5 FILLER_338_2226 ();
 b15zdnd11an1n16x5 FILLER_338_2258 ();
 b15zdnd00an1n02x5 FILLER_338_2274 ();
 b15zdnd11an1n64x5 FILLER_339_0 ();
 b15zdnd11an1n64x5 FILLER_339_64 ();
 b15zdnd11an1n64x5 FILLER_339_128 ();
 b15zdnd11an1n64x5 FILLER_339_192 ();
 b15zdnd11an1n64x5 FILLER_339_256 ();
 b15zdnd00an1n02x5 FILLER_339_320 ();
 b15zdnd11an1n64x5 FILLER_339_328 ();
 b15zdnd11an1n64x5 FILLER_339_392 ();
 b15zdnd11an1n16x5 FILLER_339_456 ();
 b15zdnd00an1n02x5 FILLER_339_472 ();
 b15zdnd00an1n01x5 FILLER_339_474 ();
 b15zdnd11an1n64x5 FILLER_339_517 ();
 b15zdnd11an1n64x5 FILLER_339_581 ();
 b15zdnd11an1n64x5 FILLER_339_645 ();
 b15zdnd11an1n64x5 FILLER_339_709 ();
 b15zdnd11an1n64x5 FILLER_339_773 ();
 b15zdnd11an1n64x5 FILLER_339_837 ();
 b15zdnd11an1n64x5 FILLER_339_901 ();
 b15zdnd11an1n32x5 FILLER_339_965 ();
 b15zdnd11an1n16x5 FILLER_339_997 ();
 b15zdnd11an1n08x5 FILLER_339_1013 ();
 b15zdnd11an1n04x5 FILLER_339_1021 ();
 b15zdnd11an1n16x5 FILLER_339_1067 ();
 b15zdnd11an1n08x5 FILLER_339_1083 ();
 b15zdnd11an1n04x5 FILLER_339_1091 ();
 b15zdnd00an1n01x5 FILLER_339_1095 ();
 b15zdnd11an1n64x5 FILLER_339_1138 ();
 b15zdnd11an1n64x5 FILLER_339_1202 ();
 b15zdnd11an1n64x5 FILLER_339_1266 ();
 b15zdnd11an1n64x5 FILLER_339_1330 ();
 b15zdnd11an1n64x5 FILLER_339_1394 ();
 b15zdnd11an1n64x5 FILLER_339_1458 ();
 b15zdnd11an1n64x5 FILLER_339_1522 ();
 b15zdnd11an1n64x5 FILLER_339_1586 ();
 b15zdnd11an1n64x5 FILLER_339_1650 ();
 b15zdnd11an1n64x5 FILLER_339_1714 ();
 b15zdnd11an1n64x5 FILLER_339_1778 ();
 b15zdnd11an1n64x5 FILLER_339_1842 ();
 b15zdnd11an1n64x5 FILLER_339_1906 ();
 b15zdnd11an1n64x5 FILLER_339_1970 ();
 b15zdnd11an1n64x5 FILLER_339_2034 ();
 b15zdnd11an1n64x5 FILLER_339_2098 ();
 b15zdnd11an1n64x5 FILLER_339_2162 ();
 b15zdnd11an1n32x5 FILLER_339_2226 ();
 b15zdnd11an1n16x5 FILLER_339_2258 ();
 b15zdnd11an1n08x5 FILLER_339_2274 ();
 b15zdnd00an1n02x5 FILLER_339_2282 ();
 b15zdnd11an1n64x5 FILLER_340_8 ();
 b15zdnd11an1n64x5 FILLER_340_72 ();
 b15zdnd11an1n64x5 FILLER_340_136 ();
 b15zdnd11an1n64x5 FILLER_340_200 ();
 b15zdnd11an1n64x5 FILLER_340_264 ();
 b15zdnd11an1n64x5 FILLER_340_328 ();
 b15zdnd11an1n64x5 FILLER_340_392 ();
 b15zdnd11an1n32x5 FILLER_340_456 ();
 b15zdnd00an1n02x5 FILLER_340_488 ();
 b15zdnd11an1n64x5 FILLER_340_532 ();
 b15zdnd11an1n64x5 FILLER_340_596 ();
 b15zdnd11an1n32x5 FILLER_340_660 ();
 b15zdnd11an1n16x5 FILLER_340_692 ();
 b15zdnd11an1n08x5 FILLER_340_708 ();
 b15zdnd00an1n02x5 FILLER_340_716 ();
 b15zdnd11an1n64x5 FILLER_340_726 ();
 b15zdnd11an1n64x5 FILLER_340_790 ();
 b15zdnd11an1n64x5 FILLER_340_854 ();
 b15zdnd11an1n64x5 FILLER_340_918 ();
 b15zdnd11an1n16x5 FILLER_340_982 ();
 b15zdnd11an1n04x5 FILLER_340_998 ();
 b15zdnd00an1n01x5 FILLER_340_1002 ();
 b15zdnd11an1n64x5 FILLER_340_1045 ();
 b15zdnd11an1n32x5 FILLER_340_1109 ();
 b15zdnd11an1n08x5 FILLER_340_1141 ();
 b15zdnd11an1n04x5 FILLER_340_1149 ();
 b15zdnd00an1n01x5 FILLER_340_1153 ();
 b15zdnd11an1n64x5 FILLER_340_1196 ();
 b15zdnd11an1n64x5 FILLER_340_1260 ();
 b15zdnd11an1n64x5 FILLER_340_1324 ();
 b15zdnd11an1n64x5 FILLER_340_1388 ();
 b15zdnd11an1n64x5 FILLER_340_1452 ();
 b15zdnd11an1n64x5 FILLER_340_1516 ();
 b15zdnd11an1n64x5 FILLER_340_1580 ();
 b15zdnd11an1n64x5 FILLER_340_1644 ();
 b15zdnd11an1n64x5 FILLER_340_1708 ();
 b15zdnd11an1n64x5 FILLER_340_1772 ();
 b15zdnd11an1n64x5 FILLER_340_1836 ();
 b15zdnd11an1n64x5 FILLER_340_1900 ();
 b15zdnd11an1n64x5 FILLER_340_1964 ();
 b15zdnd11an1n64x5 FILLER_340_2028 ();
 b15zdnd11an1n32x5 FILLER_340_2092 ();
 b15zdnd11an1n16x5 FILLER_340_2124 ();
 b15zdnd11an1n08x5 FILLER_340_2140 ();
 b15zdnd11an1n04x5 FILLER_340_2148 ();
 b15zdnd00an1n02x5 FILLER_340_2152 ();
 b15zdnd11an1n64x5 FILLER_340_2162 ();
 b15zdnd11an1n32x5 FILLER_340_2226 ();
 b15zdnd11an1n16x5 FILLER_340_2258 ();
 b15zdnd00an1n02x5 FILLER_340_2274 ();
 b15zdnd11an1n64x5 FILLER_341_0 ();
 b15zdnd11an1n64x5 FILLER_341_64 ();
 b15zdnd11an1n64x5 FILLER_341_128 ();
 b15zdnd11an1n64x5 FILLER_341_192 ();
 b15zdnd11an1n64x5 FILLER_341_256 ();
 b15zdnd11an1n64x5 FILLER_341_320 ();
 b15zdnd11an1n16x5 FILLER_341_384 ();
 b15zdnd11an1n08x5 FILLER_341_400 ();
 b15zdnd11an1n04x5 FILLER_341_408 ();
 b15zdnd00an1n01x5 FILLER_341_412 ();
 b15zdnd11an1n32x5 FILLER_341_455 ();
 b15zdnd11an1n04x5 FILLER_341_487 ();
 b15zdnd00an1n01x5 FILLER_341_491 ();
 b15zdnd11an1n64x5 FILLER_341_534 ();
 b15zdnd11an1n16x5 FILLER_341_598 ();
 b15zdnd11an1n08x5 FILLER_341_614 ();
 b15zdnd00an1n02x5 FILLER_341_622 ();
 b15zdnd11an1n04x5 FILLER_341_666 ();
 b15zdnd00an1n01x5 FILLER_341_670 ();
 b15zdnd11an1n64x5 FILLER_341_713 ();
 b15zdnd11an1n64x5 FILLER_341_777 ();
 b15zdnd11an1n64x5 FILLER_341_841 ();
 b15zdnd11an1n64x5 FILLER_341_905 ();
 b15zdnd11an1n64x5 FILLER_341_969 ();
 b15zdnd11an1n16x5 FILLER_341_1033 ();
 b15zdnd11an1n08x5 FILLER_341_1049 ();
 b15zdnd11an1n04x5 FILLER_341_1057 ();
 b15zdnd11an1n64x5 FILLER_341_1103 ();
 b15zdnd11an1n64x5 FILLER_341_1167 ();
 b15zdnd11an1n64x5 FILLER_341_1231 ();
 b15zdnd11an1n64x5 FILLER_341_1295 ();
 b15zdnd11an1n64x5 FILLER_341_1359 ();
 b15zdnd11an1n64x5 FILLER_341_1423 ();
 b15zdnd11an1n64x5 FILLER_341_1487 ();
 b15zdnd11an1n64x5 FILLER_341_1551 ();
 b15zdnd11an1n64x5 FILLER_341_1615 ();
 b15zdnd11an1n64x5 FILLER_341_1679 ();
 b15zdnd11an1n64x5 FILLER_341_1743 ();
 b15zdnd11an1n64x5 FILLER_341_1807 ();
 b15zdnd11an1n64x5 FILLER_341_1871 ();
 b15zdnd11an1n64x5 FILLER_341_1935 ();
 b15zdnd11an1n64x5 FILLER_341_1999 ();
 b15zdnd11an1n64x5 FILLER_341_2063 ();
 b15zdnd11an1n64x5 FILLER_341_2127 ();
 b15zdnd11an1n64x5 FILLER_341_2191 ();
 b15zdnd11an1n16x5 FILLER_341_2255 ();
 b15zdnd11an1n08x5 FILLER_341_2271 ();
 b15zdnd11an1n04x5 FILLER_341_2279 ();
 b15zdnd00an1n01x5 FILLER_341_2283 ();
 b15zdnd11an1n64x5 FILLER_342_8 ();
 b15zdnd11an1n64x5 FILLER_342_72 ();
 b15zdnd11an1n64x5 FILLER_342_136 ();
 b15zdnd11an1n64x5 FILLER_342_200 ();
 b15zdnd11an1n64x5 FILLER_342_264 ();
 b15zdnd11an1n64x5 FILLER_342_328 ();
 b15zdnd11an1n64x5 FILLER_342_392 ();
 b15zdnd11an1n16x5 FILLER_342_456 ();
 b15zdnd11an1n04x5 FILLER_342_472 ();
 b15zdnd00an1n02x5 FILLER_342_476 ();
 b15zdnd11an1n64x5 FILLER_342_520 ();
 b15zdnd11an1n16x5 FILLER_342_584 ();
 b15zdnd11an1n08x5 FILLER_342_600 ();
 b15zdnd00an1n02x5 FILLER_342_608 ();
 b15zdnd11an1n04x5 FILLER_342_652 ();
 b15zdnd11an1n16x5 FILLER_342_698 ();
 b15zdnd11an1n04x5 FILLER_342_714 ();
 b15zdnd00an1n02x5 FILLER_342_726 ();
 b15zdnd11an1n64x5 FILLER_342_770 ();
 b15zdnd11an1n64x5 FILLER_342_834 ();
 b15zdnd11an1n64x5 FILLER_342_898 ();
 b15zdnd11an1n64x5 FILLER_342_962 ();
 b15zdnd11an1n64x5 FILLER_342_1026 ();
 b15zdnd00an1n02x5 FILLER_342_1090 ();
 b15zdnd11an1n64x5 FILLER_342_1134 ();
 b15zdnd11an1n64x5 FILLER_342_1198 ();
 b15zdnd11an1n16x5 FILLER_342_1262 ();
 b15zdnd11an1n08x5 FILLER_342_1278 ();
 b15zdnd00an1n01x5 FILLER_342_1286 ();
 b15zdnd11an1n16x5 FILLER_342_1329 ();
 b15zdnd11an1n08x5 FILLER_342_1345 ();
 b15zdnd11an1n32x5 FILLER_342_1356 ();
 b15zdnd11an1n16x5 FILLER_342_1388 ();
 b15zdnd11an1n64x5 FILLER_342_1446 ();
 b15zdnd11an1n64x5 FILLER_342_1510 ();
 b15zdnd11an1n64x5 FILLER_342_1574 ();
 b15zdnd11an1n64x5 FILLER_342_1638 ();
 b15zdnd11an1n64x5 FILLER_342_1702 ();
 b15zdnd11an1n64x5 FILLER_342_1766 ();
 b15zdnd11an1n64x5 FILLER_342_1830 ();
 b15zdnd11an1n64x5 FILLER_342_1894 ();
 b15zdnd11an1n64x5 FILLER_342_1958 ();
 b15zdnd11an1n64x5 FILLER_342_2022 ();
 b15zdnd11an1n64x5 FILLER_342_2086 ();
 b15zdnd11an1n04x5 FILLER_342_2150 ();
 b15zdnd11an1n64x5 FILLER_342_2162 ();
 b15zdnd11an1n32x5 FILLER_342_2226 ();
 b15zdnd11an1n16x5 FILLER_342_2258 ();
 b15zdnd00an1n02x5 FILLER_342_2274 ();
 b15zdnd11an1n64x5 FILLER_343_0 ();
 b15zdnd11an1n64x5 FILLER_343_64 ();
 b15zdnd11an1n64x5 FILLER_343_128 ();
 b15zdnd11an1n64x5 FILLER_343_192 ();
 b15zdnd11an1n64x5 FILLER_343_256 ();
 b15zdnd00an1n01x5 FILLER_343_320 ();
 b15zdnd11an1n16x5 FILLER_343_325 ();
 b15zdnd00an1n02x5 FILLER_343_341 ();
 b15zdnd00an1n01x5 FILLER_343_343 ();
 b15zdnd11an1n64x5 FILLER_343_386 ();
 b15zdnd11an1n16x5 FILLER_343_450 ();
 b15zdnd11an1n08x5 FILLER_343_466 ();
 b15zdnd00an1n01x5 FILLER_343_474 ();
 b15zdnd11an1n16x5 FILLER_343_517 ();
 b15zdnd11an1n04x5 FILLER_343_533 ();
 b15zdnd00an1n02x5 FILLER_343_537 ();
 b15zdnd11an1n64x5 FILLER_343_581 ();
 b15zdnd11an1n32x5 FILLER_343_645 ();
 b15zdnd11an1n16x5 FILLER_343_677 ();
 b15zdnd11an1n04x5 FILLER_343_693 ();
 b15zdnd00an1n01x5 FILLER_343_697 ();
 b15zdnd11an1n08x5 FILLER_343_740 ();
 b15zdnd00an1n02x5 FILLER_343_748 ();
 b15zdnd00an1n01x5 FILLER_343_750 ();
 b15zdnd11an1n32x5 FILLER_343_793 ();
 b15zdnd11an1n08x5 FILLER_343_825 ();
 b15zdnd00an1n02x5 FILLER_343_833 ();
 b15zdnd11an1n64x5 FILLER_343_877 ();
 b15zdnd11an1n64x5 FILLER_343_941 ();
 b15zdnd11an1n32x5 FILLER_343_1005 ();
 b15zdnd11an1n08x5 FILLER_343_1037 ();
 b15zdnd11an1n04x5 FILLER_343_1045 ();
 b15zdnd11an1n64x5 FILLER_343_1091 ();
 b15zdnd11an1n64x5 FILLER_343_1155 ();
 b15zdnd11an1n32x5 FILLER_343_1219 ();
 b15zdnd11an1n16x5 FILLER_343_1251 ();
 b15zdnd11an1n08x5 FILLER_343_1267 ();
 b15zdnd00an1n01x5 FILLER_343_1275 ();
 b15zdnd11an1n64x5 FILLER_343_1318 ();
 b15zdnd11an1n32x5 FILLER_343_1382 ();
 b15zdnd11an1n16x5 FILLER_343_1414 ();
 b15zdnd11an1n08x5 FILLER_343_1430 ();
 b15zdnd00an1n01x5 FILLER_343_1438 ();
 b15zdnd11an1n64x5 FILLER_343_1481 ();
 b15zdnd11an1n64x5 FILLER_343_1545 ();
 b15zdnd11an1n64x5 FILLER_343_1609 ();
 b15zdnd11an1n64x5 FILLER_343_1673 ();
 b15zdnd11an1n64x5 FILLER_343_1737 ();
 b15zdnd11an1n64x5 FILLER_343_1801 ();
 b15zdnd11an1n64x5 FILLER_343_1865 ();
 b15zdnd11an1n64x5 FILLER_343_1929 ();
 b15zdnd11an1n64x5 FILLER_343_1993 ();
 b15zdnd11an1n64x5 FILLER_343_2057 ();
 b15zdnd11an1n64x5 FILLER_343_2121 ();
 b15zdnd11an1n64x5 FILLER_343_2185 ();
 b15zdnd11an1n32x5 FILLER_343_2249 ();
 b15zdnd00an1n02x5 FILLER_343_2281 ();
 b15zdnd00an1n01x5 FILLER_343_2283 ();
 b15zdnd11an1n64x5 FILLER_344_8 ();
 b15zdnd11an1n64x5 FILLER_344_72 ();
 b15zdnd11an1n64x5 FILLER_344_136 ();
 b15zdnd11an1n08x5 FILLER_344_200 ();
 b15zdnd11an1n04x5 FILLER_344_208 ();
 b15zdnd11an1n64x5 FILLER_344_254 ();
 b15zdnd11an1n64x5 FILLER_344_318 ();
 b15zdnd11an1n64x5 FILLER_344_382 ();
 b15zdnd11an1n16x5 FILLER_344_446 ();
 b15zdnd11an1n04x5 FILLER_344_462 ();
 b15zdnd00an1n02x5 FILLER_344_466 ();
 b15zdnd11an1n64x5 FILLER_344_510 ();
 b15zdnd11an1n64x5 FILLER_344_574 ();
 b15zdnd11an1n16x5 FILLER_344_638 ();
 b15zdnd11an1n04x5 FILLER_344_654 ();
 b15zdnd00an1n02x5 FILLER_344_658 ();
 b15zdnd00an1n01x5 FILLER_344_660 ();
 b15zdnd11an1n08x5 FILLER_344_703 ();
 b15zdnd11an1n04x5 FILLER_344_711 ();
 b15zdnd00an1n02x5 FILLER_344_715 ();
 b15zdnd00an1n01x5 FILLER_344_717 ();
 b15zdnd00an1n02x5 FILLER_344_726 ();
 b15zdnd11an1n64x5 FILLER_344_770 ();
 b15zdnd11an1n16x5 FILLER_344_834 ();
 b15zdnd11an1n08x5 FILLER_344_850 ();
 b15zdnd00an1n02x5 FILLER_344_858 ();
 b15zdnd11an1n64x5 FILLER_344_902 ();
 b15zdnd11an1n64x5 FILLER_344_966 ();
 b15zdnd11an1n16x5 FILLER_344_1030 ();
 b15zdnd11an1n04x5 FILLER_344_1046 ();
 b15zdnd11an1n64x5 FILLER_344_1092 ();
 b15zdnd11an1n64x5 FILLER_344_1156 ();
 b15zdnd11an1n32x5 FILLER_344_1220 ();
 b15zdnd11an1n08x5 FILLER_344_1252 ();
 b15zdnd11an1n04x5 FILLER_344_1260 ();
 b15zdnd11an1n16x5 FILLER_344_1306 ();
 b15zdnd11an1n08x5 FILLER_344_1322 ();
 b15zdnd00an1n02x5 FILLER_344_1330 ();
 b15zdnd11an1n64x5 FILLER_344_1373 ();
 b15zdnd11an1n64x5 FILLER_344_1437 ();
 b15zdnd11an1n64x5 FILLER_344_1501 ();
 b15zdnd11an1n64x5 FILLER_344_1565 ();
 b15zdnd11an1n64x5 FILLER_344_1629 ();
 b15zdnd11an1n64x5 FILLER_344_1693 ();
 b15zdnd11an1n64x5 FILLER_344_1757 ();
 b15zdnd11an1n64x5 FILLER_344_1821 ();
 b15zdnd11an1n64x5 FILLER_344_1885 ();
 b15zdnd11an1n64x5 FILLER_344_1949 ();
 b15zdnd11an1n64x5 FILLER_344_2013 ();
 b15zdnd11an1n64x5 FILLER_344_2077 ();
 b15zdnd11an1n08x5 FILLER_344_2141 ();
 b15zdnd11an1n04x5 FILLER_344_2149 ();
 b15zdnd00an1n01x5 FILLER_344_2153 ();
 b15zdnd11an1n64x5 FILLER_344_2162 ();
 b15zdnd11an1n32x5 FILLER_344_2226 ();
 b15zdnd11an1n16x5 FILLER_344_2258 ();
 b15zdnd00an1n02x5 FILLER_344_2274 ();
 b15zdnd11an1n64x5 FILLER_345_0 ();
 b15zdnd11an1n64x5 FILLER_345_64 ();
 b15zdnd11an1n64x5 FILLER_345_128 ();
 b15zdnd11an1n64x5 FILLER_345_192 ();
 b15zdnd11an1n64x5 FILLER_345_256 ();
 b15zdnd11an1n32x5 FILLER_345_320 ();
 b15zdnd11an1n16x5 FILLER_345_352 ();
 b15zdnd11an1n08x5 FILLER_345_368 ();
 b15zdnd00an1n01x5 FILLER_345_376 ();
 b15zdnd11an1n32x5 FILLER_345_419 ();
 b15zdnd11an1n04x5 FILLER_345_451 ();
 b15zdnd00an1n01x5 FILLER_345_455 ();
 b15zdnd11an1n64x5 FILLER_345_498 ();
 b15zdnd11an1n64x5 FILLER_345_562 ();
 b15zdnd11an1n64x5 FILLER_345_626 ();
 b15zdnd11an1n64x5 FILLER_345_690 ();
 b15zdnd11an1n64x5 FILLER_345_754 ();
 b15zdnd11an1n64x5 FILLER_345_818 ();
 b15zdnd11an1n64x5 FILLER_345_882 ();
 b15zdnd11an1n64x5 FILLER_345_946 ();
 b15zdnd11an1n32x5 FILLER_345_1010 ();
 b15zdnd11an1n16x5 FILLER_345_1042 ();
 b15zdnd11an1n08x5 FILLER_345_1058 ();
 b15zdnd11an1n04x5 FILLER_345_1066 ();
 b15zdnd00an1n01x5 FILLER_345_1070 ();
 b15zdnd11an1n32x5 FILLER_345_1113 ();
 b15zdnd11an1n16x5 FILLER_345_1145 ();
 b15zdnd11an1n04x5 FILLER_345_1161 ();
 b15zdnd00an1n02x5 FILLER_345_1165 ();
 b15zdnd11an1n32x5 FILLER_345_1172 ();
 b15zdnd11an1n04x5 FILLER_345_1204 ();
 b15zdnd00an1n01x5 FILLER_345_1208 ();
 b15zdnd11an1n64x5 FILLER_345_1251 ();
 b15zdnd11an1n16x5 FILLER_345_1315 ();
 b15zdnd11an1n08x5 FILLER_345_1331 ();
 b15zdnd00an1n02x5 FILLER_345_1339 ();
 b15zdnd00an1n01x5 FILLER_345_1341 ();
 b15zdnd11an1n64x5 FILLER_345_1383 ();
 b15zdnd11an1n64x5 FILLER_345_1447 ();
 b15zdnd11an1n64x5 FILLER_345_1511 ();
 b15zdnd11an1n64x5 FILLER_345_1575 ();
 b15zdnd11an1n64x5 FILLER_345_1639 ();
 b15zdnd11an1n64x5 FILLER_345_1703 ();
 b15zdnd11an1n64x5 FILLER_345_1767 ();
 b15zdnd11an1n64x5 FILLER_345_1831 ();
 b15zdnd11an1n64x5 FILLER_345_1895 ();
 b15zdnd11an1n64x5 FILLER_345_1959 ();
 b15zdnd11an1n64x5 FILLER_345_2023 ();
 b15zdnd11an1n64x5 FILLER_345_2087 ();
 b15zdnd11an1n64x5 FILLER_345_2151 ();
 b15zdnd11an1n64x5 FILLER_345_2215 ();
 b15zdnd11an1n04x5 FILLER_345_2279 ();
 b15zdnd00an1n01x5 FILLER_345_2283 ();
 b15zdnd11an1n64x5 FILLER_346_8 ();
 b15zdnd11an1n64x5 FILLER_346_72 ();
 b15zdnd11an1n64x5 FILLER_346_136 ();
 b15zdnd11an1n64x5 FILLER_346_200 ();
 b15zdnd11an1n64x5 FILLER_346_264 ();
 b15zdnd00an1n01x5 FILLER_346_328 ();
 b15zdnd11an1n64x5 FILLER_346_338 ();
 b15zdnd11an1n64x5 FILLER_346_402 ();
 b15zdnd11an1n64x5 FILLER_346_466 ();
 b15zdnd11an1n64x5 FILLER_346_530 ();
 b15zdnd11an1n64x5 FILLER_346_594 ();
 b15zdnd11an1n32x5 FILLER_346_658 ();
 b15zdnd11an1n16x5 FILLER_346_690 ();
 b15zdnd11an1n08x5 FILLER_346_706 ();
 b15zdnd11an1n04x5 FILLER_346_714 ();
 b15zdnd11an1n64x5 FILLER_346_726 ();
 b15zdnd11an1n64x5 FILLER_346_790 ();
 b15zdnd11an1n64x5 FILLER_346_854 ();
 b15zdnd11an1n64x5 FILLER_346_918 ();
 b15zdnd11an1n32x5 FILLER_346_982 ();
 b15zdnd00an1n02x5 FILLER_346_1014 ();
 b15zdnd00an1n01x5 FILLER_346_1016 ();
 b15zdnd11an1n16x5 FILLER_346_1059 ();
 b15zdnd11an1n32x5 FILLER_346_1117 ();
 b15zdnd11an1n16x5 FILLER_346_1149 ();
 b15zdnd00an1n02x5 FILLER_346_1165 ();
 b15zdnd00an1n01x5 FILLER_346_1167 ();
 b15zdnd11an1n64x5 FILLER_346_1175 ();
 b15zdnd11an1n64x5 FILLER_346_1239 ();
 b15zdnd11an1n32x5 FILLER_346_1303 ();
 b15zdnd11an1n16x5 FILLER_346_1335 ();
 b15zdnd11an1n08x5 FILLER_346_1351 ();
 b15zdnd11an1n04x5 FILLER_346_1381 ();
 b15zdnd11an1n64x5 FILLER_346_1406 ();
 b15zdnd11an1n64x5 FILLER_346_1470 ();
 b15zdnd11an1n64x5 FILLER_346_1534 ();
 b15zdnd11an1n64x5 FILLER_346_1598 ();
 b15zdnd11an1n64x5 FILLER_346_1662 ();
 b15zdnd11an1n64x5 FILLER_346_1726 ();
 b15zdnd11an1n64x5 FILLER_346_1790 ();
 b15zdnd11an1n64x5 FILLER_346_1854 ();
 b15zdnd11an1n64x5 FILLER_346_1918 ();
 b15zdnd11an1n64x5 FILLER_346_1982 ();
 b15zdnd11an1n64x5 FILLER_346_2046 ();
 b15zdnd11an1n32x5 FILLER_346_2110 ();
 b15zdnd11an1n08x5 FILLER_346_2142 ();
 b15zdnd11an1n04x5 FILLER_346_2150 ();
 b15zdnd11an1n64x5 FILLER_346_2162 ();
 b15zdnd11an1n32x5 FILLER_346_2226 ();
 b15zdnd11an1n16x5 FILLER_346_2258 ();
 b15zdnd00an1n02x5 FILLER_346_2274 ();
 b15zdnd11an1n64x5 FILLER_347_0 ();
 b15zdnd11an1n64x5 FILLER_347_64 ();
 b15zdnd11an1n64x5 FILLER_347_128 ();
 b15zdnd11an1n64x5 FILLER_347_192 ();
 b15zdnd11an1n64x5 FILLER_347_256 ();
 b15zdnd11an1n08x5 FILLER_347_320 ();
 b15zdnd11an1n04x5 FILLER_347_328 ();
 b15zdnd00an1n02x5 FILLER_347_332 ();
 b15zdnd11an1n64x5 FILLER_347_343 ();
 b15zdnd11an1n64x5 FILLER_347_407 ();
 b15zdnd11an1n32x5 FILLER_347_471 ();
 b15zdnd11an1n16x5 FILLER_347_503 ();
 b15zdnd00an1n02x5 FILLER_347_519 ();
 b15zdnd11an1n64x5 FILLER_347_563 ();
 b15zdnd11an1n64x5 FILLER_347_627 ();
 b15zdnd11an1n64x5 FILLER_347_691 ();
 b15zdnd11an1n64x5 FILLER_347_755 ();
 b15zdnd11an1n32x5 FILLER_347_819 ();
 b15zdnd11an1n04x5 FILLER_347_851 ();
 b15zdnd00an1n02x5 FILLER_347_855 ();
 b15zdnd00an1n01x5 FILLER_347_857 ();
 b15zdnd11an1n64x5 FILLER_347_900 ();
 b15zdnd11an1n64x5 FILLER_347_964 ();
 b15zdnd11an1n64x5 FILLER_347_1028 ();
 b15zdnd11an1n08x5 FILLER_347_1092 ();
 b15zdnd00an1n02x5 FILLER_347_1100 ();
 b15zdnd00an1n01x5 FILLER_347_1102 ();
 b15zdnd11an1n16x5 FILLER_347_1145 ();
 b15zdnd00an1n02x5 FILLER_347_1161 ();
 b15zdnd00an1n01x5 FILLER_347_1163 ();
 b15zdnd11an1n04x5 FILLER_347_1188 ();
 b15zdnd00an1n02x5 FILLER_347_1192 ();
 b15zdnd11an1n16x5 FILLER_347_1204 ();
 b15zdnd11an1n04x5 FILLER_347_1225 ();
 b15zdnd00an1n01x5 FILLER_347_1229 ();
 b15zdnd11an1n64x5 FILLER_347_1234 ();
 b15zdnd11an1n64x5 FILLER_347_1298 ();
 b15zdnd11an1n64x5 FILLER_347_1362 ();
 b15zdnd11an1n64x5 FILLER_347_1426 ();
 b15zdnd11an1n64x5 FILLER_347_1490 ();
 b15zdnd11an1n64x5 FILLER_347_1554 ();
 b15zdnd11an1n64x5 FILLER_347_1618 ();
 b15zdnd11an1n64x5 FILLER_347_1682 ();
 b15zdnd11an1n64x5 FILLER_347_1746 ();
 b15zdnd11an1n64x5 FILLER_347_1810 ();
 b15zdnd11an1n64x5 FILLER_347_1874 ();
 b15zdnd11an1n64x5 FILLER_347_1938 ();
 b15zdnd11an1n64x5 FILLER_347_2002 ();
 b15zdnd11an1n64x5 FILLER_347_2066 ();
 b15zdnd11an1n64x5 FILLER_347_2130 ();
 b15zdnd11an1n64x5 FILLER_347_2194 ();
 b15zdnd11an1n16x5 FILLER_347_2258 ();
 b15zdnd11an1n08x5 FILLER_347_2274 ();
 b15zdnd00an1n02x5 FILLER_347_2282 ();
 b15zdnd11an1n64x5 FILLER_348_8 ();
 b15zdnd11an1n64x5 FILLER_348_72 ();
 b15zdnd11an1n64x5 FILLER_348_136 ();
 b15zdnd11an1n64x5 FILLER_348_200 ();
 b15zdnd11an1n64x5 FILLER_348_264 ();
 b15zdnd11an1n64x5 FILLER_348_328 ();
 b15zdnd11an1n32x5 FILLER_348_392 ();
 b15zdnd11an1n16x5 FILLER_348_424 ();
 b15zdnd11an1n08x5 FILLER_348_440 ();
 b15zdnd11an1n64x5 FILLER_348_493 ();
 b15zdnd11an1n64x5 FILLER_348_557 ();
 b15zdnd11an1n64x5 FILLER_348_621 ();
 b15zdnd11an1n32x5 FILLER_348_685 ();
 b15zdnd00an1n01x5 FILLER_348_717 ();
 b15zdnd11an1n64x5 FILLER_348_726 ();
 b15zdnd11an1n64x5 FILLER_348_790 ();
 b15zdnd11an1n64x5 FILLER_348_854 ();
 b15zdnd11an1n64x5 FILLER_348_918 ();
 b15zdnd11an1n64x5 FILLER_348_982 ();
 b15zdnd11an1n64x5 FILLER_348_1046 ();
 b15zdnd11an1n16x5 FILLER_348_1110 ();
 b15zdnd11an1n08x5 FILLER_348_1126 ();
 b15zdnd00an1n01x5 FILLER_348_1134 ();
 b15zdnd11an1n08x5 FILLER_348_1177 ();
 b15zdnd11an1n04x5 FILLER_348_1185 ();
 b15zdnd00an1n02x5 FILLER_348_1189 ();
 b15zdnd00an1n01x5 FILLER_348_1191 ();
 b15zdnd11an1n32x5 FILLER_348_1199 ();
 b15zdnd11an1n08x5 FILLER_348_1231 ();
 b15zdnd11an1n64x5 FILLER_348_1245 ();
 b15zdnd11an1n32x5 FILLER_348_1309 ();
 b15zdnd11an1n16x5 FILLER_348_1341 ();
 b15zdnd11an1n04x5 FILLER_348_1357 ();
 b15zdnd00an1n01x5 FILLER_348_1361 ();
 b15zdnd11an1n64x5 FILLER_348_1385 ();
 b15zdnd11an1n64x5 FILLER_348_1449 ();
 b15zdnd11an1n64x5 FILLER_348_1513 ();
 b15zdnd11an1n64x5 FILLER_348_1577 ();
 b15zdnd11an1n64x5 FILLER_348_1641 ();
 b15zdnd11an1n64x5 FILLER_348_1705 ();
 b15zdnd11an1n64x5 FILLER_348_1769 ();
 b15zdnd11an1n64x5 FILLER_348_1833 ();
 b15zdnd11an1n64x5 FILLER_348_1897 ();
 b15zdnd11an1n64x5 FILLER_348_1961 ();
 b15zdnd11an1n64x5 FILLER_348_2025 ();
 b15zdnd11an1n64x5 FILLER_348_2089 ();
 b15zdnd00an1n01x5 FILLER_348_2153 ();
 b15zdnd11an1n64x5 FILLER_348_2162 ();
 b15zdnd11an1n32x5 FILLER_348_2226 ();
 b15zdnd11an1n16x5 FILLER_348_2258 ();
 b15zdnd00an1n02x5 FILLER_348_2274 ();
 b15zdnd11an1n64x5 FILLER_349_0 ();
 b15zdnd11an1n64x5 FILLER_349_64 ();
 b15zdnd11an1n64x5 FILLER_349_128 ();
 b15zdnd11an1n64x5 FILLER_349_192 ();
 b15zdnd11an1n32x5 FILLER_349_256 ();
 b15zdnd11an1n08x5 FILLER_349_288 ();
 b15zdnd11an1n04x5 FILLER_349_296 ();
 b15zdnd00an1n02x5 FILLER_349_300 ();
 b15zdnd00an1n01x5 FILLER_349_302 ();
 b15zdnd11an1n04x5 FILLER_349_326 ();
 b15zdnd11an1n08x5 FILLER_349_346 ();
 b15zdnd00an1n02x5 FILLER_349_354 ();
 b15zdnd11an1n32x5 FILLER_349_379 ();
 b15zdnd11an1n16x5 FILLER_349_411 ();
 b15zdnd11an1n08x5 FILLER_349_427 ();
 b15zdnd00an1n02x5 FILLER_349_435 ();
 b15zdnd00an1n01x5 FILLER_349_437 ();
 b15zdnd11an1n16x5 FILLER_349_443 ();
 b15zdnd11an1n08x5 FILLER_349_459 ();
 b15zdnd00an1n02x5 FILLER_349_467 ();
 b15zdnd00an1n01x5 FILLER_349_469 ();
 b15zdnd11an1n04x5 FILLER_349_480 ();
 b15zdnd11an1n04x5 FILLER_349_494 ();
 b15zdnd11an1n16x5 FILLER_349_502 ();
 b15zdnd11an1n04x5 FILLER_349_518 ();
 b15zdnd00an1n01x5 FILLER_349_522 ();
 b15zdnd11an1n64x5 FILLER_349_529 ();
 b15zdnd11an1n64x5 FILLER_349_593 ();
 b15zdnd11an1n64x5 FILLER_349_657 ();
 b15zdnd11an1n64x5 FILLER_349_721 ();
 b15zdnd11an1n64x5 FILLER_349_785 ();
 b15zdnd11an1n64x5 FILLER_349_849 ();
 b15zdnd11an1n64x5 FILLER_349_913 ();
 b15zdnd11an1n08x5 FILLER_349_977 ();
 b15zdnd00an1n02x5 FILLER_349_985 ();
 b15zdnd00an1n01x5 FILLER_349_987 ();
 b15zdnd11an1n64x5 FILLER_349_1030 ();
 b15zdnd11an1n04x5 FILLER_349_1094 ();
 b15zdnd00an1n02x5 FILLER_349_1098 ();
 b15zdnd00an1n01x5 FILLER_349_1100 ();
 b15zdnd11an1n08x5 FILLER_349_1143 ();
 b15zdnd11an1n04x5 FILLER_349_1151 ();
 b15zdnd00an1n02x5 FILLER_349_1155 ();
 b15zdnd11an1n32x5 FILLER_349_1167 ();
 b15zdnd11an1n16x5 FILLER_349_1199 ();
 b15zdnd11an1n08x5 FILLER_349_1215 ();
 b15zdnd11an1n04x5 FILLER_349_1223 ();
 b15zdnd00an1n02x5 FILLER_349_1227 ();
 b15zdnd00an1n01x5 FILLER_349_1229 ();
 b15zdnd11an1n64x5 FILLER_349_1250 ();
 b15zdnd11an1n64x5 FILLER_349_1314 ();
 b15zdnd11an1n64x5 FILLER_349_1378 ();
 b15zdnd11an1n64x5 FILLER_349_1442 ();
 b15zdnd11an1n64x5 FILLER_349_1506 ();
 b15zdnd11an1n64x5 FILLER_349_1570 ();
 b15zdnd11an1n64x5 FILLER_349_1634 ();
 b15zdnd11an1n64x5 FILLER_349_1698 ();
 b15zdnd11an1n64x5 FILLER_349_1762 ();
 b15zdnd11an1n64x5 FILLER_349_1826 ();
 b15zdnd11an1n64x5 FILLER_349_1890 ();
 b15zdnd11an1n64x5 FILLER_349_1954 ();
 b15zdnd11an1n64x5 FILLER_349_2018 ();
 b15zdnd11an1n64x5 FILLER_349_2082 ();
 b15zdnd11an1n64x5 FILLER_349_2146 ();
 b15zdnd11an1n64x5 FILLER_349_2210 ();
 b15zdnd11an1n08x5 FILLER_349_2274 ();
 b15zdnd00an1n02x5 FILLER_349_2282 ();
 b15zdnd11an1n64x5 FILLER_350_8 ();
 b15zdnd11an1n64x5 FILLER_350_72 ();
 b15zdnd11an1n64x5 FILLER_350_136 ();
 b15zdnd11an1n64x5 FILLER_350_200 ();
 b15zdnd11an1n16x5 FILLER_350_264 ();
 b15zdnd11an1n08x5 FILLER_350_280 ();
 b15zdnd00an1n01x5 FILLER_350_288 ();
 b15zdnd11an1n04x5 FILLER_350_307 ();
 b15zdnd11an1n32x5 FILLER_350_317 ();
 b15zdnd11an1n08x5 FILLER_350_349 ();
 b15zdnd11an1n04x5 FILLER_350_357 ();
 b15zdnd11an1n16x5 FILLER_350_403 ();
 b15zdnd00an1n01x5 FILLER_350_419 ();
 b15zdnd11an1n04x5 FILLER_350_451 ();
 b15zdnd11an1n08x5 FILLER_350_480 ();
 b15zdnd11an1n04x5 FILLER_350_488 ();
 b15zdnd00an1n01x5 FILLER_350_492 ();
 b15zdnd11an1n04x5 FILLER_350_517 ();
 b15zdnd11an1n64x5 FILLER_350_526 ();
 b15zdnd11an1n64x5 FILLER_350_590 ();
 b15zdnd11an1n64x5 FILLER_350_654 ();
 b15zdnd11an1n64x5 FILLER_350_726 ();
 b15zdnd11an1n64x5 FILLER_350_790 ();
 b15zdnd11an1n64x5 FILLER_350_854 ();
 b15zdnd11an1n64x5 FILLER_350_918 ();
 b15zdnd11an1n64x5 FILLER_350_982 ();
 b15zdnd11an1n64x5 FILLER_350_1046 ();
 b15zdnd11an1n16x5 FILLER_350_1110 ();
 b15zdnd11an1n04x5 FILLER_350_1126 ();
 b15zdnd11an1n04x5 FILLER_350_1142 ();
 b15zdnd11an1n04x5 FILLER_350_1150 ();
 b15zdnd00an1n01x5 FILLER_350_1154 ();
 b15zdnd11an1n64x5 FILLER_350_1170 ();
 b15zdnd11an1n64x5 FILLER_350_1234 ();
 b15zdnd11an1n64x5 FILLER_350_1298 ();
 b15zdnd11an1n64x5 FILLER_350_1362 ();
 b15zdnd11an1n64x5 FILLER_350_1426 ();
 b15zdnd11an1n64x5 FILLER_350_1490 ();
 b15zdnd11an1n64x5 FILLER_350_1554 ();
 b15zdnd11an1n64x5 FILLER_350_1618 ();
 b15zdnd11an1n64x5 FILLER_350_1682 ();
 b15zdnd11an1n64x5 FILLER_350_1746 ();
 b15zdnd11an1n64x5 FILLER_350_1810 ();
 b15zdnd11an1n64x5 FILLER_350_1874 ();
 b15zdnd11an1n64x5 FILLER_350_1938 ();
 b15zdnd11an1n64x5 FILLER_350_2002 ();
 b15zdnd11an1n64x5 FILLER_350_2066 ();
 b15zdnd11an1n16x5 FILLER_350_2130 ();
 b15zdnd11an1n08x5 FILLER_350_2146 ();
 b15zdnd11an1n64x5 FILLER_350_2162 ();
 b15zdnd11an1n32x5 FILLER_350_2226 ();
 b15zdnd11an1n16x5 FILLER_350_2258 ();
 b15zdnd00an1n02x5 FILLER_350_2274 ();
 b15zdnd11an1n64x5 FILLER_351_0 ();
 b15zdnd11an1n64x5 FILLER_351_64 ();
 b15zdnd11an1n64x5 FILLER_351_128 ();
 b15zdnd11an1n64x5 FILLER_351_192 ();
 b15zdnd11an1n64x5 FILLER_351_256 ();
 b15zdnd11an1n16x5 FILLER_351_320 ();
 b15zdnd11an1n04x5 FILLER_351_336 ();
 b15zdnd11an1n64x5 FILLER_351_372 ();
 b15zdnd11an1n16x5 FILLER_351_436 ();
 b15zdnd11an1n08x5 FILLER_351_452 ();
 b15zdnd00an1n02x5 FILLER_351_460 ();
 b15zdnd11an1n04x5 FILLER_351_489 ();
 b15zdnd00an1n01x5 FILLER_351_493 ();
 b15zdnd11an1n04x5 FILLER_351_508 ();
 b15zdnd11an1n64x5 FILLER_351_537 ();
 b15zdnd11an1n64x5 FILLER_351_601 ();
 b15zdnd11an1n64x5 FILLER_351_665 ();
 b15zdnd11an1n64x5 FILLER_351_729 ();
 b15zdnd11an1n64x5 FILLER_351_793 ();
 b15zdnd11an1n64x5 FILLER_351_857 ();
 b15zdnd11an1n64x5 FILLER_351_921 ();
 b15zdnd11an1n32x5 FILLER_351_985 ();
 b15zdnd11an1n16x5 FILLER_351_1017 ();
 b15zdnd11an1n04x5 FILLER_351_1033 ();
 b15zdnd00an1n02x5 FILLER_351_1037 ();
 b15zdnd00an1n01x5 FILLER_351_1039 ();
 b15zdnd11an1n32x5 FILLER_351_1082 ();
 b15zdnd00an1n02x5 FILLER_351_1114 ();
 b15zdnd11an1n04x5 FILLER_351_1121 ();
 b15zdnd11an1n16x5 FILLER_351_1143 ();
 b15zdnd00an1n01x5 FILLER_351_1159 ();
 b15zdnd11an1n64x5 FILLER_351_1202 ();
 b15zdnd11an1n64x5 FILLER_351_1266 ();
 b15zdnd11an1n64x5 FILLER_351_1330 ();
 b15zdnd11an1n64x5 FILLER_351_1394 ();
 b15zdnd11an1n64x5 FILLER_351_1458 ();
 b15zdnd11an1n64x5 FILLER_351_1522 ();
 b15zdnd11an1n64x5 FILLER_351_1586 ();
 b15zdnd11an1n64x5 FILLER_351_1650 ();
 b15zdnd11an1n64x5 FILLER_351_1714 ();
 b15zdnd11an1n64x5 FILLER_351_1778 ();
 b15zdnd11an1n64x5 FILLER_351_1842 ();
 b15zdnd11an1n64x5 FILLER_351_1906 ();
 b15zdnd11an1n64x5 FILLER_351_1970 ();
 b15zdnd11an1n64x5 FILLER_351_2034 ();
 b15zdnd11an1n64x5 FILLER_351_2098 ();
 b15zdnd11an1n64x5 FILLER_351_2162 ();
 b15zdnd11an1n32x5 FILLER_351_2226 ();
 b15zdnd11an1n16x5 FILLER_351_2258 ();
 b15zdnd11an1n08x5 FILLER_351_2274 ();
 b15zdnd00an1n02x5 FILLER_351_2282 ();
 b15zdnd11an1n64x5 FILLER_352_8 ();
 b15zdnd11an1n64x5 FILLER_352_72 ();
 b15zdnd11an1n64x5 FILLER_352_136 ();
 b15zdnd11an1n64x5 FILLER_352_200 ();
 b15zdnd11an1n64x5 FILLER_352_264 ();
 b15zdnd11an1n16x5 FILLER_352_328 ();
 b15zdnd11an1n04x5 FILLER_352_344 ();
 b15zdnd00an1n02x5 FILLER_352_348 ();
 b15zdnd00an1n01x5 FILLER_352_350 ();
 b15zdnd11an1n64x5 FILLER_352_393 ();
 b15zdnd11an1n04x5 FILLER_352_457 ();
 b15zdnd00an1n02x5 FILLER_352_461 ();
 b15zdnd00an1n01x5 FILLER_352_463 ();
 b15zdnd11an1n04x5 FILLER_352_469 ();
 b15zdnd11an1n04x5 FILLER_352_481 ();
 b15zdnd11an1n08x5 FILLER_352_489 ();
 b15zdnd11an1n04x5 FILLER_352_497 ();
 b15zdnd11an1n64x5 FILLER_352_543 ();
 b15zdnd11an1n64x5 FILLER_352_607 ();
 b15zdnd11an1n32x5 FILLER_352_671 ();
 b15zdnd11an1n08x5 FILLER_352_703 ();
 b15zdnd11an1n04x5 FILLER_352_711 ();
 b15zdnd00an1n02x5 FILLER_352_715 ();
 b15zdnd00an1n01x5 FILLER_352_717 ();
 b15zdnd11an1n64x5 FILLER_352_726 ();
 b15zdnd11an1n64x5 FILLER_352_790 ();
 b15zdnd11an1n64x5 FILLER_352_854 ();
 b15zdnd11an1n64x5 FILLER_352_918 ();
 b15zdnd11an1n32x5 FILLER_352_982 ();
 b15zdnd11an1n16x5 FILLER_352_1014 ();
 b15zdnd00an1n02x5 FILLER_352_1030 ();
 b15zdnd11an1n64x5 FILLER_352_1050 ();
 b15zdnd11an1n08x5 FILLER_352_1114 ();
 b15zdnd00an1n02x5 FILLER_352_1122 ();
 b15zdnd11an1n64x5 FILLER_352_1155 ();
 b15zdnd11an1n64x5 FILLER_352_1219 ();
 b15zdnd11an1n64x5 FILLER_352_1283 ();
 b15zdnd11an1n64x5 FILLER_352_1347 ();
 b15zdnd11an1n16x5 FILLER_352_1411 ();
 b15zdnd11an1n04x5 FILLER_352_1427 ();
 b15zdnd11an1n64x5 FILLER_352_1444 ();
 b15zdnd11an1n64x5 FILLER_352_1508 ();
 b15zdnd11an1n64x5 FILLER_352_1572 ();
 b15zdnd11an1n64x5 FILLER_352_1636 ();
 b15zdnd11an1n64x5 FILLER_352_1700 ();
 b15zdnd11an1n64x5 FILLER_352_1764 ();
 b15zdnd11an1n64x5 FILLER_352_1828 ();
 b15zdnd11an1n64x5 FILLER_352_1892 ();
 b15zdnd11an1n64x5 FILLER_352_1956 ();
 b15zdnd11an1n64x5 FILLER_352_2020 ();
 b15zdnd11an1n64x5 FILLER_352_2084 ();
 b15zdnd11an1n04x5 FILLER_352_2148 ();
 b15zdnd00an1n02x5 FILLER_352_2152 ();
 b15zdnd11an1n64x5 FILLER_352_2162 ();
 b15zdnd11an1n32x5 FILLER_352_2226 ();
 b15zdnd11an1n16x5 FILLER_352_2258 ();
 b15zdnd00an1n02x5 FILLER_352_2274 ();
 b15zdnd11an1n64x5 FILLER_353_0 ();
 b15zdnd11an1n64x5 FILLER_353_64 ();
 b15zdnd11an1n64x5 FILLER_353_128 ();
 b15zdnd11an1n64x5 FILLER_353_192 ();
 b15zdnd11an1n64x5 FILLER_353_256 ();
 b15zdnd11an1n08x5 FILLER_353_320 ();
 b15zdnd11an1n04x5 FILLER_353_328 ();
 b15zdnd00an1n02x5 FILLER_353_332 ();
 b15zdnd00an1n01x5 FILLER_353_334 ();
 b15zdnd11an1n04x5 FILLER_353_351 ();
 b15zdnd11an1n04x5 FILLER_353_367 ();
 b15zdnd11an1n04x5 FILLER_353_375 ();
 b15zdnd00an1n02x5 FILLER_353_379 ();
 b15zdnd00an1n01x5 FILLER_353_381 ();
 b15zdnd11an1n32x5 FILLER_353_410 ();
 b15zdnd11an1n08x5 FILLER_353_442 ();
 b15zdnd00an1n01x5 FILLER_353_450 ();
 b15zdnd11an1n04x5 FILLER_353_458 ();
 b15zdnd00an1n02x5 FILLER_353_462 ();
 b15zdnd00an1n01x5 FILLER_353_464 ();
 b15zdnd11an1n04x5 FILLER_353_507 ();
 b15zdnd11an1n64x5 FILLER_353_553 ();
 b15zdnd11an1n32x5 FILLER_353_617 ();
 b15zdnd11an1n08x5 FILLER_353_649 ();
 b15zdnd11an1n04x5 FILLER_353_657 ();
 b15zdnd00an1n02x5 FILLER_353_661 ();
 b15zdnd11an1n16x5 FILLER_353_675 ();
 b15zdnd11an1n04x5 FILLER_353_691 ();
 b15zdnd11an1n64x5 FILLER_353_707 ();
 b15zdnd11an1n64x5 FILLER_353_771 ();
 b15zdnd11an1n64x5 FILLER_353_835 ();
 b15zdnd11an1n64x5 FILLER_353_899 ();
 b15zdnd11an1n32x5 FILLER_353_963 ();
 b15zdnd11an1n16x5 FILLER_353_995 ();
 b15zdnd00an1n01x5 FILLER_353_1011 ();
 b15zdnd11an1n64x5 FILLER_353_1054 ();
 b15zdnd11an1n08x5 FILLER_353_1118 ();
 b15zdnd11an1n04x5 FILLER_353_1126 ();
 b15zdnd00an1n01x5 FILLER_353_1130 ();
 b15zdnd11an1n16x5 FILLER_353_1145 ();
 b15zdnd00an1n02x5 FILLER_353_1161 ();
 b15zdnd11an1n64x5 FILLER_353_1168 ();
 b15zdnd11an1n64x5 FILLER_353_1232 ();
 b15zdnd11an1n64x5 FILLER_353_1296 ();
 b15zdnd11an1n16x5 FILLER_353_1360 ();
 b15zdnd11an1n04x5 FILLER_353_1376 ();
 b15zdnd00an1n02x5 FILLER_353_1380 ();
 b15zdnd00an1n01x5 FILLER_353_1382 ();
 b15zdnd11an1n16x5 FILLER_353_1424 ();
 b15zdnd11an1n08x5 FILLER_353_1440 ();
 b15zdnd11an1n64x5 FILLER_353_1466 ();
 b15zdnd11an1n64x5 FILLER_353_1530 ();
 b15zdnd11an1n64x5 FILLER_353_1594 ();
 b15zdnd11an1n64x5 FILLER_353_1658 ();
 b15zdnd11an1n64x5 FILLER_353_1722 ();
 b15zdnd11an1n64x5 FILLER_353_1786 ();
 b15zdnd11an1n64x5 FILLER_353_1850 ();
 b15zdnd11an1n64x5 FILLER_353_1914 ();
 b15zdnd11an1n64x5 FILLER_353_1978 ();
 b15zdnd11an1n64x5 FILLER_353_2042 ();
 b15zdnd11an1n64x5 FILLER_353_2106 ();
 b15zdnd11an1n64x5 FILLER_353_2170 ();
 b15zdnd11an1n32x5 FILLER_353_2234 ();
 b15zdnd11an1n16x5 FILLER_353_2266 ();
 b15zdnd00an1n02x5 FILLER_353_2282 ();
 b15zdnd11an1n64x5 FILLER_354_8 ();
 b15zdnd11an1n64x5 FILLER_354_72 ();
 b15zdnd11an1n64x5 FILLER_354_136 ();
 b15zdnd11an1n64x5 FILLER_354_200 ();
 b15zdnd11an1n64x5 FILLER_354_264 ();
 b15zdnd11an1n16x5 FILLER_354_328 ();
 b15zdnd00an1n02x5 FILLER_354_344 ();
 b15zdnd00an1n01x5 FILLER_354_346 ();
 b15zdnd11an1n64x5 FILLER_354_389 ();
 b15zdnd11an1n16x5 FILLER_354_453 ();
 b15zdnd11an1n08x5 FILLER_354_469 ();
 b15zdnd11an1n04x5 FILLER_354_477 ();
 b15zdnd00an1n02x5 FILLER_354_481 ();
 b15zdnd00an1n01x5 FILLER_354_483 ();
 b15zdnd11an1n08x5 FILLER_354_526 ();
 b15zdnd00an1n02x5 FILLER_354_534 ();
 b15zdnd11an1n64x5 FILLER_354_539 ();
 b15zdnd11an1n04x5 FILLER_354_603 ();
 b15zdnd00an1n01x5 FILLER_354_607 ();
 b15zdnd11an1n32x5 FILLER_354_620 ();
 b15zdnd00an1n01x5 FILLER_354_652 ();
 b15zdnd11an1n16x5 FILLER_354_665 ();
 b15zdnd11an1n08x5 FILLER_354_681 ();
 b15zdnd11an1n04x5 FILLER_354_689 ();
 b15zdnd11an1n04x5 FILLER_354_712 ();
 b15zdnd00an1n02x5 FILLER_354_716 ();
 b15zdnd11an1n64x5 FILLER_354_726 ();
 b15zdnd11an1n08x5 FILLER_354_790 ();
 b15zdnd11an1n04x5 FILLER_354_798 ();
 b15zdnd00an1n02x5 FILLER_354_802 ();
 b15zdnd00an1n01x5 FILLER_354_804 ();
 b15zdnd11an1n64x5 FILLER_354_811 ();
 b15zdnd11an1n32x5 FILLER_354_875 ();
 b15zdnd11an1n16x5 FILLER_354_907 ();
 b15zdnd11an1n08x5 FILLER_354_923 ();
 b15zdnd11an1n32x5 FILLER_354_973 ();
 b15zdnd11an1n16x5 FILLER_354_1005 ();
 b15zdnd11an1n04x5 FILLER_354_1021 ();
 b15zdnd11an1n32x5 FILLER_354_1067 ();
 b15zdnd11an1n16x5 FILLER_354_1099 ();
 b15zdnd00an1n02x5 FILLER_354_1115 ();
 b15zdnd00an1n01x5 FILLER_354_1117 ();
 b15zdnd11an1n04x5 FILLER_354_1123 ();
 b15zdnd11an1n64x5 FILLER_354_1169 ();
 b15zdnd11an1n32x5 FILLER_354_1233 ();
 b15zdnd11an1n16x5 FILLER_354_1265 ();
 b15zdnd11an1n08x5 FILLER_354_1281 ();
 b15zdnd11an1n04x5 FILLER_354_1289 ();
 b15zdnd11an1n64x5 FILLER_354_1335 ();
 b15zdnd11an1n32x5 FILLER_354_1399 ();
 b15zdnd11an1n16x5 FILLER_354_1431 ();
 b15zdnd11an1n08x5 FILLER_354_1447 ();
 b15zdnd11an1n04x5 FILLER_354_1455 ();
 b15zdnd00an1n02x5 FILLER_354_1459 ();
 b15zdnd00an1n01x5 FILLER_354_1461 ();
 b15zdnd11an1n64x5 FILLER_354_1483 ();
 b15zdnd11an1n64x5 FILLER_354_1547 ();
 b15zdnd11an1n64x5 FILLER_354_1611 ();
 b15zdnd11an1n64x5 FILLER_354_1675 ();
 b15zdnd11an1n64x5 FILLER_354_1739 ();
 b15zdnd11an1n64x5 FILLER_354_1803 ();
 b15zdnd11an1n64x5 FILLER_354_1867 ();
 b15zdnd11an1n64x5 FILLER_354_1931 ();
 b15zdnd11an1n64x5 FILLER_354_1995 ();
 b15zdnd11an1n64x5 FILLER_354_2059 ();
 b15zdnd11an1n16x5 FILLER_354_2123 ();
 b15zdnd11an1n08x5 FILLER_354_2139 ();
 b15zdnd11an1n04x5 FILLER_354_2147 ();
 b15zdnd00an1n02x5 FILLER_354_2151 ();
 b15zdnd00an1n01x5 FILLER_354_2153 ();
 b15zdnd11an1n64x5 FILLER_354_2162 ();
 b15zdnd11an1n32x5 FILLER_354_2226 ();
 b15zdnd11an1n16x5 FILLER_354_2258 ();
 b15zdnd00an1n02x5 FILLER_354_2274 ();
 b15zdnd11an1n64x5 FILLER_355_0 ();
 b15zdnd11an1n64x5 FILLER_355_64 ();
 b15zdnd11an1n64x5 FILLER_355_128 ();
 b15zdnd11an1n64x5 FILLER_355_192 ();
 b15zdnd11an1n64x5 FILLER_355_256 ();
 b15zdnd11an1n08x5 FILLER_355_320 ();
 b15zdnd11an1n04x5 FILLER_355_328 ();
 b15zdnd00an1n02x5 FILLER_355_332 ();
 b15zdnd00an1n01x5 FILLER_355_334 ();
 b15zdnd11an1n04x5 FILLER_355_338 ();
 b15zdnd11an1n08x5 FILLER_355_352 ();
 b15zdnd00an1n02x5 FILLER_355_360 ();
 b15zdnd11an1n64x5 FILLER_355_383 ();
 b15zdnd11an1n16x5 FILLER_355_447 ();
 b15zdnd00an1n02x5 FILLER_355_463 ();
 b15zdnd00an1n01x5 FILLER_355_465 ();
 b15zdnd11an1n16x5 FILLER_355_493 ();
 b15zdnd11an1n04x5 FILLER_355_509 ();
 b15zdnd11an1n08x5 FILLER_355_527 ();
 b15zdnd00an1n01x5 FILLER_355_535 ();
 b15zdnd11an1n32x5 FILLER_355_551 ();
 b15zdnd11an1n08x5 FILLER_355_583 ();
 b15zdnd11an1n16x5 FILLER_355_600 ();
 b15zdnd00an1n01x5 FILLER_355_616 ();
 b15zdnd11an1n32x5 FILLER_355_629 ();
 b15zdnd11an1n16x5 FILLER_355_661 ();
 b15zdnd00an1n02x5 FILLER_355_677 ();
 b15zdnd11an1n04x5 FILLER_355_702 ();
 b15zdnd11an1n04x5 FILLER_355_709 ();
 b15zdnd11an1n64x5 FILLER_355_725 ();
 b15zdnd11an1n04x5 FILLER_355_789 ();
 b15zdnd11an1n64x5 FILLER_355_810 ();
 b15zdnd11an1n08x5 FILLER_355_874 ();
 b15zdnd00an1n02x5 FILLER_355_882 ();
 b15zdnd00an1n01x5 FILLER_355_884 ();
 b15zdnd11an1n08x5 FILLER_355_903 ();
 b15zdnd00an1n02x5 FILLER_355_911 ();
 b15zdnd00an1n01x5 FILLER_355_913 ();
 b15zdnd11an1n64x5 FILLER_355_932 ();
 b15zdnd00an1n02x5 FILLER_355_996 ();
 b15zdnd00an1n01x5 FILLER_355_998 ();
 b15zdnd11an1n04x5 FILLER_355_1041 ();
 b15zdnd11an1n64x5 FILLER_355_1050 ();
 b15zdnd11an1n64x5 FILLER_355_1114 ();
 b15zdnd11an1n64x5 FILLER_355_1178 ();
 b15zdnd11an1n64x5 FILLER_355_1242 ();
 b15zdnd11an1n64x5 FILLER_355_1306 ();
 b15zdnd11an1n32x5 FILLER_355_1370 ();
 b15zdnd11an1n08x5 FILLER_355_1402 ();
 b15zdnd00an1n02x5 FILLER_355_1410 ();
 b15zdnd00an1n01x5 FILLER_355_1412 ();
 b15zdnd11an1n64x5 FILLER_355_1465 ();
 b15zdnd11an1n64x5 FILLER_355_1529 ();
 b15zdnd11an1n64x5 FILLER_355_1593 ();
 b15zdnd11an1n64x5 FILLER_355_1657 ();
 b15zdnd11an1n64x5 FILLER_355_1721 ();
 b15zdnd11an1n64x5 FILLER_355_1785 ();
 b15zdnd11an1n64x5 FILLER_355_1849 ();
 b15zdnd11an1n64x5 FILLER_355_1913 ();
 b15zdnd11an1n64x5 FILLER_355_1977 ();
 b15zdnd11an1n64x5 FILLER_355_2041 ();
 b15zdnd11an1n64x5 FILLER_355_2105 ();
 b15zdnd11an1n64x5 FILLER_355_2169 ();
 b15zdnd11an1n32x5 FILLER_355_2233 ();
 b15zdnd11an1n16x5 FILLER_355_2265 ();
 b15zdnd00an1n02x5 FILLER_355_2281 ();
 b15zdnd00an1n01x5 FILLER_355_2283 ();
 b15zdnd11an1n64x5 FILLER_356_8 ();
 b15zdnd11an1n64x5 FILLER_356_72 ();
 b15zdnd11an1n64x5 FILLER_356_136 ();
 b15zdnd11an1n64x5 FILLER_356_200 ();
 b15zdnd11an1n64x5 FILLER_356_264 ();
 b15zdnd11an1n08x5 FILLER_356_328 ();
 b15zdnd11an1n04x5 FILLER_356_336 ();
 b15zdnd00an1n02x5 FILLER_356_340 ();
 b15zdnd00an1n01x5 FILLER_356_342 ();
 b15zdnd11an1n64x5 FILLER_356_351 ();
 b15zdnd11an1n64x5 FILLER_356_415 ();
 b15zdnd11an1n64x5 FILLER_356_479 ();
 b15zdnd11an1n08x5 FILLER_356_543 ();
 b15zdnd11an1n04x5 FILLER_356_551 ();
 b15zdnd00an1n02x5 FILLER_356_555 ();
 b15zdnd00an1n01x5 FILLER_356_557 ();
 b15zdnd11an1n64x5 FILLER_356_564 ();
 b15zdnd11an1n32x5 FILLER_356_628 ();
 b15zdnd11an1n16x5 FILLER_356_660 ();
 b15zdnd11an1n08x5 FILLER_356_676 ();
 b15zdnd00an1n02x5 FILLER_356_684 ();
 b15zdnd00an1n01x5 FILLER_356_686 ();
 b15zdnd11an1n04x5 FILLER_356_696 ();
 b15zdnd11an1n04x5 FILLER_356_712 ();
 b15zdnd00an1n02x5 FILLER_356_716 ();
 b15zdnd11an1n32x5 FILLER_356_726 ();
 b15zdnd11an1n16x5 FILLER_356_758 ();
 b15zdnd11an1n08x5 FILLER_356_774 ();
 b15zdnd11an1n04x5 FILLER_356_782 ();
 b15zdnd11an1n08x5 FILLER_356_790 ();
 b15zdnd11an1n04x5 FILLER_356_798 ();
 b15zdnd00an1n02x5 FILLER_356_802 ();
 b15zdnd11an1n04x5 FILLER_356_811 ();
 b15zdnd00an1n02x5 FILLER_356_815 ();
 b15zdnd00an1n01x5 FILLER_356_817 ();
 b15zdnd11an1n04x5 FILLER_356_830 ();
 b15zdnd11an1n08x5 FILLER_356_849 ();
 b15zdnd11an1n04x5 FILLER_356_857 ();
 b15zdnd00an1n02x5 FILLER_356_861 ();
 b15zdnd11an1n16x5 FILLER_356_887 ();
 b15zdnd11an1n08x5 FILLER_356_903 ();
 b15zdnd00an1n01x5 FILLER_356_911 ();
 b15zdnd11an1n32x5 FILLER_356_930 ();
 b15zdnd11an1n16x5 FILLER_356_962 ();
 b15zdnd00an1n02x5 FILLER_356_978 ();
 b15zdnd00an1n01x5 FILLER_356_980 ();
 b15zdnd11an1n16x5 FILLER_356_1023 ();
 b15zdnd11an1n08x5 FILLER_356_1039 ();
 b15zdnd11an1n04x5 FILLER_356_1047 ();
 b15zdnd00an1n02x5 FILLER_356_1051 ();
 b15zdnd00an1n01x5 FILLER_356_1053 ();
 b15zdnd11an1n64x5 FILLER_356_1068 ();
 b15zdnd00an1n01x5 FILLER_356_1132 ();
 b15zdnd11an1n64x5 FILLER_356_1150 ();
 b15zdnd11an1n16x5 FILLER_356_1214 ();
 b15zdnd11an1n08x5 FILLER_356_1230 ();
 b15zdnd00an1n01x5 FILLER_356_1238 ();
 b15zdnd11an1n64x5 FILLER_356_1264 ();
 b15zdnd11an1n64x5 FILLER_356_1328 ();
 b15zdnd11an1n64x5 FILLER_356_1392 ();
 b15zdnd11an1n64x5 FILLER_356_1456 ();
 b15zdnd11an1n64x5 FILLER_356_1520 ();
 b15zdnd11an1n64x5 FILLER_356_1584 ();
 b15zdnd11an1n64x5 FILLER_356_1648 ();
 b15zdnd11an1n64x5 FILLER_356_1712 ();
 b15zdnd11an1n64x5 FILLER_356_1776 ();
 b15zdnd11an1n64x5 FILLER_356_1840 ();
 b15zdnd11an1n64x5 FILLER_356_1904 ();
 b15zdnd11an1n64x5 FILLER_356_1968 ();
 b15zdnd11an1n64x5 FILLER_356_2032 ();
 b15zdnd11an1n32x5 FILLER_356_2096 ();
 b15zdnd11an1n16x5 FILLER_356_2128 ();
 b15zdnd11an1n08x5 FILLER_356_2144 ();
 b15zdnd00an1n02x5 FILLER_356_2152 ();
 b15zdnd11an1n64x5 FILLER_356_2162 ();
 b15zdnd11an1n32x5 FILLER_356_2226 ();
 b15zdnd11an1n16x5 FILLER_356_2258 ();
 b15zdnd00an1n02x5 FILLER_356_2274 ();
 b15zdnd11an1n64x5 FILLER_357_0 ();
 b15zdnd11an1n64x5 FILLER_357_64 ();
 b15zdnd11an1n64x5 FILLER_357_128 ();
 b15zdnd11an1n64x5 FILLER_357_192 ();
 b15zdnd11an1n64x5 FILLER_357_256 ();
 b15zdnd11an1n32x5 FILLER_357_320 ();
 b15zdnd11an1n16x5 FILLER_357_352 ();
 b15zdnd11an1n64x5 FILLER_357_387 ();
 b15zdnd11an1n64x5 FILLER_357_451 ();
 b15zdnd11an1n32x5 FILLER_357_515 ();
 b15zdnd11an1n16x5 FILLER_357_547 ();
 b15zdnd11an1n08x5 FILLER_357_563 ();
 b15zdnd11an1n04x5 FILLER_357_571 ();
 b15zdnd11an1n16x5 FILLER_357_580 ();
 b15zdnd11an1n04x5 FILLER_357_596 ();
 b15zdnd11an1n64x5 FILLER_357_618 ();
 b15zdnd11an1n64x5 FILLER_357_682 ();
 b15zdnd11an1n32x5 FILLER_357_746 ();
 b15zdnd11an1n16x5 FILLER_357_778 ();
 b15zdnd11an1n04x5 FILLER_357_794 ();
 b15zdnd00an1n01x5 FILLER_357_798 ();
 b15zdnd11an1n04x5 FILLER_357_813 ();
 b15zdnd11an1n64x5 FILLER_357_859 ();
 b15zdnd11an1n04x5 FILLER_357_923 ();
 b15zdnd00an1n02x5 FILLER_357_927 ();
 b15zdnd11an1n32x5 FILLER_357_939 ();
 b15zdnd11an1n04x5 FILLER_357_971 ();
 b15zdnd11an1n16x5 FILLER_357_993 ();
 b15zdnd00an1n01x5 FILLER_357_1009 ();
 b15zdnd11an1n08x5 FILLER_357_1050 ();
 b15zdnd00an1n01x5 FILLER_357_1058 ();
 b15zdnd11an1n64x5 FILLER_357_1079 ();
 b15zdnd11an1n64x5 FILLER_357_1143 ();
 b15zdnd11an1n64x5 FILLER_357_1207 ();
 b15zdnd11an1n64x5 FILLER_357_1271 ();
 b15zdnd11an1n64x5 FILLER_357_1335 ();
 b15zdnd11an1n16x5 FILLER_357_1399 ();
 b15zdnd11an1n08x5 FILLER_357_1415 ();
 b15zdnd00an1n02x5 FILLER_357_1423 ();
 b15zdnd00an1n01x5 FILLER_357_1425 ();
 b15zdnd11an1n04x5 FILLER_357_1436 ();
 b15zdnd11an1n64x5 FILLER_357_1492 ();
 b15zdnd11an1n64x5 FILLER_357_1556 ();
 b15zdnd11an1n64x5 FILLER_357_1620 ();
 b15zdnd11an1n64x5 FILLER_357_1684 ();
 b15zdnd11an1n64x5 FILLER_357_1748 ();
 b15zdnd11an1n64x5 FILLER_357_1812 ();
 b15zdnd11an1n64x5 FILLER_357_1876 ();
 b15zdnd11an1n64x5 FILLER_357_1940 ();
 b15zdnd11an1n64x5 FILLER_357_2004 ();
 b15zdnd11an1n64x5 FILLER_357_2068 ();
 b15zdnd11an1n64x5 FILLER_357_2132 ();
 b15zdnd11an1n64x5 FILLER_357_2196 ();
 b15zdnd11an1n16x5 FILLER_357_2260 ();
 b15zdnd11an1n08x5 FILLER_357_2276 ();
 b15zdnd11an1n64x5 FILLER_358_8 ();
 b15zdnd11an1n64x5 FILLER_358_72 ();
 b15zdnd11an1n64x5 FILLER_358_136 ();
 b15zdnd11an1n64x5 FILLER_358_200 ();
 b15zdnd11an1n64x5 FILLER_358_264 ();
 b15zdnd11an1n64x5 FILLER_358_328 ();
 b15zdnd11an1n64x5 FILLER_358_392 ();
 b15zdnd11an1n64x5 FILLER_358_456 ();
 b15zdnd11an1n32x5 FILLER_358_520 ();
 b15zdnd00an1n01x5 FILLER_358_552 ();
 b15zdnd11an1n64x5 FILLER_358_565 ();
 b15zdnd11an1n64x5 FILLER_358_629 ();
 b15zdnd11an1n16x5 FILLER_358_693 ();
 b15zdnd11an1n08x5 FILLER_358_709 ();
 b15zdnd00an1n01x5 FILLER_358_717 ();
 b15zdnd11an1n32x5 FILLER_358_726 ();
 b15zdnd11an1n16x5 FILLER_358_758 ();
 b15zdnd11an1n08x5 FILLER_358_774 ();
 b15zdnd11an1n04x5 FILLER_358_782 ();
 b15zdnd00an1n02x5 FILLER_358_786 ();
 b15zdnd11an1n04x5 FILLER_358_792 ();
 b15zdnd11an1n16x5 FILLER_358_816 ();
 b15zdnd11an1n04x5 FILLER_358_832 ();
 b15zdnd00an1n02x5 FILLER_358_836 ();
 b15zdnd11an1n32x5 FILLER_358_853 ();
 b15zdnd11an1n16x5 FILLER_358_885 ();
 b15zdnd11an1n08x5 FILLER_358_901 ();
 b15zdnd11an1n04x5 FILLER_358_909 ();
 b15zdnd00an1n02x5 FILLER_358_913 ();
 b15zdnd00an1n01x5 FILLER_358_915 ();
 b15zdnd11an1n08x5 FILLER_358_925 ();
 b15zdnd00an1n02x5 FILLER_358_933 ();
 b15zdnd00an1n01x5 FILLER_358_935 ();
 b15zdnd11an1n16x5 FILLER_358_978 ();
 b15zdnd11an1n04x5 FILLER_358_994 ();
 b15zdnd11an1n04x5 FILLER_358_1023 ();
 b15zdnd11an1n16x5 FILLER_358_1032 ();
 b15zdnd11an1n64x5 FILLER_358_1053 ();
 b15zdnd11an1n64x5 FILLER_358_1117 ();
 b15zdnd11an1n64x5 FILLER_358_1181 ();
 b15zdnd11an1n64x5 FILLER_358_1245 ();
 b15zdnd11an1n64x5 FILLER_358_1309 ();
 b15zdnd11an1n64x5 FILLER_358_1373 ();
 b15zdnd11an1n64x5 FILLER_358_1437 ();
 b15zdnd11an1n64x5 FILLER_358_1501 ();
 b15zdnd11an1n64x5 FILLER_358_1565 ();
 b15zdnd11an1n64x5 FILLER_358_1629 ();
 b15zdnd11an1n64x5 FILLER_358_1693 ();
 b15zdnd11an1n64x5 FILLER_358_1757 ();
 b15zdnd11an1n64x5 FILLER_358_1821 ();
 b15zdnd11an1n64x5 FILLER_358_1885 ();
 b15zdnd11an1n64x5 FILLER_358_1949 ();
 b15zdnd11an1n64x5 FILLER_358_2013 ();
 b15zdnd11an1n64x5 FILLER_358_2077 ();
 b15zdnd11an1n08x5 FILLER_358_2141 ();
 b15zdnd11an1n04x5 FILLER_358_2149 ();
 b15zdnd00an1n01x5 FILLER_358_2153 ();
 b15zdnd11an1n64x5 FILLER_358_2162 ();
 b15zdnd11an1n32x5 FILLER_358_2226 ();
 b15zdnd11an1n16x5 FILLER_358_2258 ();
 b15zdnd00an1n02x5 FILLER_358_2274 ();
 b15zdnd11an1n64x5 FILLER_359_0 ();
 b15zdnd11an1n64x5 FILLER_359_64 ();
 b15zdnd11an1n64x5 FILLER_359_128 ();
 b15zdnd11an1n64x5 FILLER_359_192 ();
 b15zdnd11an1n64x5 FILLER_359_256 ();
 b15zdnd11an1n64x5 FILLER_359_320 ();
 b15zdnd11an1n64x5 FILLER_359_384 ();
 b15zdnd11an1n64x5 FILLER_359_448 ();
 b15zdnd11an1n64x5 FILLER_359_512 ();
 b15zdnd11an1n64x5 FILLER_359_576 ();
 b15zdnd11an1n64x5 FILLER_359_640 ();
 b15zdnd11an1n64x5 FILLER_359_704 ();
 b15zdnd11an1n64x5 FILLER_359_768 ();
 b15zdnd11an1n64x5 FILLER_359_832 ();
 b15zdnd11an1n16x5 FILLER_359_896 ();
 b15zdnd00an1n02x5 FILLER_359_912 ();
 b15zdnd11an1n32x5 FILLER_359_926 ();
 b15zdnd11an1n16x5 FILLER_359_958 ();
 b15zdnd00an1n02x5 FILLER_359_974 ();
 b15zdnd11an1n16x5 FILLER_359_994 ();
 b15zdnd11an1n04x5 FILLER_359_1010 ();
 b15zdnd00an1n02x5 FILLER_359_1014 ();
 b15zdnd00an1n01x5 FILLER_359_1016 ();
 b15zdnd11an1n64x5 FILLER_359_1041 ();
 b15zdnd11an1n32x5 FILLER_359_1105 ();
 b15zdnd11an1n04x5 FILLER_359_1137 ();
 b15zdnd00an1n01x5 FILLER_359_1141 ();
 b15zdnd11an1n64x5 FILLER_359_1162 ();
 b15zdnd11an1n64x5 FILLER_359_1226 ();
 b15zdnd11an1n64x5 FILLER_359_1290 ();
 b15zdnd11an1n64x5 FILLER_359_1354 ();
 b15zdnd11an1n64x5 FILLER_359_1418 ();
 b15zdnd11an1n64x5 FILLER_359_1482 ();
 b15zdnd11an1n64x5 FILLER_359_1546 ();
 b15zdnd11an1n64x5 FILLER_359_1610 ();
 b15zdnd11an1n64x5 FILLER_359_1674 ();
 b15zdnd11an1n64x5 FILLER_359_1738 ();
 b15zdnd11an1n64x5 FILLER_359_1802 ();
 b15zdnd11an1n64x5 FILLER_359_1866 ();
 b15zdnd11an1n64x5 FILLER_359_1930 ();
 b15zdnd11an1n64x5 FILLER_359_1994 ();
 b15zdnd11an1n64x5 FILLER_359_2058 ();
 b15zdnd11an1n64x5 FILLER_359_2122 ();
 b15zdnd11an1n64x5 FILLER_359_2186 ();
 b15zdnd11an1n32x5 FILLER_359_2250 ();
 b15zdnd00an1n02x5 FILLER_359_2282 ();
 b15zdnd11an1n64x5 FILLER_360_8 ();
 b15zdnd11an1n64x5 FILLER_360_72 ();
 b15zdnd11an1n64x5 FILLER_360_136 ();
 b15zdnd11an1n64x5 FILLER_360_200 ();
 b15zdnd11an1n64x5 FILLER_360_264 ();
 b15zdnd11an1n64x5 FILLER_360_328 ();
 b15zdnd11an1n64x5 FILLER_360_392 ();
 b15zdnd11an1n64x5 FILLER_360_456 ();
 b15zdnd11an1n08x5 FILLER_360_520 ();
 b15zdnd00an1n01x5 FILLER_360_528 ();
 b15zdnd11an1n64x5 FILLER_360_571 ();
 b15zdnd11an1n64x5 FILLER_360_635 ();
 b15zdnd11an1n16x5 FILLER_360_699 ();
 b15zdnd00an1n02x5 FILLER_360_715 ();
 b15zdnd00an1n01x5 FILLER_360_717 ();
 b15zdnd11an1n64x5 FILLER_360_726 ();
 b15zdnd11an1n64x5 FILLER_360_790 ();
 b15zdnd11an1n64x5 FILLER_360_854 ();
 b15zdnd11an1n64x5 FILLER_360_918 ();
 b15zdnd11an1n64x5 FILLER_360_982 ();
 b15zdnd11an1n64x5 FILLER_360_1046 ();
 b15zdnd11an1n64x5 FILLER_360_1110 ();
 b15zdnd11an1n64x5 FILLER_360_1174 ();
 b15zdnd11an1n64x5 FILLER_360_1238 ();
 b15zdnd11an1n64x5 FILLER_360_1302 ();
 b15zdnd11an1n64x5 FILLER_360_1366 ();
 b15zdnd11an1n64x5 FILLER_360_1430 ();
 b15zdnd11an1n64x5 FILLER_360_1494 ();
 b15zdnd11an1n64x5 FILLER_360_1558 ();
 b15zdnd11an1n64x5 FILLER_360_1622 ();
 b15zdnd11an1n64x5 FILLER_360_1686 ();
 b15zdnd11an1n64x5 FILLER_360_1750 ();
 b15zdnd11an1n64x5 FILLER_360_1814 ();
 b15zdnd11an1n64x5 FILLER_360_1878 ();
 b15zdnd11an1n64x5 FILLER_360_1942 ();
 b15zdnd11an1n64x5 FILLER_360_2006 ();
 b15zdnd11an1n64x5 FILLER_360_2070 ();
 b15zdnd11an1n16x5 FILLER_360_2134 ();
 b15zdnd11an1n04x5 FILLER_360_2150 ();
 b15zdnd11an1n64x5 FILLER_360_2162 ();
 b15zdnd11an1n32x5 FILLER_360_2226 ();
 b15zdnd11an1n16x5 FILLER_360_2258 ();
 b15zdnd00an1n02x5 FILLER_360_2274 ();
 b15zdnd11an1n64x5 FILLER_361_0 ();
 b15zdnd11an1n64x5 FILLER_361_64 ();
 b15zdnd11an1n64x5 FILLER_361_128 ();
 b15zdnd11an1n64x5 FILLER_361_192 ();
 b15zdnd11an1n64x5 FILLER_361_256 ();
 b15zdnd11an1n32x5 FILLER_361_320 ();
 b15zdnd00an1n02x5 FILLER_361_352 ();
 b15zdnd11an1n64x5 FILLER_361_374 ();
 b15zdnd11an1n64x5 FILLER_361_438 ();
 b15zdnd11an1n64x5 FILLER_361_502 ();
 b15zdnd11an1n64x5 FILLER_361_566 ();
 b15zdnd11an1n64x5 FILLER_361_630 ();
 b15zdnd11an1n64x5 FILLER_361_694 ();
 b15zdnd11an1n16x5 FILLER_361_758 ();
 b15zdnd11an1n08x5 FILLER_361_774 ();
 b15zdnd00an1n02x5 FILLER_361_782 ();
 b15zdnd00an1n01x5 FILLER_361_784 ();
 b15zdnd11an1n04x5 FILLER_361_789 ();
 b15zdnd11an1n64x5 FILLER_361_813 ();
 b15zdnd11an1n64x5 FILLER_361_877 ();
 b15zdnd11an1n64x5 FILLER_361_941 ();
 b15zdnd11an1n08x5 FILLER_361_1005 ();
 b15zdnd00an1n02x5 FILLER_361_1013 ();
 b15zdnd00an1n01x5 FILLER_361_1015 ();
 b15zdnd11an1n64x5 FILLER_361_1033 ();
 b15zdnd11an1n16x5 FILLER_361_1097 ();
 b15zdnd11an1n08x5 FILLER_361_1113 ();
 b15zdnd00an1n01x5 FILLER_361_1121 ();
 b15zdnd11an1n04x5 FILLER_361_1147 ();
 b15zdnd11an1n64x5 FILLER_361_1155 ();
 b15zdnd11an1n64x5 FILLER_361_1219 ();
 b15zdnd11an1n64x5 FILLER_361_1283 ();
 b15zdnd11an1n64x5 FILLER_361_1347 ();
 b15zdnd11an1n64x5 FILLER_361_1411 ();
 b15zdnd11an1n64x5 FILLER_361_1475 ();
 b15zdnd11an1n64x5 FILLER_361_1539 ();
 b15zdnd11an1n64x5 FILLER_361_1603 ();
 b15zdnd11an1n64x5 FILLER_361_1667 ();
 b15zdnd11an1n64x5 FILLER_361_1731 ();
 b15zdnd11an1n64x5 FILLER_361_1795 ();
 b15zdnd11an1n64x5 FILLER_361_1859 ();
 b15zdnd11an1n64x5 FILLER_361_1923 ();
 b15zdnd11an1n64x5 FILLER_361_1987 ();
 b15zdnd11an1n64x5 FILLER_361_2051 ();
 b15zdnd11an1n64x5 FILLER_361_2115 ();
 b15zdnd11an1n64x5 FILLER_361_2179 ();
 b15zdnd11an1n32x5 FILLER_361_2243 ();
 b15zdnd11an1n08x5 FILLER_361_2275 ();
 b15zdnd00an1n01x5 FILLER_361_2283 ();
 b15zdnd11an1n64x5 FILLER_362_8 ();
 b15zdnd11an1n64x5 FILLER_362_72 ();
 b15zdnd11an1n64x5 FILLER_362_136 ();
 b15zdnd11an1n64x5 FILLER_362_200 ();
 b15zdnd11an1n64x5 FILLER_362_264 ();
 b15zdnd11an1n64x5 FILLER_362_328 ();
 b15zdnd11an1n64x5 FILLER_362_392 ();
 b15zdnd11an1n64x5 FILLER_362_456 ();
 b15zdnd11an1n64x5 FILLER_362_520 ();
 b15zdnd11an1n64x5 FILLER_362_584 ();
 b15zdnd11an1n64x5 FILLER_362_648 ();
 b15zdnd11an1n04x5 FILLER_362_712 ();
 b15zdnd00an1n02x5 FILLER_362_716 ();
 b15zdnd11an1n64x5 FILLER_362_726 ();
 b15zdnd11an1n64x5 FILLER_362_790 ();
 b15zdnd11an1n64x5 FILLER_362_854 ();
 b15zdnd11an1n64x5 FILLER_362_918 ();
 b15zdnd11an1n64x5 FILLER_362_982 ();
 b15zdnd11an1n32x5 FILLER_362_1046 ();
 b15zdnd11an1n16x5 FILLER_362_1078 ();
 b15zdnd00an1n02x5 FILLER_362_1094 ();
 b15zdnd11an1n64x5 FILLER_362_1136 ();
 b15zdnd11an1n32x5 FILLER_362_1200 ();
 b15zdnd00an1n01x5 FILLER_362_1232 ();
 b15zdnd11an1n08x5 FILLER_362_1237 ();
 b15zdnd11an1n04x5 FILLER_362_1245 ();
 b15zdnd00an1n01x5 FILLER_362_1249 ();
 b15zdnd11an1n64x5 FILLER_362_1254 ();
 b15zdnd11an1n64x5 FILLER_362_1318 ();
 b15zdnd11an1n64x5 FILLER_362_1382 ();
 b15zdnd11an1n64x5 FILLER_362_1446 ();
 b15zdnd11an1n64x5 FILLER_362_1510 ();
 b15zdnd11an1n64x5 FILLER_362_1574 ();
 b15zdnd11an1n64x5 FILLER_362_1638 ();
 b15zdnd11an1n64x5 FILLER_362_1702 ();
 b15zdnd11an1n64x5 FILLER_362_1766 ();
 b15zdnd11an1n64x5 FILLER_362_1830 ();
 b15zdnd11an1n64x5 FILLER_362_1894 ();
 b15zdnd11an1n64x5 FILLER_362_1958 ();
 b15zdnd11an1n64x5 FILLER_362_2022 ();
 b15zdnd11an1n64x5 FILLER_362_2086 ();
 b15zdnd11an1n04x5 FILLER_362_2150 ();
 b15zdnd11an1n64x5 FILLER_362_2162 ();
 b15zdnd11an1n32x5 FILLER_362_2226 ();
 b15zdnd11an1n16x5 FILLER_362_2258 ();
 b15zdnd00an1n02x5 FILLER_362_2274 ();
 b15zdnd11an1n64x5 FILLER_363_0 ();
 b15zdnd11an1n64x5 FILLER_363_64 ();
 b15zdnd11an1n64x5 FILLER_363_128 ();
 b15zdnd11an1n64x5 FILLER_363_192 ();
 b15zdnd11an1n64x5 FILLER_363_256 ();
 b15zdnd11an1n64x5 FILLER_363_320 ();
 b15zdnd11an1n64x5 FILLER_363_384 ();
 b15zdnd11an1n64x5 FILLER_363_448 ();
 b15zdnd11an1n64x5 FILLER_363_512 ();
 b15zdnd11an1n64x5 FILLER_363_576 ();
 b15zdnd11an1n64x5 FILLER_363_640 ();
 b15zdnd11an1n64x5 FILLER_363_704 ();
 b15zdnd11an1n64x5 FILLER_363_768 ();
 b15zdnd11an1n64x5 FILLER_363_832 ();
 b15zdnd11an1n64x5 FILLER_363_896 ();
 b15zdnd11an1n64x5 FILLER_363_960 ();
 b15zdnd11an1n04x5 FILLER_363_1024 ();
 b15zdnd00an1n02x5 FILLER_363_1028 ();
 b15zdnd11an1n64x5 FILLER_363_1050 ();
 b15zdnd11an1n64x5 FILLER_363_1114 ();
 b15zdnd11an1n08x5 FILLER_363_1178 ();
 b15zdnd11an1n04x5 FILLER_363_1186 ();
 b15zdnd00an1n02x5 FILLER_363_1190 ();
 b15zdnd00an1n01x5 FILLER_363_1192 ();
 b15zdnd11an1n16x5 FILLER_363_1198 ();
 b15zdnd11an1n04x5 FILLER_363_1214 ();
 b15zdnd11an1n04x5 FILLER_363_1238 ();
 b15zdnd00an1n01x5 FILLER_363_1242 ();
 b15zdnd11an1n64x5 FILLER_363_1285 ();
 b15zdnd11an1n64x5 FILLER_363_1349 ();
 b15zdnd11an1n64x5 FILLER_363_1413 ();
 b15zdnd11an1n64x5 FILLER_363_1477 ();
 b15zdnd11an1n64x5 FILLER_363_1541 ();
 b15zdnd11an1n64x5 FILLER_363_1605 ();
 b15zdnd11an1n64x5 FILLER_363_1669 ();
 b15zdnd11an1n64x5 FILLER_363_1733 ();
 b15zdnd11an1n64x5 FILLER_363_1797 ();
 b15zdnd11an1n64x5 FILLER_363_1861 ();
 b15zdnd11an1n64x5 FILLER_363_1925 ();
 b15zdnd11an1n64x5 FILLER_363_1989 ();
 b15zdnd11an1n64x5 FILLER_363_2053 ();
 b15zdnd11an1n64x5 FILLER_363_2117 ();
 b15zdnd11an1n64x5 FILLER_363_2181 ();
 b15zdnd11an1n32x5 FILLER_363_2245 ();
 b15zdnd11an1n04x5 FILLER_363_2277 ();
 b15zdnd00an1n02x5 FILLER_363_2281 ();
 b15zdnd00an1n01x5 FILLER_363_2283 ();
 b15zdnd11an1n64x5 FILLER_364_8 ();
 b15zdnd11an1n64x5 FILLER_364_72 ();
 b15zdnd11an1n64x5 FILLER_364_136 ();
 b15zdnd11an1n64x5 FILLER_364_200 ();
 b15zdnd11an1n64x5 FILLER_364_264 ();
 b15zdnd11an1n64x5 FILLER_364_328 ();
 b15zdnd11an1n64x5 FILLER_364_392 ();
 b15zdnd11an1n64x5 FILLER_364_456 ();
 b15zdnd11an1n08x5 FILLER_364_520 ();
 b15zdnd11an1n64x5 FILLER_364_570 ();
 b15zdnd11an1n64x5 FILLER_364_634 ();
 b15zdnd11an1n16x5 FILLER_364_698 ();
 b15zdnd11an1n04x5 FILLER_364_714 ();
 b15zdnd11an1n64x5 FILLER_364_726 ();
 b15zdnd11an1n64x5 FILLER_364_790 ();
 b15zdnd11an1n64x5 FILLER_364_854 ();
 b15zdnd11an1n64x5 FILLER_364_918 ();
 b15zdnd11an1n64x5 FILLER_364_982 ();
 b15zdnd11an1n64x5 FILLER_364_1046 ();
 b15zdnd11an1n32x5 FILLER_364_1110 ();
 b15zdnd11an1n16x5 FILLER_364_1142 ();
 b15zdnd11an1n08x5 FILLER_364_1158 ();
 b15zdnd00an1n02x5 FILLER_364_1166 ();
 b15zdnd11an1n04x5 FILLER_364_1210 ();
 b15zdnd11an1n04x5 FILLER_364_1256 ();
 b15zdnd11an1n64x5 FILLER_364_1264 ();
 b15zdnd11an1n64x5 FILLER_364_1328 ();
 b15zdnd11an1n64x5 FILLER_364_1392 ();
 b15zdnd11an1n64x5 FILLER_364_1456 ();
 b15zdnd11an1n64x5 FILLER_364_1520 ();
 b15zdnd11an1n64x5 FILLER_364_1584 ();
 b15zdnd11an1n64x5 FILLER_364_1648 ();
 b15zdnd11an1n64x5 FILLER_364_1712 ();
 b15zdnd11an1n64x5 FILLER_364_1776 ();
 b15zdnd11an1n64x5 FILLER_364_1840 ();
 b15zdnd11an1n64x5 FILLER_364_1904 ();
 b15zdnd11an1n64x5 FILLER_364_1968 ();
 b15zdnd11an1n64x5 FILLER_364_2032 ();
 b15zdnd11an1n32x5 FILLER_364_2096 ();
 b15zdnd11an1n16x5 FILLER_364_2128 ();
 b15zdnd11an1n08x5 FILLER_364_2144 ();
 b15zdnd00an1n02x5 FILLER_364_2152 ();
 b15zdnd11an1n64x5 FILLER_364_2162 ();
 b15zdnd11an1n32x5 FILLER_364_2226 ();
 b15zdnd11an1n16x5 FILLER_364_2258 ();
 b15zdnd00an1n02x5 FILLER_364_2274 ();
 b15zdnd11an1n64x5 FILLER_365_0 ();
 b15zdnd11an1n64x5 FILLER_365_64 ();
 b15zdnd11an1n64x5 FILLER_365_128 ();
 b15zdnd11an1n64x5 FILLER_365_192 ();
 b15zdnd11an1n64x5 FILLER_365_256 ();
 b15zdnd11an1n64x5 FILLER_365_320 ();
 b15zdnd11an1n64x5 FILLER_365_384 ();
 b15zdnd00an1n01x5 FILLER_365_448 ();
 b15zdnd11an1n64x5 FILLER_365_452 ();
 b15zdnd11an1n16x5 FILLER_365_516 ();
 b15zdnd11an1n08x5 FILLER_365_532 ();
 b15zdnd11an1n04x5 FILLER_365_540 ();
 b15zdnd11an1n04x5 FILLER_365_586 ();
 b15zdnd00an1n02x5 FILLER_365_590 ();
 b15zdnd00an1n01x5 FILLER_365_592 ();
 b15zdnd11an1n64x5 FILLER_365_635 ();
 b15zdnd11an1n64x5 FILLER_365_699 ();
 b15zdnd11an1n64x5 FILLER_365_763 ();
 b15zdnd11an1n64x5 FILLER_365_827 ();
 b15zdnd11an1n64x5 FILLER_365_891 ();
 b15zdnd11an1n64x5 FILLER_365_955 ();
 b15zdnd11an1n64x5 FILLER_365_1019 ();
 b15zdnd11an1n64x5 FILLER_365_1083 ();
 b15zdnd00an1n02x5 FILLER_365_1147 ();
 b15zdnd11an1n16x5 FILLER_365_1191 ();
 b15zdnd00an1n02x5 FILLER_365_1207 ();
 b15zdnd11an1n04x5 FILLER_365_1223 ();
 b15zdnd11an1n08x5 FILLER_365_1239 ();
 b15zdnd00an1n02x5 FILLER_365_1247 ();
 b15zdnd11an1n04x5 FILLER_365_1269 ();
 b15zdnd00an1n01x5 FILLER_365_1273 ();
 b15zdnd11an1n64x5 FILLER_365_1305 ();
 b15zdnd11an1n64x5 FILLER_365_1369 ();
 b15zdnd11an1n64x5 FILLER_365_1433 ();
 b15zdnd11an1n64x5 FILLER_365_1497 ();
 b15zdnd11an1n64x5 FILLER_365_1561 ();
 b15zdnd11an1n64x5 FILLER_365_1625 ();
 b15zdnd11an1n64x5 FILLER_365_1689 ();
 b15zdnd11an1n64x5 FILLER_365_1753 ();
 b15zdnd11an1n64x5 FILLER_365_1817 ();
 b15zdnd11an1n64x5 FILLER_365_1881 ();
 b15zdnd11an1n64x5 FILLER_365_1945 ();
 b15zdnd11an1n64x5 FILLER_365_2009 ();
 b15zdnd11an1n64x5 FILLER_365_2073 ();
 b15zdnd11an1n64x5 FILLER_365_2137 ();
 b15zdnd11an1n64x5 FILLER_365_2201 ();
 b15zdnd11an1n16x5 FILLER_365_2265 ();
 b15zdnd00an1n02x5 FILLER_365_2281 ();
 b15zdnd00an1n01x5 FILLER_365_2283 ();
 b15zdnd11an1n64x5 FILLER_366_8 ();
 b15zdnd11an1n64x5 FILLER_366_72 ();
 b15zdnd11an1n64x5 FILLER_366_136 ();
 b15zdnd11an1n64x5 FILLER_366_200 ();
 b15zdnd11an1n64x5 FILLER_366_264 ();
 b15zdnd11an1n32x5 FILLER_366_328 ();
 b15zdnd11an1n08x5 FILLER_366_360 ();
 b15zdnd00an1n02x5 FILLER_366_368 ();
 b15zdnd11an1n64x5 FILLER_366_374 ();
 b15zdnd11an1n64x5 FILLER_366_438 ();
 b15zdnd11an1n08x5 FILLER_366_502 ();
 b15zdnd00an1n01x5 FILLER_366_510 ();
 b15zdnd11an1n16x5 FILLER_366_542 ();
 b15zdnd11an1n08x5 FILLER_366_558 ();
 b15zdnd11an1n04x5 FILLER_366_566 ();
 b15zdnd11an1n64x5 FILLER_366_612 ();
 b15zdnd11an1n32x5 FILLER_366_676 ();
 b15zdnd11an1n08x5 FILLER_366_708 ();
 b15zdnd00an1n02x5 FILLER_366_716 ();
 b15zdnd11an1n64x5 FILLER_366_726 ();
 b15zdnd11an1n64x5 FILLER_366_790 ();
 b15zdnd11an1n32x5 FILLER_366_854 ();
 b15zdnd11an1n16x5 FILLER_366_886 ();
 b15zdnd11an1n04x5 FILLER_366_902 ();
 b15zdnd00an1n02x5 FILLER_366_906 ();
 b15zdnd00an1n01x5 FILLER_366_908 ();
 b15zdnd11an1n64x5 FILLER_366_921 ();
 b15zdnd11an1n64x5 FILLER_366_985 ();
 b15zdnd11an1n64x5 FILLER_366_1049 ();
 b15zdnd11an1n08x5 FILLER_366_1113 ();
 b15zdnd11an1n04x5 FILLER_366_1121 ();
 b15zdnd00an1n02x5 FILLER_366_1125 ();
 b15zdnd11an1n16x5 FILLER_366_1169 ();
 b15zdnd00an1n01x5 FILLER_366_1185 ();
 b15zdnd11an1n04x5 FILLER_366_1210 ();
 b15zdnd11an1n08x5 FILLER_366_1229 ();
 b15zdnd11an1n04x5 FILLER_366_1237 ();
 b15zdnd11an1n04x5 FILLER_366_1261 ();
 b15zdnd11an1n64x5 FILLER_366_1269 ();
 b15zdnd11an1n64x5 FILLER_366_1333 ();
 b15zdnd11an1n64x5 FILLER_366_1397 ();
 b15zdnd11an1n64x5 FILLER_366_1461 ();
 b15zdnd11an1n64x5 FILLER_366_1525 ();
 b15zdnd11an1n64x5 FILLER_366_1589 ();
 b15zdnd11an1n64x5 FILLER_366_1653 ();
 b15zdnd11an1n64x5 FILLER_366_1717 ();
 b15zdnd11an1n64x5 FILLER_366_1781 ();
 b15zdnd11an1n64x5 FILLER_366_1845 ();
 b15zdnd11an1n64x5 FILLER_366_1909 ();
 b15zdnd11an1n64x5 FILLER_366_1973 ();
 b15zdnd11an1n64x5 FILLER_366_2037 ();
 b15zdnd11an1n32x5 FILLER_366_2101 ();
 b15zdnd11an1n16x5 FILLER_366_2133 ();
 b15zdnd11an1n04x5 FILLER_366_2149 ();
 b15zdnd00an1n01x5 FILLER_366_2153 ();
 b15zdnd11an1n64x5 FILLER_366_2162 ();
 b15zdnd11an1n32x5 FILLER_366_2226 ();
 b15zdnd11an1n16x5 FILLER_366_2258 ();
 b15zdnd00an1n02x5 FILLER_366_2274 ();
 b15zdnd11an1n64x5 FILLER_367_0 ();
 b15zdnd11an1n64x5 FILLER_367_64 ();
 b15zdnd11an1n64x5 FILLER_367_128 ();
 b15zdnd11an1n64x5 FILLER_367_192 ();
 b15zdnd11an1n64x5 FILLER_367_256 ();
 b15zdnd11an1n32x5 FILLER_367_320 ();
 b15zdnd11an1n16x5 FILLER_367_352 ();
 b15zdnd11an1n04x5 FILLER_367_368 ();
 b15zdnd00an1n01x5 FILLER_367_372 ();
 b15zdnd11an1n64x5 FILLER_367_383 ();
 b15zdnd11an1n64x5 FILLER_367_447 ();
 b15zdnd11an1n64x5 FILLER_367_511 ();
 b15zdnd11an1n32x5 FILLER_367_575 ();
 b15zdnd11an1n64x5 FILLER_367_649 ();
 b15zdnd11an1n64x5 FILLER_367_713 ();
 b15zdnd11an1n32x5 FILLER_367_777 ();
 b15zdnd11an1n16x5 FILLER_367_809 ();
 b15zdnd11an1n04x5 FILLER_367_825 ();
 b15zdnd00an1n02x5 FILLER_367_829 ();
 b15zdnd00an1n01x5 FILLER_367_831 ();
 b15zdnd11an1n64x5 FILLER_367_874 ();
 b15zdnd11an1n64x5 FILLER_367_938 ();
 b15zdnd11an1n64x5 FILLER_367_1002 ();
 b15zdnd11an1n64x5 FILLER_367_1066 ();
 b15zdnd11an1n32x5 FILLER_367_1130 ();
 b15zdnd11an1n64x5 FILLER_367_1204 ();
 b15zdnd11an1n64x5 FILLER_367_1268 ();
 b15zdnd11an1n64x5 FILLER_367_1332 ();
 b15zdnd11an1n64x5 FILLER_367_1396 ();
 b15zdnd11an1n64x5 FILLER_367_1460 ();
 b15zdnd11an1n64x5 FILLER_367_1524 ();
 b15zdnd11an1n64x5 FILLER_367_1588 ();
 b15zdnd11an1n64x5 FILLER_367_1652 ();
 b15zdnd11an1n64x5 FILLER_367_1716 ();
 b15zdnd11an1n64x5 FILLER_367_1780 ();
 b15zdnd11an1n64x5 FILLER_367_1844 ();
 b15zdnd11an1n64x5 FILLER_367_1908 ();
 b15zdnd11an1n64x5 FILLER_367_1972 ();
 b15zdnd11an1n64x5 FILLER_367_2036 ();
 b15zdnd11an1n64x5 FILLER_367_2100 ();
 b15zdnd11an1n64x5 FILLER_367_2164 ();
 b15zdnd11an1n32x5 FILLER_367_2228 ();
 b15zdnd11an1n16x5 FILLER_367_2260 ();
 b15zdnd11an1n08x5 FILLER_367_2276 ();
 b15zdnd11an1n64x5 FILLER_368_8 ();
 b15zdnd11an1n64x5 FILLER_368_72 ();
 b15zdnd11an1n64x5 FILLER_368_136 ();
 b15zdnd11an1n64x5 FILLER_368_200 ();
 b15zdnd11an1n64x5 FILLER_368_264 ();
 b15zdnd11an1n64x5 FILLER_368_328 ();
 b15zdnd11an1n64x5 FILLER_368_392 ();
 b15zdnd11an1n64x5 FILLER_368_456 ();
 b15zdnd11an1n04x5 FILLER_368_520 ();
 b15zdnd00an1n02x5 FILLER_368_524 ();
 b15zdnd11an1n64x5 FILLER_368_568 ();
 b15zdnd11an1n64x5 FILLER_368_632 ();
 b15zdnd11an1n16x5 FILLER_368_696 ();
 b15zdnd11an1n04x5 FILLER_368_712 ();
 b15zdnd00an1n02x5 FILLER_368_716 ();
 b15zdnd11an1n64x5 FILLER_368_726 ();
 b15zdnd11an1n08x5 FILLER_368_790 ();
 b15zdnd00an1n02x5 FILLER_368_798 ();
 b15zdnd11an1n64x5 FILLER_368_842 ();
 b15zdnd11an1n64x5 FILLER_368_906 ();
 b15zdnd11an1n08x5 FILLER_368_970 ();
 b15zdnd00an1n01x5 FILLER_368_978 ();
 b15zdnd11an1n64x5 FILLER_368_1021 ();
 b15zdnd11an1n08x5 FILLER_368_1085 ();
 b15zdnd11an1n04x5 FILLER_368_1093 ();
 b15zdnd00an1n02x5 FILLER_368_1097 ();
 b15zdnd00an1n01x5 FILLER_368_1099 ();
 b15zdnd11an1n16x5 FILLER_368_1125 ();
 b15zdnd00an1n02x5 FILLER_368_1141 ();
 b15zdnd00an1n01x5 FILLER_368_1143 ();
 b15zdnd11an1n04x5 FILLER_368_1148 ();
 b15zdnd11an1n64x5 FILLER_368_1194 ();
 b15zdnd11an1n64x5 FILLER_368_1258 ();
 b15zdnd11an1n64x5 FILLER_368_1322 ();
 b15zdnd11an1n64x5 FILLER_368_1386 ();
 b15zdnd11an1n64x5 FILLER_368_1450 ();
 b15zdnd11an1n64x5 FILLER_368_1514 ();
 b15zdnd11an1n64x5 FILLER_368_1578 ();
 b15zdnd11an1n64x5 FILLER_368_1642 ();
 b15zdnd11an1n64x5 FILLER_368_1706 ();
 b15zdnd11an1n64x5 FILLER_368_1770 ();
 b15zdnd11an1n64x5 FILLER_368_1834 ();
 b15zdnd11an1n64x5 FILLER_368_1898 ();
 b15zdnd11an1n64x5 FILLER_368_1962 ();
 b15zdnd11an1n64x5 FILLER_368_2026 ();
 b15zdnd11an1n64x5 FILLER_368_2090 ();
 b15zdnd11an1n64x5 FILLER_368_2162 ();
 b15zdnd11an1n32x5 FILLER_368_2226 ();
 b15zdnd11an1n16x5 FILLER_368_2258 ();
 b15zdnd00an1n02x5 FILLER_368_2274 ();
 b15zdnd11an1n64x5 FILLER_369_0 ();
 b15zdnd11an1n64x5 FILLER_369_64 ();
 b15zdnd11an1n64x5 FILLER_369_128 ();
 b15zdnd11an1n64x5 FILLER_369_192 ();
 b15zdnd11an1n64x5 FILLER_369_256 ();
 b15zdnd11an1n64x5 FILLER_369_320 ();
 b15zdnd11an1n64x5 FILLER_369_384 ();
 b15zdnd11an1n32x5 FILLER_369_448 ();
 b15zdnd11an1n16x5 FILLER_369_480 ();
 b15zdnd11an1n08x5 FILLER_369_496 ();
 b15zdnd11an1n04x5 FILLER_369_504 ();
 b15zdnd00an1n01x5 FILLER_369_508 ();
 b15zdnd11an1n64x5 FILLER_369_551 ();
 b15zdnd11an1n64x5 FILLER_369_615 ();
 b15zdnd11an1n64x5 FILLER_369_679 ();
 b15zdnd11an1n32x5 FILLER_369_743 ();
 b15zdnd11an1n16x5 FILLER_369_775 ();
 b15zdnd11an1n04x5 FILLER_369_791 ();
 b15zdnd00an1n02x5 FILLER_369_795 ();
 b15zdnd11an1n64x5 FILLER_369_839 ();
 b15zdnd00an1n02x5 FILLER_369_903 ();
 b15zdnd00an1n01x5 FILLER_369_905 ();
 b15zdnd11an1n64x5 FILLER_369_948 ();
 b15zdnd11an1n08x5 FILLER_369_1012 ();
 b15zdnd00an1n02x5 FILLER_369_1020 ();
 b15zdnd00an1n01x5 FILLER_369_1022 ();
 b15zdnd11an1n64x5 FILLER_369_1065 ();
 b15zdnd11an1n08x5 FILLER_369_1129 ();
 b15zdnd00an1n02x5 FILLER_369_1137 ();
 b15zdnd11an1n64x5 FILLER_369_1181 ();
 b15zdnd11an1n64x5 FILLER_369_1245 ();
 b15zdnd11an1n64x5 FILLER_369_1309 ();
 b15zdnd11an1n64x5 FILLER_369_1373 ();
 b15zdnd11an1n64x5 FILLER_369_1437 ();
 b15zdnd11an1n64x5 FILLER_369_1501 ();
 b15zdnd11an1n64x5 FILLER_369_1565 ();
 b15zdnd11an1n64x5 FILLER_369_1629 ();
 b15zdnd11an1n64x5 FILLER_369_1693 ();
 b15zdnd11an1n64x5 FILLER_369_1757 ();
 b15zdnd11an1n64x5 FILLER_369_1821 ();
 b15zdnd11an1n64x5 FILLER_369_1885 ();
 b15zdnd11an1n64x5 FILLER_369_1949 ();
 b15zdnd11an1n64x5 FILLER_369_2013 ();
 b15zdnd11an1n64x5 FILLER_369_2077 ();
 b15zdnd11an1n64x5 FILLER_369_2141 ();
 b15zdnd11an1n64x5 FILLER_369_2205 ();
 b15zdnd11an1n08x5 FILLER_369_2269 ();
 b15zdnd11an1n04x5 FILLER_369_2277 ();
 b15zdnd00an1n02x5 FILLER_369_2281 ();
 b15zdnd00an1n01x5 FILLER_369_2283 ();
 b15zdnd11an1n64x5 FILLER_370_8 ();
 b15zdnd11an1n64x5 FILLER_370_72 ();
 b15zdnd11an1n64x5 FILLER_370_136 ();
 b15zdnd11an1n64x5 FILLER_370_200 ();
 b15zdnd11an1n64x5 FILLER_370_264 ();
 b15zdnd11an1n64x5 FILLER_370_328 ();
 b15zdnd11an1n32x5 FILLER_370_392 ();
 b15zdnd11an1n08x5 FILLER_370_424 ();
 b15zdnd11an1n32x5 FILLER_370_474 ();
 b15zdnd11an1n16x5 FILLER_370_506 ();
 b15zdnd11an1n08x5 FILLER_370_522 ();
 b15zdnd00an1n02x5 FILLER_370_530 ();
 b15zdnd00an1n01x5 FILLER_370_532 ();
 b15zdnd11an1n64x5 FILLER_370_537 ();
 b15zdnd11an1n64x5 FILLER_370_601 ();
 b15zdnd11an1n32x5 FILLER_370_665 ();
 b15zdnd11an1n16x5 FILLER_370_697 ();
 b15zdnd11an1n04x5 FILLER_370_713 ();
 b15zdnd00an1n01x5 FILLER_370_717 ();
 b15zdnd00an1n02x5 FILLER_370_726 ();
 b15zdnd11an1n64x5 FILLER_370_770 ();
 b15zdnd11an1n64x5 FILLER_370_834 ();
 b15zdnd11an1n64x5 FILLER_370_898 ();
 b15zdnd11an1n64x5 FILLER_370_962 ();
 b15zdnd11an1n64x5 FILLER_370_1026 ();
 b15zdnd11an1n16x5 FILLER_370_1090 ();
 b15zdnd11an1n04x5 FILLER_370_1106 ();
 b15zdnd00an1n01x5 FILLER_370_1110 ();
 b15zdnd11an1n08x5 FILLER_370_1131 ();
 b15zdnd11an1n04x5 FILLER_370_1139 ();
 b15zdnd00an1n02x5 FILLER_370_1143 ();
 b15zdnd11an1n64x5 FILLER_370_1187 ();
 b15zdnd11an1n64x5 FILLER_370_1251 ();
 b15zdnd11an1n64x5 FILLER_370_1315 ();
 b15zdnd11an1n64x5 FILLER_370_1379 ();
 b15zdnd11an1n64x5 FILLER_370_1443 ();
 b15zdnd11an1n64x5 FILLER_370_1507 ();
 b15zdnd11an1n64x5 FILLER_370_1571 ();
 b15zdnd11an1n64x5 FILLER_370_1635 ();
 b15zdnd11an1n64x5 FILLER_370_1699 ();
 b15zdnd11an1n64x5 FILLER_370_1763 ();
 b15zdnd11an1n64x5 FILLER_370_1827 ();
 b15zdnd11an1n64x5 FILLER_370_1891 ();
 b15zdnd11an1n64x5 FILLER_370_1955 ();
 b15zdnd11an1n64x5 FILLER_370_2019 ();
 b15zdnd11an1n64x5 FILLER_370_2083 ();
 b15zdnd11an1n04x5 FILLER_370_2147 ();
 b15zdnd00an1n02x5 FILLER_370_2151 ();
 b15zdnd00an1n01x5 FILLER_370_2153 ();
 b15zdnd11an1n64x5 FILLER_370_2162 ();
 b15zdnd11an1n32x5 FILLER_370_2226 ();
 b15zdnd11an1n16x5 FILLER_370_2258 ();
 b15zdnd00an1n02x5 FILLER_370_2274 ();
 b15zdnd11an1n64x5 FILLER_371_0 ();
 b15zdnd11an1n64x5 FILLER_371_64 ();
 b15zdnd11an1n64x5 FILLER_371_128 ();
 b15zdnd11an1n64x5 FILLER_371_192 ();
 b15zdnd11an1n64x5 FILLER_371_256 ();
 b15zdnd11an1n64x5 FILLER_371_320 ();
 b15zdnd11an1n64x5 FILLER_371_384 ();
 b15zdnd11an1n64x5 FILLER_371_448 ();
 b15zdnd11an1n64x5 FILLER_371_512 ();
 b15zdnd11an1n64x5 FILLER_371_576 ();
 b15zdnd11an1n32x5 FILLER_371_640 ();
 b15zdnd11an1n16x5 FILLER_371_714 ();
 b15zdnd11an1n08x5 FILLER_371_730 ();
 b15zdnd00an1n02x5 FILLER_371_738 ();
 b15zdnd00an1n01x5 FILLER_371_740 ();
 b15zdnd11an1n16x5 FILLER_371_783 ();
 b15zdnd11an1n64x5 FILLER_371_841 ();
 b15zdnd11an1n64x5 FILLER_371_905 ();
 b15zdnd11an1n64x5 FILLER_371_969 ();
 b15zdnd11an1n64x5 FILLER_371_1033 ();
 b15zdnd11an1n04x5 FILLER_371_1097 ();
 b15zdnd00an1n02x5 FILLER_371_1101 ();
 b15zdnd11an1n08x5 FILLER_371_1134 ();
 b15zdnd11an1n04x5 FILLER_371_1142 ();
 b15zdnd00an1n02x5 FILLER_371_1146 ();
 b15zdnd11an1n64x5 FILLER_371_1190 ();
 b15zdnd11an1n64x5 FILLER_371_1254 ();
 b15zdnd11an1n64x5 FILLER_371_1318 ();
 b15zdnd11an1n64x5 FILLER_371_1382 ();
 b15zdnd11an1n64x5 FILLER_371_1446 ();
 b15zdnd11an1n64x5 FILLER_371_1510 ();
 b15zdnd11an1n64x5 FILLER_371_1574 ();
 b15zdnd11an1n64x5 FILLER_371_1638 ();
 b15zdnd11an1n64x5 FILLER_371_1702 ();
 b15zdnd11an1n64x5 FILLER_371_1766 ();
 b15zdnd11an1n64x5 FILLER_371_1830 ();
 b15zdnd11an1n64x5 FILLER_371_1894 ();
 b15zdnd11an1n64x5 FILLER_371_1958 ();
 b15zdnd11an1n64x5 FILLER_371_2022 ();
 b15zdnd11an1n64x5 FILLER_371_2086 ();
 b15zdnd11an1n64x5 FILLER_371_2150 ();
 b15zdnd11an1n64x5 FILLER_371_2214 ();
 b15zdnd11an1n04x5 FILLER_371_2278 ();
 b15zdnd00an1n02x5 FILLER_371_2282 ();
 b15zdnd11an1n64x5 FILLER_372_8 ();
 b15zdnd11an1n64x5 FILLER_372_72 ();
 b15zdnd11an1n64x5 FILLER_372_136 ();
 b15zdnd11an1n64x5 FILLER_372_200 ();
 b15zdnd11an1n64x5 FILLER_372_264 ();
 b15zdnd11an1n64x5 FILLER_372_328 ();
 b15zdnd11an1n64x5 FILLER_372_392 ();
 b15zdnd11an1n64x5 FILLER_372_456 ();
 b15zdnd11an1n32x5 FILLER_372_520 ();
 b15zdnd11an1n16x5 FILLER_372_594 ();
 b15zdnd11an1n08x5 FILLER_372_610 ();
 b15zdnd11an1n04x5 FILLER_372_660 ();
 b15zdnd11an1n08x5 FILLER_372_706 ();
 b15zdnd11an1n04x5 FILLER_372_714 ();
 b15zdnd11an1n64x5 FILLER_372_726 ();
 b15zdnd11an1n64x5 FILLER_372_790 ();
 b15zdnd11an1n64x5 FILLER_372_854 ();
 b15zdnd11an1n64x5 FILLER_372_918 ();
 b15zdnd11an1n64x5 FILLER_372_982 ();
 b15zdnd11an1n64x5 FILLER_372_1046 ();
 b15zdnd11an1n64x5 FILLER_372_1110 ();
 b15zdnd11an1n32x5 FILLER_372_1174 ();
 b15zdnd11an1n16x5 FILLER_372_1206 ();
 b15zdnd11an1n08x5 FILLER_372_1222 ();
 b15zdnd11an1n04x5 FILLER_372_1230 ();
 b15zdnd00an1n02x5 FILLER_372_1234 ();
 b15zdnd00an1n01x5 FILLER_372_1236 ();
 b15zdnd11an1n64x5 FILLER_372_1279 ();
 b15zdnd11an1n64x5 FILLER_372_1343 ();
 b15zdnd11an1n64x5 FILLER_372_1407 ();
 b15zdnd11an1n64x5 FILLER_372_1471 ();
 b15zdnd11an1n64x5 FILLER_372_1535 ();
 b15zdnd11an1n64x5 FILLER_372_1599 ();
 b15zdnd11an1n64x5 FILLER_372_1663 ();
 b15zdnd11an1n64x5 FILLER_372_1727 ();
 b15zdnd11an1n64x5 FILLER_372_1791 ();
 b15zdnd11an1n64x5 FILLER_372_1855 ();
 b15zdnd11an1n64x5 FILLER_372_1919 ();
 b15zdnd11an1n64x5 FILLER_372_1983 ();
 b15zdnd11an1n64x5 FILLER_372_2047 ();
 b15zdnd11an1n32x5 FILLER_372_2111 ();
 b15zdnd11an1n08x5 FILLER_372_2143 ();
 b15zdnd00an1n02x5 FILLER_372_2151 ();
 b15zdnd00an1n01x5 FILLER_372_2153 ();
 b15zdnd11an1n64x5 FILLER_372_2162 ();
 b15zdnd11an1n32x5 FILLER_372_2226 ();
 b15zdnd11an1n16x5 FILLER_372_2258 ();
 b15zdnd00an1n02x5 FILLER_372_2274 ();
 b15zdnd11an1n64x5 FILLER_373_0 ();
 b15zdnd11an1n64x5 FILLER_373_64 ();
 b15zdnd11an1n64x5 FILLER_373_128 ();
 b15zdnd11an1n64x5 FILLER_373_192 ();
 b15zdnd11an1n64x5 FILLER_373_256 ();
 b15zdnd11an1n64x5 FILLER_373_320 ();
 b15zdnd11an1n64x5 FILLER_373_384 ();
 b15zdnd11an1n64x5 FILLER_373_448 ();
 b15zdnd11an1n64x5 FILLER_373_512 ();
 b15zdnd11an1n32x5 FILLER_373_576 ();
 b15zdnd11an1n16x5 FILLER_373_608 ();
 b15zdnd00an1n02x5 FILLER_373_624 ();
 b15zdnd00an1n01x5 FILLER_373_626 ();
 b15zdnd11an1n32x5 FILLER_373_669 ();
 b15zdnd11an1n04x5 FILLER_373_701 ();
 b15zdnd11an1n04x5 FILLER_373_747 ();
 b15zdnd11an1n32x5 FILLER_373_793 ();
 b15zdnd11an1n08x5 FILLER_373_825 ();
 b15zdnd11an1n04x5 FILLER_373_833 ();
 b15zdnd00an1n02x5 FILLER_373_837 ();
 b15zdnd11an1n64x5 FILLER_373_881 ();
 b15zdnd11an1n08x5 FILLER_373_945 ();
 b15zdnd11an1n04x5 FILLER_373_953 ();
 b15zdnd00an1n02x5 FILLER_373_957 ();
 b15zdnd00an1n01x5 FILLER_373_959 ();
 b15zdnd11an1n64x5 FILLER_373_977 ();
 b15zdnd11an1n64x5 FILLER_373_1041 ();
 b15zdnd11an1n64x5 FILLER_373_1105 ();
 b15zdnd11an1n32x5 FILLER_373_1169 ();
 b15zdnd11an1n16x5 FILLER_373_1201 ();
 b15zdnd11an1n04x5 FILLER_373_1217 ();
 b15zdnd00an1n02x5 FILLER_373_1221 ();
 b15zdnd00an1n01x5 FILLER_373_1223 ();
 b15zdnd11an1n04x5 FILLER_373_1266 ();
 b15zdnd11an1n64x5 FILLER_373_1312 ();
 b15zdnd11an1n64x5 FILLER_373_1376 ();
 b15zdnd11an1n64x5 FILLER_373_1440 ();
 b15zdnd11an1n64x5 FILLER_373_1504 ();
 b15zdnd11an1n64x5 FILLER_373_1568 ();
 b15zdnd11an1n64x5 FILLER_373_1632 ();
 b15zdnd11an1n64x5 FILLER_373_1696 ();
 b15zdnd11an1n64x5 FILLER_373_1760 ();
 b15zdnd11an1n64x5 FILLER_373_1824 ();
 b15zdnd11an1n64x5 FILLER_373_1888 ();
 b15zdnd11an1n64x5 FILLER_373_1952 ();
 b15zdnd11an1n64x5 FILLER_373_2016 ();
 b15zdnd11an1n64x5 FILLER_373_2080 ();
 b15zdnd11an1n64x5 FILLER_373_2144 ();
 b15zdnd11an1n64x5 FILLER_373_2208 ();
 b15zdnd11an1n08x5 FILLER_373_2272 ();
 b15zdnd11an1n04x5 FILLER_373_2280 ();
 b15zdnd11an1n64x5 FILLER_374_8 ();
 b15zdnd11an1n64x5 FILLER_374_72 ();
 b15zdnd11an1n64x5 FILLER_374_136 ();
 b15zdnd11an1n64x5 FILLER_374_200 ();
 b15zdnd11an1n64x5 FILLER_374_264 ();
 b15zdnd11an1n64x5 FILLER_374_328 ();
 b15zdnd11an1n64x5 FILLER_374_392 ();
 b15zdnd11an1n64x5 FILLER_374_456 ();
 b15zdnd11an1n16x5 FILLER_374_520 ();
 b15zdnd11an1n04x5 FILLER_374_536 ();
 b15zdnd00an1n02x5 FILLER_374_540 ();
 b15zdnd11an1n32x5 FILLER_374_568 ();
 b15zdnd11an1n08x5 FILLER_374_600 ();
 b15zdnd00an1n01x5 FILLER_374_608 ();
 b15zdnd11an1n64x5 FILLER_374_613 ();
 b15zdnd11an1n32x5 FILLER_374_677 ();
 b15zdnd11an1n08x5 FILLER_374_709 ();
 b15zdnd00an1n01x5 FILLER_374_717 ();
 b15zdnd11an1n32x5 FILLER_374_726 ();
 b15zdnd11an1n04x5 FILLER_374_758 ();
 b15zdnd00an1n02x5 FILLER_374_762 ();
 b15zdnd11an1n64x5 FILLER_374_795 ();
 b15zdnd11an1n64x5 FILLER_374_859 ();
 b15zdnd11an1n64x5 FILLER_374_923 ();
 b15zdnd11an1n08x5 FILLER_374_987 ();
 b15zdnd11an1n32x5 FILLER_374_999 ();
 b15zdnd11an1n08x5 FILLER_374_1031 ();
 b15zdnd11an1n64x5 FILLER_374_1054 ();
 b15zdnd11an1n64x5 FILLER_374_1118 ();
 b15zdnd11an1n64x5 FILLER_374_1182 ();
 b15zdnd11an1n64x5 FILLER_374_1246 ();
 b15zdnd11an1n64x5 FILLER_374_1310 ();
 b15zdnd11an1n64x5 FILLER_374_1374 ();
 b15zdnd11an1n64x5 FILLER_374_1438 ();
 b15zdnd11an1n64x5 FILLER_374_1502 ();
 b15zdnd11an1n64x5 FILLER_374_1566 ();
 b15zdnd11an1n64x5 FILLER_374_1630 ();
 b15zdnd11an1n64x5 FILLER_374_1694 ();
 b15zdnd11an1n64x5 FILLER_374_1758 ();
 b15zdnd11an1n64x5 FILLER_374_1822 ();
 b15zdnd11an1n64x5 FILLER_374_1886 ();
 b15zdnd11an1n64x5 FILLER_374_1950 ();
 b15zdnd11an1n64x5 FILLER_374_2014 ();
 b15zdnd11an1n64x5 FILLER_374_2078 ();
 b15zdnd11an1n08x5 FILLER_374_2142 ();
 b15zdnd11an1n04x5 FILLER_374_2150 ();
 b15zdnd11an1n64x5 FILLER_374_2162 ();
 b15zdnd11an1n32x5 FILLER_374_2226 ();
 b15zdnd11an1n16x5 FILLER_374_2258 ();
 b15zdnd00an1n02x5 FILLER_374_2274 ();
 b15zdnd11an1n64x5 FILLER_375_0 ();
 b15zdnd11an1n64x5 FILLER_375_64 ();
 b15zdnd11an1n64x5 FILLER_375_128 ();
 b15zdnd11an1n64x5 FILLER_375_192 ();
 b15zdnd11an1n64x5 FILLER_375_256 ();
 b15zdnd11an1n64x5 FILLER_375_320 ();
 b15zdnd11an1n64x5 FILLER_375_384 ();
 b15zdnd11an1n64x5 FILLER_375_448 ();
 b15zdnd11an1n16x5 FILLER_375_512 ();
 b15zdnd11an1n08x5 FILLER_375_528 ();
 b15zdnd00an1n01x5 FILLER_375_536 ();
 b15zdnd11an1n04x5 FILLER_375_540 ();
 b15zdnd11an1n04x5 FILLER_375_558 ();
 b15zdnd11an1n16x5 FILLER_375_566 ();
 b15zdnd11an1n08x5 FILLER_375_582 ();
 b15zdnd11an1n04x5 FILLER_375_590 ();
 b15zdnd00an1n02x5 FILLER_375_594 ();
 b15zdnd11an1n04x5 FILLER_375_604 ();
 b15zdnd11an1n64x5 FILLER_375_650 ();
 b15zdnd11an1n32x5 FILLER_375_714 ();
 b15zdnd11an1n16x5 FILLER_375_746 ();
 b15zdnd11an1n08x5 FILLER_375_762 ();
 b15zdnd11an1n04x5 FILLER_375_770 ();
 b15zdnd00an1n02x5 FILLER_375_774 ();
 b15zdnd00an1n01x5 FILLER_375_776 ();
 b15zdnd11an1n16x5 FILLER_375_789 ();
 b15zdnd11an1n04x5 FILLER_375_805 ();
 b15zdnd00an1n02x5 FILLER_375_809 ();
 b15zdnd00an1n01x5 FILLER_375_811 ();
 b15zdnd11an1n64x5 FILLER_375_827 ();
 b15zdnd11an1n08x5 FILLER_375_891 ();
 b15zdnd00an1n01x5 FILLER_375_899 ();
 b15zdnd11an1n16x5 FILLER_375_905 ();
 b15zdnd11an1n04x5 FILLER_375_921 ();
 b15zdnd00an1n01x5 FILLER_375_925 ();
 b15zdnd11an1n08x5 FILLER_375_930 ();
 b15zdnd11an1n04x5 FILLER_375_950 ();
 b15zdnd00an1n01x5 FILLER_375_954 ();
 b15zdnd11an1n64x5 FILLER_375_958 ();
 b15zdnd11an1n08x5 FILLER_375_1022 ();
 b15zdnd11an1n04x5 FILLER_375_1030 ();
 b15zdnd00an1n02x5 FILLER_375_1034 ();
 b15zdnd11an1n64x5 FILLER_375_1053 ();
 b15zdnd11an1n16x5 FILLER_375_1117 ();
 b15zdnd00an1n01x5 FILLER_375_1133 ();
 b15zdnd11an1n64x5 FILLER_375_1176 ();
 b15zdnd11an1n64x5 FILLER_375_1240 ();
 b15zdnd11an1n64x5 FILLER_375_1304 ();
 b15zdnd11an1n64x5 FILLER_375_1368 ();
 b15zdnd11an1n64x5 FILLER_375_1432 ();
 b15zdnd11an1n64x5 FILLER_375_1496 ();
 b15zdnd11an1n64x5 FILLER_375_1560 ();
 b15zdnd11an1n64x5 FILLER_375_1624 ();
 b15zdnd11an1n64x5 FILLER_375_1688 ();
 b15zdnd11an1n64x5 FILLER_375_1752 ();
 b15zdnd11an1n64x5 FILLER_375_1816 ();
 b15zdnd11an1n64x5 FILLER_375_1880 ();
 b15zdnd11an1n64x5 FILLER_375_1944 ();
 b15zdnd11an1n64x5 FILLER_375_2008 ();
 b15zdnd11an1n64x5 FILLER_375_2072 ();
 b15zdnd11an1n64x5 FILLER_375_2136 ();
 b15zdnd11an1n64x5 FILLER_375_2200 ();
 b15zdnd11an1n16x5 FILLER_375_2264 ();
 b15zdnd11an1n04x5 FILLER_375_2280 ();
 b15zdnd11an1n16x5 FILLER_376_8 ();
 b15zdnd00an1n02x5 FILLER_376_24 ();
 b15zdnd11an1n64x5 FILLER_376_32 ();
 b15zdnd11an1n64x5 FILLER_376_96 ();
 b15zdnd11an1n64x5 FILLER_376_160 ();
 b15zdnd11an1n64x5 FILLER_376_224 ();
 b15zdnd11an1n64x5 FILLER_376_288 ();
 b15zdnd11an1n64x5 FILLER_376_352 ();
 b15zdnd11an1n64x5 FILLER_376_416 ();
 b15zdnd11an1n32x5 FILLER_376_480 ();
 b15zdnd11an1n16x5 FILLER_376_512 ();
 b15zdnd11an1n04x5 FILLER_376_528 ();
 b15zdnd00an1n02x5 FILLER_376_532 ();
 b15zdnd00an1n01x5 FILLER_376_534 ();
 b15zdnd11an1n04x5 FILLER_376_538 ();
 b15zdnd00an1n01x5 FILLER_376_542 ();
 b15zdnd11an1n04x5 FILLER_376_558 ();
 b15zdnd11an1n08x5 FILLER_376_567 ();
 b15zdnd00an1n01x5 FILLER_376_575 ();
 b15zdnd11an1n32x5 FILLER_376_581 ();
 b15zdnd11an1n16x5 FILLER_376_613 ();
 b15zdnd11an1n08x5 FILLER_376_629 ();
 b15zdnd00an1n02x5 FILLER_376_637 ();
 b15zdnd11an1n32x5 FILLER_376_659 ();
 b15zdnd11an1n16x5 FILLER_376_691 ();
 b15zdnd11an1n08x5 FILLER_376_707 ();
 b15zdnd00an1n02x5 FILLER_376_715 ();
 b15zdnd00an1n01x5 FILLER_376_717 ();
 b15zdnd11an1n32x5 FILLER_376_726 ();
 b15zdnd11an1n16x5 FILLER_376_758 ();
 b15zdnd11an1n08x5 FILLER_376_774 ();
 b15zdnd11an1n04x5 FILLER_376_782 ();
 b15zdnd00an1n01x5 FILLER_376_786 ();
 b15zdnd11an1n08x5 FILLER_376_792 ();
 b15zdnd11an1n04x5 FILLER_376_810 ();
 b15zdnd11an1n64x5 FILLER_376_819 ();
 b15zdnd11an1n16x5 FILLER_376_883 ();
 b15zdnd00an1n02x5 FILLER_376_899 ();
 b15zdnd00an1n01x5 FILLER_376_901 ();
 b15zdnd11an1n04x5 FILLER_376_919 ();
 b15zdnd11an1n32x5 FILLER_376_965 ();
 b15zdnd11an1n08x5 FILLER_376_997 ();
 b15zdnd11an1n04x5 FILLER_376_1005 ();
 b15zdnd00an1n02x5 FILLER_376_1009 ();
 b15zdnd00an1n01x5 FILLER_376_1011 ();
 b15zdnd11an1n04x5 FILLER_376_1017 ();
 b15zdnd00an1n02x5 FILLER_376_1021 ();
 b15zdnd11an1n04x5 FILLER_376_1030 ();
 b15zdnd11an1n04x5 FILLER_376_1038 ();
 b15zdnd11an1n64x5 FILLER_376_1054 ();
 b15zdnd11an1n64x5 FILLER_376_1118 ();
 b15zdnd11an1n64x5 FILLER_376_1182 ();
 b15zdnd11an1n64x5 FILLER_376_1246 ();
 b15zdnd11an1n64x5 FILLER_376_1310 ();
 b15zdnd11an1n64x5 FILLER_376_1374 ();
 b15zdnd11an1n64x5 FILLER_376_1438 ();
 b15zdnd11an1n64x5 FILLER_376_1502 ();
 b15zdnd11an1n64x5 FILLER_376_1566 ();
 b15zdnd11an1n64x5 FILLER_376_1630 ();
 b15zdnd11an1n64x5 FILLER_376_1694 ();
 b15zdnd11an1n64x5 FILLER_376_1758 ();
 b15zdnd11an1n64x5 FILLER_376_1822 ();
 b15zdnd11an1n64x5 FILLER_376_1886 ();
 b15zdnd11an1n64x5 FILLER_376_1950 ();
 b15zdnd11an1n64x5 FILLER_376_2014 ();
 b15zdnd11an1n64x5 FILLER_376_2078 ();
 b15zdnd11an1n08x5 FILLER_376_2142 ();
 b15zdnd11an1n04x5 FILLER_376_2150 ();
 b15zdnd11an1n64x5 FILLER_376_2162 ();
 b15zdnd11an1n32x5 FILLER_376_2226 ();
 b15zdnd11an1n16x5 FILLER_376_2258 ();
 b15zdnd00an1n02x5 FILLER_376_2274 ();
 b15zdnd11an1n08x5 FILLER_377_0 ();
 b15zdnd11an1n64x5 FILLER_377_50 ();
 b15zdnd11an1n64x5 FILLER_377_114 ();
 b15zdnd11an1n64x5 FILLER_377_178 ();
 b15zdnd11an1n64x5 FILLER_377_242 ();
 b15zdnd11an1n64x5 FILLER_377_306 ();
 b15zdnd11an1n64x5 FILLER_377_370 ();
 b15zdnd11an1n64x5 FILLER_377_434 ();
 b15zdnd11an1n32x5 FILLER_377_498 ();
 b15zdnd11an1n08x5 FILLER_377_530 ();
 b15zdnd11an1n04x5 FILLER_377_538 ();
 b15zdnd00an1n02x5 FILLER_377_542 ();
 b15zdnd11an1n04x5 FILLER_377_551 ();
 b15zdnd11an1n64x5 FILLER_377_597 ();
 b15zdnd11an1n64x5 FILLER_377_661 ();
 b15zdnd11an1n32x5 FILLER_377_725 ();
 b15zdnd11an1n16x5 FILLER_377_757 ();
 b15zdnd11an1n08x5 FILLER_377_787 ();
 b15zdnd11an1n04x5 FILLER_377_795 ();
 b15zdnd00an1n02x5 FILLER_377_799 ();
 b15zdnd00an1n01x5 FILLER_377_801 ();
 b15zdnd11an1n04x5 FILLER_377_806 ();
 b15zdnd00an1n01x5 FILLER_377_810 ();
 b15zdnd11an1n16x5 FILLER_377_822 ();
 b15zdnd11an1n08x5 FILLER_377_838 ();
 b15zdnd00an1n02x5 FILLER_377_846 ();
 b15zdnd11an1n16x5 FILLER_377_853 ();
 b15zdnd11an1n08x5 FILLER_377_869 ();
 b15zdnd11an1n08x5 FILLER_377_884 ();
 b15zdnd11an1n04x5 FILLER_377_892 ();
 b15zdnd00an1n02x5 FILLER_377_896 ();
 b15zdnd00an1n01x5 FILLER_377_898 ();
 b15zdnd11an1n04x5 FILLER_377_909 ();
 b15zdnd11an1n32x5 FILLER_377_916 ();
 b15zdnd11an1n08x5 FILLER_377_948 ();
 b15zdnd11an1n04x5 FILLER_377_956 ();
 b15zdnd00an1n02x5 FILLER_377_960 ();
 b15zdnd00an1n01x5 FILLER_377_962 ();
 b15zdnd11an1n08x5 FILLER_377_968 ();
 b15zdnd11an1n04x5 FILLER_377_976 ();
 b15zdnd00an1n02x5 FILLER_377_980 ();
 b15zdnd11an1n08x5 FILLER_377_1024 ();
 b15zdnd11an1n04x5 FILLER_377_1032 ();
 b15zdnd00an1n02x5 FILLER_377_1036 ();
 b15zdnd11an1n04x5 FILLER_377_1043 ();
 b15zdnd11an1n04x5 FILLER_377_1064 ();
 b15zdnd11an1n64x5 FILLER_377_1072 ();
 b15zdnd11an1n64x5 FILLER_377_1136 ();
 b15zdnd11an1n64x5 FILLER_377_1200 ();
 b15zdnd11an1n64x5 FILLER_377_1264 ();
 b15zdnd11an1n64x5 FILLER_377_1328 ();
 b15zdnd11an1n64x5 FILLER_377_1392 ();
 b15zdnd11an1n64x5 FILLER_377_1456 ();
 b15zdnd11an1n64x5 FILLER_377_1520 ();
 b15zdnd11an1n64x5 FILLER_377_1584 ();
 b15zdnd11an1n64x5 FILLER_377_1648 ();
 b15zdnd11an1n64x5 FILLER_377_1712 ();
 b15zdnd11an1n64x5 FILLER_377_1776 ();
 b15zdnd11an1n64x5 FILLER_377_1840 ();
 b15zdnd11an1n64x5 FILLER_377_1904 ();
 b15zdnd11an1n64x5 FILLER_377_1968 ();
 b15zdnd11an1n64x5 FILLER_377_2032 ();
 b15zdnd11an1n64x5 FILLER_377_2096 ();
 b15zdnd11an1n64x5 FILLER_377_2160 ();
 b15zdnd11an1n32x5 FILLER_377_2224 ();
 b15zdnd11an1n16x5 FILLER_377_2256 ();
 b15zdnd11an1n08x5 FILLER_377_2272 ();
 b15zdnd11an1n04x5 FILLER_377_2280 ();
 b15zdnd11an1n64x5 FILLER_378_8 ();
 b15zdnd11an1n64x5 FILLER_378_72 ();
 b15zdnd11an1n64x5 FILLER_378_136 ();
 b15zdnd11an1n64x5 FILLER_378_200 ();
 b15zdnd11an1n64x5 FILLER_378_264 ();
 b15zdnd11an1n64x5 FILLER_378_328 ();
 b15zdnd11an1n64x5 FILLER_378_392 ();
 b15zdnd11an1n64x5 FILLER_378_456 ();
 b15zdnd11an1n32x5 FILLER_378_520 ();
 b15zdnd11an1n08x5 FILLER_378_552 ();
 b15zdnd11an1n64x5 FILLER_378_573 ();
 b15zdnd11an1n32x5 FILLER_378_637 ();
 b15zdnd11an1n16x5 FILLER_378_669 ();
 b15zdnd11an1n04x5 FILLER_378_685 ();
 b15zdnd00an1n02x5 FILLER_378_689 ();
 b15zdnd11an1n08x5 FILLER_378_695 ();
 b15zdnd00an1n01x5 FILLER_378_703 ();
 b15zdnd11an1n08x5 FILLER_378_710 ();
 b15zdnd00an1n02x5 FILLER_378_726 ();
 b15zdnd11an1n04x5 FILLER_378_770 ();
 b15zdnd11an1n04x5 FILLER_378_791 ();
 b15zdnd00an1n02x5 FILLER_378_795 ();
 b15zdnd11an1n04x5 FILLER_378_805 ();
 b15zdnd11an1n16x5 FILLER_378_819 ();
 b15zdnd11an1n08x5 FILLER_378_835 ();
 b15zdnd11an1n04x5 FILLER_378_843 ();
 b15zdnd11an1n08x5 FILLER_378_857 ();
 b15zdnd11an1n04x5 FILLER_378_907 ();
 b15zdnd11an1n16x5 FILLER_378_921 ();
 b15zdnd11an1n08x5 FILLER_378_937 ();
 b15zdnd11an1n04x5 FILLER_378_945 ();
 b15zdnd00an1n01x5 FILLER_378_949 ();
 b15zdnd11an1n16x5 FILLER_378_992 ();
 b15zdnd11an1n04x5 FILLER_378_1050 ();
 b15zdnd00an1n01x5 FILLER_378_1054 ();
 b15zdnd11an1n32x5 FILLER_378_1097 ();
 b15zdnd11an1n16x5 FILLER_378_1129 ();
 b15zdnd00an1n02x5 FILLER_378_1145 ();
 b15zdnd00an1n01x5 FILLER_378_1147 ();
 b15zdnd11an1n64x5 FILLER_378_1153 ();
 b15zdnd11an1n64x5 FILLER_378_1217 ();
 b15zdnd11an1n64x5 FILLER_378_1281 ();
 b15zdnd11an1n64x5 FILLER_378_1345 ();
 b15zdnd11an1n64x5 FILLER_378_1409 ();
 b15zdnd11an1n64x5 FILLER_378_1473 ();
 b15zdnd11an1n64x5 FILLER_378_1537 ();
 b15zdnd11an1n64x5 FILLER_378_1601 ();
 b15zdnd11an1n64x5 FILLER_378_1665 ();
 b15zdnd11an1n64x5 FILLER_378_1729 ();
 b15zdnd11an1n64x5 FILLER_378_1793 ();
 b15zdnd11an1n64x5 FILLER_378_1857 ();
 b15zdnd11an1n64x5 FILLER_378_1921 ();
 b15zdnd11an1n64x5 FILLER_378_1985 ();
 b15zdnd11an1n64x5 FILLER_378_2049 ();
 b15zdnd11an1n32x5 FILLER_378_2113 ();
 b15zdnd11an1n08x5 FILLER_378_2145 ();
 b15zdnd00an1n01x5 FILLER_378_2153 ();
 b15zdnd11an1n64x5 FILLER_378_2162 ();
 b15zdnd11an1n32x5 FILLER_378_2226 ();
 b15zdnd11an1n16x5 FILLER_378_2258 ();
 b15zdnd00an1n02x5 FILLER_378_2274 ();
 b15zdnd11an1n64x5 FILLER_379_0 ();
 b15zdnd11an1n64x5 FILLER_379_64 ();
 b15zdnd11an1n64x5 FILLER_379_128 ();
 b15zdnd11an1n64x5 FILLER_379_192 ();
 b15zdnd11an1n64x5 FILLER_379_256 ();
 b15zdnd11an1n64x5 FILLER_379_320 ();
 b15zdnd11an1n64x5 FILLER_379_384 ();
 b15zdnd11an1n64x5 FILLER_379_448 ();
 b15zdnd11an1n32x5 FILLER_379_512 ();
 b15zdnd11an1n08x5 FILLER_379_544 ();
 b15zdnd00an1n01x5 FILLER_379_552 ();
 b15zdnd11an1n04x5 FILLER_379_562 ();
 b15zdnd11an1n64x5 FILLER_379_576 ();
 b15zdnd11an1n64x5 FILLER_379_640 ();
 b15zdnd11an1n64x5 FILLER_379_704 ();
 b15zdnd11an1n04x5 FILLER_379_768 ();
 b15zdnd00an1n02x5 FILLER_379_772 ();
 b15zdnd11an1n04x5 FILLER_379_778 ();
 b15zdnd11an1n16x5 FILLER_379_796 ();
 b15zdnd11an1n16x5 FILLER_379_820 ();
 b15zdnd00an1n02x5 FILLER_379_836 ();
 b15zdnd11an1n32x5 FILLER_379_880 ();
 b15zdnd11an1n16x5 FILLER_379_912 ();
 b15zdnd11an1n04x5 FILLER_379_928 ();
 b15zdnd00an1n01x5 FILLER_379_932 ();
 b15zdnd11an1n32x5 FILLER_379_975 ();
 b15zdnd11an1n04x5 FILLER_379_1007 ();
 b15zdnd00an1n02x5 FILLER_379_1011 ();
 b15zdnd00an1n01x5 FILLER_379_1013 ();
 b15zdnd11an1n16x5 FILLER_379_1021 ();
 b15zdnd11an1n04x5 FILLER_379_1037 ();
 b15zdnd00an1n01x5 FILLER_379_1041 ();
 b15zdnd11an1n04x5 FILLER_379_1045 ();
 b15zdnd11an1n32x5 FILLER_379_1091 ();
 b15zdnd11an1n04x5 FILLER_379_1123 ();
 b15zdnd11an1n64x5 FILLER_379_1169 ();
 b15zdnd11an1n64x5 FILLER_379_1233 ();
 b15zdnd11an1n64x5 FILLER_379_1297 ();
 b15zdnd11an1n64x5 FILLER_379_1361 ();
 b15zdnd11an1n64x5 FILLER_379_1425 ();
 b15zdnd11an1n64x5 FILLER_379_1489 ();
 b15zdnd11an1n64x5 FILLER_379_1553 ();
 b15zdnd11an1n64x5 FILLER_379_1617 ();
 b15zdnd11an1n64x5 FILLER_379_1681 ();
 b15zdnd11an1n64x5 FILLER_379_1745 ();
 b15zdnd11an1n64x5 FILLER_379_1809 ();
 b15zdnd11an1n64x5 FILLER_379_1873 ();
 b15zdnd11an1n64x5 FILLER_379_1937 ();
 b15zdnd11an1n64x5 FILLER_379_2001 ();
 b15zdnd11an1n64x5 FILLER_379_2065 ();
 b15zdnd11an1n64x5 FILLER_379_2129 ();
 b15zdnd11an1n64x5 FILLER_379_2193 ();
 b15zdnd11an1n16x5 FILLER_379_2257 ();
 b15zdnd11an1n08x5 FILLER_379_2273 ();
 b15zdnd00an1n02x5 FILLER_379_2281 ();
 b15zdnd00an1n01x5 FILLER_379_2283 ();
 b15zdnd11an1n64x5 FILLER_380_8 ();
 b15zdnd11an1n64x5 FILLER_380_72 ();
 b15zdnd11an1n64x5 FILLER_380_136 ();
 b15zdnd11an1n64x5 FILLER_380_200 ();
 b15zdnd11an1n64x5 FILLER_380_264 ();
 b15zdnd11an1n32x5 FILLER_380_328 ();
 b15zdnd11an1n04x5 FILLER_380_360 ();
 b15zdnd11an1n64x5 FILLER_380_384 ();
 b15zdnd11an1n64x5 FILLER_380_448 ();
 b15zdnd11an1n64x5 FILLER_380_512 ();
 b15zdnd11an1n16x5 FILLER_380_576 ();
 b15zdnd11an1n08x5 FILLER_380_592 ();
 b15zdnd11an1n04x5 FILLER_380_600 ();
 b15zdnd11an1n64x5 FILLER_380_607 ();
 b15zdnd11an1n32x5 FILLER_380_671 ();
 b15zdnd11an1n08x5 FILLER_380_703 ();
 b15zdnd11an1n04x5 FILLER_380_711 ();
 b15zdnd00an1n02x5 FILLER_380_715 ();
 b15zdnd00an1n01x5 FILLER_380_717 ();
 b15zdnd11an1n64x5 FILLER_380_726 ();
 b15zdnd11an1n64x5 FILLER_380_790 ();
 b15zdnd11an1n08x5 FILLER_380_854 ();
 b15zdnd11an1n04x5 FILLER_380_862 ();
 b15zdnd00an1n02x5 FILLER_380_866 ();
 b15zdnd00an1n01x5 FILLER_380_868 ();
 b15zdnd11an1n64x5 FILLER_380_874 ();
 b15zdnd00an1n02x5 FILLER_380_938 ();
 b15zdnd00an1n01x5 FILLER_380_940 ();
 b15zdnd11an1n16x5 FILLER_380_946 ();
 b15zdnd00an1n02x5 FILLER_380_962 ();
 b15zdnd00an1n01x5 FILLER_380_964 ();
 b15zdnd11an1n64x5 FILLER_380_972 ();
 b15zdnd11an1n08x5 FILLER_380_1036 ();
 b15zdnd11an1n04x5 FILLER_380_1044 ();
 b15zdnd00an1n01x5 FILLER_380_1048 ();
 b15zdnd11an1n08x5 FILLER_380_1054 ();
 b15zdnd11an1n16x5 FILLER_380_1104 ();
 b15zdnd11an1n08x5 FILLER_380_1120 ();
 b15zdnd11an1n04x5 FILLER_380_1128 ();
 b15zdnd11an1n04x5 FILLER_380_1137 ();
 b15zdnd11an1n08x5 FILLER_380_1146 ();
 b15zdnd00an1n01x5 FILLER_380_1154 ();
 b15zdnd11an1n16x5 FILLER_380_1162 ();
 b15zdnd00an1n01x5 FILLER_380_1178 ();
 b15zdnd11an1n08x5 FILLER_380_1189 ();
 b15zdnd00an1n02x5 FILLER_380_1197 ();
 b15zdnd00an1n01x5 FILLER_380_1199 ();
 b15zdnd11an1n04x5 FILLER_380_1205 ();
 b15zdnd11an1n16x5 FILLER_380_1219 ();
 b15zdnd00an1n02x5 FILLER_380_1235 ();
 b15zdnd11an1n04x5 FILLER_380_1242 ();
 b15zdnd00an1n02x5 FILLER_380_1246 ();
 b15zdnd00an1n01x5 FILLER_380_1248 ();
 b15zdnd11an1n04x5 FILLER_380_1256 ();
 b15zdnd11an1n64x5 FILLER_380_1265 ();
 b15zdnd11an1n64x5 FILLER_380_1329 ();
 b15zdnd11an1n64x5 FILLER_380_1393 ();
 b15zdnd11an1n64x5 FILLER_380_1457 ();
 b15zdnd11an1n64x5 FILLER_380_1521 ();
 b15zdnd11an1n64x5 FILLER_380_1585 ();
 b15zdnd11an1n64x5 FILLER_380_1649 ();
 b15zdnd11an1n64x5 FILLER_380_1713 ();
 b15zdnd11an1n64x5 FILLER_380_1777 ();
 b15zdnd11an1n64x5 FILLER_380_1841 ();
 b15zdnd11an1n64x5 FILLER_380_1905 ();
 b15zdnd11an1n64x5 FILLER_380_1969 ();
 b15zdnd11an1n64x5 FILLER_380_2033 ();
 b15zdnd11an1n32x5 FILLER_380_2097 ();
 b15zdnd11an1n16x5 FILLER_380_2129 ();
 b15zdnd11an1n08x5 FILLER_380_2145 ();
 b15zdnd00an1n01x5 FILLER_380_2153 ();
 b15zdnd11an1n64x5 FILLER_380_2162 ();
 b15zdnd11an1n32x5 FILLER_380_2226 ();
 b15zdnd11an1n16x5 FILLER_380_2258 ();
 b15zdnd00an1n02x5 FILLER_380_2274 ();
 b15zdnd11an1n64x5 FILLER_381_0 ();
 b15zdnd11an1n64x5 FILLER_381_64 ();
 b15zdnd11an1n64x5 FILLER_381_128 ();
 b15zdnd11an1n64x5 FILLER_381_192 ();
 b15zdnd11an1n64x5 FILLER_381_256 ();
 b15zdnd11an1n32x5 FILLER_381_320 ();
 b15zdnd11an1n08x5 FILLER_381_352 ();
 b15zdnd11an1n04x5 FILLER_381_360 ();
 b15zdnd11an1n64x5 FILLER_381_376 ();
 b15zdnd11an1n64x5 FILLER_381_440 ();
 b15zdnd11an1n16x5 FILLER_381_504 ();
 b15zdnd11an1n08x5 FILLER_381_520 ();
 b15zdnd00an1n01x5 FILLER_381_528 ();
 b15zdnd11an1n64x5 FILLER_381_533 ();
 b15zdnd11an1n04x5 FILLER_381_597 ();
 b15zdnd00an1n01x5 FILLER_381_601 ();
 b15zdnd11an1n64x5 FILLER_381_644 ();
 b15zdnd11an1n08x5 FILLER_381_708 ();
 b15zdnd00an1n01x5 FILLER_381_716 ();
 b15zdnd11an1n32x5 FILLER_381_759 ();
 b15zdnd11an1n04x5 FILLER_381_791 ();
 b15zdnd11an1n04x5 FILLER_381_805 ();
 b15zdnd11an1n64x5 FILLER_381_816 ();
 b15zdnd11an1n32x5 FILLER_381_880 ();
 b15zdnd11an1n04x5 FILLER_381_912 ();
 b15zdnd00an1n01x5 FILLER_381_916 ();
 b15zdnd11an1n08x5 FILLER_381_924 ();
 b15zdnd00an1n02x5 FILLER_381_932 ();
 b15zdnd00an1n01x5 FILLER_381_934 ();
 b15zdnd11an1n16x5 FILLER_381_942 ();
 b15zdnd11an1n04x5 FILLER_381_958 ();
 b15zdnd11an1n64x5 FILLER_381_969 ();
 b15zdnd11an1n04x5 FILLER_381_1033 ();
 b15zdnd00an1n01x5 FILLER_381_1037 ();
 b15zdnd11an1n04x5 FILLER_381_1046 ();
 b15zdnd00an1n02x5 FILLER_381_1050 ();
 b15zdnd11an1n04x5 FILLER_381_1057 ();
 b15zdnd11an1n04x5 FILLER_381_1068 ();
 b15zdnd11an1n04x5 FILLER_381_1079 ();
 b15zdnd00an1n02x5 FILLER_381_1083 ();
 b15zdnd11an1n16x5 FILLER_381_1096 ();
 b15zdnd11an1n04x5 FILLER_381_1112 ();
 b15zdnd00an1n02x5 FILLER_381_1116 ();
 b15zdnd11an1n16x5 FILLER_381_1125 ();
 b15zdnd11an1n04x5 FILLER_381_1141 ();
 b15zdnd00an1n02x5 FILLER_381_1145 ();
 b15zdnd00an1n01x5 FILLER_381_1147 ();
 b15zdnd11an1n08x5 FILLER_381_1153 ();
 b15zdnd00an1n02x5 FILLER_381_1161 ();
 b15zdnd00an1n01x5 FILLER_381_1163 ();
 b15zdnd11an1n16x5 FILLER_381_1169 ();
 b15zdnd11an1n08x5 FILLER_381_1185 ();
 b15zdnd11an1n04x5 FILLER_381_1193 ();
 b15zdnd11an1n16x5 FILLER_381_1204 ();
 b15zdnd00an1n02x5 FILLER_381_1220 ();
 b15zdnd11an1n04x5 FILLER_381_1232 ();
 b15zdnd11an1n08x5 FILLER_381_1243 ();
 b15zdnd11an1n04x5 FILLER_381_1256 ();
 b15zdnd11an1n64x5 FILLER_381_1267 ();
 b15zdnd11an1n64x5 FILLER_381_1331 ();
 b15zdnd11an1n64x5 FILLER_381_1395 ();
 b15zdnd11an1n64x5 FILLER_381_1459 ();
 b15zdnd11an1n64x5 FILLER_381_1523 ();
 b15zdnd11an1n64x5 FILLER_381_1587 ();
 b15zdnd11an1n64x5 FILLER_381_1651 ();
 b15zdnd11an1n64x5 FILLER_381_1715 ();
 b15zdnd11an1n64x5 FILLER_381_1779 ();
 b15zdnd11an1n64x5 FILLER_381_1843 ();
 b15zdnd11an1n64x5 FILLER_381_1907 ();
 b15zdnd11an1n64x5 FILLER_381_1971 ();
 b15zdnd11an1n64x5 FILLER_381_2035 ();
 b15zdnd11an1n64x5 FILLER_381_2099 ();
 b15zdnd11an1n64x5 FILLER_381_2163 ();
 b15zdnd11an1n32x5 FILLER_381_2227 ();
 b15zdnd11an1n16x5 FILLER_381_2259 ();
 b15zdnd11an1n08x5 FILLER_381_2275 ();
 b15zdnd00an1n01x5 FILLER_381_2283 ();
 b15zdnd11an1n64x5 FILLER_382_8 ();
 b15zdnd11an1n64x5 FILLER_382_72 ();
 b15zdnd11an1n64x5 FILLER_382_136 ();
 b15zdnd11an1n64x5 FILLER_382_200 ();
 b15zdnd11an1n64x5 FILLER_382_264 ();
 b15zdnd11an1n16x5 FILLER_382_328 ();
 b15zdnd11an1n08x5 FILLER_382_344 ();
 b15zdnd11an1n04x5 FILLER_382_352 ();
 b15zdnd00an1n01x5 FILLER_382_356 ();
 b15zdnd11an1n16x5 FILLER_382_361 ();
 b15zdnd00an1n02x5 FILLER_382_377 ();
 b15zdnd11an1n64x5 FILLER_382_387 ();
 b15zdnd11an1n64x5 FILLER_382_451 ();
 b15zdnd11an1n16x5 FILLER_382_515 ();
 b15zdnd11an1n32x5 FILLER_382_537 ();
 b15zdnd00an1n01x5 FILLER_382_569 ();
 b15zdnd11an1n04x5 FILLER_382_612 ();
 b15zdnd11an1n32x5 FILLER_382_658 ();
 b15zdnd11an1n16x5 FILLER_382_690 ();
 b15zdnd11an1n08x5 FILLER_382_706 ();
 b15zdnd11an1n04x5 FILLER_382_714 ();
 b15zdnd11an1n08x5 FILLER_382_726 ();
 b15zdnd00an1n01x5 FILLER_382_734 ();
 b15zdnd11an1n64x5 FILLER_382_741 ();
 b15zdnd11an1n64x5 FILLER_382_805 ();
 b15zdnd11an1n64x5 FILLER_382_869 ();
 b15zdnd11an1n64x5 FILLER_382_933 ();
 b15zdnd11an1n64x5 FILLER_382_997 ();
 b15zdnd11an1n64x5 FILLER_382_1061 ();
 b15zdnd11an1n64x5 FILLER_382_1125 ();
 b15zdnd11an1n64x5 FILLER_382_1189 ();
 b15zdnd11an1n64x5 FILLER_382_1253 ();
 b15zdnd11an1n64x5 FILLER_382_1317 ();
 b15zdnd11an1n64x5 FILLER_382_1381 ();
 b15zdnd11an1n64x5 FILLER_382_1445 ();
 b15zdnd11an1n64x5 FILLER_382_1509 ();
 b15zdnd11an1n64x5 FILLER_382_1573 ();
 b15zdnd11an1n64x5 FILLER_382_1637 ();
 b15zdnd11an1n64x5 FILLER_382_1701 ();
 b15zdnd11an1n64x5 FILLER_382_1765 ();
 b15zdnd11an1n64x5 FILLER_382_1829 ();
 b15zdnd11an1n64x5 FILLER_382_1893 ();
 b15zdnd11an1n64x5 FILLER_382_1957 ();
 b15zdnd11an1n64x5 FILLER_382_2021 ();
 b15zdnd11an1n64x5 FILLER_382_2085 ();
 b15zdnd11an1n04x5 FILLER_382_2149 ();
 b15zdnd00an1n01x5 FILLER_382_2153 ();
 b15zdnd11an1n64x5 FILLER_382_2162 ();
 b15zdnd11an1n32x5 FILLER_382_2226 ();
 b15zdnd11an1n16x5 FILLER_382_2258 ();
 b15zdnd00an1n02x5 FILLER_382_2274 ();
 b15zdnd11an1n64x5 FILLER_383_0 ();
 b15zdnd11an1n64x5 FILLER_383_64 ();
 b15zdnd11an1n64x5 FILLER_383_128 ();
 b15zdnd11an1n64x5 FILLER_383_192 ();
 b15zdnd11an1n64x5 FILLER_383_256 ();
 b15zdnd11an1n32x5 FILLER_383_320 ();
 b15zdnd11an1n08x5 FILLER_383_352 ();
 b15zdnd11an1n04x5 FILLER_383_360 ();
 b15zdnd00an1n02x5 FILLER_383_364 ();
 b15zdnd00an1n01x5 FILLER_383_366 ();
 b15zdnd11an1n04x5 FILLER_383_373 ();
 b15zdnd11an1n64x5 FILLER_383_383 ();
 b15zdnd11an1n64x5 FILLER_383_447 ();
 b15zdnd11an1n32x5 FILLER_383_511 ();
 b15zdnd11an1n08x5 FILLER_383_543 ();
 b15zdnd11an1n04x5 FILLER_383_551 ();
 b15zdnd00an1n01x5 FILLER_383_555 ();
 b15zdnd11an1n04x5 FILLER_383_598 ();
 b15zdnd11an1n32x5 FILLER_383_644 ();
 b15zdnd11an1n16x5 FILLER_383_676 ();
 b15zdnd11an1n08x5 FILLER_383_692 ();
 b15zdnd00an1n01x5 FILLER_383_700 ();
 b15zdnd11an1n64x5 FILLER_383_743 ();
 b15zdnd11an1n32x5 FILLER_383_807 ();
 b15zdnd00an1n02x5 FILLER_383_839 ();
 b15zdnd00an1n01x5 FILLER_383_841 ();
 b15zdnd11an1n04x5 FILLER_383_884 ();
 b15zdnd00an1n02x5 FILLER_383_888 ();
 b15zdnd11an1n64x5 FILLER_383_932 ();
 b15zdnd11an1n64x5 FILLER_383_996 ();
 b15zdnd11an1n64x5 FILLER_383_1060 ();
 b15zdnd11an1n64x5 FILLER_383_1124 ();
 b15zdnd11an1n64x5 FILLER_383_1188 ();
 b15zdnd11an1n64x5 FILLER_383_1252 ();
 b15zdnd11an1n64x5 FILLER_383_1316 ();
 b15zdnd11an1n64x5 FILLER_383_1380 ();
 b15zdnd11an1n64x5 FILLER_383_1444 ();
 b15zdnd11an1n64x5 FILLER_383_1508 ();
 b15zdnd11an1n64x5 FILLER_383_1572 ();
 b15zdnd11an1n64x5 FILLER_383_1636 ();
 b15zdnd11an1n64x5 FILLER_383_1700 ();
 b15zdnd11an1n64x5 FILLER_383_1764 ();
 b15zdnd11an1n64x5 FILLER_383_1828 ();
 b15zdnd11an1n64x5 FILLER_383_1892 ();
 b15zdnd11an1n64x5 FILLER_383_1956 ();
 b15zdnd11an1n64x5 FILLER_383_2020 ();
 b15zdnd11an1n64x5 FILLER_383_2084 ();
 b15zdnd11an1n64x5 FILLER_383_2148 ();
 b15zdnd11an1n64x5 FILLER_383_2212 ();
 b15zdnd11an1n08x5 FILLER_383_2276 ();
 b15zdnd11an1n64x5 FILLER_384_8 ();
 b15zdnd11an1n64x5 FILLER_384_72 ();
 b15zdnd11an1n64x5 FILLER_384_136 ();
 b15zdnd11an1n64x5 FILLER_384_200 ();
 b15zdnd11an1n64x5 FILLER_384_264 ();
 b15zdnd11an1n64x5 FILLER_384_328 ();
 b15zdnd11an1n64x5 FILLER_384_392 ();
 b15zdnd11an1n64x5 FILLER_384_456 ();
 b15zdnd11an1n64x5 FILLER_384_520 ();
 b15zdnd00an1n01x5 FILLER_384_584 ();
 b15zdnd11an1n04x5 FILLER_384_627 ();
 b15zdnd11an1n64x5 FILLER_384_635 ();
 b15zdnd11an1n16x5 FILLER_384_699 ();
 b15zdnd00an1n02x5 FILLER_384_715 ();
 b15zdnd00an1n01x5 FILLER_384_717 ();
 b15zdnd00an1n02x5 FILLER_384_726 ();
 b15zdnd11an1n32x5 FILLER_384_770 ();
 b15zdnd11an1n08x5 FILLER_384_802 ();
 b15zdnd11an1n04x5 FILLER_384_810 ();
 b15zdnd11an1n04x5 FILLER_384_856 ();
 b15zdnd00an1n02x5 FILLER_384_860 ();
 b15zdnd00an1n01x5 FILLER_384_862 ();
 b15zdnd11an1n04x5 FILLER_384_905 ();
 b15zdnd11an1n64x5 FILLER_384_951 ();
 b15zdnd11an1n64x5 FILLER_384_1015 ();
 b15zdnd11an1n64x5 FILLER_384_1079 ();
 b15zdnd11an1n64x5 FILLER_384_1143 ();
 b15zdnd11an1n64x5 FILLER_384_1207 ();
 b15zdnd11an1n64x5 FILLER_384_1271 ();
 b15zdnd11an1n64x5 FILLER_384_1335 ();
 b15zdnd11an1n64x5 FILLER_384_1399 ();
 b15zdnd11an1n64x5 FILLER_384_1463 ();
 b15zdnd11an1n64x5 FILLER_384_1527 ();
 b15zdnd11an1n64x5 FILLER_384_1591 ();
 b15zdnd11an1n64x5 FILLER_384_1655 ();
 b15zdnd11an1n64x5 FILLER_384_1719 ();
 b15zdnd11an1n64x5 FILLER_384_1783 ();
 b15zdnd11an1n64x5 FILLER_384_1847 ();
 b15zdnd11an1n64x5 FILLER_384_1911 ();
 b15zdnd11an1n64x5 FILLER_384_1975 ();
 b15zdnd11an1n64x5 FILLER_384_2039 ();
 b15zdnd11an1n32x5 FILLER_384_2103 ();
 b15zdnd11an1n16x5 FILLER_384_2135 ();
 b15zdnd00an1n02x5 FILLER_384_2151 ();
 b15zdnd00an1n01x5 FILLER_384_2153 ();
 b15zdnd11an1n64x5 FILLER_384_2162 ();
 b15zdnd11an1n32x5 FILLER_384_2226 ();
 b15zdnd11an1n16x5 FILLER_384_2258 ();
 b15zdnd00an1n02x5 FILLER_384_2274 ();
 b15zdnd11an1n64x5 FILLER_385_0 ();
 b15zdnd11an1n64x5 FILLER_385_64 ();
 b15zdnd11an1n64x5 FILLER_385_128 ();
 b15zdnd11an1n64x5 FILLER_385_192 ();
 b15zdnd11an1n64x5 FILLER_385_256 ();
 b15zdnd11an1n32x5 FILLER_385_320 ();
 b15zdnd11an1n16x5 FILLER_385_352 ();
 b15zdnd00an1n01x5 FILLER_385_368 ();
 b15zdnd11an1n64x5 FILLER_385_373 ();
 b15zdnd11an1n64x5 FILLER_385_437 ();
 b15zdnd11an1n16x5 FILLER_385_501 ();
 b15zdnd11an1n08x5 FILLER_385_517 ();
 b15zdnd11an1n04x5 FILLER_385_525 ();
 b15zdnd00an1n02x5 FILLER_385_529 ();
 b15zdnd00an1n01x5 FILLER_385_531 ();
 b15zdnd11an1n04x5 FILLER_385_574 ();
 b15zdnd00an1n02x5 FILLER_385_578 ();
 b15zdnd00an1n01x5 FILLER_385_580 ();
 b15zdnd11an1n08x5 FILLER_385_623 ();
 b15zdnd00an1n01x5 FILLER_385_631 ();
 b15zdnd11an1n04x5 FILLER_385_638 ();
 b15zdnd11an1n64x5 FILLER_385_648 ();
 b15zdnd11an1n16x5 FILLER_385_712 ();
 b15zdnd11an1n08x5 FILLER_385_728 ();
 b15zdnd00an1n02x5 FILLER_385_736 ();
 b15zdnd00an1n01x5 FILLER_385_738 ();
 b15zdnd11an1n32x5 FILLER_385_781 ();
 b15zdnd00an1n02x5 FILLER_385_813 ();
 b15zdnd11an1n16x5 FILLER_385_857 ();
 b15zdnd11an1n04x5 FILLER_385_873 ();
 b15zdnd11an1n04x5 FILLER_385_919 ();
 b15zdnd11an1n16x5 FILLER_385_965 ();
 b15zdnd00an1n02x5 FILLER_385_981 ();
 b15zdnd11an1n64x5 FILLER_385_1025 ();
 b15zdnd11an1n64x5 FILLER_385_1089 ();
 b15zdnd11an1n16x5 FILLER_385_1195 ();
 b15zdnd00an1n01x5 FILLER_385_1211 ();
 b15zdnd11an1n64x5 FILLER_385_1254 ();
 b15zdnd11an1n64x5 FILLER_385_1318 ();
 b15zdnd11an1n64x5 FILLER_385_1382 ();
 b15zdnd11an1n64x5 FILLER_385_1446 ();
 b15zdnd11an1n64x5 FILLER_385_1510 ();
 b15zdnd11an1n64x5 FILLER_385_1574 ();
 b15zdnd11an1n64x5 FILLER_385_1638 ();
 b15zdnd11an1n64x5 FILLER_385_1702 ();
 b15zdnd11an1n64x5 FILLER_385_1766 ();
 b15zdnd11an1n64x5 FILLER_385_1830 ();
 b15zdnd11an1n64x5 FILLER_385_1894 ();
 b15zdnd11an1n64x5 FILLER_385_1958 ();
 b15zdnd11an1n64x5 FILLER_385_2022 ();
 b15zdnd11an1n64x5 FILLER_385_2086 ();
 b15zdnd11an1n64x5 FILLER_385_2150 ();
 b15zdnd11an1n64x5 FILLER_385_2214 ();
 b15zdnd11an1n04x5 FILLER_385_2278 ();
 b15zdnd00an1n02x5 FILLER_385_2282 ();
 b15zdnd11an1n64x5 FILLER_386_8 ();
 b15zdnd11an1n64x5 FILLER_386_72 ();
 b15zdnd11an1n64x5 FILLER_386_136 ();
 b15zdnd11an1n64x5 FILLER_386_200 ();
 b15zdnd11an1n64x5 FILLER_386_264 ();
 b15zdnd11an1n32x5 FILLER_386_328 ();
 b15zdnd00an1n01x5 FILLER_386_360 ();
 b15zdnd11an1n04x5 FILLER_386_365 ();
 b15zdnd11an1n04x5 FILLER_386_373 ();
 b15zdnd11an1n64x5 FILLER_386_381 ();
 b15zdnd11an1n64x5 FILLER_386_445 ();
 b15zdnd11an1n16x5 FILLER_386_509 ();
 b15zdnd11an1n08x5 FILLER_386_525 ();
 b15zdnd11an1n04x5 FILLER_386_533 ();
 b15zdnd00an1n02x5 FILLER_386_537 ();
 b15zdnd11an1n08x5 FILLER_386_581 ();
 b15zdnd00an1n01x5 FILLER_386_589 ();
 b15zdnd11an1n04x5 FILLER_386_594 ();
 b15zdnd11an1n04x5 FILLER_386_640 ();
 b15zdnd11an1n08x5 FILLER_386_650 ();
 b15zdnd00an1n02x5 FILLER_386_658 ();
 b15zdnd00an1n01x5 FILLER_386_660 ();
 b15zdnd11an1n04x5 FILLER_386_665 ();
 b15zdnd11an1n04x5 FILLER_386_673 ();
 b15zdnd11an1n32x5 FILLER_386_681 ();
 b15zdnd11an1n04x5 FILLER_386_713 ();
 b15zdnd00an1n01x5 FILLER_386_717 ();
 b15zdnd11an1n16x5 FILLER_386_726 ();
 b15zdnd11an1n64x5 FILLER_386_784 ();
 b15zdnd11an1n64x5 FILLER_386_848 ();
 b15zdnd11an1n64x5 FILLER_386_912 ();
 b15zdnd11an1n64x5 FILLER_386_976 ();
 b15zdnd11an1n64x5 FILLER_386_1040 ();
 b15zdnd11an1n64x5 FILLER_386_1104 ();
 b15zdnd11an1n64x5 FILLER_386_1168 ();
 b15zdnd11an1n64x5 FILLER_386_1232 ();
 b15zdnd11an1n64x5 FILLER_386_1296 ();
 b15zdnd11an1n64x5 FILLER_386_1360 ();
 b15zdnd11an1n64x5 FILLER_386_1424 ();
 b15zdnd11an1n64x5 FILLER_386_1488 ();
 b15zdnd11an1n64x5 FILLER_386_1552 ();
 b15zdnd11an1n64x5 FILLER_386_1616 ();
 b15zdnd11an1n64x5 FILLER_386_1680 ();
 b15zdnd11an1n64x5 FILLER_386_1744 ();
 b15zdnd11an1n64x5 FILLER_386_1808 ();
 b15zdnd11an1n64x5 FILLER_386_1872 ();
 b15zdnd11an1n64x5 FILLER_386_1936 ();
 b15zdnd11an1n64x5 FILLER_386_2000 ();
 b15zdnd11an1n64x5 FILLER_386_2064 ();
 b15zdnd11an1n16x5 FILLER_386_2128 ();
 b15zdnd11an1n08x5 FILLER_386_2144 ();
 b15zdnd00an1n02x5 FILLER_386_2152 ();
 b15zdnd11an1n64x5 FILLER_386_2162 ();
 b15zdnd11an1n32x5 FILLER_386_2226 ();
 b15zdnd11an1n16x5 FILLER_386_2258 ();
 b15zdnd00an1n02x5 FILLER_386_2274 ();
 b15zdnd11an1n64x5 FILLER_387_0 ();
 b15zdnd11an1n64x5 FILLER_387_64 ();
 b15zdnd11an1n64x5 FILLER_387_128 ();
 b15zdnd11an1n64x5 FILLER_387_192 ();
 b15zdnd11an1n64x5 FILLER_387_256 ();
 b15zdnd11an1n32x5 FILLER_387_320 ();
 b15zdnd11an1n08x5 FILLER_387_352 ();
 b15zdnd00an1n01x5 FILLER_387_360 ();
 b15zdnd11an1n04x5 FILLER_387_365 ();
 b15zdnd11an1n04x5 FILLER_387_373 ();
 b15zdnd00an1n02x5 FILLER_387_377 ();
 b15zdnd00an1n01x5 FILLER_387_379 ();
 b15zdnd11an1n64x5 FILLER_387_384 ();
 b15zdnd11an1n64x5 FILLER_387_448 ();
 b15zdnd11an1n16x5 FILLER_387_512 ();
 b15zdnd11an1n08x5 FILLER_387_528 ();
 b15zdnd00an1n02x5 FILLER_387_536 ();
 b15zdnd00an1n01x5 FILLER_387_538 ();
 b15zdnd11an1n04x5 FILLER_387_581 ();
 b15zdnd00an1n02x5 FILLER_387_585 ();
 b15zdnd11an1n04x5 FILLER_387_591 ();
 b15zdnd11an1n04x5 FILLER_387_599 ();
 b15zdnd11an1n04x5 FILLER_387_607 ();
 b15zdnd11an1n08x5 FILLER_387_653 ();
 b15zdnd00an1n02x5 FILLER_387_661 ();
 b15zdnd00an1n01x5 FILLER_387_663 ();
 b15zdnd11an1n16x5 FILLER_387_706 ();
 b15zdnd11an1n08x5 FILLER_387_722 ();
 b15zdnd11an1n04x5 FILLER_387_730 ();
 b15zdnd00an1n01x5 FILLER_387_734 ();
 b15zdnd11an1n04x5 FILLER_387_739 ();
 b15zdnd11an1n04x5 FILLER_387_785 ();
 b15zdnd11an1n04x5 FILLER_387_795 ();
 b15zdnd11an1n08x5 FILLER_387_803 ();
 b15zdnd00an1n02x5 FILLER_387_811 ();
 b15zdnd00an1n01x5 FILLER_387_813 ();
 b15zdnd11an1n64x5 FILLER_387_818 ();
 b15zdnd11an1n64x5 FILLER_387_882 ();
 b15zdnd11an1n64x5 FILLER_387_946 ();
 b15zdnd11an1n64x5 FILLER_387_1010 ();
 b15zdnd11an1n64x5 FILLER_387_1074 ();
 b15zdnd11an1n64x5 FILLER_387_1138 ();
 b15zdnd11an1n32x5 FILLER_387_1202 ();
 b15zdnd11an1n16x5 FILLER_387_1234 ();
 b15zdnd11an1n08x5 FILLER_387_1250 ();
 b15zdnd00an1n02x5 FILLER_387_1258 ();
 b15zdnd00an1n01x5 FILLER_387_1260 ();
 b15zdnd11an1n64x5 FILLER_387_1265 ();
 b15zdnd11an1n64x5 FILLER_387_1329 ();
 b15zdnd11an1n64x5 FILLER_387_1393 ();
 b15zdnd11an1n64x5 FILLER_387_1457 ();
 b15zdnd11an1n64x5 FILLER_387_1521 ();
 b15zdnd11an1n64x5 FILLER_387_1585 ();
 b15zdnd11an1n64x5 FILLER_387_1649 ();
 b15zdnd11an1n64x5 FILLER_387_1713 ();
 b15zdnd11an1n64x5 FILLER_387_1777 ();
 b15zdnd11an1n64x5 FILLER_387_1841 ();
 b15zdnd11an1n64x5 FILLER_387_1905 ();
 b15zdnd11an1n64x5 FILLER_387_1969 ();
 b15zdnd11an1n64x5 FILLER_387_2033 ();
 b15zdnd11an1n64x5 FILLER_387_2097 ();
 b15zdnd11an1n64x5 FILLER_387_2161 ();
 b15zdnd11an1n32x5 FILLER_387_2225 ();
 b15zdnd11an1n16x5 FILLER_387_2257 ();
 b15zdnd11an1n08x5 FILLER_387_2273 ();
 b15zdnd00an1n02x5 FILLER_387_2281 ();
 b15zdnd00an1n01x5 FILLER_387_2283 ();
 b15zdnd11an1n64x5 FILLER_388_8 ();
 b15zdnd11an1n64x5 FILLER_388_72 ();
 b15zdnd11an1n64x5 FILLER_388_136 ();
 b15zdnd11an1n64x5 FILLER_388_200 ();
 b15zdnd11an1n64x5 FILLER_388_264 ();
 b15zdnd11an1n16x5 FILLER_388_328 ();
 b15zdnd11an1n08x5 FILLER_388_344 ();
 b15zdnd11an1n04x5 FILLER_388_352 ();
 b15zdnd00an1n02x5 FILLER_388_356 ();
 b15zdnd00an1n01x5 FILLER_388_358 ();
 b15zdnd11an1n04x5 FILLER_388_364 ();
 b15zdnd11an1n04x5 FILLER_388_372 ();
 b15zdnd11an1n04x5 FILLER_388_380 ();
 b15zdnd11an1n16x5 FILLER_388_388 ();
 b15zdnd00an1n01x5 FILLER_388_404 ();
 b15zdnd11an1n64x5 FILLER_388_410 ();
 b15zdnd11an1n16x5 FILLER_388_474 ();
 b15zdnd00an1n02x5 FILLER_388_490 ();
 b15zdnd11an1n32x5 FILLER_388_496 ();
 b15zdnd11an1n04x5 FILLER_388_528 ();
 b15zdnd11an1n16x5 FILLER_388_536 ();
 b15zdnd00an1n02x5 FILLER_388_552 ();
 b15zdnd00an1n01x5 FILLER_388_554 ();
 b15zdnd11an1n04x5 FILLER_388_559 ();
 b15zdnd11an1n04x5 FILLER_388_567 ();
 b15zdnd11an1n04x5 FILLER_388_613 ();
 b15zdnd11an1n04x5 FILLER_388_659 ();
 b15zdnd00an1n02x5 FILLER_388_663 ();
 b15zdnd00an1n01x5 FILLER_388_665 ();
 b15zdnd11an1n04x5 FILLER_388_708 ();
 b15zdnd00an1n02x5 FILLER_388_716 ();
 b15zdnd11an1n08x5 FILLER_388_726 ();
 b15zdnd00an1n02x5 FILLER_388_734 ();
 b15zdnd11an1n04x5 FILLER_388_740 ();
 b15zdnd11an1n04x5 FILLER_388_748 ();
 b15zdnd11an1n04x5 FILLER_388_757 ();
 b15zdnd11an1n04x5 FILLER_388_767 ();
 b15zdnd11an1n08x5 FILLER_388_813 ();
 b15zdnd00an1n02x5 FILLER_388_821 ();
 b15zdnd11an1n04x5 FILLER_388_827 ();
 b15zdnd11an1n16x5 FILLER_388_835 ();
 b15zdnd11an1n08x5 FILLER_388_851 ();
 b15zdnd11an1n04x5 FILLER_388_859 ();
 b15zdnd11an1n04x5 FILLER_388_867 ();
 b15zdnd11an1n64x5 FILLER_388_875 ();
 b15zdnd11an1n04x5 FILLER_388_939 ();
 b15zdnd00an1n01x5 FILLER_388_943 ();
 b15zdnd11an1n32x5 FILLER_388_948 ();
 b15zdnd11an1n16x5 FILLER_388_980 ();
 b15zdnd11an1n16x5 FILLER_388_1000 ();
 b15zdnd11an1n08x5 FILLER_388_1016 ();
 b15zdnd00an1n02x5 FILLER_388_1024 ();
 b15zdnd00an1n01x5 FILLER_388_1026 ();
 b15zdnd11an1n16x5 FILLER_388_1031 ();
 b15zdnd11an1n64x5 FILLER_388_1051 ();
 b15zdnd11an1n16x5 FILLER_388_1115 ();
 b15zdnd11an1n08x5 FILLER_388_1131 ();
 b15zdnd11an1n04x5 FILLER_388_1139 ();
 b15zdnd00an1n02x5 FILLER_388_1143 ();
 b15zdnd00an1n01x5 FILLER_388_1145 ();
 b15zdnd11an1n16x5 FILLER_388_1150 ();
 b15zdnd00an1n02x5 FILLER_388_1166 ();
 b15zdnd11an1n64x5 FILLER_388_1172 ();
 b15zdnd11an1n04x5 FILLER_388_1236 ();
 b15zdnd00an1n02x5 FILLER_388_1240 ();
 b15zdnd00an1n01x5 FILLER_388_1242 ();
 b15zdnd11an1n08x5 FILLER_388_1247 ();
 b15zdnd00an1n01x5 FILLER_388_1255 ();
 b15zdnd11an1n04x5 FILLER_388_1260 ();
 b15zdnd11an1n04x5 FILLER_388_1268 ();
 b15zdnd11an1n64x5 FILLER_388_1276 ();
 b15zdnd11an1n64x5 FILLER_388_1340 ();
 b15zdnd11an1n64x5 FILLER_388_1404 ();
 b15zdnd11an1n64x5 FILLER_388_1468 ();
 b15zdnd11an1n64x5 FILLER_388_1532 ();
 b15zdnd11an1n64x5 FILLER_388_1596 ();
 b15zdnd11an1n64x5 FILLER_388_1660 ();
 b15zdnd11an1n64x5 FILLER_388_1724 ();
 b15zdnd11an1n64x5 FILLER_388_1788 ();
 b15zdnd11an1n64x5 FILLER_388_1852 ();
 b15zdnd11an1n64x5 FILLER_388_1916 ();
 b15zdnd11an1n64x5 FILLER_388_1980 ();
 b15zdnd11an1n64x5 FILLER_388_2044 ();
 b15zdnd11an1n32x5 FILLER_388_2108 ();
 b15zdnd11an1n08x5 FILLER_388_2140 ();
 b15zdnd11an1n04x5 FILLER_388_2148 ();
 b15zdnd00an1n02x5 FILLER_388_2152 ();
 b15zdnd11an1n64x5 FILLER_388_2162 ();
 b15zdnd11an1n32x5 FILLER_388_2226 ();
 b15zdnd11an1n16x5 FILLER_388_2258 ();
 b15zdnd00an1n02x5 FILLER_388_2274 ();
 b15zdnd11an1n64x5 FILLER_389_0 ();
 b15zdnd11an1n64x5 FILLER_389_64 ();
 b15zdnd11an1n64x5 FILLER_389_128 ();
 b15zdnd11an1n64x5 FILLER_389_192 ();
 b15zdnd11an1n64x5 FILLER_389_256 ();
 b15zdnd11an1n16x5 FILLER_389_320 ();
 b15zdnd11an1n04x5 FILLER_389_336 ();
 b15zdnd00an1n02x5 FILLER_389_340 ();
 b15zdnd11an1n08x5 FILLER_389_348 ();
 b15zdnd11an1n04x5 FILLER_389_360 ();
 b15zdnd00an1n01x5 FILLER_389_364 ();
 b15zdnd11an1n08x5 FILLER_389_369 ();
 b15zdnd00an1n01x5 FILLER_389_377 ();
 b15zdnd11an1n04x5 FILLER_389_382 ();
 b15zdnd11an1n64x5 FILLER_389_390 ();
 b15zdnd11an1n32x5 FILLER_389_454 ();
 b15zdnd11an1n04x5 FILLER_389_486 ();
 b15zdnd00an1n02x5 FILLER_389_490 ();
 b15zdnd00an1n01x5 FILLER_389_492 ();
 b15zdnd11an1n32x5 FILLER_389_501 ();
 b15zdnd11an1n04x5 FILLER_389_533 ();
 b15zdnd00an1n02x5 FILLER_389_537 ();
 b15zdnd00an1n01x5 FILLER_389_539 ();
 b15zdnd11an1n08x5 FILLER_389_544 ();
 b15zdnd11an1n04x5 FILLER_389_552 ();
 b15zdnd11an1n04x5 FILLER_389_560 ();
 b15zdnd11an1n04x5 FILLER_389_568 ();
 b15zdnd11an1n04x5 FILLER_389_614 ();
 b15zdnd11an1n04x5 FILLER_389_660 ();
 b15zdnd11an1n08x5 FILLER_389_670 ();
 b15zdnd11an1n04x5 FILLER_389_720 ();
 b15zdnd00an1n01x5 FILLER_389_724 ();
 b15zdnd11an1n04x5 FILLER_389_729 ();
 b15zdnd11an1n04x5 FILLER_389_737 ();
 b15zdnd11an1n04x5 FILLER_389_746 ();
 b15zdnd11an1n04x5 FILLER_389_792 ();
 b15zdnd11an1n04x5 FILLER_389_838 ();
 b15zdnd11an1n32x5 FILLER_389_846 ();
 b15zdnd11an1n08x5 FILLER_389_878 ();
 b15zdnd00an1n02x5 FILLER_389_886 ();
 b15zdnd11an1n08x5 FILLER_389_892 ();
 b15zdnd11an1n04x5 FILLER_389_904 ();
 b15zdnd11an1n08x5 FILLER_389_912 ();
 b15zdnd00an1n01x5 FILLER_389_920 ();
 b15zdnd11an1n16x5 FILLER_389_925 ();
 b15zdnd00an1n02x5 FILLER_389_941 ();
 b15zdnd11an1n08x5 FILLER_389_947 ();
 b15zdnd11an1n04x5 FILLER_389_955 ();
 b15zdnd00an1n01x5 FILLER_389_959 ();
 b15zdnd11an1n04x5 FILLER_389_964 ();
 b15zdnd11an1n32x5 FILLER_389_972 ();
 b15zdnd00an1n02x5 FILLER_389_1004 ();
 b15zdnd11an1n32x5 FILLER_389_1010 ();
 b15zdnd11an1n08x5 FILLER_389_1042 ();
 b15zdnd00an1n01x5 FILLER_389_1050 ();
 b15zdnd11an1n16x5 FILLER_389_1055 ();
 b15zdnd11an1n08x5 FILLER_389_1071 ();
 b15zdnd11an1n16x5 FILLER_389_1083 ();
 b15zdnd11an1n04x5 FILLER_389_1099 ();
 b15zdnd00an1n02x5 FILLER_389_1103 ();
 b15zdnd11an1n16x5 FILLER_389_1109 ();
 b15zdnd11an1n08x5 FILLER_389_1125 ();
 b15zdnd11an1n04x5 FILLER_389_1133 ();
 b15zdnd11an1n04x5 FILLER_389_1141 ();
 b15zdnd11an1n04x5 FILLER_389_1149 ();
 b15zdnd11an1n04x5 FILLER_389_1157 ();
 b15zdnd11an1n32x5 FILLER_389_1165 ();
 b15zdnd11an1n04x5 FILLER_389_1197 ();
 b15zdnd11an1n08x5 FILLER_389_1205 ();
 b15zdnd11an1n04x5 FILLER_389_1213 ();
 b15zdnd00an1n01x5 FILLER_389_1217 ();
 b15zdnd11an1n16x5 FILLER_389_1222 ();
 b15zdnd00an1n02x5 FILLER_389_1238 ();
 b15zdnd00an1n01x5 FILLER_389_1240 ();
 b15zdnd11an1n04x5 FILLER_389_1245 ();
 b15zdnd11an1n04x5 FILLER_389_1253 ();
 b15zdnd11an1n04x5 FILLER_389_1261 ();
 b15zdnd00an1n02x5 FILLER_389_1265 ();
 b15zdnd00an1n01x5 FILLER_389_1267 ();
 b15zdnd11an1n04x5 FILLER_389_1272 ();
 b15zdnd00an1n02x5 FILLER_389_1276 ();
 b15zdnd11an1n64x5 FILLER_389_1282 ();
 b15zdnd11an1n64x5 FILLER_389_1346 ();
 b15zdnd11an1n64x5 FILLER_389_1410 ();
 b15zdnd11an1n64x5 FILLER_389_1474 ();
 b15zdnd11an1n64x5 FILLER_389_1538 ();
 b15zdnd11an1n64x5 FILLER_389_1602 ();
 b15zdnd11an1n64x5 FILLER_389_1666 ();
 b15zdnd11an1n64x5 FILLER_389_1730 ();
 b15zdnd11an1n64x5 FILLER_389_1794 ();
 b15zdnd11an1n64x5 FILLER_389_1858 ();
 b15zdnd11an1n64x5 FILLER_389_1922 ();
 b15zdnd11an1n64x5 FILLER_389_1986 ();
 b15zdnd11an1n64x5 FILLER_389_2050 ();
 b15zdnd11an1n64x5 FILLER_389_2114 ();
 b15zdnd11an1n64x5 FILLER_389_2178 ();
 b15zdnd11an1n32x5 FILLER_389_2242 ();
 b15zdnd11an1n08x5 FILLER_389_2274 ();
 b15zdnd00an1n02x5 FILLER_389_2282 ();
endmodule
