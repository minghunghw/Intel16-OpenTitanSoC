module Noise_injection_block_Stuck (
    RANDOM,
    S,
    VB,
    IOUT
);

input RANDOM;
input [15:0] S;
input [3:0] VB;
output IOUT;

endmodule