module xbar_west (

);

endmodule