module b15ztpn00an1d03x5();
endmodule

module b15ztpn00an1n08x5();
endmodule

module b15zdnd00an1n01x5();
endmodule

module b15zdnd00an1n02x5();
endmodule

module b15zdnd11an1n04x5();
endmodule

module b15zdnd11an1n08x5();
endmodule

module b15zdnd11an1n16x5();
endmodule

module b15zdnd11an1n32x5();
endmodule

module b15zdnd11an1n64x5();
endmodule