module gpio (clk_i,
    rst_ni,
    alert_rx_i,
    alert_tx_o,
    cio_gpio_en_o,
    cio_gpio_i,
    cio_gpio_o,
    intr_gpio_o,
    tl_i,
    tl_o);
 input clk_i;
 input rst_ni;
 input [3:0] alert_rx_i;
 output [1:0] alert_tx_o;
 output [31:0] cio_gpio_en_o;
 input [31:0] cio_gpio_i;
 output [31:0] cio_gpio_o;
 output [31:0] intr_gpio_o;
 input [108:0] tl_i;
 output [65:0] tl_o;

 wire N113;
 wire N114;
 wire N115;
 wire N116;
 wire N117;
 wire N118;
 wire N119;
 wire N120;
 wire N121;
 wire N122;
 wire N123;
 wire N124;
 wire N125;
 wire N126;
 wire N127;
 wire N128;
 wire N129;
 wire N130;
 wire N131;
 wire N132;
 wire N133;
 wire N134;
 wire N135;
 wire N136;
 wire N137;
 wire N138;
 wire N139;
 wire N140;
 wire N141;
 wire N142;
 wire N143;
 wire N144;
 wire N145;
 wire N146;
 wire N38;
 wire N39;
 wire N40;
 wire N41;
 wire N42;
 wire N43;
 wire N44;
 wire N45;
 wire N46;
 wire N47;
 wire N48;
 wire N49;
 wire N50;
 wire N51;
 wire N52;
 wire N53;
 wire N54;
 wire N55;
 wire N56;
 wire N57;
 wire N58;
 wire N59;
 wire N60;
 wire N61;
 wire N62;
 wire N63;
 wire N64;
 wire N65;
 wire N66;
 wire N67;
 wire N68;
 wire N69;
 wire N70;
 wire N71;
 wire eq_x_101_n25;
 wire eq_x_106_n25;
 wire eq_x_111_n25;
 wire eq_x_116_n25;
 wire eq_x_121_n25;
 wire eq_x_126_n25;
 wire eq_x_131_n25;
 wire eq_x_136_n25;
 wire eq_x_141_n25;
 wire eq_x_146_n25;
 wire eq_x_151_n25;
 wire eq_x_156_n25;
 wire eq_x_161_n25;
 wire eq_x_166_n25;
 wire eq_x_171_n25;
 wire eq_x_176_n25;
 wire eq_x_181_n25;
 wire eq_x_26_n25;
 wire eq_x_31_n25;
 wire eq_x_36_n25;
 wire eq_x_41_n25;
 wire eq_x_46_n25;
 wire eq_x_51_n25;
 wire eq_x_56_n25;
 wire eq_x_61_n25;
 wire eq_x_66_n25;
 wire eq_x_71_n25;
 wire eq_x_76_n25;
 wire eq_x_81_n25;
 wire eq_x_86_n25;
 wire eq_x_91_n25;
 wire eq_x_96_n25;
 wire gen_alert_tx_0__u_prim_alert_sender_ack_level;
 wire gen_alert_tx_0__u_prim_alert_sender_alert_nd;
 wire gen_alert_tx_0__u_prim_alert_sender_alert_pd;
 wire gen_alert_tx_0__u_prim_alert_sender_alert_req_trigger;
 wire gen_alert_tx_0__u_prim_alert_sender_alert_test_set_d;
 wire gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q;
 wire gen_alert_tx_0__u_prim_alert_sender_n1;
 wire gen_alert_tx_0__u_prim_alert_sender_ping_set_d;
 wire gen_alert_tx_0__u_prim_alert_sender_ping_set_q;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nd;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_intq_0_;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_intq_0_;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_intq_0_;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_intq_0_;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q;
 wire gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_n3;
 wire gen_filter_0__u_filter_filter_q;
 wire gen_filter_0__u_filter_filter_synced;
 wire gen_filter_0__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_0__u_filter_stored_value_q;
 wire gen_filter_10__u_filter_filter_q;
 wire gen_filter_10__u_filter_filter_synced;
 wire gen_filter_10__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_10__u_filter_stored_value_q;
 wire gen_filter_11__u_filter_filter_q;
 wire gen_filter_11__u_filter_filter_synced;
 wire gen_filter_11__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_11__u_filter_stored_value_q;
 wire gen_filter_12__u_filter_filter_q;
 wire gen_filter_12__u_filter_filter_synced;
 wire gen_filter_12__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_12__u_filter_stored_value_q;
 wire gen_filter_13__u_filter_filter_q;
 wire gen_filter_13__u_filter_filter_synced;
 wire gen_filter_13__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_13__u_filter_stored_value_q;
 wire gen_filter_14__u_filter_filter_q;
 wire gen_filter_14__u_filter_filter_synced;
 wire gen_filter_14__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_14__u_filter_stored_value_q;
 wire gen_filter_15__u_filter_filter_q;
 wire gen_filter_15__u_filter_filter_synced;
 wire gen_filter_15__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_15__u_filter_stored_value_q;
 wire gen_filter_16__u_filter_filter_q;
 wire gen_filter_16__u_filter_filter_synced;
 wire gen_filter_16__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_16__u_filter_stored_value_q;
 wire gen_filter_17__u_filter_filter_q;
 wire gen_filter_17__u_filter_filter_synced;
 wire gen_filter_17__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_17__u_filter_stored_value_q;
 wire gen_filter_18__u_filter_filter_q;
 wire gen_filter_18__u_filter_filter_synced;
 wire gen_filter_18__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_18__u_filter_stored_value_q;
 wire gen_filter_19__u_filter_filter_q;
 wire gen_filter_19__u_filter_filter_synced;
 wire gen_filter_19__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_19__u_filter_stored_value_q;
 wire gen_filter_1__u_filter_filter_q;
 wire gen_filter_1__u_filter_filter_synced;
 wire gen_filter_1__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_1__u_filter_stored_value_q;
 wire gen_filter_20__u_filter_filter_q;
 wire gen_filter_20__u_filter_filter_synced;
 wire gen_filter_20__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_20__u_filter_stored_value_q;
 wire gen_filter_21__u_filter_filter_q;
 wire gen_filter_21__u_filter_filter_synced;
 wire gen_filter_21__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_21__u_filter_stored_value_q;
 wire gen_filter_22__u_filter_filter_q;
 wire gen_filter_22__u_filter_filter_synced;
 wire gen_filter_22__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_22__u_filter_stored_value_q;
 wire gen_filter_23__u_filter_filter_q;
 wire gen_filter_23__u_filter_filter_synced;
 wire gen_filter_23__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_23__u_filter_stored_value_q;
 wire gen_filter_24__u_filter_filter_q;
 wire gen_filter_24__u_filter_filter_synced;
 wire gen_filter_24__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_24__u_filter_stored_value_q;
 wire gen_filter_25__u_filter_filter_q;
 wire gen_filter_25__u_filter_filter_synced;
 wire gen_filter_25__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_25__u_filter_stored_value_q;
 wire gen_filter_26__u_filter_filter_q;
 wire gen_filter_26__u_filter_filter_synced;
 wire gen_filter_26__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_26__u_filter_stored_value_q;
 wire gen_filter_27__u_filter_filter_q;
 wire gen_filter_27__u_filter_filter_synced;
 wire gen_filter_27__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_27__u_filter_stored_value_q;
 wire gen_filter_28__u_filter_filter_q;
 wire gen_filter_28__u_filter_filter_synced;
 wire gen_filter_28__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_28__u_filter_stored_value_q;
 wire gen_filter_29__u_filter_filter_q;
 wire gen_filter_29__u_filter_filter_synced;
 wire gen_filter_29__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_29__u_filter_stored_value_q;
 wire gen_filter_2__u_filter_filter_q;
 wire gen_filter_2__u_filter_filter_synced;
 wire gen_filter_2__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_2__u_filter_stored_value_q;
 wire gen_filter_30__u_filter_filter_q;
 wire gen_filter_30__u_filter_filter_synced;
 wire gen_filter_30__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_30__u_filter_stored_value_q;
 wire gen_filter_31__u_filter_filter_q;
 wire gen_filter_31__u_filter_filter_synced;
 wire gen_filter_31__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_31__u_filter_stored_value_q;
 wire gen_filter_3__u_filter_filter_q;
 wire gen_filter_3__u_filter_filter_synced;
 wire gen_filter_3__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_3__u_filter_stored_value_q;
 wire gen_filter_4__u_filter_filter_q;
 wire gen_filter_4__u_filter_filter_synced;
 wire gen_filter_4__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_4__u_filter_stored_value_q;
 wire gen_filter_5__u_filter_filter_q;
 wire gen_filter_5__u_filter_filter_synced;
 wire gen_filter_5__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_5__u_filter_stored_value_q;
 wire gen_filter_6__u_filter_filter_q;
 wire gen_filter_6__u_filter_filter_synced;
 wire gen_filter_6__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_6__u_filter_stored_value_q;
 wire gen_filter_7__u_filter_filter_q;
 wire gen_filter_7__u_filter_filter_synced;
 wire gen_filter_7__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_7__u_filter_stored_value_q;
 wire gen_filter_8__u_filter_filter_q;
 wire gen_filter_8__u_filter_filter_synced;
 wire gen_filter_8__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_8__u_filter_stored_value_q;
 wire gen_filter_9__u_filter_filter_q;
 wire gen_filter_9__u_filter_filter_synced;
 wire gen_filter_9__u_filter_gen_async_prim_flop_2sync_intq_0_;
 wire gen_filter_9__u_filter_stored_value_q;
 wire intr_hw_N1;
 wire intr_hw_N10;
 wire intr_hw_N11;
 wire intr_hw_N12;
 wire intr_hw_N13;
 wire intr_hw_N14;
 wire intr_hw_N15;
 wire intr_hw_N16;
 wire intr_hw_N17;
 wire intr_hw_N18;
 wire intr_hw_N19;
 wire intr_hw_N2;
 wire intr_hw_N20;
 wire intr_hw_N21;
 wire intr_hw_N22;
 wire intr_hw_N23;
 wire intr_hw_N24;
 wire intr_hw_N25;
 wire intr_hw_N26;
 wire intr_hw_N27;
 wire intr_hw_N28;
 wire intr_hw_N29;
 wire intr_hw_N3;
 wire intr_hw_N30;
 wire intr_hw_N31;
 wire intr_hw_N32;
 wire intr_hw_N4;
 wire intr_hw_N5;
 wire intr_hw_N6;
 wire intr_hw_N7;
 wire intr_hw_N8;
 wire intr_hw_N9;
 wire n1429;
 wire n1432;
 wire n1439;
 wire n2683;
 wire n2684;
 wire n2685;
 wire n2686;
 wire n2687;
 wire n2688;
 wire n2689;
 wire n2690;
 wire n2691;
 wire n2692;
 wire n2693;
 wire n2694;
 wire n2695;
 wire n2696;
 wire n2697;
 wire n2698;
 wire n2699;
 wire n2700;
 wire n2701;
 wire n2702;
 wire n2703;
 wire n2704;
 wire n2705;
 wire n2706;
 wire n2707;
 wire n2708;
 wire n2709;
 wire n2710;
 wire n2711;
 wire n2712;
 wire n2713;
 wire n2714;
 wire n2715;
 wire n2716;
 wire n2717;
 wire n2718;
 wire n2719;
 wire n2720;
 wire n2721;
 wire n2722;
 wire n2723;
 wire n2724;
 wire n2725;
 wire n2726;
 wire n2727;
 wire n2728;
 wire n2729;
 wire n2730;
 wire n2731;
 wire n2732;
 wire n2733;
 wire n2734;
 wire n2735;
 wire n2736;
 wire n2737;
 wire n2738;
 wire n2739;
 wire n2740;
 wire n2741;
 wire n2742;
 wire n2743;
 wire n2744;
 wire n2745;
 wire n2746;
 wire n2747;
 wire n2748;
 wire n2749;
 wire n2750;
 wire n2751;
 wire n2752;
 wire n2753;
 wire n2754;
 wire n2755;
 wire n2756;
 wire n2757;
 wire n2758;
 wire n2759;
 wire n2760;
 wire n2761;
 wire n2762;
 wire n2763;
 wire n2764;
 wire n2765;
 wire n2766;
 wire n2767;
 wire n2768;
 wire n2769;
 wire n2770;
 wire n2771;
 wire n2772;
 wire n2773;
 wire n2774;
 wire n2775;
 wire n2776;
 wire n2777;
 wire n2778;
 wire n2779;
 wire n2780;
 wire n2781;
 wire n2782;
 wire n2783;
 wire n2784;
 wire n2785;
 wire n2786;
 wire n2787;
 wire n2788;
 wire n2789;
 wire n2790;
 wire n2791;
 wire n2792;
 wire n2793;
 wire n2794;
 wire n2795;
 wire n2796;
 wire n2797;
 wire n2798;
 wire n2799;
 wire n2800;
 wire n2801;
 wire n2802;
 wire n2803;
 wire n2804;
 wire n2805;
 wire n2806;
 wire n2807;
 wire n2808;
 wire n2809;
 wire n2810;
 wire n2811;
 wire n2812;
 wire n2813;
 wire n2814;
 wire n2815;
 wire n2816;
 wire n2817;
 wire n2818;
 wire n2819;
 wire n2820;
 wire n2821;
 wire n2822;
 wire n2823;
 wire n2824;
 wire n2825;
 wire n2826;
 wire n2827;
 wire n2828;
 wire n2829;
 wire n2830;
 wire n2831;
 wire n2832;
 wire n2833;
 wire n2834;
 wire n2835;
 wire n2836;
 wire n2837;
 wire n2838;
 wire n2839;
 wire n2840;
 wire n2841;
 wire n2842;
 wire n2843;
 wire n2844;
 wire n2845;
 wire n2846;
 wire n2847;
 wire n2848;
 wire n2849;
 wire n2850;
 wire n2851;
 wire n2852;
 wire n2853;
 wire n2854;
 wire n2855;
 wire n2856;
 wire n2857;
 wire n2858;
 wire n2859;
 wire n2860;
 wire n2861;
 wire n2862;
 wire n2863;
 wire n2864;
 wire n2865;
 wire n2866;
 wire n2867;
 wire n2868;
 wire n2869;
 wire n2870;
 wire n2871;
 wire n2872;
 wire n2873;
 wire n2874;
 wire n2875;
 wire n2876;
 wire n2877;
 wire n2878;
 wire n2879;
 wire n2880;
 wire n2881;
 wire n2882;
 wire n2883;
 wire n2884;
 wire n2885;
 wire n2886;
 wire n2887;
 wire n2888;
 wire n2889;
 wire n2890;
 wire n2891;
 wire n2892;
 wire n2893;
 wire n2894;
 wire n2895;
 wire n2896;
 wire n2897;
 wire n2898;
 wire n2899;
 wire n2900;
 wire n2901;
 wire n2902;
 wire n2903;
 wire n2904;
 wire n2905;
 wire n2906;
 wire n2907;
 wire n2908;
 wire n2909;
 wire n2910;
 wire n2911;
 wire n2912;
 wire n2913;
 wire n2914;
 wire n2915;
 wire n2916;
 wire n2917;
 wire n2918;
 wire n2919;
 wire n2920;
 wire n2921;
 wire n2922;
 wire n2923;
 wire n2924;
 wire n2925;
 wire n2926;
 wire n2927;
 wire n2928;
 wire n2929;
 wire n2930;
 wire n2931;
 wire n2932;
 wire n2933;
 wire n2934;
 wire n2935;
 wire n2936;
 wire n2937;
 wire n2938;
 wire n2939;
 wire n2940;
 wire n2941;
 wire n2942;
 wire n2943;
 wire n2944;
 wire n2945;
 wire n2946;
 wire n2947;
 wire n2948;
 wire n2949;
 wire n2950;
 wire n2951;
 wire n2952;
 wire n2953;
 wire n2954;
 wire n2955;
 wire n2956;
 wire n2957;
 wire n2958;
 wire n2959;
 wire n2960;
 wire n2961;
 wire n2962;
 wire n2963;
 wire n2964;
 wire n2965;
 wire n2966;
 wire n2967;
 wire n2968;
 wire n2969;
 wire n2970;
 wire n2971;
 wire n2972;
 wire n2973;
 wire n2974;
 wire n2975;
 wire n2976;
 wire n2977;
 wire n2978;
 wire n2979;
 wire n2980;
 wire n2981;
 wire n2982;
 wire n2983;
 wire n2984;
 wire n2985;
 wire n2986;
 wire n2987;
 wire n2988;
 wire n2989;
 wire n2990;
 wire n2991;
 wire n2992;
 wire n2993;
 wire n2994;
 wire n2995;
 wire n2996;
 wire n2997;
 wire n2998;
 wire n2999;
 wire n3000;
 wire n3001;
 wire n3002;
 wire n3003;
 wire n3004;
 wire n3005;
 wire n3006;
 wire n3007;
 wire n3008;
 wire n3009;
 wire n3010;
 wire n3011;
 wire n3012;
 wire n3013;
 wire n3014;
 wire n3015;
 wire n3016;
 wire n3017;
 wire n3018;
 wire n3019;
 wire n3020;
 wire n3021;
 wire n3022;
 wire n3023;
 wire n3024;
 wire n3025;
 wire n3026;
 wire n3027;
 wire n3028;
 wire n3029;
 wire n3030;
 wire n3031;
 wire n3032;
 wire n3033;
 wire n3034;
 wire n3035;
 wire n3036;
 wire n3037;
 wire n3038;
 wire n3039;
 wire n3040;
 wire n3041;
 wire n3042;
 wire n3043;
 wire n3044;
 wire n3045;
 wire n3046;
 wire n3047;
 wire n3048;
 wire n3049;
 wire n3050;
 wire n3051;
 wire n3052;
 wire n3053;
 wire n3054;
 wire n3055;
 wire n3056;
 wire n3057;
 wire n3058;
 wire n3059;
 wire n3060;
 wire n3061;
 wire n3062;
 wire n3063;
 wire n3064;
 wire n3065;
 wire n3066;
 wire n3067;
 wire n3068;
 wire n3069;
 wire n3070;
 wire n3071;
 wire n3072;
 wire n3073;
 wire n3074;
 wire n3075;
 wire n3076;
 wire n3077;
 wire n3078;
 wire n3079;
 wire n3080;
 wire n3081;
 wire n3082;
 wire n3083;
 wire n3084;
 wire n3085;
 wire n3086;
 wire n3087;
 wire n3088;
 wire n3089;
 wire n3090;
 wire n3091;
 wire n3092;
 wire n3093;
 wire n3094;
 wire n3095;
 wire n3096;
 wire n3097;
 wire n3098;
 wire n3099;
 wire n3100;
 wire n3101;
 wire n3102;
 wire n3103;
 wire n3104;
 wire n3105;
 wire n3106;
 wire n3107;
 wire n3108;
 wire n3109;
 wire n3110;
 wire n3111;
 wire n3112;
 wire n3113;
 wire n3114;
 wire n3115;
 wire n3116;
 wire n3117;
 wire n3118;
 wire n3119;
 wire n3120;
 wire n3121;
 wire n3122;
 wire n3123;
 wire n3124;
 wire n3125;
 wire n3126;
 wire n3127;
 wire n3128;
 wire n3129;
 wire n3130;
 wire n3131;
 wire n3132;
 wire n3133;
 wire n3134;
 wire n3135;
 wire n3136;
 wire n3137;
 wire n3138;
 wire n3139;
 wire n3140;
 wire n3141;
 wire n3142;
 wire n3143;
 wire n3144;
 wire n3145;
 wire n3146;
 wire n3147;
 wire n3148;
 wire n3149;
 wire n3150;
 wire n3151;
 wire n3152;
 wire n3153;
 wire n3154;
 wire n3155;
 wire n3156;
 wire n3157;
 wire n3158;
 wire n3159;
 wire n3160;
 wire n3161;
 wire n3162;
 wire n3163;
 wire n3164;
 wire n3165;
 wire n3166;
 wire n3167;
 wire n3168;
 wire n3169;
 wire n3170;
 wire n3171;
 wire n3172;
 wire n3173;
 wire n3174;
 wire n3175;
 wire n3176;
 wire n3177;
 wire n3178;
 wire n3179;
 wire n3180;
 wire n3181;
 wire n3182;
 wire n3183;
 wire n3184;
 wire n3185;
 wire n3186;
 wire n3187;
 wire n3188;
 wire n3189;
 wire n3190;
 wire n3191;
 wire n3192;
 wire n3193;
 wire n3194;
 wire n3195;
 wire n3196;
 wire n3197;
 wire n3198;
 wire n3199;
 wire n3200;
 wire n3201;
 wire n3202;
 wire n3203;
 wire n3204;
 wire n3205;
 wire n3206;
 wire n3207;
 wire n3208;
 wire n3209;
 wire n3210;
 wire n3211;
 wire n3212;
 wire n3213;
 wire n3214;
 wire n3215;
 wire n3216;
 wire n3217;
 wire n3218;
 wire n3219;
 wire n3220;
 wire n3221;
 wire n3222;
 wire n3223;
 wire n3224;
 wire n3225;
 wire n3226;
 wire n3227;
 wire n3228;
 wire n3229;
 wire n3230;
 wire n3231;
 wire n3232;
 wire n3233;
 wire n3234;
 wire n3235;
 wire n3236;
 wire n3237;
 wire n3238;
 wire n3239;
 wire n3240;
 wire n3241;
 wire n3242;
 wire n3243;
 wire n3244;
 wire n3245;
 wire n3246;
 wire n3247;
 wire n3248;
 wire n3249;
 wire n3250;
 wire n3251;
 wire n3252;
 wire n3253;
 wire n3254;
 wire n3255;
 wire n3256;
 wire n3257;
 wire n3258;
 wire n3259;
 wire n3260;
 wire n3261;
 wire n3262;
 wire n3263;
 wire n3264;
 wire n3265;
 wire n3266;
 wire n3267;
 wire n3268;
 wire n3269;
 wire n3270;
 wire n3271;
 wire n3272;
 wire n3273;
 wire n3274;
 wire n3275;
 wire n3276;
 wire n3277;
 wire n3278;
 wire n3279;
 wire n3280;
 wire n3281;
 wire n3282;
 wire n3283;
 wire n3284;
 wire n3285;
 wire n3286;
 wire n3287;
 wire n3288;
 wire n3289;
 wire n3290;
 wire n3291;
 wire n3292;
 wire n3293;
 wire n3294;
 wire n3295;
 wire n3296;
 wire n3297;
 wire n3298;
 wire n3299;
 wire n3300;
 wire n3301;
 wire n3302;
 wire n3303;
 wire n3304;
 wire n3305;
 wire n3306;
 wire n3307;
 wire n3308;
 wire n3309;
 wire n3310;
 wire n3311;
 wire n3312;
 wire n3313;
 wire n3314;
 wire n3315;
 wire n3316;
 wire n3317;
 wire n3318;
 wire n3319;
 wire n3320;
 wire n3321;
 wire n3322;
 wire n3323;
 wire n3324;
 wire n3326;
 wire n3327;
 wire n3328;
 wire n3329;
 wire n3330;
 wire n3331;
 wire n3332;
 wire n3333;
 wire n3334;
 wire n3335;
 wire n3336;
 wire n3337;
 wire n3338;
 wire n3359;
 wire n3361;
 wire n3362;
 wire n3363;
 wire n3364;
 wire n3365;
 wire n3366;
 wire n3367;
 wire n3368;
 wire n3369;
 wire n3370;
 wire n3371;
 wire n3372;
 wire n3373;
 wire n3374;
 wire n3375;
 wire n3376;
 wire n3377;
 wire n3378;
 wire n3379;
 wire n3380;
 wire n3381;
 wire n3382;
 wire n3383;
 wire n3384;
 wire n3385;
 wire n3386;
 wire n3387;
 wire n3389;
 wire n3390;
 wire n3392;
 wire n3397;
 wire n3398;
 wire n3399;
 wire n3400;
 wire n3401;
 wire n3402;
 wire n3403;
 wire n3404;
 wire n3405;
 wire n3406;
 wire n3407;
 wire n3408;
 wire n3409;
 wire n3410;
 wire n3411;
 wire n3412;
 wire n3414;
 wire n3415;
 wire n3416;
 wire n3417;
 wire n3418;
 wire n3419;
 wire n3420;
 wire n3421;
 wire n3422;
 wire n3423;
 wire n3424;
 wire n3425;
 wire n3426;
 wire n3427;
 wire n3428;
 wire n3429;
 wire n3431;
 wire n3432;
 wire n3433;
 wire n3434;
 wire n3435;
 wire n3436;
 wire n3437;
 wire n3438;
 wire n3439;
 wire n3440;
 wire n3441;
 wire n3442;
 wire n3443;
 wire n3444;
 wire n3445;
 wire n3446;
 wire n3447;
 wire n3448;
 wire n3449;
 wire n3450;
 wire n3451;
 wire n3452;
 wire n3453;
 wire n3454;
 wire n3455;
 wire n3456;
 wire n3457;
 wire n3458;
 wire n3459;
 wire n3460;
 wire n3461;
 wire n3462;
 wire n3463;
 wire n3464;
 wire n3465;
 wire n3466;
 wire n3467;
 wire n3468;
 wire n3469;
 wire n3471;
 wire n3472;
 wire n3473;
 wire n3474;
 wire n3475;
 wire n3476;
 wire n3477;
 wire n3479;
 wire n3480;
 wire n3481;
 wire n3482;
 wire n3483;
 wire n3484;
 wire n3486;
 wire n3487;
 wire n3488;
 wire n3489;
 wire n3490;
 wire n3492;
 wire n3493;
 wire n3494;
 wire n3495;
 wire n3496;
 wire n3497;
 wire n3498;
 wire n3499;
 wire n3500;
 wire n3501;
 wire n3502;
 wire n3504;
 wire n3505;
 wire n3506;
 wire n3507;
 wire n3508;
 wire n3509;
 wire n3511;
 wire n3512;
 wire n3513;
 wire n3514;
 wire n3515;
 wire n3516;
 wire n3518;
 wire n3519;
 wire n3520;
 wire n3521;
 wire n3522;
 wire n3523;
 wire n3524;
 wire n3525;
 wire n3526;
 wire n3527;
 wire n3528;
 wire n3529;
 wire n3530;
 wire n3532;
 wire n3533;
 wire n3534;
 wire n3535;
 wire n3536;
 wire n3537;
 wire n3538;
 wire n3539;
 wire n3540;
 wire n3541;
 wire n3542;
 wire n3543;
 wire n3544;
 wire n3546;
 wire n3547;
 wire n3548;
 wire n3549;
 wire n3550;
 wire n3551;
 wire n3553;
 wire n3554;
 wire n3555;
 wire n3556;
 wire n3557;
 wire n3558;
 wire n3560;
 wire n3561;
 wire n3562;
 wire n3563;
 wire n3564;
 wire n3565;
 wire n3567;
 wire n3568;
 wire n3569;
 wire n3570;
 wire n3571;
 wire n3572;
 wire n3574;
 wire n3575;
 wire n3576;
 wire n3577;
 wire n3578;
 wire n3579;
 wire n3581;
 wire n3582;
 wire n3583;
 wire n3584;
 wire n3585;
 wire n3586;
 wire n3588;
 wire n3589;
 wire n3590;
 wire n3591;
 wire n3592;
 wire n3593;
 wire n3595;
 wire n3596;
 wire n3597;
 wire n3598;
 wire n3599;
 wire n3600;
 wire n3602;
 wire n3603;
 wire n3604;
 wire n3605;
 wire n3606;
 wire n3607;
 wire n3610;
 wire n3611;
 wire n3613;
 wire n3614;
 wire n3615;
 wire n3616;
 wire n3618;
 wire n3619;
 wire n3620;
 wire n3621;
 wire n3622;
 wire n3623;
 wire n3625;
 wire n3626;
 wire n3627;
 wire n3628;
 wire n3629;
 wire n3630;
 wire n3632;
 wire n3633;
 wire n3634;
 wire n3635;
 wire n3636;
 wire n3637;
 wire n3639;
 wire n3640;
 wire n3641;
 wire n3642;
 wire n3643;
 wire n3644;
 wire n3646;
 wire n3647;
 wire n3648;
 wire n3649;
 wire n3650;
 wire n3651;
 wire n3653;
 wire n3654;
 wire n3655;
 wire n3656;
 wire n3657;
 wire n3658;
 wire n3660;
 wire n3661;
 wire n3662;
 wire n3663;
 wire n3664;
 wire n3665;
 wire n3667;
 wire n3668;
 wire n3669;
 wire n3670;
 wire n3671;
 wire n3672;
 wire n3674;
 wire n3675;
 wire n3676;
 wire n3677;
 wire n3678;
 wire n3679;
 wire n3681;
 wire n3682;
 wire n3683;
 wire n3684;
 wire n3685;
 wire n3686;
 wire n3688;
 wire n3689;
 wire n3690;
 wire n3691;
 wire n3692;
 wire n3693;
 wire n3696;
 wire n3697;
 wire n3698;
 wire n3699;
 wire n3700;
 wire n3701;
 wire n3703;
 wire n3704;
 wire n3705;
 wire n3706;
 wire n3707;
 wire n3708;
 wire n3712;
 wire n3713;
 wire n3714;
 wire n3715;
 wire n3716;
 wire n3717;
 wire n3718;
 wire n3719;
 wire n3720;
 wire n3721;
 wire n3722;
 wire n3723;
 wire n3725;
 wire n3726;
 wire n3727;
 wire n3728;
 wire n3729;
 wire n3730;
 wire n3731;
 wire n3732;
 wire n3733;
 wire n3734;
 wire n3735;
 wire n3736;
 wire n3737;
 wire n3738;
 wire n3739;
 wire n3740;
 wire n3741;
 wire n3742;
 wire n3743;
 wire n3744;
 wire n3745;
 wire n3746;
 wire n3747;
 wire n3748;
 wire n3749;
 wire n3750;
 wire n3751;
 wire n3752;
 wire n3753;
 wire n3754;
 wire n3755;
 wire n3756;
 wire n3759;
 wire n3760;
 wire n3761;
 wire n3762;
 wire n3763;
 wire n3764;
 wire n3765;
 wire n3766;
 wire n3767;
 wire n3770;
 wire n3771;
 wire n3772;
 wire n3773;
 wire n3774;
 wire n3775;
 wire n3776;
 wire n3777;
 wire n3778;
 wire n3779;
 wire n3780;
 wire n3781;
 wire n3782;
 wire n3783;
 wire n3784;
 wire n3785;
 wire n3786;
 wire n3787;
 wire n3788;
 wire n3789;
 wire n3790;
 wire n3791;
 wire n3792;
 wire n3793;
 wire n3794;
 wire n3795;
 wire n3796;
 wire n3797;
 wire n3798;
 wire n3799;
 wire n3800;
 wire n3801;
 wire n3802;
 wire n3803;
 wire n3804;
 wire n3805;
 wire n3806;
 wire n3807;
 wire n3808;
 wire n3809;
 wire n3810;
 wire n3811;
 wire n3812;
 wire n3813;
 wire n3814;
 wire n3815;
 wire n3816;
 wire n3817;
 wire n3818;
 wire n3819;
 wire n3820;
 wire n3821;
 wire n3822;
 wire n3823;
 wire n3824;
 wire n3825;
 wire n3826;
 wire n3827;
 wire n3828;
 wire n3829;
 wire n3830;
 wire n3831;
 wire n3832;
 wire n3833;
 wire n3834;
 wire n3835;
 wire n3836;
 wire n3837;
 wire n3838;
 wire n3839;
 wire n3840;
 wire n3841;
 wire n3842;
 wire n3843;
 wire n3845;
 wire n3846;
 wire n3847;
 wire n3849;
 wire n3850;
 wire n3851;
 wire n3852;
 wire n3853;
 wire n3854;
 wire n3855;
 wire n3856;
 wire n3857;
 wire n3858;
 wire n3859;
 wire n3860;
 wire n3861;
 wire n3862;
 wire n3863;
 wire n3864;
 wire n3865;
 wire n3866;
 wire n3867;
 wire n3868;
 wire n3869;
 wire n3870;
 wire n3871;
 wire n3872;
 wire n3873;
 wire n3874;
 wire n3875;
 wire n3876;
 wire n3877;
 wire n3878;
 wire n3879;
 wire n3880;
 wire n3881;
 wire n3882;
 wire n3883;
 wire n3884;
 wire n3885;
 wire n3886;
 wire n3887;
 wire n3889;
 wire n3890;
 wire n3891;
 wire n3892;
 wire n3893;
 wire n3894;
 wire n3895;
 wire n3896;
 wire n3897;
 wire n3898;
 wire n3899;
 wire n3900;
 wire n3901;
 wire n3902;
 wire n3903;
 wire n3904;
 wire n3905;
 wire n3906;
 wire n3907;
 wire n3908;
 wire n3909;
 wire n3911;
 wire n3912;
 wire n3913;
 wire n3915;
 wire n3916;
 wire n3917;
 wire n3918;
 wire n3920;
 wire n3921;
 wire n3922;
 wire n3924;
 wire n3925;
 wire n3926;
 wire n3927;
 wire n3931;
 wire n3932;
 wire n3933;
 wire n3935;
 wire n3936;
 wire n3937;
 wire n3938;
 wire n3939;
 wire n3940;
 wire n3941;
 wire n3942;
 wire n3943;
 wire n3944;
 wire n3945;
 wire n3946;
 wire n3947;
 wire n3948;
 wire n3949;
 wire n3950;
 wire n3951;
 wire n3952;
 wire n3953;
 wire n3954;
 wire n3955;
 wire n3958;
 wire n3959;
 wire n3960;
 wire n3961;
 wire n3966;
 wire n3967;
 wire n3968;
 wire n3970;
 wire n3971;
 wire n3972;
 wire n3973;
 wire n3981;
 wire n3982;
 wire n3983;
 wire n3984;
 wire n3986;
 wire n3989;
 wire n3990;
 wire n3991;
 wire n3992;
 wire n3993;
 wire n3994;
 wire n3995;
 wire n3996;
 wire n4067;
 wire n4068;
 wire n4069;
 wire n4070;
 wire n4071;
 wire n4072;
 wire n4073;
 wire n4074;
 wire n4075;
 wire n4076;
 wire n4077;
 wire n4078;
 wire n4079;
 wire n4080;
 wire n4081;
 wire n4082;
 wire n4083;
 wire n4084;
 wire n4085;
 wire n4086;
 wire n4087;
 wire n4088;
 wire n4089;
 wire n4090;
 wire n4091;
 wire n4092;
 wire n4093;
 wire n4094;
 wire n4095;
 wire n4096;
 wire net96;
 wire net95;
 wire net94;
 wire net93;
 wire net92;
 wire net91;
 wire net90;
 wire net89;
 wire net88;
 wire net87;
 wire net85;
 wire net83;
 wire net82;
 wire net81;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire net75;
 wire net74;
 wire net73;
 wire net72;
 wire n4123;
 wire n4124;
 wire n4125;
 wire n4126;
 wire n4127;
 wire n4128;
 wire n4129;
 wire n4130;
 wire net71;
 wire net70;
 wire net69;
 wire net68;
 wire net67;
 wire net66;
 wire net65;
 wire net64;
 wire net63;
 wire net62;
 wire net61;
 wire net60;
 wire net59;
 wire net58;
 wire net57;
 wire net56;
 wire net55;
 wire net54;
 wire net53;
 wire net52;
 wire net51;
 wire net50;
 wire net49;
 wire net48;
 wire net47;
 wire net46;
 wire net45;
 wire net44;
 wire net43;
 wire net42;
 wire net41;
 wire net40;
 wire net39;
 wire net38;
 wire net37;
 wire net36;
 wire net35;
 wire net34;
 wire net33;
 wire net32;
 wire net31;
 wire net30;
 wire net29;
 wire net28;
 wire net27;
 wire net26;
 wire net25;
 wire net24;
 wire net23;
 wire net22;
 wire net21;
 wire net20;
 wire net19;
 wire net18;
 wire net17;
 wire net16;
 wire net15;
 wire net14;
 wire net13;
 wire net12;
 wire net11;
 wire net10;
 wire net9;
 wire net8;
 wire net7;
 wire net6;
 wire net5;
 wire net4;
 wire net3;
 wire net2;
 wire net1;
 wire net86;
 wire net84;
 wire net2034;
 wire net2040;
 wire net2045;
 wire net2050;
 wire clknet_leaf_0_clk_i;
 wire reg2hw_ctrl_en_input_filter__q__0_;
 wire reg2hw_ctrl_en_input_filter__q__10_;
 wire reg2hw_ctrl_en_input_filter__q__11_;
 wire reg2hw_ctrl_en_input_filter__q__12_;
 wire reg2hw_ctrl_en_input_filter__q__13_;
 wire reg2hw_ctrl_en_input_filter__q__14_;
 wire reg2hw_ctrl_en_input_filter__q__15_;
 wire reg2hw_ctrl_en_input_filter__q__16_;
 wire reg2hw_ctrl_en_input_filter__q__17_;
 wire reg2hw_ctrl_en_input_filter__q__18_;
 wire reg2hw_ctrl_en_input_filter__q__19_;
 wire reg2hw_ctrl_en_input_filter__q__1_;
 wire reg2hw_ctrl_en_input_filter__q__20_;
 wire reg2hw_ctrl_en_input_filter__q__21_;
 wire reg2hw_ctrl_en_input_filter__q__22_;
 wire reg2hw_ctrl_en_input_filter__q__23_;
 wire reg2hw_ctrl_en_input_filter__q__24_;
 wire reg2hw_ctrl_en_input_filter__q__25_;
 wire reg2hw_ctrl_en_input_filter__q__26_;
 wire reg2hw_ctrl_en_input_filter__q__27_;
 wire reg2hw_ctrl_en_input_filter__q__28_;
 wire reg2hw_ctrl_en_input_filter__q__29_;
 wire reg2hw_ctrl_en_input_filter__q__2_;
 wire reg2hw_ctrl_en_input_filter__q__30_;
 wire reg2hw_ctrl_en_input_filter__q__31_;
 wire reg2hw_ctrl_en_input_filter__q__3_;
 wire reg2hw_ctrl_en_input_filter__q__4_;
 wire reg2hw_ctrl_en_input_filter__q__5_;
 wire reg2hw_ctrl_en_input_filter__q__6_;
 wire reg2hw_ctrl_en_input_filter__q__7_;
 wire reg2hw_ctrl_en_input_filter__q__8_;
 wire reg2hw_ctrl_en_input_filter__q__9_;
 wire reg2hw_intr_ctrl_en_falling__q__0_;
 wire reg2hw_intr_ctrl_en_falling__q__10_;
 wire reg2hw_intr_ctrl_en_falling__q__11_;
 wire reg2hw_intr_ctrl_en_falling__q__12_;
 wire reg2hw_intr_ctrl_en_falling__q__13_;
 wire reg2hw_intr_ctrl_en_falling__q__14_;
 wire reg2hw_intr_ctrl_en_falling__q__15_;
 wire reg2hw_intr_ctrl_en_falling__q__16_;
 wire reg2hw_intr_ctrl_en_falling__q__17_;
 wire reg2hw_intr_ctrl_en_falling__q__18_;
 wire reg2hw_intr_ctrl_en_falling__q__19_;
 wire reg2hw_intr_ctrl_en_falling__q__1_;
 wire reg2hw_intr_ctrl_en_falling__q__20_;
 wire reg2hw_intr_ctrl_en_falling__q__21_;
 wire reg2hw_intr_ctrl_en_falling__q__22_;
 wire reg2hw_intr_ctrl_en_falling__q__23_;
 wire reg2hw_intr_ctrl_en_falling__q__24_;
 wire reg2hw_intr_ctrl_en_falling__q__25_;
 wire reg2hw_intr_ctrl_en_falling__q__26_;
 wire reg2hw_intr_ctrl_en_falling__q__27_;
 wire reg2hw_intr_ctrl_en_falling__q__28_;
 wire reg2hw_intr_ctrl_en_falling__q__29_;
 wire reg2hw_intr_ctrl_en_falling__q__2_;
 wire reg2hw_intr_ctrl_en_falling__q__30_;
 wire reg2hw_intr_ctrl_en_falling__q__31_;
 wire reg2hw_intr_ctrl_en_falling__q__3_;
 wire reg2hw_intr_ctrl_en_falling__q__4_;
 wire reg2hw_intr_ctrl_en_falling__q__5_;
 wire reg2hw_intr_ctrl_en_falling__q__6_;
 wire reg2hw_intr_ctrl_en_falling__q__7_;
 wire reg2hw_intr_ctrl_en_falling__q__8_;
 wire reg2hw_intr_ctrl_en_falling__q__9_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__0_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__10_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__11_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__12_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__13_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__14_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__15_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__16_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__17_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__18_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__19_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__1_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__20_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__21_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__22_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__23_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__24_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__25_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__26_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__27_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__28_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__29_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__2_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__30_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__31_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__3_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__4_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__5_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__6_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__7_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__8_;
 wire reg2hw_intr_ctrl_en_lvlhigh__q__9_;
 wire reg2hw_intr_ctrl_en_lvllow__q__0_;
 wire reg2hw_intr_ctrl_en_lvllow__q__10_;
 wire reg2hw_intr_ctrl_en_lvllow__q__11_;
 wire reg2hw_intr_ctrl_en_lvllow__q__12_;
 wire reg2hw_intr_ctrl_en_lvllow__q__13_;
 wire reg2hw_intr_ctrl_en_lvllow__q__14_;
 wire reg2hw_intr_ctrl_en_lvllow__q__15_;
 wire reg2hw_intr_ctrl_en_lvllow__q__16_;
 wire reg2hw_intr_ctrl_en_lvllow__q__17_;
 wire reg2hw_intr_ctrl_en_lvllow__q__18_;
 wire reg2hw_intr_ctrl_en_lvllow__q__19_;
 wire reg2hw_intr_ctrl_en_lvllow__q__1_;
 wire reg2hw_intr_ctrl_en_lvllow__q__20_;
 wire reg2hw_intr_ctrl_en_lvllow__q__21_;
 wire reg2hw_intr_ctrl_en_lvllow__q__22_;
 wire reg2hw_intr_ctrl_en_lvllow__q__23_;
 wire reg2hw_intr_ctrl_en_lvllow__q__24_;
 wire reg2hw_intr_ctrl_en_lvllow__q__25_;
 wire reg2hw_intr_ctrl_en_lvllow__q__26_;
 wire reg2hw_intr_ctrl_en_lvllow__q__27_;
 wire reg2hw_intr_ctrl_en_lvllow__q__28_;
 wire reg2hw_intr_ctrl_en_lvllow__q__29_;
 wire reg2hw_intr_ctrl_en_lvllow__q__2_;
 wire reg2hw_intr_ctrl_en_lvllow__q__30_;
 wire reg2hw_intr_ctrl_en_lvllow__q__31_;
 wire reg2hw_intr_ctrl_en_lvllow__q__3_;
 wire reg2hw_intr_ctrl_en_lvllow__q__4_;
 wire reg2hw_intr_ctrl_en_lvllow__q__5_;
 wire reg2hw_intr_ctrl_en_lvllow__q__6_;
 wire reg2hw_intr_ctrl_en_lvllow__q__7_;
 wire reg2hw_intr_ctrl_en_lvllow__q__8_;
 wire reg2hw_intr_ctrl_en_lvllow__q__9_;
 wire reg2hw_intr_ctrl_en_rising__q__0_;
 wire reg2hw_intr_ctrl_en_rising__q__10_;
 wire reg2hw_intr_ctrl_en_rising__q__11_;
 wire reg2hw_intr_ctrl_en_rising__q__12_;
 wire reg2hw_intr_ctrl_en_rising__q__13_;
 wire reg2hw_intr_ctrl_en_rising__q__14_;
 wire reg2hw_intr_ctrl_en_rising__q__15_;
 wire reg2hw_intr_ctrl_en_rising__q__16_;
 wire reg2hw_intr_ctrl_en_rising__q__17_;
 wire reg2hw_intr_ctrl_en_rising__q__18_;
 wire reg2hw_intr_ctrl_en_rising__q__19_;
 wire reg2hw_intr_ctrl_en_rising__q__1_;
 wire reg2hw_intr_ctrl_en_rising__q__20_;
 wire reg2hw_intr_ctrl_en_rising__q__21_;
 wire reg2hw_intr_ctrl_en_rising__q__22_;
 wire reg2hw_intr_ctrl_en_rising__q__23_;
 wire reg2hw_intr_ctrl_en_rising__q__24_;
 wire reg2hw_intr_ctrl_en_rising__q__25_;
 wire reg2hw_intr_ctrl_en_rising__q__26_;
 wire reg2hw_intr_ctrl_en_rising__q__27_;
 wire reg2hw_intr_ctrl_en_rising__q__28_;
 wire reg2hw_intr_ctrl_en_rising__q__29_;
 wire reg2hw_intr_ctrl_en_rising__q__2_;
 wire reg2hw_intr_ctrl_en_rising__q__30_;
 wire reg2hw_intr_ctrl_en_rising__q__31_;
 wire reg2hw_intr_ctrl_en_rising__q__3_;
 wire reg2hw_intr_ctrl_en_rising__q__4_;
 wire reg2hw_intr_ctrl_en_rising__q__5_;
 wire reg2hw_intr_ctrl_en_rising__q__6_;
 wire reg2hw_intr_ctrl_en_rising__q__7_;
 wire reg2hw_intr_ctrl_en_rising__q__8_;
 wire reg2hw_intr_ctrl_en_rising__q__9_;
 wire reg2hw_intr_enable__q__0_;
 wire reg2hw_intr_enable__q__10_;
 wire reg2hw_intr_enable__q__11_;
 wire reg2hw_intr_enable__q__12_;
 wire reg2hw_intr_enable__q__13_;
 wire reg2hw_intr_enable__q__14_;
 wire reg2hw_intr_enable__q__15_;
 wire reg2hw_intr_enable__q__16_;
 wire reg2hw_intr_enable__q__17_;
 wire reg2hw_intr_enable__q__18_;
 wire reg2hw_intr_enable__q__19_;
 wire reg2hw_intr_enable__q__1_;
 wire reg2hw_intr_enable__q__20_;
 wire reg2hw_intr_enable__q__21_;
 wire reg2hw_intr_enable__q__22_;
 wire reg2hw_intr_enable__q__23_;
 wire reg2hw_intr_enable__q__24_;
 wire reg2hw_intr_enable__q__25_;
 wire reg2hw_intr_enable__q__26_;
 wire reg2hw_intr_enable__q__27_;
 wire reg2hw_intr_enable__q__28_;
 wire reg2hw_intr_enable__q__29_;
 wire reg2hw_intr_enable__q__2_;
 wire reg2hw_intr_enable__q__30_;
 wire reg2hw_intr_enable__q__31_;
 wire reg2hw_intr_enable__q__3_;
 wire reg2hw_intr_enable__q__4_;
 wire reg2hw_intr_enable__q__5_;
 wire reg2hw_intr_enable__q__6_;
 wire reg2hw_intr_enable__q__7_;
 wire reg2hw_intr_enable__q__8_;
 wire reg2hw_intr_enable__q__9_;
 wire reg2hw_intr_state__q__0_;
 wire reg2hw_intr_state__q__10_;
 wire reg2hw_intr_state__q__11_;
 wire reg2hw_intr_state__q__12_;
 wire reg2hw_intr_state__q__13_;
 wire reg2hw_intr_state__q__14_;
 wire reg2hw_intr_state__q__15_;
 wire reg2hw_intr_state__q__16_;
 wire reg2hw_intr_state__q__17_;
 wire reg2hw_intr_state__q__18_;
 wire reg2hw_intr_state__q__19_;
 wire reg2hw_intr_state__q__1_;
 wire reg2hw_intr_state__q__20_;
 wire reg2hw_intr_state__q__21_;
 wire reg2hw_intr_state__q__22_;
 wire reg2hw_intr_state__q__23_;
 wire reg2hw_intr_state__q__24_;
 wire reg2hw_intr_state__q__25_;
 wire reg2hw_intr_state__q__26_;
 wire reg2hw_intr_state__q__27_;
 wire reg2hw_intr_state__q__28_;
 wire reg2hw_intr_state__q__29_;
 wire reg2hw_intr_state__q__2_;
 wire reg2hw_intr_state__q__30_;
 wire reg2hw_intr_state__q__31_;
 wire reg2hw_intr_state__q__3_;
 wire reg2hw_intr_state__q__4_;
 wire reg2hw_intr_state__q__5_;
 wire reg2hw_intr_state__q__6_;
 wire reg2hw_intr_state__q__7_;
 wire reg2hw_intr_state__q__8_;
 wire reg2hw_intr_state__q__9_;
 wire u_reg_err_q;
 wire u_reg_u_ctrl_en_input_filter_net2067;
 wire u_reg_u_ctrl_en_input_filter_net2073;
 wire u_reg_u_intr_ctrl_en_falling_net2067;
 wire u_reg_u_intr_ctrl_en_falling_net2073;
 wire u_reg_u_intr_ctrl_en_lvlhigh_net2067;
 wire u_reg_u_intr_ctrl_en_lvlhigh_net2073;
 wire u_reg_u_intr_ctrl_en_lvllow_net2067;
 wire u_reg_u_intr_ctrl_en_lvllow_net2073;
 wire u_reg_u_intr_ctrl_en_rising_net2067;
 wire u_reg_u_intr_ctrl_en_rising_net2073;
 wire u_reg_u_intr_enable_net2067;
 wire u_reg_u_intr_enable_net2073;
 wire u_reg_u_intr_state_n1;
 wire u_reg_u_intr_state_net2090;
 wire u_reg_u_intr_state_net2096;
 wire u_reg_u_reg_if_N14;
 wire u_reg_u_reg_if_N15;
 wire u_reg_u_reg_if_N16;
 wire u_reg_u_reg_if_N17;
 wire u_reg_u_reg_if_N18;
 wire u_reg_u_reg_if_N19;
 wire u_reg_u_reg_if_N20;
 wire u_reg_u_reg_if_N21;
 wire u_reg_u_reg_if_N22;
 wire u_reg_u_reg_if_N23;
 wire u_reg_u_reg_if_N24;
 wire u_reg_u_reg_if_N25;
 wire u_reg_u_reg_if_N26;
 wire u_reg_u_reg_if_N27;
 wire u_reg_u_reg_if_N28;
 wire u_reg_u_reg_if_N29;
 wire u_reg_u_reg_if_N30;
 wire u_reg_u_reg_if_N31;
 wire u_reg_u_reg_if_N32;
 wire u_reg_u_reg_if_N33;
 wire u_reg_u_reg_if_N34;
 wire u_reg_u_reg_if_N35;
 wire u_reg_u_reg_if_N36;
 wire u_reg_u_reg_if_N37;
 wire u_reg_u_reg_if_N38;
 wire u_reg_u_reg_if_N39;
 wire u_reg_u_reg_if_N40;
 wire u_reg_u_reg_if_N41;
 wire u_reg_u_reg_if_N42;
 wire u_reg_u_reg_if_N43;
 wire u_reg_u_reg_if_N44;
 wire u_reg_u_reg_if_N45;
 wire u_reg_u_reg_if_N46;
 wire u_reg_u_reg_if_N7;
 wire u_reg_u_reg_if_a_ack;
 wire u_reg_u_reg_if_net2113;
 wire u_reg_u_reg_if_net2119;
 wire u_reg_u_reg_if_net2124;
 wire u_reg_u_reg_if_rd_req;
 wire net1606;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire clknet_leaf_1_clk_i;
 wire clknet_leaf_2_clk_i;
 wire clknet_leaf_3_clk_i;
 wire clknet_leaf_4_clk_i;
 wire clknet_leaf_5_clk_i;
 wire clknet_leaf_6_clk_i;
 wire clknet_leaf_7_clk_i;
 wire clknet_leaf_8_clk_i;
 wire clknet_leaf_9_clk_i;
 wire clknet_leaf_10_clk_i;
 wire clknet_leaf_11_clk_i;
 wire clknet_0_clk_i;
 wire clknet_1_0__leaf_clk_i;
 wire clknet_1_1__leaf_clk_i;
 wire clknet_0_u_reg_u_reg_if_net2113;
 wire clknet_1_0__leaf_u_reg_u_reg_if_net2113;
 wire clknet_1_1__leaf_u_reg_u_reg_if_net2113;
 wire clknet_0_u_reg_u_reg_if_net2119;
 wire clknet_1_0__leaf_u_reg_u_reg_if_net2119;
 wire clknet_1_1__leaf_u_reg_u_reg_if_net2119;
 wire clknet_0_u_reg_u_reg_if_net2124;
 wire clknet_1_0__leaf_u_reg_u_reg_if_net2124;
 wire clknet_1_1__leaf_u_reg_u_reg_if_net2124;
 wire clknet_0_u_reg_u_intr_state_net2090;
 wire clknet_1_0__leaf_u_reg_u_intr_state_net2090;
 wire clknet_1_1__leaf_u_reg_u_intr_state_net2090;
 wire clknet_0_u_reg_u_intr_state_net2096;
 wire clknet_1_0__leaf_u_reg_u_intr_state_net2096;
 wire clknet_1_1__leaf_u_reg_u_intr_state_net2096;
 wire clknet_0_u_reg_u_intr_enable_net2067;
 wire clknet_1_0__leaf_u_reg_u_intr_enable_net2067;
 wire clknet_1_1__leaf_u_reg_u_intr_enable_net2067;
 wire clknet_0_u_reg_u_intr_enable_net2073;
 wire clknet_1_0__leaf_u_reg_u_intr_enable_net2073;
 wire clknet_1_1__leaf_u_reg_u_intr_enable_net2073;
 wire clknet_0_u_reg_u_intr_ctrl_en_rising_net2067;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2067;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2067;
 wire clknet_0_u_reg_u_intr_ctrl_en_rising_net2073;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2073;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2073;
 wire clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2067;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2067;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2067;
 wire clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2073;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2073;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2073;
 wire clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2067;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2067;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2067;
 wire clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2073;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2073;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2073;
 wire clknet_0_u_reg_u_intr_ctrl_en_falling_net2067;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2067;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2067;
 wire clknet_0_u_reg_u_intr_ctrl_en_falling_net2073;
 wire clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2073;
 wire clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2073;
 wire clknet_0_u_reg_u_ctrl_en_input_filter_net2067;
 wire clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2067;
 wire clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2067;
 wire clknet_0_u_reg_u_ctrl_en_input_filter_net2073;
 wire clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2073;
 wire clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2073;
 wire clknet_0_net2034;
 wire clknet_1_0__leaf_net2034;
 wire clknet_1_1__leaf_net2034;
 wire clknet_0_net2040;
 wire clknet_1_0__leaf_net2040;
 wire clknet_1_1__leaf_net2040;
 wire clknet_0_net2045;
 wire clknet_1_0__leaf_net2045;
 wire clknet_1_1__leaf_net2045;
 wire clknet_0_net2050;
 wire clknet_1_0__leaf_net2050;
 wire clknet_1_1__leaf_net2050;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire [31:0] data_in_q;
 wire [2:0] gen_alert_tx_0__u_prim_alert_sender_state_d;
 wire [2:0] gen_alert_tx_0__u_prim_alert_sender_state_q;
 wire [1:0] gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d;
 wire [1:0] gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q;
 wire [1:0] gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d;
 wire [1:0] gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q;
 wire [3:0] gen_filter_0__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_0__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_10__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_10__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_11__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_11__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_12__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_12__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_13__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_13__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_14__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_14__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_15__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_15__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_16__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_16__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_17__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_17__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_18__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_18__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_19__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_19__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_1__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_1__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_20__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_20__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_21__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_21__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_22__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_22__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_23__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_23__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_24__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_24__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_25__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_25__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_26__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_26__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_27__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_27__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_28__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_28__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_29__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_29__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_2__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_2__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_30__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_30__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_31__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_31__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_3__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_3__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_4__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_4__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_5__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_5__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_6__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_6__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_7__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_7__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_8__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_8__u_filter_diff_ctr_q;
 wire [3:0] gen_filter_9__u_filter_diff_ctr_d;
 wire [3:0] gen_filter_9__u_filter_diff_ctr_q;
 wire [31:0] u_reg_data_in_qs;
 wire [31:0] u_reg_u_ctrl_en_input_filter_wr_data;
 wire [31:0] u_reg_u_data_in_wr_data;
 wire [31:0] u_reg_u_intr_ctrl_en_falling_wr_data;
 wire [31:0] u_reg_u_intr_ctrl_en_lvlhigh_wr_data;
 wire [31:0] u_reg_u_intr_ctrl_en_lvllow_wr_data;
 wire [31:0] u_reg_u_intr_ctrl_en_rising_wr_data;
 wire [31:0] u_reg_u_intr_enable_wr_data;
 wire [31:0] u_reg_u_intr_state_wr_data;

 b15bfn000al1n02x5 U3240 (.a(net2026),
    .o(net241));
 b15bfn000an1n02x5 U3241 (.a(net2055),
    .o(net243));
 b15inv000as1n80x5 U3242 (.a(net55),
    .o1(n4067));
 b15inv000as1n80x5 U3243 (.a(net832),
    .o1(n4068));
 b15inv000as1n64x5 U3244 (.a(net831),
    .o1(n4069));
 b15and002an1n08x5 U3245 (.a(net2482),
    .b(reg2hw_intr_enable__q__9_),
    .o(intr_hw_N23));
 b15and002an1n08x5 U3246 (.a(reg2hw_intr_state__q__10_),
    .b(reg2hw_intr_enable__q__10_),
    .o(intr_hw_N22));
 b15and002an1n24x5 U3247 (.a(reg2hw_intr_state__q__2_),
    .b(reg2hw_intr_enable__q__2_),
    .o(intr_hw_N30));
 b15and002as1n08x5 U3248 (.a(reg2hw_intr_state__q__8_),
    .b(net2484),
    .o(intr_hw_N24));
 b15and002ar1n02x5 U3249 (.a(reg2hw_intr_state__q__12_),
    .b(reg2hw_intr_enable__q__12_),
    .o(intr_hw_N20));
 b15and002ah1n04x5 U3250 (.a(reg2hw_intr_state__q__26_),
    .b(reg2hw_intr_enable__q__26_),
    .o(intr_hw_N6));
 b15and002ah1n04x5 U3251 (.a(net519),
    .b(reg2hw_intr_enable__q__4_),
    .o(intr_hw_N28));
 b15and002ar1n08x5 U3252 (.a(reg2hw_intr_state__q__15_),
    .b(reg2hw_intr_enable__q__15_),
    .o(intr_hw_N17));
 b15and002al1n16x5 U3253 (.a(reg2hw_intr_state__q__3_),
    .b(reg2hw_intr_enable__q__3_),
    .o(intr_hw_N29));
 b15and002al1n16x5 U3254 (.a(net517),
    .b(reg2hw_intr_enable__q__5_),
    .o(intr_hw_N27));
 b15and002as1n08x5 U3255 (.a(net526),
    .b(net542),
    .o(intr_hw_N32));
 b15and002an1n02x5 U3256 (.a(net512),
    .b(net2519),
    .o(intr_hw_N25));
 b15and002an1n08x5 U3257 (.a(net514),
    .b(reg2hw_intr_enable__q__6_),
    .o(intr_hw_N26));
 b15and002aq1n02x5 U3258 (.a(reg2hw_intr_state__q__14_),
    .b(net536),
    .o(intr_hw_N18));
 b15and002an1n02x5 U3259 (.a(reg2hw_intr_state__q__13_),
    .b(reg2hw_intr_enable__q__13_),
    .o(intr_hw_N19));
 b15and002aq1n16x5 U3260 (.a(net524),
    .b(net541),
    .o(intr_hw_N31));
 b15and002an1n08x5 U3261 (.a(net537),
    .b(reg2hw_intr_state__q__11_),
    .o(intr_hw_N21));
 b15inv040as1n12x5 U3262 (.a(net2495),
    .o1(n3947));
 b15nonb02as1n16x5 U3263 (.a(net531),
    .b(n3947),
    .out0(intr_hw_N7));
 b15inv000as1n80x5 U3264 (.a(net830),
    .o1(n4070));
 b15inv000ah1n80x5 U3265 (.a(net829),
    .o1(n4071));
 b15inv040as1n60x5 U3266 (.a(net62),
    .o1(n4072));
 b15inv000as1n48x5 U3267 (.a(net63),
    .o1(n4073));
 b15inv000an1n80x5 U3268 (.a(net64),
    .o1(n4074));
 b15inv040as1n60x5 U3269 (.a(net65),
    .o1(n4075));
 b15inv040aq1n60x5 U3270 (.a(net66),
    .o1(n4076));
 b15inv020as1n64x5 U3271 (.a(net67),
    .o1(n4077));
 b15inv000as1n48x5 U3272 (.a(net68),
    .o1(n4078));
 b15inv040as1n48x5 U3273 (.a(net70),
    .o1(n4079));
 b15inv040as1n60x5 U3274 (.a(net71),
    .o1(n4080));
 b15inv000as1n80x5 U3275 (.a(net73),
    .o1(n4081));
 b15inv040as1n16x5 U3276 (.a(net828),
    .o1(n4082));
 b15inv000as1n24x5 U3277 (.a(net75),
    .o1(n4083));
 b15inv000as1n80x5 U3278 (.a(net826),
    .o1(n4084));
 b15inv040as1n48x5 U3279 (.a(net77),
    .o1(n4085));
 b15inv000as1n28x5 U3280 (.a(net78),
    .o1(n4086));
 b15inv020an1n16x5 U3281 (.a(net79),
    .o1(n4087));
 b15inv000as1n80x5 U3282 (.a(net80),
    .o1(n4088));
 b15inv020aq1n16x5 U3283 (.a(net823),
    .o1(n4089));
 b15inv040as1n40x5 U3284 (.a(net822),
    .o1(n4090));
 b15inv000as1n16x5 U3285 (.a(net84),
    .o1(n4091));
 b15inv000aq1n16x5 U3286 (.a(net85),
    .o1(n4092));
 b15inv000as1n20x5 U3287 (.a(net821),
    .o1(n4093));
 b15inv000as1n80x5 U3288 (.a(net87),
    .o1(n4094));
 b15inv000an1n24x5 U3289 (.a(net88),
    .o1(n4095));
 b15inv000ah1n24x5 U3290 (.a(net89),
    .o1(n4096));
 b15ztpn00an1n08x5 PHY_97 ();
 b15ztpn00an1n08x5 PHY_96 ();
 b15ztpn00an1n08x5 PHY_95 ();
 b15ztpn00an1n08x5 PHY_94 ();
 b15ztpn00an1n08x5 PHY_93 ();
 b15ztpn00an1n08x5 PHY_92 ();
 b15ztpn00an1n08x5 PHY_91 ();
 b15ztpn00an1n08x5 PHY_90 ();
 b15ztpn00an1n08x5 PHY_89 ();
 b15ztpn00an1n08x5 PHY_88 ();
 b15ztpn00an1n08x5 PHY_87 ();
 b15ztpn00an1n08x5 PHY_86 ();
 b15ztpn00an1n08x5 PHY_85 ();
 b15ztpn00an1n08x5 PHY_84 ();
 b15ztpn00an1n08x5 PHY_83 ();
 b15ztpn00an1n08x5 PHY_82 ();
 b15ztpn00an1n08x5 PHY_81 ();
 b15ztpn00an1n08x5 PHY_80 ();
 b15ztpn00an1n08x5 PHY_79 ();
 b15ztpn00an1n08x5 PHY_78 ();
 b15ztpn00an1n08x5 PHY_77 ();
 b15ztpn00an1n08x5 PHY_76 ();
 b15ztpn00an1n08x5 PHY_75 ();
 b15ztpn00an1n08x5 PHY_74 ();
 b15ztpn00an1n08x5 PHY_73 ();
 b15inv000as1n80x5 U3317 (.a(net435),
    .o1(n4123));
 b15inv000an1n24x5 U3318 (.a(net346),
    .o1(n4124));
 b15inv000ar1n24x5 U3319 (.a(net344),
    .o1(n4125));
 b15inv000as1n08x5 U3320 (.a(net350),
    .o1(n4126));
 b15inv000ar1n20x5 U3321 (.a(net351),
    .o1(n4127));
 b15inv000aq1n24x5 U3322 (.a(net353),
    .o1(n4128));
 b15inv000ar1n28x5 U3323 (.a(net357),
    .o1(n4129));
 b15inv000al1n10x5 U3324 (.a(n3497),
    .o1(n4130));
 b15inv000ar1n03x5 U3325 (.a(net1606),
    .o1(tl_o[48]));
 b15inv000ar1n03x5 U3327 (.a(net1607),
    .o1(tl_o[59]));
 b15inv000ar1n03x5 U3329 (.a(net1608),
    .o1(tl_o[60]));
 b15inv000ar1n03x5 U3331 (.a(net1609),
    .o1(tl_o[61]));
 b15ztpn00an1n08x5 PHY_72 ();
 b15ztpn00an1n08x5 PHY_71 ();
 b15ztpn00an1n08x5 PHY_70 ();
 b15ztpn00an1n08x5 PHY_69 ();
 b15ztpn00an1n08x5 PHY_68 ();
 b15inv020aq1n10x5 U3340 (.a(reg2hw_intr_state__q__17_),
    .o1(n3890));
 b15nonb02ah1n06x5 U3341 (.a(reg2hw_intr_enable__q__17_),
    .b(n3890),
    .out0(intr_hw_N15));
 b15inv000ah1n06x5 U3342 (.a(reg2hw_intr_state__q__16_),
    .o1(n3882));
 b15nonb02al1n08x5 U3343 (.a(reg2hw_intr_enable__q__16_),
    .b(n3882),
    .out0(intr_hw_N16));
 b15inv040as1n06x5 U3344 (.a(reg2hw_intr_state__q__22_),
    .o1(n3921));
 b15nonb02an1n03x5 U3345 (.a(net532),
    .b(n3921),
    .out0(intr_hw_N10));
 b15inv000an1n16x5 U3346 (.a(reg2hw_intr_state__q__19_),
    .o1(n3327));
 b15nonb02al1n08x5 U3347 (.a(reg2hw_intr_enable__q__19_),
    .b(n3327),
    .out0(intr_hw_N13));
 b15inv020ah1n04x5 U3348 (.a(reg2hw_intr_state__q__21_),
    .o1(n3912));
 b15nonb02as1n02x5 U3349 (.a(net533),
    .b(n3912),
    .out0(intr_hw_N11));
 b15qgbin1an1n05x5 U3350 (.a(reg2hw_intr_state__q__23_),
    .o1(n3932));
 b15nonb02as1n06x5 U3351 (.a(reg2hw_intr_enable__q__23_),
    .b(n3932),
    .out0(intr_hw_N9));
 b15inv040as1n03x5 U3352 (.a(reg2hw_intr_state__q__20_),
    .o1(n3904));
 b15nonb02ah1n04x5 U3353 (.a(net534),
    .b(n3904),
    .out0(intr_hw_N12));
 b15inv040an1n08x5 U3354 (.a(reg2hw_intr_state__q__24_),
    .o1(n3940));
 b15nonb02aq1n12x5 U3355 (.a(reg2hw_intr_enable__q__24_),
    .b(n3940),
    .out0(intr_hw_N8));
 b15inv000an1n06x5 U3356 (.a(reg2hw_intr_state__q__29_),
    .o1(n3984));
 b15nonb02aq1n16x5 U3357 (.a(reg2hw_intr_enable__q__29_),
    .b(n3984),
    .out0(intr_hw_N3));
 b15inv020ah1n08x5 U3358 (.a(reg2hw_intr_state__q__27_),
    .o1(n3305));
 b15nonb02ah1n08x5 U3359 (.a(reg2hw_intr_enable__q__27_),
    .b(n3305),
    .out0(intr_hw_N5));
 b15inv040as1n12x5 U3360 (.a(reg2hw_intr_state__q__28_),
    .o1(n3967));
 b15nonb02an1n03x5 U3361 (.a(reg2hw_intr_enable__q__28_),
    .b(n3967),
    .out0(intr_hw_N4));
 b15inv000as1n10x5 U3362 (.a(reg2hw_intr_state__q__31_),
    .o1(n3319));
 b15nonb02aq1n12x5 U3363 (.a(reg2hw_intr_enable__q__31_),
    .b(n3319),
    .out0(intr_hw_N1));
 b15inv000ar1n20x5 U3364 (.a(reg2hw_intr_state__q__18_),
    .o1(n3897));
 b15nonb02an1n02x5 U3365 (.a(net535),
    .b(n3897),
    .out0(intr_hw_N14));
 b15inv020ah1n08x5 U3366 (.a(reg2hw_intr_state__q__30_),
    .o1(n3312));
 b15nonb02as1n08x5 U3367 (.a(reg2hw_intr_enable__q__30_),
    .b(n3312),
    .out0(intr_hw_N2));
 b15ztpn00an1n08x5 PHY_67 ();
 b15ztpn00an1n08x5 PHY_66 ();
 b15ztpn00an1n08x5 PHY_65 ();
 b15ztpn00an1n08x5 PHY_64 ();
 b15inv000aq1n02x5 U3372 (.a(net2406),
    .o1(n2821));
 b15nand03aq1n03x5 U3373 (.a(gen_filter_5__u_filter_diff_ctr_q[0]),
    .b(gen_filter_5__u_filter_diff_ctr_q[1]),
    .c(gen_filter_5__u_filter_diff_ctr_q[2]),
    .o1(n2731));
 b15xor002aq1n08x5 U3374 (.a(net2415),
    .b(net741),
    .out0(n2819));
 b15aoi012ar1n02x5 U3375 (.a(n2819),
    .b(n2821),
    .c(net2448),
    .o1(gen_filter_5__u_filter_diff_ctr_d[3]));
 b15inv040al1n02x5 U3376 (.a(net2477),
    .o1(n2779));
 b15nandp3al1n03x5 U3377 (.a(gen_filter_14__u_filter_diff_ctr_q[0]),
    .b(gen_filter_14__u_filter_diff_ctr_q[1]),
    .c(net2462),
    .o1(n2732));
 b15xor002ar1n16x5 U3378 (.a(gen_filter_14__u_filter_filter_q),
    .b(gen_filter_14__u_filter_filter_synced),
    .out0(n2777));
 b15aoi012an1n02x5 U3379 (.a(n2777),
    .b(n2779),
    .c(n2732),
    .o1(gen_filter_14__u_filter_diff_ctr_d[3]));
 b15inv000al1n02x5 U3380 (.a(gen_filter_31__u_filter_diff_ctr_q[3]),
    .o1(n2828));
 b15nandp3ar1n03x5 U3381 (.a(gen_filter_31__u_filter_diff_ctr_q[0]),
    .b(gen_filter_31__u_filter_diff_ctr_q[1]),
    .c(net2630),
    .o1(n2737));
 b15xor002an1n16x5 U3382 (.a(gen_filter_31__u_filter_filter_q),
    .b(net746),
    .out0(n2826));
 b15aoi012ar1n02x5 U3383 (.a(n2826),
    .b(n2828),
    .c(n2737),
    .o1(gen_filter_31__u_filter_diff_ctr_d[3]));
 b15inv000ar1n03x5 U3384 (.a(gen_filter_28__u_filter_diff_ctr_q[3]),
    .o1(n2786));
 b15nandp3ah1n03x5 U3385 (.a(gen_filter_28__u_filter_diff_ctr_q[0]),
    .b(gen_filter_28__u_filter_diff_ctr_q[1]),
    .c(net2543),
    .o1(n2735));
 b15xor002an1n12x5 U3386 (.a(net2454),
    .b(gen_filter_28__u_filter_filter_synced),
    .out0(n2784));
 b15aoi012aq1n02x5 U3387 (.a(n2784),
    .b(n2786),
    .c(n2735),
    .o1(gen_filter_28__u_filter_diff_ctr_d[3]));
 b15inv000al1n02x5 U3388 (.a(gen_filter_26__u_filter_diff_ctr_q[3]),
    .o1(n2793));
 b15nand03al1n06x5 U3389 (.a(gen_filter_26__u_filter_diff_ctr_q[0]),
    .b(gen_filter_26__u_filter_diff_ctr_q[1]),
    .c(gen_filter_26__u_filter_diff_ctr_q[2]),
    .o1(n2734));
 b15xor002as1n08x5 U3390 (.a(net2479),
    .b(gen_filter_26__u_filter_filter_synced),
    .out0(n2791));
 b15aoi012as1n02x5 U3391 (.a(n2791),
    .b(n2793),
    .c(n2734),
    .o1(gen_filter_26__u_filter_diff_ctr_d[3]));
 b15inv000al1n03x5 U3392 (.a(net2633),
    .o1(n2814));
 b15nand03ah1n06x5 U3393 (.a(gen_filter_19__u_filter_diff_ctr_q[0]),
    .b(gen_filter_19__u_filter_diff_ctr_q[1]),
    .c(net2367),
    .o1(n2739));
 b15xor002as1n06x5 U3394 (.a(net2358),
    .b(gen_filter_19__u_filter_filter_synced),
    .out0(n2812));
 b15aoi012al1n02x5 U3395 (.a(n2812),
    .b(n2814),
    .c(n2739),
    .o1(gen_filter_19__u_filter_diff_ctr_d[3]));
 b15inv020an1n03x5 U3396 (.a(gen_filter_8__u_filter_diff_ctr_q[3]),
    .o1(n2765));
 b15nandp3ah1n03x5 U3397 (.a(gen_filter_8__u_filter_diff_ctr_q[0]),
    .b(gen_filter_8__u_filter_diff_ctr_q[1]),
    .c(net2492),
    .o1(n2733));
 b15xor002an1n16x5 U3398 (.a(gen_filter_8__u_filter_filter_q),
    .b(net740),
    .out0(n2763));
 b15aoi012ar1n04x5 U3399 (.a(n2763),
    .b(n2765),
    .c(n2733),
    .o1(gen_filter_8__u_filter_diff_ctr_d[3]));
 b15inv000an1n02x5 U3400 (.a(gen_filter_13__u_filter_diff_ctr_q[3]),
    .o1(n2772));
 b15nandp3al1n04x5 U3401 (.a(net2329),
    .b(gen_filter_13__u_filter_diff_ctr_q[1]),
    .c(net2363),
    .o1(n2738));
 b15xor002an1n12x5 U3402 (.a(net2378),
    .b(gen_filter_13__u_filter_filter_synced),
    .out0(n2770));
 b15aoi012an1n02x5 U3403 (.a(n2770),
    .b(n2772),
    .c(n2738),
    .o1(gen_filter_13__u_filter_diff_ctr_d[3]));
 b15inv000aq1n02x5 U3404 (.a(gen_filter_9__u_filter_diff_ctr_q[3]),
    .o1(n2800));
 b15nand03an1n06x5 U3405 (.a(gen_filter_9__u_filter_diff_ctr_q[0]),
    .b(gen_filter_9__u_filter_diff_ctr_q[1]),
    .c(gen_filter_9__u_filter_diff_ctr_q[2]),
    .o1(n2730));
 b15xor002al1n12x5 U3406 (.a(net2490),
    .b(gen_filter_9__u_filter_filter_synced),
    .out0(n2798));
 b15aoi012ah1n02x5 U3407 (.a(n2798),
    .b(n2800),
    .c(n2730),
    .o1(gen_filter_9__u_filter_diff_ctr_d[3]));
 b15inv000an1n02x5 U3408 (.a(gen_filter_0__u_filter_diff_ctr_q[3]),
    .o1(n2807));
 b15nandp3al1n04x5 U3409 (.a(gen_filter_0__u_filter_diff_ctr_q[0]),
    .b(gen_filter_0__u_filter_diff_ctr_q[1]),
    .c(gen_filter_0__u_filter_diff_ctr_q[2]),
    .o1(n2736));
 b15xor002aq1n08x5 U3410 (.a(net2386),
    .b(gen_filter_0__u_filter_filter_synced),
    .out0(n2805));
 b15aoi012ar1n02x5 U3411 (.a(n2805),
    .b(net2413),
    .c(n2736),
    .o1(gen_filter_0__u_filter_diff_ctr_d[3]));
 b15xor002aq1n16x5 U3412 (.a(net752),
    .b(net2379),
    .out0(n2706));
 b15and002ah1n02x5 U3413 (.a(net2334),
    .b(net2383),
    .o(n2704));
 b15nandp3al1n04x5 U3414 (.a(net2334),
    .b(gen_filter_22__u_filter_diff_ctr_q[1]),
    .c(gen_filter_22__u_filter_diff_ctr_q[2]),
    .o1(n2684));
 b15oai022ar1n02x5 U3415 (.a(n2704),
    .b(gen_filter_22__u_filter_diff_ctr_q[2]),
    .c(gen_filter_22__u_filter_diff_ctr_q[3]),
    .d(net2335),
    .o1(n2683));
 b15norp02ar1n02x5 U3416 (.a(net2380),
    .b(net2384),
    .o1(gen_filter_22__u_filter_diff_ctr_d[2]));
 b15and003aq1n03x5 U3417 (.a(gen_filter_25__u_filter_diff_ctr_q[0]),
    .b(gen_filter_25__u_filter_diff_ctr_q[1]),
    .c(net2432),
    .o(n2719));
 b15inv000as1n06x5 U3418 (.a(net748),
    .o1(n3490));
 b15xor002aq1n08x5 U3419 (.a(n3490),
    .b(gen_filter_25__u_filter_filter_q),
    .out0(n2717));
 b15inv040aq1n04x5 U3420 (.a(n2717),
    .o1(n2748));
 b15oab012ar1n02x5 U3421 (.a(n2748),
    .b(gen_filter_25__u_filter_diff_ctr_q[3]),
    .c(n2719),
    .out0(gen_filter_25__u_filter_diff_ctr_d[3]));
 b15nand03an1n08x5 U3422 (.a(gen_filter_22__u_filter_diff_ctr_q[3]),
    .b(gen_filter_22__u_filter_diff_ctr_q[1]),
    .c(gen_filter_22__u_filter_diff_ctr_q[2]),
    .o1(n2705));
 b15aoi012ar1n02x5 U3423 (.a(n2706),
    .b(net2334),
    .c(n2705),
    .o1(gen_filter_22__u_filter_diff_ctr_d[0]));
 b15inv000al1n02x5 U3424 (.a(gen_filter_22__u_filter_diff_ctr_q[3]),
    .o1(n2685));
 b15aoi012ar1n02x5 U3425 (.a(n2706),
    .b(n2685),
    .c(net2335),
    .o1(gen_filter_22__u_filter_diff_ctr_d[3]));
 b15and003aq1n04x5 U3426 (.a(gen_filter_16__u_filter_diff_ctr_q[0]),
    .b(gen_filter_16__u_filter_diff_ctr_q[1]),
    .c(net2331),
    .o(n2855));
 b15xor002an1n16x5 U3427 (.a(net2427),
    .b(gen_filter_16__u_filter_filter_synced),
    .out0(n2856));
 b15oab012al1n02x5 U3428 (.a(n2856),
    .b(net2368),
    .c(n2855),
    .out0(gen_filter_16__u_filter_diff_ctr_d[3]));
 b15and003ah1n03x5 U3429 (.a(gen_filter_2__u_filter_diff_ctr_q[0]),
    .b(net2396),
    .c(net2512),
    .o(n2839));
 b15xor002an1n16x5 U3430 (.a(gen_filter_2__u_filter_filter_q),
    .b(gen_filter_2__u_filter_filter_synced),
    .out0(n2840));
 b15oab012ar1n02x5 U3431 (.a(n2840),
    .b(net2404),
    .c(n2839),
    .out0(gen_filter_2__u_filter_diff_ctr_d[3]));
 b15and003al1n04x5 U3432 (.a(gen_filter_11__u_filter_diff_ctr_q[0]),
    .b(gen_filter_11__u_filter_diff_ctr_q[1]),
    .c(gen_filter_11__u_filter_diff_ctr_q[2]),
    .o(n2847));
 b15xor002as1n06x5 U3433 (.a(net2372),
    .b(gen_filter_11__u_filter_filter_synced),
    .out0(n2848));
 b15oab012ar1n02x5 U3434 (.a(n2848),
    .b(gen_filter_11__u_filter_diff_ctr_q[3]),
    .c(n2847),
    .out0(gen_filter_11__u_filter_diff_ctr_d[3]));
 b15and003ah1n04x5 U3435 (.a(gen_filter_27__u_filter_diff_ctr_q[0]),
    .b(gen_filter_27__u_filter_diff_ctr_q[1]),
    .c(gen_filter_27__u_filter_diff_ctr_q[2]),
    .o(n2831));
 b15xor002ah1n16x5 U3436 (.a(net2449),
    .b(gen_filter_27__u_filter_filter_synced),
    .out0(n2832));
 b15oab012ar1n02x5 U3437 (.a(n2832),
    .b(net2440),
    .c(n2831),
    .out0(gen_filter_27__u_filter_diff_ctr_d[3]));
 b15and003aq1n03x5 U3438 (.a(gen_filter_12__u_filter_diff_ctr_q[0]),
    .b(gen_filter_12__u_filter_diff_ctr_q[1]),
    .c(net2637),
    .o(n2863));
 b15xor002ah1n08x5 U3439 (.a(net2326),
    .b(gen_filter_12__u_filter_filter_synced),
    .out0(n2864));
 b15oab012al1n02x5 U3440 (.a(net2327),
    .b(net2344),
    .c(n2863),
    .out0(gen_filter_12__u_filter_diff_ctr_d[3]));
 b15and003ah1n03x5 U3441 (.a(net2476),
    .b(gen_filter_30__u_filter_diff_ctr_q[0]),
    .c(gen_filter_30__u_filter_diff_ctr_q[1]),
    .o(n2949));
 b15xor002as1n08x5 U3442 (.a(net2365),
    .b(gen_filter_30__u_filter_filter_synced),
    .out0(n2952));
 b15oab012al1n03x5 U3443 (.a(n2952),
    .b(net2409),
    .c(n2949),
    .out0(gen_filter_30__u_filter_diff_ctr_d[3]));
 b15and003ar1n03x5 U3444 (.a(net2487),
    .b(gen_filter_1__u_filter_diff_ctr_q[0]),
    .c(gen_filter_1__u_filter_diff_ctr_q[1]),
    .o(n2943));
 b15xor002al1n12x5 U3445 (.a(gen_filter_1__u_filter_filter_q),
    .b(gen_filter_1__u_filter_filter_synced),
    .out0(n2946));
 b15oab012ar1n02x5 U3446 (.a(n2946),
    .b(net2424),
    .c(n2943),
    .out0(gen_filter_1__u_filter_diff_ctr_d[3]));
 b15and003al1n04x5 U3447 (.a(gen_filter_4__u_filter_diff_ctr_q[0]),
    .b(gen_filter_4__u_filter_diff_ctr_q[1]),
    .c(net2503),
    .o(n2750));
 b15xor002as1n12x5 U3448 (.a(gen_filter_4__u_filter_filter_synced),
    .b(net2531),
    .out0(n2752));
 b15oab012al1n04x5 U3449 (.a(n2752),
    .b(gen_filter_4__u_filter_diff_ctr_q[3]),
    .c(n2750),
    .out0(gen_filter_4__u_filter_diff_ctr_d[3]));
 b15and003ar1n04x5 U3450 (.a(net2391),
    .b(gen_filter_29__u_filter_diff_ctr_q[1]),
    .c(gen_filter_29__u_filter_diff_ctr_q[2]),
    .o(n2713));
 b15xor002as1n08x5 U3451 (.a(net747),
    .b(net2410),
    .out0(n2755));
 b15oab012ar1n02x5 U3452 (.a(n2755),
    .b(net2442),
    .c(n2713),
    .out0(gen_filter_29__u_filter_diff_ctr_d[3]));
 b15and003aq1n04x5 U3453 (.a(net2375),
    .b(gen_filter_23__u_filter_diff_ctr_q[0]),
    .c(gen_filter_23__u_filter_diff_ctr_q[1]),
    .o(n2729));
 b15xor002ah1n12x5 U3454 (.a(net749),
    .b(net2528),
    .out0(n2913));
 b15oab012ar1n02x5 U3455 (.a(n2913),
    .b(gen_filter_23__u_filter_diff_ctr_q[3]),
    .c(n2729),
    .out0(gen_filter_23__u_filter_diff_ctr_d[3]));
 b15and003ah1n02x5 U3456 (.a(net2452),
    .b(gen_filter_20__u_filter_diff_ctr_q[0]),
    .c(gen_filter_20__u_filter_diff_ctr_q[1]),
    .o(n2725));
 b15xor002an1n16x5 U3457 (.a(net754),
    .b(gen_filter_20__u_filter_filter_q),
    .out0(n2919));
 b15oab012ar1n02x5 U3458 (.a(n2919),
    .b(net2435),
    .c(n2725),
    .out0(gen_filter_20__u_filter_diff_ctr_d[3]));
 b15and003al1n04x5 U3459 (.a(gen_filter_15__u_filter_diff_ctr_q[0]),
    .b(gen_filter_15__u_filter_diff_ctr_q[1]),
    .c(net2515),
    .o(n2712));
 b15inv000ah1n10x5 U3460 (.a(gen_filter_15__u_filter_filter_synced),
    .o1(n3540));
 b15xor002aq1n08x5 U3461 (.a(n3540),
    .b(gen_filter_15__u_filter_filter_q),
    .out0(n2710));
 b15inv000aq1n06x5 U3462 (.a(n2710),
    .o1(n2925));
 b15oab012ar1n04x5 U3463 (.a(n2925),
    .b(gen_filter_15__u_filter_diff_ctr_q[3]),
    .c(n2712),
    .out0(gen_filter_15__u_filter_diff_ctr_d[3]));
 b15and003ah1n03x5 U3464 (.a(gen_filter_21__u_filter_diff_ctr_q[0]),
    .b(gen_filter_21__u_filter_diff_ctr_q[1]),
    .c(net2467),
    .o(n2709));
 b15inv040as1n08x5 U3465 (.a(gen_filter_21__u_filter_filter_synced),
    .o1(n3619));
 b15xor002ah1n06x5 U3466 (.a(n3619),
    .b(net2527),
    .out0(n2707));
 b15inv000al1n04x5 U3467 (.a(n2707),
    .o1(n2931));
 b15oab012ah1n02x5 U3468 (.a(n2931),
    .b(net2552),
    .c(n2709),
    .out0(gen_filter_21__u_filter_diff_ctr_d[3]));
 b15inv000aq1n08x5 U3469 (.a(net2400),
    .o1(n2893));
 b15nandp3al1n12x5 U3470 (.o1(n2891),
    .a(gen_filter_6__u_filter_diff_ctr_q[0]),
    .b(gen_filter_6__u_filter_diff_ctr_q[1]),
    .c(gen_filter_6__u_filter_diff_ctr_q[2]));
 b15xor002as1n08x5 U3471 (.a(gen_filter_6__u_filter_filter_synced),
    .b(net2398),
    .out0(n2890));
 b15aoi012ar1n06x5 U3472 (.a(n2890),
    .b(n2893),
    .c(n2891),
    .o1(gen_filter_6__u_filter_diff_ctr_d[3]));
 b15inv000ah1n05x5 U3473 (.a(gen_filter_4__u_filter_diff_ctr_q[3]),
    .o1(n3993));
 b15aoi012an1n08x5 U3474 (.a(net2503),
    .b(gen_filter_4__u_filter_diff_ctr_q[1]),
    .c(gen_filter_4__u_filter_diff_ctr_q[0]),
    .o1(n3994));
 b15aoi112al1n03x5 U3475 (.a(n2752),
    .b(n3994),
    .c(n2750),
    .d(n3993),
    .o1(gen_filter_4__u_filter_diff_ctr_d[2]));
 b15inv020aq1n10x5 U3476 (.a(net2360),
    .o1(n2905));
 b15nandp3as1n08x5 U3477 (.a(gen_filter_17__u_filter_diff_ctr_q[0]),
    .b(gen_filter_17__u_filter_diff_ctr_q[1]),
    .c(net2388),
    .o1(n2903));
 b15xor002as1n08x5 U3478 (.a(gen_filter_17__u_filter_filter_synced),
    .b(net2351),
    .out0(n2902));
 b15aoi012an1n02x5 U3479 (.a(n2902),
    .b(n2905),
    .c(net2389),
    .o1(gen_filter_17__u_filter_diff_ctr_d[3]));
 b15inv020ah1n12x5 U3480 (.a(net2546),
    .o1(n2875));
 b15nand03aq1n16x5 U3481 (.a(gen_filter_7__u_filter_diff_ctr_q[0]),
    .b(gen_filter_7__u_filter_diff_ctr_q[1]),
    .c(gen_filter_7__u_filter_diff_ctr_q[2]),
    .o1(n2873));
 b15xor002al1n16x5 U3482 (.a(gen_filter_7__u_filter_filter_synced),
    .b(net2537),
    .out0(n2872));
 b15aoi012al1n04x5 U3483 (.a(n2872),
    .b(n2875),
    .c(n2873),
    .o1(gen_filter_7__u_filter_diff_ctr_d[3]));
 b15inv020ah1n10x5 U3484 (.a(net2323),
    .o1(n2911));
 b15nand03al1n16x5 U3485 (.a(gen_filter_24__u_filter_diff_ctr_q[0]),
    .b(gen_filter_24__u_filter_diff_ctr_q[1]),
    .c(gen_filter_24__u_filter_diff_ctr_q[2]),
    .o1(n2909));
 b15xor002an1n16x5 U3486 (.a(gen_filter_24__u_filter_filter_synced),
    .b(net2319),
    .out0(n2908));
 b15aoi012ah1n02x5 U3487 (.a(n2908),
    .b(n2911),
    .c(n2909),
    .o1(gen_filter_24__u_filter_diff_ctr_d[3]));
 b15inv040al1n10x5 U3488 (.a(net2511),
    .o1(n2887));
 b15nandp3an1n16x5 U3489 (.a(gen_filter_3__u_filter_diff_ctr_q[0]),
    .b(gen_filter_3__u_filter_diff_ctr_q[1]),
    .c(gen_filter_3__u_filter_diff_ctr_q[2]),
    .o1(n2885));
 b15xor002as1n12x5 U3490 (.a(net744),
    .b(net2485),
    .out0(n2884));
 b15aoi012ar1n06x5 U3491 (.a(n2884),
    .b(n2887),
    .c(n2885),
    .o1(gen_filter_3__u_filter_diff_ctr_d[3]));
 b15inv000al1n10x5 U3492 (.a(net2393),
    .o1(n2881));
 b15nandp3ar1n16x5 U3493 (.a(gen_filter_10__u_filter_diff_ctr_q[0]),
    .b(gen_filter_10__u_filter_diff_ctr_q[1]),
    .c(gen_filter_10__u_filter_diff_ctr_q[2]),
    .o1(n2879));
 b15xor002as1n16x5 U3494 (.a(gen_filter_10__u_filter_filter_synced),
    .b(gen_filter_10__u_filter_filter_q),
    .out0(n2878));
 b15aoi012ar1n02x5 U3495 (.a(n2878),
    .b(n2881),
    .c(n2879),
    .o1(gen_filter_10__u_filter_diff_ctr_d[3]));
 b15inv040an1n05x5 U3496 (.a(net2353),
    .o1(n2899));
 b15nandp3ar1n12x5 U3497 (.o1(n2897),
    .a(gen_filter_18__u_filter_diff_ctr_q[0]),
    .b(gen_filter_18__u_filter_diff_ctr_q[1]),
    .c(gen_filter_18__u_filter_diff_ctr_q[2]));
 b15xor002aq1n16x5 U3498 (.a(gen_filter_18__u_filter_filter_synced),
    .b(gen_filter_18__u_filter_filter_q),
    .out0(n2896));
 b15aoi012ar1n02x5 U3499 (.a(n2896),
    .b(n2899),
    .c(n2897),
    .o1(gen_filter_18__u_filter_diff_ctr_d[3]));
 b15inv000al1n02x5 U3500 (.a(gen_filter_29__u_filter_diff_ctr_q[3]),
    .o1(n2687));
 b15aoi012al1n02x5 U3501 (.a(gen_filter_29__u_filter_diff_ctr_q[2]),
    .b(gen_filter_29__u_filter_diff_ctr_q[1]),
    .c(net2391),
    .o1(n2686));
 b15aoi112aq1n02x5 U3502 (.a(n2755),
    .b(n2686),
    .c(n2713),
    .d(n2687),
    .o1(gen_filter_29__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3503 (.a(n2879),
    .o1(n2689));
 b15aoi012al1n02x5 U3504 (.a(gen_filter_10__u_filter_diff_ctr_q[2]),
    .b(gen_filter_10__u_filter_diff_ctr_q[1]),
    .c(gen_filter_10__u_filter_diff_ctr_q[0]),
    .o1(n2688));
 b15aoi112ah1n03x5 U3505 (.a(n2688),
    .b(n2878),
    .c(n2689),
    .d(n2881),
    .o1(gen_filter_10__u_filter_diff_ctr_d[2]));
 b15inv000aq1n02x5 U3506 (.a(n2909),
    .o1(n2691));
 b15aoi012as1n02x5 U3507 (.a(gen_filter_24__u_filter_diff_ctr_q[2]),
    .b(gen_filter_24__u_filter_diff_ctr_q[1]),
    .c(gen_filter_24__u_filter_diff_ctr_q[0]),
    .o1(n2690));
 b15aoi112ar1n06x5 U3508 (.a(n2690),
    .b(n2908),
    .c(n2691),
    .d(n2911),
    .o1(gen_filter_24__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3509 (.a(n2891),
    .o1(n2693));
 b15aoi012ar1n02x5 U3510 (.a(net2417),
    .b(gen_filter_6__u_filter_diff_ctr_q[1]),
    .c(gen_filter_6__u_filter_diff_ctr_q[0]),
    .o1(n2692));
 b15aoi112an1n02x5 U3511 (.a(net2418),
    .b(n2890),
    .c(n2693),
    .d(n2893),
    .o1(gen_filter_6__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3512 (.a(n2903),
    .o1(n2695));
 b15aoi012ah1n02x5 U3513 (.a(gen_filter_17__u_filter_diff_ctr_q[2]),
    .b(gen_filter_17__u_filter_diff_ctr_q[1]),
    .c(gen_filter_17__u_filter_diff_ctr_q[0]),
    .o1(n2694));
 b15aoi112ah1n04x5 U3514 (.a(n2694),
    .b(n2902),
    .c(n2695),
    .d(n2905),
    .o1(gen_filter_17__u_filter_diff_ctr_d[2]));
 b15inv000an1n02x5 U3515 (.a(n2873),
    .o1(n2697));
 b15aoi012as1n02x5 U3516 (.a(net2556),
    .b(net2558),
    .c(gen_filter_7__u_filter_diff_ctr_q[0]),
    .o1(n2696));
 b15aoi112an1n04x5 U3517 (.a(n2696),
    .b(n2872),
    .c(n2697),
    .d(n2875),
    .o1(gen_filter_7__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3518 (.a(n2897),
    .o1(n2699));
 b15aoi012ar1n02x5 U3519 (.a(gen_filter_18__u_filter_diff_ctr_q[2]),
    .b(gen_filter_18__u_filter_diff_ctr_q[1]),
    .c(gen_filter_18__u_filter_diff_ctr_q[0]),
    .o1(n2698));
 b15aoi112al1n02x5 U3520 (.a(n2698),
    .b(n2896),
    .c(n2699),
    .d(n2899),
    .o1(gen_filter_18__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3521 (.a(n2885),
    .o1(n2701));
 b15aoi012al1n02x5 U3522 (.a(gen_filter_3__u_filter_diff_ctr_q[2]),
    .b(gen_filter_3__u_filter_diff_ctr_q[1]),
    .c(gen_filter_3__u_filter_diff_ctr_q[0]),
    .o1(n2700));
 b15aoi112aq1n03x5 U3523 (.a(n2700),
    .b(n2884),
    .c(n2701),
    .d(n2887),
    .o1(gen_filter_3__u_filter_diff_ctr_d[2]));
 b15nandp2al1n02x5 U3524 (.a(gen_filter_22__u_filter_diff_ctr_q[3]),
    .b(gen_filter_22__u_filter_diff_ctr_q[2]),
    .o1(n2703));
 b15norp02ar1n02x5 U3525 (.a(net2510),
    .b(gen_filter_22__u_filter_diff_ctr_q[1]),
    .o1(n2702));
 b15aoi112al1n02x5 U3526 (.a(n2706),
    .b(n2702),
    .c(n2704),
    .d(n2703),
    .o1(gen_filter_22__u_filter_diff_ctr_d[1]));
 b15norp02ar1n08x5 U3527 (.a(n2706),
    .b(n2705),
    .o1(eq_x_71_n25));
 b15inv020ar1n04x5 U3528 (.a(net2381),
    .o1(n2846));
 b15aoi012aq1n04x5 U3529 (.a(net2566),
    .b(gen_filter_11__u_filter_diff_ctr_q[1]),
    .c(gen_filter_11__u_filter_diff_ctr_q[0]),
    .o1(n2853));
 b15aoi112as1n02x5 U3530 (.a(n2853),
    .b(n2848),
    .c(n2847),
    .d(n2846),
    .o1(gen_filter_11__u_filter_diff_ctr_d[2]));
 b15inv000an1n02x5 U3531 (.a(gen_filter_12__u_filter_diff_ctr_q[3]),
    .o1(n2862));
 b15aoi012aq1n04x5 U3532 (.a(net2551),
    .b(gen_filter_12__u_filter_diff_ctr_q[1]),
    .c(gen_filter_12__u_filter_diff_ctr_q[0]),
    .o1(n2869));
 b15aoi112as1n02x5 U3533 (.a(n2869),
    .b(net2327),
    .c(n2863),
    .d(n2862),
    .o1(gen_filter_12__u_filter_diff_ctr_d[2]));
 b15inv020ah1n03x5 U3534 (.a(net2368),
    .o1(n2854));
 b15aoi012as1n04x5 U3535 (.a(net2331),
    .b(gen_filter_16__u_filter_diff_ctr_q[1]),
    .c(gen_filter_16__u_filter_diff_ctr_q[0]),
    .o1(n2861));
 b15aoi112ar1n04x5 U3536 (.a(net2332),
    .b(n2856),
    .c(n2855),
    .d(n2854),
    .o1(gen_filter_16__u_filter_diff_ctr_d[2]));
 b15inv020ah1n03x5 U3537 (.a(net2404),
    .o1(n2838));
 b15aoi012aq1n06x5 U3538 (.a(net2512),
    .b(gen_filter_2__u_filter_diff_ctr_q[1]),
    .c(gen_filter_2__u_filter_diff_ctr_q[0]),
    .o1(n2845));
 b15aoi112ar1n04x5 U3539 (.a(net2513),
    .b(n2840),
    .c(n2839),
    .d(n2838),
    .o1(gen_filter_2__u_filter_diff_ctr_d[2]));
 b15inv040aq1n03x5 U3540 (.a(net2440),
    .o1(n2830));
 b15aoi012ar1n08x5 U3541 (.a(gen_filter_27__u_filter_diff_ctr_q[2]),
    .b(gen_filter_27__u_filter_diff_ctr_q[1]),
    .c(gen_filter_27__u_filter_diff_ctr_q[0]),
    .o1(n2837));
 b15aoi112an1n04x5 U3542 (.a(n2837),
    .b(n2832),
    .c(n2831),
    .d(n2830),
    .o1(gen_filter_27__u_filter_diff_ctr_d[2]));
 b15nandp2as1n05x5 U3543 (.a(net2435),
    .b(n2725),
    .o1(n2923));
 b15aoi012an1n02x5 U3544 (.a(n2919),
    .b(net2420),
    .c(n2923),
    .o1(gen_filter_20__u_filter_diff_ctr_d[0]));
 b15nandp2as1n08x5 U3545 (.a(gen_filter_23__u_filter_diff_ctr_q[3]),
    .b(n2729),
    .o1(n2917));
 b15aoi012aq1n12x5 U3546 (.a(n2913),
    .b(gen_filter_23__u_filter_diff_ctr_q[0]),
    .c(n2917),
    .o1(gen_filter_23__u_filter_diff_ctr_d[0]));
 b15nand02ah1n08x5 U3547 (.a(gen_filter_15__u_filter_diff_ctr_q[3]),
    .b(n2712),
    .o1(n2929));
 b15aoi012al1n02x5 U3548 (.a(n2925),
    .b(gen_filter_15__u_filter_diff_ctr_q[0]),
    .c(n2929),
    .o1(gen_filter_15__u_filter_diff_ctr_d[0]));
 b15nand02al1n08x5 U3549 (.a(gen_filter_21__u_filter_diff_ctr_q[3]),
    .b(n2709),
    .o1(n2935));
 b15aoi012aq1n04x5 U3550 (.a(n2931),
    .b(gen_filter_21__u_filter_diff_ctr_q[0]),
    .c(n2935),
    .o1(gen_filter_21__u_filter_diff_ctr_d[0]));
 b15inv000al1n02x5 U3551 (.a(gen_filter_21__u_filter_diff_ctr_q[3]),
    .o1(n2708));
 b15aoai13an1n06x5 U3552 (.a(n2707),
    .b(net2467),
    .c(gen_filter_21__u_filter_diff_ctr_q[1]),
    .d(gen_filter_21__u_filter_diff_ctr_q[0]),
    .o1(n2934));
 b15aoi012al1n02x5 U3553 (.a(n2934),
    .b(net2468),
    .c(n2708),
    .o1(gen_filter_21__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3554 (.a(gen_filter_15__u_filter_diff_ctr_q[3]),
    .o1(n2711));
 b15aoai13an1n08x5 U3555 (.a(n2710),
    .b(net2515),
    .c(gen_filter_15__u_filter_diff_ctr_q[1]),
    .d(gen_filter_15__u_filter_diff_ctr_q[0]),
    .o1(n2928));
 b15aoi012an1n02x5 U3556 (.a(n2928),
    .b(n2712),
    .c(n2711),
    .o1(gen_filter_15__u_filter_diff_ctr_d[2]));
 b15nand02ar1n02x5 U3557 (.a(net2639),
    .b(gen_filter_29__u_filter_diff_ctr_q[1]),
    .o1(n2715));
 b15nand02aq1n04x5 U3558 (.a(gen_filter_29__u_filter_diff_ctr_q[3]),
    .b(n2713),
    .o1(n2756));
 b15inv000al1n02x5 U3559 (.a(n2756),
    .o1(n2714));
 b15oaoi13ar1n02x3 U3560 (.a(n2714),
    .b(n2715),
    .c(gen_filter_29__u_filter_diff_ctr_q[0]),
    .d(gen_filter_29__u_filter_diff_ctr_q[1]),
    .o1(n2716));
 b15norp02ar1n03x5 U3561 (.a(n2716),
    .b(n2755),
    .o1(gen_filter_29__u_filter_diff_ctr_d[1]));
 b15inv000al1n02x5 U3562 (.a(gen_filter_25__u_filter_diff_ctr_q[3]),
    .o1(n2718));
 b15aoai13ah1n06x5 U3563 (.a(n2717),
    .b(net2432),
    .c(gen_filter_25__u_filter_diff_ctr_q[1]),
    .d(gen_filter_25__u_filter_diff_ctr_q[0]),
    .o1(n3995));
 b15aoi012ar1n02x5 U3564 (.a(net2433),
    .b(n2719),
    .c(n2718),
    .o1(gen_filter_25__u_filter_diff_ctr_d[2]));
 b15inv040ar1n06x5 U3565 (.a(net2082),
    .o1(net237));
 b15nand02as1n16x5 U3566 (.a(net44),
    .b(net237),
    .o1(n2744));
 b15aob012an1n04x5 U3567 (.a(n2744),
    .b(net2081),
    .c(net38),
    .out0(u_reg_u_reg_if_N7));
 b15nand02al1n02x5 U3568 (.a(gen_filter_25__u_filter_diff_ctr_q[0]),
    .b(gen_filter_25__u_filter_diff_ctr_q[1]),
    .o1(n2721));
 b15nand02al1n06x5 U3569 (.a(gen_filter_25__u_filter_diff_ctr_q[3]),
    .b(n2719),
    .o1(n2749));
 b15inv000al1n02x5 U3570 (.a(n2749),
    .o1(n2720));
 b15oaoi13an1n04x5 U3571 (.a(n2720),
    .b(n2721),
    .c(gen_filter_25__u_filter_diff_ctr_q[0]),
    .d(gen_filter_25__u_filter_diff_ctr_q[1]),
    .o1(n3996));
 b15norp02ar1n03x5 U3572 (.a(n2748),
    .b(n3996),
    .o1(gen_filter_25__u_filter_diff_ctr_d[1]));
 b15inv000al1n02x5 U3573 (.a(gen_filter_20__u_filter_diff_ctr_q[2]),
    .o1(n2722));
 b15nandp2ah1n02x5 U3574 (.a(gen_filter_20__u_filter_diff_ctr_q[0]),
    .b(gen_filter_20__u_filter_diff_ctr_q[1]),
    .o1(n2918));
 b15aoi012an1n02x5 U3575 (.a(n2919),
    .b(n2722),
    .c(n2918),
    .o1(n2723));
 b15inv000al1n02x5 U3576 (.a(n2723),
    .o1(n2724));
 b15nandp2aq1n04x5 U3577 (.a(n2723),
    .b(net2435),
    .o1(n2922));
 b15oai012ar1n02x5 U3578 (.a(n2922),
    .b(net2453),
    .c(n2724),
    .o1(gen_filter_20__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3579 (.a(net2375),
    .o1(n2726));
 b15nand02aq1n04x5 U3580 (.a(gen_filter_23__u_filter_diff_ctr_q[0]),
    .b(gen_filter_23__u_filter_diff_ctr_q[1]),
    .o1(n2912));
 b15aoi012as1n02x5 U3581 (.a(n2913),
    .b(n2726),
    .c(n2912),
    .o1(n2727));
 b15inv000al1n02x5 U3582 (.a(n2727),
    .o1(n2728));
 b15nand02as1n06x5 U3583 (.a(n2727),
    .b(gen_filter_23__u_filter_diff_ctr_q[3]),
    .o1(n2916));
 b15oai012as1n02x5 U3584 (.a(n2916),
    .b(net2376),
    .c(n2728),
    .o1(gen_filter_23__u_filter_diff_ctr_d[2]));
 b15inv000as1n03x5 U3585 (.a(n2798),
    .o1(n2795));
 b15aoai13ar1n04x5 U3586 (.a(n2795),
    .b(gen_filter_9__u_filter_diff_ctr_q[2]),
    .c(gen_filter_9__u_filter_diff_ctr_q[1]),
    .d(gen_filter_9__u_filter_diff_ctr_q[0]),
    .o1(n2799));
 b15oab012ar1n02x5 U3587 (.a(n2799),
    .b(gen_filter_9__u_filter_diff_ctr_q[3]),
    .c(n2730),
    .out0(gen_filter_9__u_filter_diff_ctr_d[2]));
 b15inv000an1n04x5 U3588 (.a(n2819),
    .o1(n2816));
 b15aoai13ar1n06x5 U3589 (.a(n2816),
    .b(net2447),
    .c(gen_filter_5__u_filter_diff_ctr_q[1]),
    .d(gen_filter_5__u_filter_diff_ctr_q[0]),
    .o1(n2820));
 b15oab012ar1n02x5 U3590 (.a(n2820),
    .b(net2406),
    .c(net2448),
    .out0(gen_filter_5__u_filter_diff_ctr_d[2]));
 b15inv000ar1n05x5 U3591 (.a(n2777),
    .o1(n2774));
 b15aoai13as1n03x5 U3592 (.a(n2774),
    .b(net2462),
    .c(gen_filter_14__u_filter_diff_ctr_q[1]),
    .d(gen_filter_14__u_filter_diff_ctr_q[0]),
    .o1(n2778));
 b15oab012al1n02x5 U3593 (.a(n2778),
    .b(net2477),
    .c(n2732),
    .out0(gen_filter_14__u_filter_diff_ctr_d[2]));
 b15inv040aq1n03x5 U3594 (.a(n2763),
    .o1(n2760));
 b15aoai13as1n02x5 U3595 (.a(n2760),
    .b(net2492),
    .c(gen_filter_8__u_filter_diff_ctr_q[1]),
    .d(gen_filter_8__u_filter_diff_ctr_q[0]),
    .o1(n2764));
 b15oab012an1n03x5 U3596 (.a(n2764),
    .b(net2534),
    .c(n2733),
    .out0(gen_filter_8__u_filter_diff_ctr_d[2]));
 b15inv000ar1n05x5 U3597 (.a(n2791),
    .o1(n2788));
 b15aoai13ah1n03x5 U3598 (.a(n2788),
    .b(gen_filter_26__u_filter_diff_ctr_q[2]),
    .c(gen_filter_26__u_filter_diff_ctr_q[1]),
    .d(gen_filter_26__u_filter_diff_ctr_q[0]),
    .o1(n2792));
 b15oab012an1n02x5 U3599 (.a(n2792),
    .b(net2522),
    .c(n2734),
    .out0(gen_filter_26__u_filter_diff_ctr_d[2]));
 b15inv020ah1n03x5 U3600 (.a(n2784),
    .o1(n2781));
 b15aoai13ar1n04x5 U3601 (.a(n2781),
    .b(net2543),
    .c(gen_filter_28__u_filter_diff_ctr_q[1]),
    .d(gen_filter_28__u_filter_diff_ctr_q[0]),
    .o1(n2785));
 b15oab012ar1n02x5 U3602 (.a(n2785),
    .b(net2550),
    .c(n2735),
    .out0(gen_filter_28__u_filter_diff_ctr_d[2]));
 b15inv040al1n04x5 U3603 (.a(n2805),
    .o1(n2802));
 b15aoai13al1n06x5 U3604 (.a(n2802),
    .b(gen_filter_0__u_filter_diff_ctr_q[2]),
    .c(gen_filter_0__u_filter_diff_ctr_q[1]),
    .d(gen_filter_0__u_filter_diff_ctr_q[0]),
    .o1(n2806));
 b15oab012as1n02x5 U3605 (.a(n2806),
    .b(net2412),
    .c(net2507),
    .out0(gen_filter_0__u_filter_diff_ctr_d[2]));
 b15inv040ah1n04x5 U3606 (.a(n2826),
    .o1(n2823));
 b15aoai13ah1n02x5 U3607 (.a(n2823),
    .b(net2535),
    .c(gen_filter_31__u_filter_diff_ctr_q[1]),
    .d(gen_filter_31__u_filter_diff_ctr_q[0]),
    .o1(n2827));
 b15oab012ar1n02x5 U3608 (.a(n2827),
    .b(gen_filter_31__u_filter_diff_ctr_q[3]),
    .c(n2737),
    .out0(gen_filter_31__u_filter_diff_ctr_d[2]));
 b15inv040as1n02x5 U3609 (.a(n2770),
    .o1(n2767));
 b15aoai13al1n03x5 U3610 (.a(n2767),
    .b(net2363),
    .c(gen_filter_13__u_filter_diff_ctr_q[1]),
    .d(net2329),
    .o1(n2771));
 b15oab012aq1n02x5 U3611 (.a(n2771),
    .b(gen_filter_13__u_filter_diff_ctr_q[3]),
    .c(n2738),
    .out0(gen_filter_13__u_filter_diff_ctr_d[2]));
 b15inv000ah1n03x5 U3612 (.a(n2812),
    .o1(n2809));
 b15aoai13ah1n03x5 U3613 (.a(n2809),
    .b(net2367),
    .c(gen_filter_19__u_filter_diff_ctr_q[1]),
    .d(gen_filter_19__u_filter_diff_ctr_q[0]),
    .o1(n2813));
 b15oab012ar1n02x5 U3614 (.a(n2813),
    .b(net2474),
    .c(n2739),
    .out0(gen_filter_19__u_filter_diff_ctr_d[2]));
 b15inv040an1n06x5 U3615 (.a(net2041),
    .o1(n2936));
 b15inv000as1n03x5 U3616 (.a(net2012),
    .o1(n2937));
 b15aoi022al1n06x5 U3617 (.a(net2012),
    .b(net2007),
    .c(n2936),
    .d(n2937),
    .o1(net239));
 b15nor002an1n03x5 U3618 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .b(net2489),
    .o1(n2743));
 b15inv000al1n02x5 U3619 (.a(n2743),
    .o1(n2741));
 b15nandp3an1n02x5 U3620 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq),
    .c(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq),
    .o1(n2740));
 b15oai013ar1n06x5 U3621 (.a(n2740),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq),
    .c(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq),
    .d(n2741),
    .o1(n2742));
 b15nor003ar1n06x5 U3622 (.a(net2317),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[1]),
    .c(n2742),
    .o1(n2964));
 b15aoi012an1n08x5 U3623 (.a(n2743),
    .b(net2374),
    .c(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .o1(n2965));
 b15nonb02ar1n02x3 U3624 (.a(n2964),
    .b(n2965),
    .out0(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[0]));
 b15inv000as1n48x5 U3625 (.a(n2744),
    .o1(u_reg_u_reg_if_a_ack));
 b15qgbin1an1n15x5 U3626 (.a(net2054),
    .o1(n2938));
 b15nor002as1n08x5 U3627 (.a(net409),
    .b(n2938),
    .o1(n1429));
 b15norp02ar1n02x5 U3628 (.a(u_reg_u_reg_if_a_ack),
    .b(n2936),
    .o1(n1432));
 b15inv040as1n05x5 U3629 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd),
    .o1(n2746));
 b15inv000aq1n12x5 U3630 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd),
    .o1(n2747));
 b15aoi022an1n16x5 U3631 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd),
    .c(n2746),
    .d(n2747),
    .o1(n2967));
 b15nanb02al1n12x5 U3632 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .b(n2967),
    .out0(n2973));
 b15nandp2ar1n02x5 U3633 (.a(n2973),
    .b(net2394),
    .o1(n2745));
 b15oai012al1n04x5 U3634 (.a(n2745),
    .b(n2973),
    .c(n2747),
    .o1(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_n3));
 b15xor002ar1n16x5 U3635 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq),
    .b(n2746),
    .out0(n2972));
 b15xor002an1n12x5 U3636 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq),
    .b(n2747),
    .out0(n2971));
 b15aoi112al1n06x5 U3637 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[0]),
    .c(n2972),
    .d(n2971),
    .o1(n2966));
 b15nonb02al1n02x5 U3638 (.a(n2966),
    .b(n2967),
    .out0(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[0]));
 b15aoi012as1n04x5 U3639 (.a(n2748),
    .b(net2509),
    .c(n2749),
    .o1(gen_filter_25__u_filter_diff_ctr_d[0]));
 b15nand02al1n08x5 U3640 (.a(gen_filter_4__u_filter_diff_ctr_q[3]),
    .b(n2750),
    .o1(n2754));
 b15aoi012aq1n06x5 U3641 (.a(n2752),
    .b(gen_filter_4__u_filter_diff_ctr_q[0]),
    .c(n2754),
    .o1(gen_filter_4__u_filter_diff_ctr_d[0]));
 b15nand02al1n02x5 U3642 (.a(gen_filter_4__u_filter_diff_ctr_q[0]),
    .b(gen_filter_4__u_filter_diff_ctr_q[1]),
    .o1(n2751));
 b15oai012al1n06x5 U3643 (.a(n2751),
    .b(gen_filter_4__u_filter_diff_ctr_q[0]),
    .c(gen_filter_4__u_filter_diff_ctr_q[1]),
    .o1(n2753));
 b15aoi012al1n08x5 U3644 (.a(n2752),
    .b(n2754),
    .c(n2753),
    .o1(gen_filter_4__u_filter_diff_ctr_d[1]));
 b15aoi012as1n04x5 U3645 (.a(n2755),
    .b(net2391),
    .c(n2756),
    .o1(gen_filter_29__u_filter_diff_ctr_d[0]));
 b15nandp3ah1n02x5 U3646 (.a(net2471),
    .b(gen_filter_29__u_filter_diff_ctr_q[2]),
    .c(gen_filter_29__u_filter_diff_ctr_q[3]),
    .o1(n2757));
 b15nonb02as1n04x5 U3647 (.a(gen_filter_29__u_filter_diff_ctr_d[0]),
    .b(net2472),
    .out0(eq_x_36_n25));
 b15inv020ar1n04x5 U3648 (.a(n2952),
    .o1(n2948));
 b15aoai13as1n04x5 U3649 (.a(n2948),
    .b(net2476),
    .c(gen_filter_30__u_filter_diff_ctr_q[0]),
    .d(gen_filter_30__u_filter_diff_ctr_q[1]),
    .o1(n2758));
 b15nonb02al1n06x5 U3650 (.a(gen_filter_30__u_filter_diff_ctr_q[3]),
    .b(n2758),
    .out0(n2953));
 b15oabi12an1n03x5 U3651 (.a(n2953),
    .b(n2949),
    .c(n2758),
    .out0(gen_filter_30__u_filter_diff_ctr_d[2]));
 b15inv000al1n02x5 U3652 (.a(n2946),
    .o1(n2942));
 b15aoai13ar1n03x5 U3653 (.a(n2942),
    .b(net2487),
    .c(gen_filter_1__u_filter_diff_ctr_q[0]),
    .d(gen_filter_1__u_filter_diff_ctr_q[1]),
    .o1(n2759));
 b15nonb02ah1n02x5 U3654 (.a(net2424),
    .b(n2759),
    .out0(n2947));
 b15oabi12aq1n02x5 U3655 (.a(n2947),
    .b(n2943),
    .c(n2759),
    .out0(gen_filter_1__u_filter_diff_ctr_d[2]));
 b15oai012aq1n04x5 U3656 (.a(n2760),
    .b(gen_filter_8__u_filter_diff_ctr_q[0]),
    .c(gen_filter_8__u_filter_diff_ctr_q[1]),
    .o1(n2761));
 b15nand04ah1n08x5 U3657 (.a(gen_filter_8__u_filter_diff_ctr_q[1]),
    .b(gen_filter_8__u_filter_diff_ctr_q[3]),
    .c(net2492),
    .d(n2760),
    .o1(n2762));
 b15aoai13as1n06x5 U3658 (.a(net2493),
    .b(n2761),
    .c(gen_filter_8__u_filter_diff_ctr_q[1]),
    .d(gen_filter_8__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_8__u_filter_diff_ctr_d[1]));
 b15oai012ar1n12x5 U3659 (.a(net2493),
    .b(gen_filter_8__u_filter_diff_ctr_q[0]),
    .c(n2763),
    .o1(gen_filter_8__u_filter_diff_ctr_d[0]));
 b15nor002aq1n02x5 U3660 (.a(n2765),
    .b(n2764),
    .o1(n2766));
 b15and003ah1n03x5 U3661 (.a(n2766),
    .b(gen_filter_8__u_filter_diff_ctr_d[1]),
    .c(gen_filter_8__u_filter_diff_ctr_d[0]),
    .o(eq_x_141_n25));
 b15oai012ah1n02x5 U3662 (.a(n2767),
    .b(net2329),
    .c(gen_filter_13__u_filter_diff_ctr_q[1]),
    .o1(n2768));
 b15nand04as1n06x5 U3663 (.a(gen_filter_13__u_filter_diff_ctr_q[1]),
    .b(gen_filter_13__u_filter_diff_ctr_q[3]),
    .c(gen_filter_13__u_filter_diff_ctr_q[2]),
    .d(n2767),
    .o1(n2769));
 b15aoai13an1n06x5 U3664 (.a(n2769),
    .b(n2768),
    .c(gen_filter_13__u_filter_diff_ctr_q[1]),
    .d(net2329),
    .o1(gen_filter_13__u_filter_diff_ctr_d[1]));
 b15oai012an1n08x5 U3665 (.a(n2769),
    .b(net2627),
    .c(n2770),
    .o1(gen_filter_13__u_filter_diff_ctr_d[0]));
 b15norp02al1n02x5 U3666 (.a(n2772),
    .b(n2771),
    .o1(n2773));
 b15and003al1n04x5 U3667 (.a(n2773),
    .b(gen_filter_13__u_filter_diff_ctr_d[1]),
    .c(gen_filter_13__u_filter_diff_ctr_d[0]),
    .o(eq_x_116_n25));
 b15oai012an1n04x5 U3668 (.a(n2774),
    .b(gen_filter_14__u_filter_diff_ctr_q[0]),
    .c(gen_filter_14__u_filter_diff_ctr_q[1]),
    .o1(n2775));
 b15nand04aq1n08x5 U3669 (.a(gen_filter_14__u_filter_diff_ctr_q[1]),
    .b(gen_filter_14__u_filter_diff_ctr_q[3]),
    .c(net2462),
    .d(n2774),
    .o1(n2776));
 b15aoai13al1n08x5 U3670 (.a(net2463),
    .b(n2775),
    .c(gen_filter_14__u_filter_diff_ctr_q[1]),
    .d(gen_filter_14__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_14__u_filter_diff_ctr_d[1]));
 b15oai012ah1n06x5 U3671 (.a(net2463),
    .b(gen_filter_14__u_filter_diff_ctr_q[0]),
    .c(n2777),
    .o1(gen_filter_14__u_filter_diff_ctr_d[0]));
 b15norp02ar1n02x5 U3672 (.a(n2779),
    .b(n2778),
    .o1(n2780));
 b15and003aq1n04x5 U3673 (.a(n2780),
    .b(gen_filter_14__u_filter_diff_ctr_d[1]),
    .c(gen_filter_14__u_filter_diff_ctr_d[0]),
    .o(eq_x_111_n25));
 b15oai012ar1n02x5 U3674 (.a(n2781),
    .b(gen_filter_28__u_filter_diff_ctr_q[0]),
    .c(gen_filter_28__u_filter_diff_ctr_q[1]),
    .o1(n2782));
 b15nand04as1n06x5 U3675 (.a(gen_filter_28__u_filter_diff_ctr_q[1]),
    .b(gen_filter_28__u_filter_diff_ctr_q[3]),
    .c(net2543),
    .d(n2781),
    .o1(n2783));
 b15aoai13ar1n03x5 U3676 (.a(net2544),
    .b(n2782),
    .c(gen_filter_28__u_filter_diff_ctr_q[1]),
    .d(gen_filter_28__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_28__u_filter_diff_ctr_d[1]));
 b15oai012aq1n12x5 U3677 (.a(net2544),
    .b(gen_filter_28__u_filter_diff_ctr_q[0]),
    .c(n2784),
    .o1(gen_filter_28__u_filter_diff_ctr_d[0]));
 b15norp02aq1n02x5 U3678 (.a(n2786),
    .b(n2785),
    .o1(n2787));
 b15and003al1n04x5 U3679 (.a(n2787),
    .b(gen_filter_28__u_filter_diff_ctr_d[1]),
    .c(gen_filter_28__u_filter_diff_ctr_d[0]),
    .o(eq_x_41_n25));
 b15oai012as1n02x5 U3680 (.a(n2788),
    .b(gen_filter_26__u_filter_diff_ctr_q[0]),
    .c(gen_filter_26__u_filter_diff_ctr_q[1]),
    .o1(n2789));
 b15nand04ah1n06x5 U3681 (.a(gen_filter_26__u_filter_diff_ctr_q[1]),
    .b(net2522),
    .c(gen_filter_26__u_filter_diff_ctr_q[2]),
    .d(n2788),
    .o1(n2790));
 b15aoai13al1n06x5 U3682 (.a(net2523),
    .b(n2789),
    .c(gen_filter_26__u_filter_diff_ctr_q[1]),
    .d(gen_filter_26__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_26__u_filter_diff_ctr_d[1]));
 b15oai012ar1n06x5 U3683 (.a(net2523),
    .b(net2553),
    .c(n2791),
    .o1(gen_filter_26__u_filter_diff_ctr_d[0]));
 b15norp02ar1n02x5 U3684 (.a(n2793),
    .b(n2792),
    .o1(n2794));
 b15and003al1n04x5 U3685 (.a(n2794),
    .b(gen_filter_26__u_filter_diff_ctr_d[1]),
    .c(gen_filter_26__u_filter_diff_ctr_d[0]),
    .o(eq_x_51_n25));
 b15oai012al1n02x5 U3686 (.a(n2795),
    .b(gen_filter_9__u_filter_diff_ctr_q[0]),
    .c(gen_filter_9__u_filter_diff_ctr_q[1]),
    .o1(n2796));
 b15nand04ar1n12x5 U3687 (.a(gen_filter_9__u_filter_diff_ctr_q[1]),
    .b(gen_filter_9__u_filter_diff_ctr_q[3]),
    .c(gen_filter_9__u_filter_diff_ctr_q[2]),
    .d(n2795),
    .o1(n2797));
 b15aoai13al1n04x5 U3688 (.a(n2797),
    .b(n2796),
    .c(gen_filter_9__u_filter_diff_ctr_q[1]),
    .d(gen_filter_9__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_9__u_filter_diff_ctr_d[1]));
 b15oai012aq1n08x5 U3689 (.a(n2797),
    .b(gen_filter_9__u_filter_diff_ctr_q[0]),
    .c(n2798),
    .o1(gen_filter_9__u_filter_diff_ctr_d[0]));
 b15norp02al1n02x5 U3690 (.a(n2800),
    .b(n2799),
    .o1(n2801));
 b15and003an1n04x5 U3691 (.a(n2801),
    .b(gen_filter_9__u_filter_diff_ctr_d[1]),
    .c(gen_filter_9__u_filter_diff_ctr_d[0]),
    .o(eq_x_136_n25));
 b15oai012an1n04x5 U3692 (.a(n2802),
    .b(gen_filter_0__u_filter_diff_ctr_q[0]),
    .c(gen_filter_0__u_filter_diff_ctr_q[1]),
    .o1(n2803));
 b15nand04ah1n08x5 U3693 (.a(gen_filter_0__u_filter_diff_ctr_q[1]),
    .b(net2412),
    .c(net2506),
    .d(n2802),
    .o1(n2804));
 b15aoai13al1n08x5 U3694 (.a(n2804),
    .b(n2803),
    .c(gen_filter_0__u_filter_diff_ctr_q[1]),
    .d(gen_filter_0__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_0__u_filter_diff_ctr_d[1]));
 b15oai012ah1n06x5 U3695 (.a(n2804),
    .b(gen_filter_0__u_filter_diff_ctr_q[0]),
    .c(n2805),
    .o1(gen_filter_0__u_filter_diff_ctr_d[0]));
 b15nor002ar1n03x5 U3696 (.a(n2807),
    .b(n2806),
    .o1(n2808));
 b15and003aq1n04x5 U3697 (.a(n2808),
    .b(gen_filter_0__u_filter_diff_ctr_d[1]),
    .c(gen_filter_0__u_filter_diff_ctr_d[0]),
    .o(eq_x_181_n25));
 b15oai012ah1n03x5 U3698 (.a(n2809),
    .b(gen_filter_19__u_filter_diff_ctr_q[0]),
    .c(gen_filter_19__u_filter_diff_ctr_q[1]),
    .o1(n2810));
 b15nand04an1n08x5 U3699 (.a(gen_filter_19__u_filter_diff_ctr_q[1]),
    .b(net2474),
    .c(net2367),
    .d(n2809),
    .o1(n2811));
 b15aoai13ah1n06x5 U3700 (.a(n2811),
    .b(n2810),
    .c(gen_filter_19__u_filter_diff_ctr_q[1]),
    .d(gen_filter_19__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_19__u_filter_diff_ctr_d[1]));
 b15oai012ah1n04x5 U3701 (.a(n2811),
    .b(gen_filter_19__u_filter_diff_ctr_q[0]),
    .c(n2812),
    .o1(gen_filter_19__u_filter_diff_ctr_d[0]));
 b15norp02an1n02x5 U3702 (.a(n2814),
    .b(n2813),
    .o1(n2815));
 b15and003aq1n03x5 U3703 (.a(n2815),
    .b(gen_filter_19__u_filter_diff_ctr_d[1]),
    .c(gen_filter_19__u_filter_diff_ctr_d[0]),
    .o(eq_x_86_n25));
 b15oai012aq1n02x5 U3704 (.a(n2816),
    .b(gen_filter_5__u_filter_diff_ctr_q[0]),
    .c(gen_filter_5__u_filter_diff_ctr_q[1]),
    .o1(n2817));
 b15nand04an1n08x5 U3705 (.a(gen_filter_5__u_filter_diff_ctr_q[1]),
    .b(net2406),
    .c(gen_filter_5__u_filter_diff_ctr_q[2]),
    .d(n2816),
    .o1(n2818));
 b15aoai13as1n04x5 U3706 (.a(net2407),
    .b(n2817),
    .c(gen_filter_5__u_filter_diff_ctr_q[1]),
    .d(gen_filter_5__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_5__u_filter_diff_ctr_d[1]));
 b15oai012ah1n06x5 U3707 (.a(net2407),
    .b(gen_filter_5__u_filter_diff_ctr_q[0]),
    .c(n2819),
    .o1(gen_filter_5__u_filter_diff_ctr_d[0]));
 b15nor002ah1n02x5 U3708 (.a(n2821),
    .b(n2820),
    .o1(n2822));
 b15and003an1n12x5 U3709 (.a(n2822),
    .b(gen_filter_5__u_filter_diff_ctr_d[1]),
    .c(gen_filter_5__u_filter_diff_ctr_d[0]),
    .o(eq_x_156_n25));
 b15oai012an1n04x5 U3710 (.a(n2823),
    .b(gen_filter_31__u_filter_diff_ctr_q[0]),
    .c(gen_filter_31__u_filter_diff_ctr_q[1]),
    .o1(n2824));
 b15nand04ah1n12x5 U3711 (.a(gen_filter_31__u_filter_diff_ctr_q[1]),
    .b(net2561),
    .c(net2535),
    .d(n2823),
    .o1(n2825));
 b15aoai13al1n08x5 U3712 (.a(n2825),
    .b(n2824),
    .c(gen_filter_31__u_filter_diff_ctr_q[1]),
    .d(gen_filter_31__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_31__u_filter_diff_ctr_d[1]));
 b15oai012ar1n12x5 U3713 (.a(n2825),
    .b(gen_filter_31__u_filter_diff_ctr_q[0]),
    .c(n2826),
    .o1(gen_filter_31__u_filter_diff_ctr_d[0]));
 b15nor002as1n02x5 U3714 (.a(n2828),
    .b(n2827),
    .o1(n2829));
 b15and003as1n04x5 U3715 (.a(n2829),
    .b(gen_filter_31__u_filter_diff_ctr_d[1]),
    .c(gen_filter_31__u_filter_diff_ctr_d[0]),
    .o(eq_x_26_n25));
 b15norp02an1n04x5 U3716 (.a(n2830),
    .b(n2832),
    .o1(n2835));
 b15nandp2ah1n03x5 U3717 (.a(n2835),
    .b(n2831),
    .o1(n2833));
 b15oai012aq1n06x5 U3718 (.a(n2833),
    .b(net2526),
    .c(n2832),
    .o1(gen_filter_27__u_filter_diff_ctr_d[0]));
 b15oabi12an1n02x5 U3719 (.a(n2832),
    .b(gen_filter_27__u_filter_diff_ctr_q[0]),
    .c(gen_filter_27__u_filter_diff_ctr_q[1]),
    .out0(n2834));
 b15aoai13as1n04x5 U3720 (.a(n2833),
    .b(n2834),
    .c(net2458),
    .d(gen_filter_27__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_27__u_filter_diff_ctr_d[1]));
 b15nand03ar1n06x5 U3721 (.a(n2835),
    .b(gen_filter_27__u_filter_diff_ctr_d[0]),
    .c(gen_filter_27__u_filter_diff_ctr_d[1]),
    .o1(n2836));
 b15nor002an1n04x5 U3722 (.a(n2837),
    .b(n2836),
    .o1(eq_x_46_n25));
 b15norp02aq1n03x5 U3723 (.a(n2838),
    .b(n2840),
    .o1(n2843));
 b15nand02ah1n03x5 U3724 (.a(n2843),
    .b(n2839),
    .o1(n2841));
 b15oai012ah1n03x5 U3725 (.a(n2841),
    .b(net2430),
    .c(n2840),
    .o1(gen_filter_2__u_filter_diff_ctr_d[0]));
 b15oabi12al1n02x5 U3726 (.a(n2840),
    .b(gen_filter_2__u_filter_diff_ctr_q[0]),
    .c(gen_filter_2__u_filter_diff_ctr_q[1]),
    .out0(n2842));
 b15aoai13ah1n03x5 U3727 (.a(n2841),
    .b(n2842),
    .c(net2396),
    .d(gen_filter_2__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_2__u_filter_diff_ctr_d[1]));
 b15nandp3aq1n04x5 U3728 (.a(n2843),
    .b(gen_filter_2__u_filter_diff_ctr_d[0]),
    .c(gen_filter_2__u_filter_diff_ctr_d[1]),
    .o1(n2844));
 b15norp02al1n12x5 U3729 (.a(n2845),
    .b(n2844),
    .o1(eq_x_171_n25));
 b15norp02aq1n03x5 U3730 (.a(n2846),
    .b(n2848),
    .o1(n2851));
 b15nandp2al1n03x5 U3731 (.a(n2851),
    .b(n2847),
    .o1(n2849));
 b15oai012aq1n04x5 U3732 (.a(n2849),
    .b(net2426),
    .c(n2848),
    .o1(gen_filter_11__u_filter_diff_ctr_d[0]));
 b15oabi12ar1n04x5 U3733 (.a(n2848),
    .b(gen_filter_11__u_filter_diff_ctr_q[0]),
    .c(gen_filter_11__u_filter_diff_ctr_q[1]),
    .out0(n2850));
 b15aoai13ar1n06x5 U3734 (.a(n2849),
    .b(n2850),
    .c(net2554),
    .d(gen_filter_11__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_11__u_filter_diff_ctr_d[1]));
 b15nandp3al1n04x5 U3735 (.a(n2851),
    .b(gen_filter_11__u_filter_diff_ctr_d[0]),
    .c(gen_filter_11__u_filter_diff_ctr_d[1]),
    .o1(n2852));
 b15nor002ar1n06x5 U3736 (.a(n2853),
    .b(n2852),
    .o1(eq_x_126_n25));
 b15norp02an1n03x5 U3737 (.a(n2854),
    .b(n2856),
    .o1(n2859));
 b15nandp2al1n04x5 U3738 (.a(n2859),
    .b(n2855),
    .o1(n2857));
 b15oai012ah1n06x5 U3739 (.a(n2857),
    .b(net2517),
    .c(n2856),
    .o1(gen_filter_16__u_filter_diff_ctr_d[0]));
 b15oabi12al1n02x5 U3740 (.a(n2856),
    .b(gen_filter_16__u_filter_diff_ctr_q[0]),
    .c(gen_filter_16__u_filter_diff_ctr_q[1]),
    .out0(n2858));
 b15aoai13aq1n04x5 U3741 (.a(n2857),
    .b(n2858),
    .c(net2460),
    .d(gen_filter_16__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_16__u_filter_diff_ctr_d[1]));
 b15nand03ah1n04x5 U3742 (.a(n2859),
    .b(gen_filter_16__u_filter_diff_ctr_d[0]),
    .c(gen_filter_16__u_filter_diff_ctr_d[1]),
    .o1(n2860));
 b15nor002al1n06x5 U3743 (.a(net2332),
    .b(n2860),
    .o1(eq_x_101_n25));
 b15nor002an1n03x5 U3744 (.a(n2862),
    .b(n2864),
    .o1(n2867));
 b15nandp2aq1n04x5 U3745 (.a(n2867),
    .b(n2863),
    .o1(n2865));
 b15oai012al1n06x5 U3746 (.a(n2865),
    .b(net2350),
    .c(net2327),
    .o1(gen_filter_12__u_filter_diff_ctr_d[0]));
 b15oabi12ar1n03x5 U3747 (.a(n2864),
    .b(gen_filter_12__u_filter_diff_ctr_q[0]),
    .c(gen_filter_12__u_filter_diff_ctr_q[1]),
    .out0(n2866));
 b15aoai13ah1n04x5 U3748 (.a(n2865),
    .b(n2866),
    .c(net2497),
    .d(net2350),
    .o1(gen_filter_12__u_filter_diff_ctr_d[1]));
 b15nandp3al1n03x5 U3749 (.a(n2867),
    .b(gen_filter_12__u_filter_diff_ctr_d[0]),
    .c(gen_filter_12__u_filter_diff_ctr_d[1]),
    .o1(n2868));
 b15norp02aq1n03x5 U3750 (.a(n2869),
    .b(n2868),
    .o1(eq_x_121_n25));
 b15nand02al1n02x5 U3751 (.a(gen_filter_7__u_filter_diff_ctr_q[0]),
    .b(gen_filter_7__u_filter_diff_ctr_q[1]),
    .o1(n2870));
 b15oai012ar1n06x5 U3752 (.a(n2870),
    .b(gen_filter_7__u_filter_diff_ctr_q[0]),
    .c(gen_filter_7__u_filter_diff_ctr_q[1]),
    .o1(n2871));
 b15oaoi13as1n04x5 U3753 (.a(n2872),
    .b(n2871),
    .c(n2875),
    .d(n2873),
    .o1(gen_filter_7__u_filter_diff_ctr_d[1]));
 b15oaoi13al1n08x5 U3754 (.a(n2872),
    .b(gen_filter_7__u_filter_diff_ctr_q[0]),
    .c(n2875),
    .d(n2873),
    .o1(gen_filter_7__u_filter_diff_ctr_d[0]));
 b15nand03ar1n06x5 U3755 (.a(gen_filter_7__u_filter_diff_ctr_q[2]),
    .b(gen_filter_7__u_filter_diff_ctr_d[1]),
    .c(gen_filter_7__u_filter_diff_ctr_d[0]),
    .o1(n2874));
 b15nor002as1n04x5 U3756 (.a(n2875),
    .b(n2874),
    .o1(eq_x_146_n25));
 b15nand02ar1n02x5 U3757 (.a(gen_filter_10__u_filter_diff_ctr_q[0]),
    .b(gen_filter_10__u_filter_diff_ctr_q[1]),
    .o1(n2876));
 b15oai012ah1n03x5 U3758 (.a(n2876),
    .b(gen_filter_10__u_filter_diff_ctr_q[0]),
    .c(gen_filter_10__u_filter_diff_ctr_q[1]),
    .o1(n2877));
 b15oaoi13al1n08x5 U3759 (.a(n2878),
    .b(n2877),
    .c(n2881),
    .d(n2879),
    .o1(gen_filter_10__u_filter_diff_ctr_d[1]));
 b15oaoi13al1n04x5 U3760 (.a(n2878),
    .b(gen_filter_10__u_filter_diff_ctr_q[0]),
    .c(n2881),
    .d(n2879),
    .o1(gen_filter_10__u_filter_diff_ctr_d[0]));
 b15nandp3ar1n04x5 U3761 (.a(gen_filter_10__u_filter_diff_ctr_q[2]),
    .b(gen_filter_10__u_filter_diff_ctr_d[1]),
    .c(gen_filter_10__u_filter_diff_ctr_d[0]),
    .o1(n2880));
 b15norp02al1n08x5 U3762 (.a(n2881),
    .b(n2880),
    .o1(eq_x_131_n25));
 b15nandp2al1n02x5 U3763 (.a(gen_filter_3__u_filter_diff_ctr_q[0]),
    .b(gen_filter_3__u_filter_diff_ctr_q[1]),
    .o1(n2882));
 b15oai012ar1n06x5 U3764 (.a(n2882),
    .b(gen_filter_3__u_filter_diff_ctr_q[0]),
    .c(gen_filter_3__u_filter_diff_ctr_q[1]),
    .o1(n2883));
 b15oaoi13ah1n04x5 U3765 (.a(n2884),
    .b(n2883),
    .c(n2887),
    .d(n2885),
    .o1(gen_filter_3__u_filter_diff_ctr_d[1]));
 b15oaoi13an1n08x5 U3766 (.a(n2884),
    .b(gen_filter_3__u_filter_diff_ctr_q[0]),
    .c(n2887),
    .d(n2885),
    .o1(gen_filter_3__u_filter_diff_ctr_d[0]));
 b15nandp3ar1n02x5 U3767 (.a(gen_filter_3__u_filter_diff_ctr_q[2]),
    .b(gen_filter_3__u_filter_diff_ctr_d[1]),
    .c(gen_filter_3__u_filter_diff_ctr_d[0]),
    .o1(n2886));
 b15norp02ar1n03x5 U3768 (.a(n2887),
    .b(n2886),
    .o1(eq_x_166_n25));
 b15nand02ar1n02x5 U3769 (.a(gen_filter_6__u_filter_diff_ctr_q[0]),
    .b(gen_filter_6__u_filter_diff_ctr_q[1]),
    .o1(n2888));
 b15oai012an1n02x5 U3770 (.a(n2888),
    .b(gen_filter_6__u_filter_diff_ctr_q[0]),
    .c(gen_filter_6__u_filter_diff_ctr_q[1]),
    .o1(n2889));
 b15oaoi13ar1n04x5 U3771 (.a(n2890),
    .b(n2889),
    .c(n2893),
    .d(n2891),
    .o1(gen_filter_6__u_filter_diff_ctr_d[1]));
 b15oaoi13aq1n04x5 U3772 (.a(n2890),
    .b(gen_filter_6__u_filter_diff_ctr_q[0]),
    .c(n2893),
    .d(n2891),
    .o1(gen_filter_6__u_filter_diff_ctr_d[0]));
 b15nand03ah1n03x5 U3773 (.a(gen_filter_6__u_filter_diff_ctr_q[2]),
    .b(gen_filter_6__u_filter_diff_ctr_d[1]),
    .c(gen_filter_6__u_filter_diff_ctr_d[0]),
    .o1(n2892));
 b15norp02al1n02x5 U3774 (.a(n2893),
    .b(n2892),
    .o1(eq_x_151_n25));
 b15nand02ar1n02x5 U3775 (.a(gen_filter_18__u_filter_diff_ctr_q[0]),
    .b(gen_filter_18__u_filter_diff_ctr_q[1]),
    .o1(n2894));
 b15oai012al1n02x5 U3776 (.a(n2894),
    .b(gen_filter_18__u_filter_diff_ctr_q[0]),
    .c(gen_filter_18__u_filter_diff_ctr_q[1]),
    .o1(n2895));
 b15oaoi13ah1n03x5 U3777 (.a(n2896),
    .b(n2895),
    .c(n2899),
    .d(n2897),
    .o1(gen_filter_18__u_filter_diff_ctr_d[1]));
 b15oaoi13ah1n03x5 U3778 (.a(n2896),
    .b(net2357),
    .c(n2899),
    .d(n2897),
    .o1(gen_filter_18__u_filter_diff_ctr_d[0]));
 b15nand03al1n02x5 U3779 (.a(gen_filter_18__u_filter_diff_ctr_q[2]),
    .b(gen_filter_18__u_filter_diff_ctr_d[1]),
    .c(gen_filter_18__u_filter_diff_ctr_d[0]),
    .o1(n2898));
 b15norp02ar1n03x5 U3780 (.a(n2899),
    .b(n2898),
    .o1(eq_x_91_n25));
 b15nand02ar1n02x5 U3781 (.a(gen_filter_17__u_filter_diff_ctr_q[0]),
    .b(gen_filter_17__u_filter_diff_ctr_q[1]),
    .o1(n2900));
 b15oai012an1n03x5 U3782 (.a(n2900),
    .b(gen_filter_17__u_filter_diff_ctr_q[0]),
    .c(gen_filter_17__u_filter_diff_ctr_q[1]),
    .o1(n2901));
 b15oaoi13ah1n04x5 U3783 (.a(n2902),
    .b(n2901),
    .c(n2905),
    .d(n2903),
    .o1(gen_filter_17__u_filter_diff_ctr_d[1]));
 b15oaoi13as1n04x5 U3784 (.a(n2902),
    .b(net2473),
    .c(n2905),
    .d(n2903),
    .o1(gen_filter_17__u_filter_diff_ctr_d[0]));
 b15nand03aq1n03x5 U3785 (.a(gen_filter_17__u_filter_diff_ctr_q[2]),
    .b(gen_filter_17__u_filter_diff_ctr_d[1]),
    .c(gen_filter_17__u_filter_diff_ctr_d[0]),
    .o1(n2904));
 b15nor002an1n04x5 U3786 (.a(n2905),
    .b(n2904),
    .o1(eq_x_96_n25));
 b15nand02ar1n02x5 U3787 (.a(gen_filter_24__u_filter_diff_ctr_q[0]),
    .b(gen_filter_24__u_filter_diff_ctr_q[1]),
    .o1(n2906));
 b15oai012an1n04x5 U3788 (.a(n2906),
    .b(gen_filter_24__u_filter_diff_ctr_q[0]),
    .c(gen_filter_24__u_filter_diff_ctr_q[1]),
    .o1(n2907));
 b15oaoi13aq1n04x5 U3789 (.a(n2908),
    .b(n2907),
    .c(n2911),
    .d(n2909),
    .o1(gen_filter_24__u_filter_diff_ctr_d[1]));
 b15oaoi13ah1n08x5 U3790 (.a(n2908),
    .b(gen_filter_24__u_filter_diff_ctr_q[0]),
    .c(n2911),
    .d(n2909),
    .o1(gen_filter_24__u_filter_diff_ctr_d[0]));
 b15nandp3ar1n03x5 U3791 (.a(gen_filter_24__u_filter_diff_ctr_q[2]),
    .b(gen_filter_24__u_filter_diff_ctr_d[1]),
    .c(gen_filter_24__u_filter_diff_ctr_d[0]),
    .o1(n2910));
 b15nor002an1n04x5 U3792 (.a(n2911),
    .b(n2910),
    .o1(eq_x_61_n25));
 b15oai012an1n03x5 U3793 (.a(n2912),
    .b(gen_filter_23__u_filter_diff_ctr_q[0]),
    .c(gen_filter_23__u_filter_diff_ctr_q[1]),
    .o1(n2914));
 b15aoi012an1n04x5 U3794 (.a(n2913),
    .b(n2917),
    .c(n2914),
    .o1(gen_filter_23__u_filter_diff_ctr_d[1]));
 b15inv020ah1n03x5 U3795 (.a(gen_filter_23__u_filter_diff_ctr_d[1]),
    .o1(n2915));
 b15aoi112as1n08x5 U3796 (.a(n2916),
    .b(n2915),
    .c(gen_filter_23__u_filter_diff_ctr_q[0]),
    .d(n2917),
    .o1(eq_x_66_n25));
 b15oai012an1n04x5 U3797 (.a(n2918),
    .b(gen_filter_20__u_filter_diff_ctr_q[0]),
    .c(gen_filter_20__u_filter_diff_ctr_q[1]),
    .o1(n2920));
 b15aoi012ar1n06x5 U3798 (.a(n2919),
    .b(net2436),
    .c(n2920),
    .o1(gen_filter_20__u_filter_diff_ctr_d[1]));
 b15inv040ar1n02x5 U3799 (.a(gen_filter_20__u_filter_diff_ctr_d[1]),
    .o1(n2921));
 b15aoi112ah1n04x5 U3800 (.a(n2922),
    .b(n2921),
    .c(net2420),
    .d(n2923),
    .o1(eq_x_81_n25));
 b15nand02ar1n02x5 U3801 (.a(gen_filter_15__u_filter_diff_ctr_q[0]),
    .b(gen_filter_15__u_filter_diff_ctr_q[1]),
    .o1(n2924));
 b15oai012al1n03x5 U3802 (.a(n2924),
    .b(gen_filter_15__u_filter_diff_ctr_q[0]),
    .c(gen_filter_15__u_filter_diff_ctr_q[1]),
    .o1(n2926));
 b15aoi012aq1n04x5 U3803 (.a(n2925),
    .b(n2929),
    .c(n2926),
    .o1(gen_filter_15__u_filter_diff_ctr_d[1]));
 b15nandp2al1n04x5 U3804 (.a(gen_filter_15__u_filter_diff_ctr_q[3]),
    .b(gen_filter_15__u_filter_diff_ctr_d[1]),
    .o1(n2927));
 b15aoi112as1n08x5 U3805 (.a(n2928),
    .b(n2927),
    .c(gen_filter_15__u_filter_diff_ctr_q[0]),
    .d(n2929),
    .o1(eq_x_106_n25));
 b15nand02ar1n02x5 U3806 (.a(gen_filter_21__u_filter_diff_ctr_q[0]),
    .b(gen_filter_21__u_filter_diff_ctr_q[1]),
    .o1(n2930));
 b15oai012ah1n02x5 U3807 (.a(n2930),
    .b(gen_filter_21__u_filter_diff_ctr_q[0]),
    .c(gen_filter_21__u_filter_diff_ctr_q[1]),
    .o1(n2932));
 b15aoi012ar1n04x5 U3808 (.a(n2931),
    .b(n2935),
    .c(n2932),
    .o1(gen_filter_21__u_filter_diff_ctr_d[1]));
 b15nand02al1n03x5 U3809 (.a(gen_filter_21__u_filter_diff_ctr_q[3]),
    .b(gen_filter_21__u_filter_diff_ctr_d[1]),
    .o1(n2933));
 b15aoi112ah1n04x5 U3810 (.a(n2934),
    .b(n2933),
    .c(gen_filter_21__u_filter_diff_ctr_q[0]),
    .d(n2935),
    .o1(eq_x_76_n25));
 b15aboi22al1n12x5 U3811 (.a(net2030),
    .b(net2041),
    .c(net2030),
    .d(n2936),
    .out0(net240));
 b15inv000as1n05x5 U3812 (.a(net2122),
    .o1(net242));
 b15aboi22aq1n04x5 U3813 (.a(net2026),
    .b(n2937),
    .c(net2026),
    .d(net2012),
    .out0(n2940));
 b15aoi022ah1n16x5 U3814 (.a(net2055),
    .b(net242),
    .c(net291),
    .d(n2938),
    .o1(n2939));
 b15xor002as1n03x5 U3815 (.a(n2940),
    .b(net2056),
    .out0(n2941));
 b15xor002an1n03x5 U3816 (.a(net2057),
    .b(net2042),
    .out0(net298));
 b15xor002al1n03x5 U3817 (.a(net2076),
    .b(net2057),
    .out0(net238));
 b15oai012ah1n02x5 U3818 (.a(n2942),
    .b(gen_filter_1__u_filter_diff_ctr_q[0]),
    .c(net2450),
    .o1(n2944));
 b15nand02as1n03x5 U3819 (.a(n2947),
    .b(n2943),
    .o1(n2945));
 b15aoai13al1n06x5 U3820 (.a(n2945),
    .b(n2944),
    .c(net2450),
    .d(gen_filter_1__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_1__u_filter_diff_ctr_d[1]));
 b15oai012al1n06x5 U3821 (.a(n2945),
    .b(net2499),
    .c(n2946),
    .o1(gen_filter_1__u_filter_diff_ctr_d[0]));
 b15and003an1n04x5 U3822 (.a(n2947),
    .b(gen_filter_1__u_filter_diff_ctr_d[1]),
    .c(gen_filter_1__u_filter_diff_ctr_d[0]),
    .o(eq_x_176_n25));
 b15oai012aq1n03x5 U3823 (.a(n2948),
    .b(gen_filter_30__u_filter_diff_ctr_q[0]),
    .c(gen_filter_30__u_filter_diff_ctr_q[1]),
    .o1(n2950));
 b15nand02as1n06x5 U3824 (.a(n2953),
    .b(n2949),
    .o1(n2951));
 b15aoai13aq1n08x5 U3825 (.a(n2951),
    .b(n2950),
    .c(gen_filter_30__u_filter_diff_ctr_q[1]),
    .d(gen_filter_30__u_filter_diff_ctr_q[0]),
    .o1(gen_filter_30__u_filter_diff_ctr_d[1]));
 b15oai012ar1n16x5 U3826 (.a(n2951),
    .b(gen_filter_30__u_filter_diff_ctr_q[0]),
    .c(n2952),
    .o1(gen_filter_30__u_filter_diff_ctr_d[0]));
 b15and003an1n03x5 U3827 (.a(n2953),
    .b(gen_filter_30__u_filter_diff_ctr_d[1]),
    .c(gen_filter_30__u_filter_diff_ctr_d[0]),
    .o(eq_x_31_n25));
 b15inv040ah1n16x5 U3828 (.a(net2166),
    .o1(n3037));
 b15aboi22aq1n16x5 U3829 (.a(net2214),
    .b(n3037),
    .c(net2166),
    .d(net2214),
    .out0(n2957));
 b15inv000ah1n16x5 U3830 (.a(net476),
    .o1(n3042));
 b15inv000as1n10x5 U3831 (.a(net268),
    .o1(n2988));
 b15aoi022an1n48x5 U3832 (.a(net268),
    .b(n3042),
    .c(net2157),
    .d(n2988),
    .o1(n3025));
 b15inv000aq1n12x5 U3833 (.a(net253),
    .o1(n2977));
 b15inv040as1n08x5 U3834 (.a(net266),
    .o1(n2982));
 b15aoi022al1n24x5 U3835 (.a(net266),
    .b(n2977),
    .c(net2180),
    .d(n2982),
    .o1(n2954));
 b15qgbxo2an1n10x5 U3836 (.a(n3025),
    .b(n2954),
    .out0(n2955));
 b15inv000ah1n10x5 U3837 (.a(net484),
    .o1(n3021));
 b15inv000al1n20x5 U3838 (.a(net471),
    .o1(n2987));
 b15aoi022ar1n32x5 U3839 (.a(net472),
    .b(net483),
    .c(n3021),
    .d(n2987),
    .o1(n3001));
 b15xor002aq1n08x5 U3840 (.a(n2955),
    .b(n3001),
    .out0(n2956));
 b15xor002an1n12x5 U3841 (.a(net2215),
    .b(n2956),
    .out0(n2960));
 b15inv000ar1n28x5 U3842 (.a(net2146),
    .o1(n2989));
 b15inv000ar1n24x5 U3843 (.a(net2143),
    .o1(n3038));
 b15aoi022as1n48x5 U3844 (.a(net2144),
    .b(net502),
    .c(n2989),
    .d(n3038),
    .o1(n3056));
 b15inv040al1n12x5 U3845 (.a(net498),
    .o1(n3014));
 b15inv000as1n20x5 U3846 (.a(net2175),
    .o1(n3000));
 b15aoi022al1n32x5 U3847 (.a(net482),
    .b(net498),
    .c(n3014),
    .d(net458),
    .o1(n2958));
 b15xor002as1n12x5 U3848 (.a(n3056),
    .b(n2958),
    .out0(n2959));
 b15xor002ah1n16x5 U3849 (.a(net2216),
    .b(n2959),
    .out0(net297));
 b15nanb02as1n12x5 U3850 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[1]),
    .b(n2965),
    .out0(n2963));
 b15inv020ar1n08x5 U3851 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .o1(n2962));
 b15nandp2al1n08x5 U3852 (.a(n2963),
    .b(net2438),
    .o1(n2961));
 b15oai012an1n32x5 U3853 (.a(n2961),
    .b(n2963),
    .c(n2962),
    .o1(gen_alert_tx_0__u_prim_alert_sender_ack_level));
 b15nandp2ar1n08x5 U3854 (.a(net2317),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[1]),
    .o1(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39));
 b15nonb03an1n06x5 U3855 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39),
    .b(n2965),
    .c(n2964),
    .out0(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[1]));
 b15nand02as1n06x5 U3856 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[0]),
    .b(net2564),
    .o1(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39));
 b15nonb03ar1n08x5 U3857 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39),
    .b(n2967),
    .c(n2966),
    .out0(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[1]));
 b15inv020ar1n08x5 U3858 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .o1(n3367));
 b15nandp2ar1n05x5 U3859 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .b(n3367),
    .o1(n2969));
 b15qgbno2an1n05x5 U3860 (.o1(n3365),
    .a(n3367),
    .b(gen_alert_tx_0__u_prim_alert_sender_state_q[2]));
 b15inv000al1n02x5 U3861 (.a(gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .o1(n2968));
 b15obai22ah1n06x5 U3862 (.a(n2969),
    .b(n3365),
    .c(n2968),
    .d(net2636),
    .out0(n2970));
 b15inv020as1n08x5 U3863 (.a(net2525),
    .o1(n3435));
 b15nor003ar1n12x5 U3864 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .b(gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .c(n3435),
    .o1(n3434));
 b15orn002ah1n12x5 U3865 (.a(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[1]),
    .b(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[1]),
    .o(n3439));
 b15aoi112as1n04x5 U3866 (.a(n3434),
    .b(n3439),
    .c(n2969),
    .d(n2970),
    .o1(gen_alert_tx_0__u_prim_alert_sender_state_d[2]));
 b15nor002as1n04x5 U3867 (.a(n2970),
    .b(net2636),
    .o1(n3438));
 b15nor002aq1n04x5 U3868 (.a(n2972),
    .b(n2971),
    .o1(n2975));
 b15inv000aq1n02x5 U3869 (.a(n2973),
    .o1(n2974));
 b15oaoi13al1n08x5 U3870 (.a(net2443),
    .b(n2974),
    .c(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[0]),
    .d(n2975),
    .o1(n3364));
 b15aoi112an1n02x5 U3871 (.a(n3364),
    .b(n3439),
    .c(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .d(n3438),
    .o1(gen_alert_tx_0__u_prim_alert_sender_ping_set_d));
 b15inv020as1n12x5 U3872 (.a(net466),
    .o1(n3048));
 b15inv020an1n16x5 U3873 (.a(net262),
    .o1(n3030));
 b15aoi022an1n16x5 U3874 (.a(net2205),
    .b(net465),
    .c(n3048),
    .d(n3030),
    .o1(n2976));
 b15xor002as1n16x5 U3875 (.a(net507),
    .b(n2976),
    .out0(n2993));
 b15inv000aq1n20x5 U3876 (.a(net491),
    .o1(n3015));
 b15aboi22ah1n24x5 U3877 (.a(net495),
    .b(net253),
    .c(net495),
    .d(n2977),
    .out0(n2978));
 b15xor002as1n16x5 U3878 (.a(net504),
    .b(n2978),
    .out0(n3046));
 b15xor002ah1n08x5 U3879 (.a(n3015),
    .b(n3046),
    .out0(n2980));
 b15inv000ah1n16x5 U3880 (.a(net473),
    .o1(n2998));
 b15aoi022as1n48x5 U3881 (.a(net462),
    .b(net474),
    .c(n2998),
    .d(n3037),
    .o1(n2979));
 b15xor002al1n16x5 U3882 (.a(n2980),
    .b(n2979),
    .out0(n2981));
 b15xor002as1n12x5 U3883 (.a(n2993),
    .b(n2981),
    .out0(n2986));
 b15inv040as1n08x5 U3884 (.a(net497),
    .o1(n3041));
 b15aoi022ah1n32x5 U3885 (.a(net266),
    .b(net2134),
    .c(n3041),
    .d(n2982),
    .o1(n2984));
 b15inv040ah1n05x5 U3886 (.a(net494),
    .o1(n3029));
 b15inv000as1n05x5 U3887 (.a(net265),
    .o1(n3020));
 b15aoi022aq1n16x5 U3888 (.a(net265),
    .b(net494),
    .c(net457),
    .d(n3020),
    .o1(n2983));
 b15xor002as1n16x5 U3889 (.a(n2984),
    .b(n2983),
    .out0(n2985));
 b15xor002as1n16x5 U3890 (.a(n2985),
    .b(net2276),
    .out0(n3003));
 b15xor002as1n06x5 U3891 (.a(n2986),
    .b(n3003),
    .out0(net280));
 b15aoi022an1n16x5 U3892 (.a(net471),
    .b(net268),
    .c(n2988),
    .d(n2987),
    .o1(n2997));
 b15inv020ah1n32x5 U3893 (.a(net2141),
    .o1(n3012));
 b15aoi022ah1n48x5 U3894 (.a(net501),
    .b(net503),
    .c(n2989),
    .d(n3012),
    .o1(n2991));
 b15inv040al1n10x5 U3895 (.a(net459),
    .o1(n3016));
 b15aboi22as1n24x5 U3896 (.a(net277),
    .b(n3016),
    .c(net277),
    .d(net460),
    .out0(n2990));
 b15xor002al1n16x5 U3897 (.a(n2991),
    .b(n2990),
    .out0(n2995));
 b15inv020ar1n32x5 U3898 (.a(net510),
    .o1(n3047));
 b15inv040as1n04x5 U3899 (.a(net468),
    .o1(n3007));
 b15aoi022as1n48x5 U3900 (.a(net469),
    .b(net511),
    .c(n3047),
    .d(net456),
    .o1(n3028));
 b15inv020as1n16x5 U3901 (.a(net488),
    .o1(n3043));
 b15aboi22aq1n24x5 U3902 (.a(n3028),
    .b(n3043),
    .c(net272),
    .d(n3028),
    .out0(n2992));
 b15xor002as1n16x5 U3903 (.a(n2993),
    .b(n2992),
    .out0(n2994));
 b15xor002as1n16x5 U3904 (.a(n2995),
    .b(n2994),
    .out0(n2996));
 b15xor002ar1n16x5 U3905 (.a(n2997),
    .b(n2996),
    .out0(n2999));
 b15inv000ah1n10x5 U3906 (.a(net269),
    .o1(n3008));
 b15aoi022al1n32x5 U3907 (.a(net2136),
    .b(net2115),
    .c(n2998),
    .d(n3008),
    .o1(n3013));
 b15xor002aq1n06x5 U3908 (.a(n2999),
    .b(net2137),
    .out0(net295));
 b15aboi22as1n24x5 U3909 (.a(net263),
    .b(net480),
    .c(net263),
    .d(net458),
    .out0(n3035));
 b15xor002as1n08x5 U3910 (.a(n3001),
    .b(net464),
    .out0(n3005));
 b15inv040ah1n24x5 U3911 (.a(net486),
    .o1(n3011));
 b15aoi022an1n48x5 U3912 (.a(net489),
    .b(net487),
    .c(n3011),
    .d(n3043),
    .o1(n3002));
 b15xor002as1n16x5 U3913 (.a(n3003),
    .b(n3002),
    .out0(n3004));
 b15xor002ah1n12x5 U3914 (.a(n3005),
    .b(n3004),
    .out0(n3006));
 b15xor002an1n16x5 U3915 (.a(n3035),
    .b(n3006),
    .out0(n3010));
 b15aoi022an1n32x5 U3916 (.a(net2177),
    .b(net2136),
    .c(n3008),
    .d(net456),
    .o1(n3009));
 b15xor002aq1n16x5 U3917 (.a(n3010),
    .b(net2178),
    .out0(net270));
 b15aoi022as1n48x5 U3918 (.a(net485),
    .b(net499),
    .c(n3012),
    .d(n3011),
    .o1(n3053));
 b15xor002as1n06x5 U3919 (.a(net2137),
    .b(n3053),
    .out0(n3024));
 b15aoi022as1n12x5 U3920 (.a(net2129),
    .b(net490),
    .c(n3015),
    .d(n3014),
    .o1(n3018));
 b15inv040aq1n05x5 U3921 (.a(net478),
    .o1(n3044));
 b15aoi022ah1n08x5 U3922 (.a(net459),
    .b(net478),
    .c(n3044),
    .d(n3016),
    .o1(n3017));
 b15xor002ah1n12x5 U3923 (.a(n3018),
    .b(net407),
    .out0(n3019));
 b15xor002as1n16x5 U3924 (.a(n3019),
    .b(net464),
    .out0(n3032));
 b15aoi022as1n12x5 U3925 (.a(net265),
    .b(net483),
    .c(n3021),
    .d(n3020),
    .o1(n3022));
 b15xor002an1n16x5 U3926 (.a(n3032),
    .b(n3022),
    .out0(n3023));
 b15qgbxo2an1n10x5 U3927 (.a(n3024),
    .b(n3023),
    .out0(n3026));
 b15xor002an1n16x5 U3928 (.a(n3026),
    .b(n3025),
    .out0(n3027));
 b15xor002an1n12x5 U3929 (.a(n3027),
    .b(net2182),
    .out0(net296));
 b15xor002aq1n08x5 U3930 (.a(net504),
    .b(n3028),
    .out0(n3034));
 b15aoi022as1n48x5 U3931 (.a(net492),
    .b(net496),
    .c(n3030),
    .d(net457),
    .o1(n3031));
 b15xor002ah1n12x5 U3932 (.a(n3032),
    .b(n3031),
    .out0(n3033));
 b15xor002an1n16x5 U3933 (.a(n3034),
    .b(n3033),
    .out0(n3036));
 b15xor002an1n12x5 U3934 (.a(n3036),
    .b(n3035),
    .out0(n3040));
 b15aoi022an1n48x5 U3935 (.a(net2167),
    .b(net505),
    .c(n3038),
    .d(n3037),
    .o1(n3039));
 b15xor002as1n16x5 U3936 (.a(n3040),
    .b(net2201),
    .out0(net290));
 b15aoi022as1n32x5 U3937 (.a(net2133),
    .b(net2156),
    .c(n3042),
    .d(n3041),
    .o1(n3052));
 b15aoi022an1n16x5 U3938 (.a(net488),
    .b(n3044),
    .c(net478),
    .d(n3043),
    .o1(n3045));
 b15xor002an1n12x5 U3939 (.a(n3046),
    .b(n3045),
    .out0(n3050));
 b15aoi022aq1n16x5 U3940 (.a(net509),
    .b(net465),
    .c(n3048),
    .d(n3047),
    .o1(n3049));
 b15xor002as1n16x5 U3941 (.a(n3050),
    .b(n3049),
    .out0(n3051));
 b15xor002as1n03x5 U3942 (.a(n3052),
    .b(n3051),
    .out0(n3054));
 b15xor002as1n08x5 U3943 (.a(n3054),
    .b(n3053),
    .out0(n3055));
 b15xor002as1n16x5 U3944 (.a(n3056),
    .b(n3055),
    .out0(n3057));
 b15xor002as1n06x5 U3945 (.a(n3057),
    .b(net2292),
    .out0(net259));
 b15inv040aq1n06x5 U3946 (.a(net96),
    .o1(n3159));
 b15norp02aq1n12x5 U3947 (.a(net95),
    .b(n3159),
    .o1(n3074));
 b15norp02ar1n02x5 U3948 (.a(net91),
    .b(net90),
    .o1(n3058));
 b15nandp2aq1n02x5 U3949 (.a(n3074),
    .b(n3058),
    .o1(n3061));
 b15inv000an1n06x5 U3950 (.a(net93),
    .o1(n3264));
 b15inv000an1n06x5 U3951 (.a(net95),
    .o1(n3194));
 b15nor002ah1n06x5 U3952 (.a(n3194),
    .b(net96),
    .o1(n3075));
 b15aboi22aq1n02x5 U3953 (.a(n3075),
    .b(net91),
    .c(net90),
    .d(net95),
    .out0(n3059));
 b15inv000al1n10x5 U3954 (.a(net92),
    .o1(n3265));
 b15oai112ah1n06x5 U3955 (.a(n3059),
    .b(n3265),
    .c(net96),
    .d(n3264),
    .o1(n3060));
 b15oai022an1n08x5 U3956 (.a(n3061),
    .b(net93),
    .c(n3074),
    .d(n3060),
    .o1(n3285));
 b15inv000ar1n06x5 U3957 (.a(net39),
    .o1(n3271));
 b15nanb02ah1n08x5 U3958 (.a(net40),
    .b(n3271),
    .out0(n3284));
 b15inv000an1n08x5 U3959 (.a(net91),
    .o1(n3145));
 b15norp03ah1n12x5 U3960 (.a(n3145),
    .b(n3265),
    .c(n3264),
    .o1(n3279));
 b15nor002ah1n24x5 U3961 (.a(net100),
    .b(net99),
    .o1(n3484));
 b15inv000ah1n24x5 U3962 (.a(n3484),
    .o1(n3300));
 b15nandp2an1n48x5 U3963 (.a(net97),
    .b(net98),
    .o1(n3361));
 b15norp02ar1n16x5 U3964 (.a(n3300),
    .b(n3361),
    .o1(n3286));
 b15qgbin1an1n15x5 U3965 (.a(net43),
    .o1(n3280));
 b15nand02as1n24x5 U3966 (.a(u_reg_u_reg_if_a_ack),
    .b(n3280),
    .o1(n3297));
 b15oaoi13al1n04x5 U3967 (.a(n3297),
    .b(net90),
    .c(n3279),
    .d(n3286),
    .o1(n3275));
 b15xor002an1n12x5 U3968 (.a(net104),
    .b(net107),
    .out0(n3063));
 b15xor002as1n08x5 U3969 (.a(net103),
    .b(net106),
    .out0(n3062));
 b15xor002as1n16x5 U3970 (.a(n3063),
    .b(n3062),
    .out0(n3118));
 b15xor002an1n06x5 U3971 (.a(net45),
    .b(net118),
    .out0(n3065));
 b15xor002as1n16x5 U3972 (.a(net126),
    .b(net129),
    .out0(n3084));
 b15xor002ah1n06x5 U3973 (.a(net115),
    .b(n3084),
    .out0(n3064));
 b15qgbxo2an1n10x5 U3974 (.a(n3065),
    .b(n3064),
    .out0(n3066));
 b15xor002as1n08x5 U3975 (.a(n3118),
    .b(n3066),
    .out0(n3069));
 b15inv000as1n06x5 U3976 (.a(net42),
    .o1(n3267));
 b15aboi22aq1n16x5 U3977 (.a(net117),
    .b(n3267),
    .c(net42),
    .d(net117),
    .out0(n3067));
 b15xor002as1n16x5 U3978 (.a(net114),
    .b(n3067),
    .out0(n3152));
 b15inv000ah1n08x5 U3979 (.a(net51),
    .o1(n3193));
 b15inv020an1n16x5 U3980 (.a(net50),
    .o1(n3177));
 b15aoi022al1n32x5 U3981 (.a(net50),
    .b(net51),
    .c(n3193),
    .d(n3177),
    .o1(n3080));
 b15xor002aq1n08x5 U3982 (.a(n3152),
    .b(n3080),
    .out0(n3068));
 b15xor002as1n06x5 U3983 (.a(n3069),
    .b(n3068),
    .out0(n3070));
 b15xor002as1n12x5 U3984 (.a(net119),
    .b(n3070),
    .out0(n3072));
 b15xor002as1n16x5 U3985 (.a(net128),
    .b(net125),
    .out0(n3148));
 b15xor002as1n16x5 U3986 (.a(n3148),
    .b(net90),
    .out0(n3085));
 b15xor002an1n12x5 U3987 (.a(n3085),
    .b(net120),
    .out0(n3071));
 b15xor002an1n16x5 U3988 (.a(n3072),
    .b(n3071),
    .out0(n3261));
 b15oai012al1n06x5 U3989 (.a(net43),
    .b(n3075),
    .c(n3074),
    .o1(n3073));
 b15oai013as1n12x5 U3990 (.a(n3073),
    .b(n3075),
    .c(net43),
    .d(n3074),
    .o1(n3260));
 b15norp02ar1n02x5 U3991 (.a(net91),
    .b(net92),
    .o1(n3076));
 b15aoi012aq1n04x5 U3992 (.a(n3076),
    .b(net92),
    .c(net91),
    .o1(n3252));
 b15aboi22an1n12x5 U3993 (.a(net101),
    .b(n3267),
    .c(net42),
    .d(net101),
    .out0(n3077));
 b15xor002as1n12x5 U3994 (.a(net127),
    .b(n3077),
    .out0(n3079));
 b15inv000as1n20x5 U3995 (.a(net98),
    .o1(n3293));
 b15nandp2al1n32x5 U3996 (.a(n3293),
    .b(net97),
    .o1(n3299));
 b15qbfin1bn1n40x5 U3997 (.a(net97),
    .o1(n3372));
 b15nand02ah1n48x5 U3998 (.a(n3372),
    .b(net98),
    .o1(n3442));
 b15and002aq1n12x5 U3999 (.a(n3299),
    .b(n3442),
    .o(n3760));
 b15inv000ah1n08x5 U4000 (.a(net52),
    .o1(n3268));
 b15inv020ah1n10x5 U4001 (.a(net53),
    .o1(n3263));
 b15aoi022aq1n32x5 U4002 (.a(net53),
    .b(net52),
    .c(n3268),
    .d(n3263),
    .o1(n3119));
 b15xor002al1n12x5 U4003 (.a(n3760),
    .b(n3119),
    .out0(n3144));
 b15xor002aq1n08x5 U4004 (.a(n3144),
    .b(net102),
    .out0(n3078));
 b15xor002ar1n12x5 U4005 (.a(n3079),
    .b(n3078),
    .out0(n3083));
 b15inv040ah1n12x5 U4006 (.a(net100),
    .o1(n3296));
 b15inv000as1n20x5 U4007 (.a(net99),
    .o1(n3291));
 b15norp02an1n24x5 U4008 (.a(n3296),
    .b(n3291),
    .o1(n3337));
 b15xnr002as1n16x5 U4009 (.a(net41),
    .b(n3080),
    .out0(n3113));
 b15oai012ah1n02x5 U4010 (.a(n3113),
    .b(n3484),
    .c(n3337),
    .o1(n3081));
 b15oai013aq1n08x5 U4011 (.a(n3081),
    .b(n3484),
    .c(n3337),
    .d(n3113),
    .o1(n3082));
 b15xor002al1n04x5 U4012 (.a(n3083),
    .b(n3082),
    .out0(n3086));
 b15xor002as1n12x5 U4013 (.a(net93),
    .b(n3084),
    .out0(n3198));
 b15xor002an1n12x5 U4014 (.a(n3198),
    .b(n3085),
    .out0(n3120));
 b15xor002ar1n03x5 U4015 (.a(n3086),
    .b(n3120),
    .out0(n3087));
 b15xor002as1n02x5 U4016 (.a(n3260),
    .b(n3087),
    .out0(n3123));
 b15ztpn00an1n08x5 PHY_63 ();
 b15inv040as1n36x5 U4018 (.a(net59),
    .o1(n3538));
 b15ztpn00an1n08x5 PHY_62 ();
 b15oai022as1n24x5 U4020 (.a(net757),
    .b(net820),
    .c(net55),
    .d(net59),
    .o1(n3208));
 b15inv040ah1n06x5 U4021 (.a(n3208),
    .o1(n3088));
 b15xor002as1n08x5 U4022 (.a(n4070),
    .b(n3088),
    .out0(n3111));
 b15ztpn00an1n08x5 PHY_61 ();
 b15ztpn00an1n08x5 PHY_60 ();
 b15aoi022ah1n24x5 U4025 (.a(net89),
    .b(net88),
    .c(net761),
    .d(net760),
    .o1(n3097));
 b15ztpn00an1n08x5 PHY_59 ();
 b15ztpn00an1n08x5 PHY_58 ();
 b15norp02as1n48x5 U4028 (.a(n4075),
    .b(net777),
    .o1(n3450));
 b15oabi12aq1n03x5 U4029 (.a(n3450),
    .b(net65),
    .c(net822),
    .out0(n3090));
 b15nand02ar1n02x5 U4030 (.a(n3090),
    .b(net94),
    .o1(n3089));
 b15oai012ah1n03x5 U4031 (.a(n3089),
    .b(net94),
    .c(n3090),
    .o1(n3091));
 b15xor002an1n04x5 U4032 (.a(net832),
    .b(n3091),
    .out0(n3094));
 b15ztpn00an1n08x5 PHY_57 ();
 b15ztpn00an1n08x5 PHY_56 ();
 b15aoi022ar1n48x5 U4035 (.a(net80),
    .b(net79),
    .c(net786),
    .d(n4088),
    .o1(n3232));
 b15ztpn00an1n08x5 PHY_55 ();
 b15inv000as1n64x5 U4037 (.a(net69),
    .o1(n3524));
 b15aoi022aq1n16x5 U4038 (.a(net69),
    .b(net68),
    .c(n4078),
    .d(n3524),
    .o1(n3092));
 b15xor002aq1n16x5 U4039 (.a(n3232),
    .b(n3092),
    .out0(n3093));
 b15xor002an1n06x5 U4040 (.a(n3094),
    .b(n3093),
    .out0(n3095));
 b15xor002aq1n08x5 U4041 (.a(n3097),
    .b(n3095),
    .out0(n3096));
 b15ztpn00an1n08x5 PHY_54 ();
 b15ztpn00an1n08x5 PHY_53 ();
 b15aoi022aq1n48x5 U4044 (.a(net73),
    .b(net60),
    .c(n4071),
    .d(n4081),
    .o1(n3220));
 b15xor002ar1n16x5 U4045 (.a(n3096),
    .b(n3220),
    .out0(n3110));
 b15ztpn00an1n08x5 PHY_52 ();
 b15ztpn00an1n08x5 PHY_51 ();
 b15aoi022aq1n16x5 U4048 (.a(net828),
    .b(net71),
    .c(n4080),
    .d(net805),
    .o1(n3128));
 b15ztpn00an1n08x5 PHY_50 ();
 b15ztpn00an1n08x5 PHY_49 ();
 b15aoi022as1n24x5 U4051 (.a(net84),
    .b(net85),
    .c(net771),
    .d(net774),
    .o1(n3231));
 b15xor002as1n08x5 U4052 (.a(n3128),
    .b(n3231),
    .out0(n3099));
 b15xor002ah1n06x5 U4053 (.a(n3097),
    .b(net826),
    .out0(n3098));
 b15xor002as1n08x5 U4054 (.a(n3099),
    .b(n3098),
    .out0(n3109));
 b15ztpn00an1n08x5 PHY_48 ();
 b15aoi022as1n12x5 U4056 (.a(net822),
    .b(net86),
    .c(net770),
    .d(net777),
    .o1(n3103));
 b15ztpn00an1n08x5 PHY_47 ();
 b15nor002as1n32x5 U4058 (.a(net757),
    .b(net795),
    .o1(n3462));
 b15oabi12al1n12x5 U4059 (.a(n3462),
    .b(net59),
    .c(net77),
    .out0(n3101));
 b15nandp2as1n04x5 U4060 (.a(n3101),
    .b(net61),
    .o1(n3100));
 b15oai012al1n24x5 U4061 (.a(n3100),
    .b(net61),
    .c(n3101),
    .o1(n3102));
 b15xor002al1n06x5 U4062 (.a(n3103),
    .b(n3102),
    .out0(n3106));
 b15ztpn00an1n08x5 PHY_46 ();
 b15ztpn00an1n08x5 PHY_45 ();
 b15aoi022al1n24x5 U4065 (.a(net825),
    .b(net62),
    .c(n4072),
    .d(net789),
    .o1(n3104));
 b15xor002as1n06x5 U4066 (.a(net80),
    .b(n3104),
    .out0(n3105));
 b15xor002an1n08x5 U4067 (.a(n3106),
    .b(n3105),
    .out0(n3108));
 b15oai022as1n06x5 U4068 (.a(n3111),
    .b(n3110),
    .c(n3108),
    .d(n3109),
    .o1(n3107));
 b15aoi122as1n08x5 U4069 (.a(n3107),
    .b(n3111),
    .c(n3110),
    .d(n3109),
    .e(n3108),
    .o1(n3112));
 b15oai012as1n04x5 U4070 (.a(n3112),
    .b(n3252),
    .c(n3123),
    .o1(n3258));
 b15xor002an1n08x5 U4071 (.a(net113),
    .b(net112),
    .out0(n3114));
 b15xor002ah1n08x5 U4072 (.a(n3114),
    .b(n3113),
    .out0(n3174));
 b15xnr002aq1n06x5 U4073 (.a(n3174),
    .b(net138),
    .out0(n3116));
 b15xor002as1n06x5 U4074 (.a(net109),
    .b(net108),
    .out0(n3147));
 b15xor002al1n04x5 U4075 (.a(net110),
    .b(n3147),
    .out0(n3115));
 b15xor002ah1n03x5 U4076 (.a(n3116),
    .b(n3115),
    .out0(n3117));
 b15xor002as1n06x5 U4077 (.a(n3118),
    .b(n3117),
    .out0(n3122));
 b15xor002al1n16x5 U4078 (.a(n3119),
    .b(net111),
    .out0(n3186));
 b15xor002as1n04x5 U4079 (.a(n3120),
    .b(n3186),
    .out0(n3121));
 b15xor002ah1n04x5 U4080 (.a(n3122),
    .b(n3121),
    .out0(n3256));
 b15inv000al1n02x5 U4081 (.a(n3123),
    .o1(n3255));
 b15ztpn00an1n08x5 PHY_44 ();
 b15ztpn00an1n08x5 PHY_43 ();
 b15aoi022aq1n16x5 U4084 (.a(net64),
    .b(net831),
    .c(n4069),
    .d(n4074),
    .o1(n3125));
 b15ztpn00an1n08x5 PHY_42 ();
 b15aoi022an1n12x5 U4086 (.a(net68),
    .b(net66),
    .c(n4076),
    .d(n4078),
    .o1(n3124));
 b15xor002an1n12x5 U4087 (.a(n3125),
    .b(n3124),
    .out0(n3143));
 b15ztpn00an1n08x5 PHY_41 ();
 b15aoi022ah1n12x5 U4089 (.a(net84),
    .b(net800),
    .c(net827),
    .d(n4091),
    .o1(n3132));
 b15ztpn00an1n08x5 PHY_40 ();
 b15aoi022ah1n12x5 U4091 (.a(net822),
    .b(net67),
    .c(n4077),
    .d(net777),
    .o1(n3127));
 b15aoi022ah1n24x5 U4092 (.a(net55),
    .b(net60),
    .c(n4071),
    .d(net820),
    .o1(n3126));
 b15xor002as1n12x5 U4093 (.a(n3127),
    .b(n3126),
    .out0(n3130));
 b15xor002an1n12x5 U4094 (.a(n3128),
    .b(net54),
    .out0(n3129));
 b15xor002ah1n08x5 U4095 (.a(n3130),
    .b(n3129),
    .out0(n3131));
 b15xor002as1n12x5 U4096 (.a(n3132),
    .b(n3131),
    .out0(n3133));
 b15ztpn00an1n08x5 PHY_39 ();
 b15norp02aq1n48x5 U4098 (.a(n3524),
    .b(net765),
    .o1(n3460));
 b15oabi12aq1n12x5 U4099 (.a(n3460),
    .b(net69),
    .c(net87),
    .out0(n3228));
 b15xor002aq1n08x5 U4100 (.a(n3133),
    .b(n3228),
    .out0(n3142));
 b15ztpn00an1n08x5 PHY_38 ();
 b15aoi022aq1n08x5 U4102 (.a(net86),
    .b(net70),
    .c(net810),
    .d(net770),
    .o1(n3139));
 b15ztpn00an1n08x5 PHY_37 ();
 b15aoi022as1n48x5 U4104 (.a(net77),
    .b(net63),
    .c(net814),
    .d(net795),
    .o1(n3219));
 b15xor002al1n12x5 U4105 (.a(n3219),
    .b(net116),
    .out0(n3137));
 b15aoi022as1n08x5 U4106 (.a(net89),
    .b(net79),
    .c(n4087),
    .d(net758),
    .o1(n3135));
 b15ztpn00an1n08x5 PHY_36 ();
 b15aoi022al1n12x5 U4108 (.a(net832),
    .b(net85),
    .c(net771),
    .d(n4068),
    .o1(n3134));
 b15xor002as1n06x5 U4109 (.a(n3135),
    .b(n3134),
    .out0(n3136));
 b15xor002al1n08x5 U4110 (.a(n3137),
    .b(n3136),
    .out0(n3138));
 b15xor002aq1n08x5 U4111 (.a(n3139),
    .b(n3138),
    .out0(n3141));
 b15nand03as1n03x5 U4112 (.a(n3143),
    .b(n3142),
    .c(n3141),
    .o1(n3140));
 b15oai013an1n12x5 U4113 (.a(n3140),
    .b(n3143),
    .c(n3142),
    .d(n3141),
    .o1(n3254));
 b15inv040aq1n02x5 U4114 (.a(n3144),
    .o1(n3176));
 b15inv000ah1n05x5 U4115 (.a(net110),
    .o1(n3160));
 b15aboi22an1n06x5 U4116 (.a(net122),
    .b(n3160),
    .c(net122),
    .d(net110),
    .out0(n3156));
 b15aoi022an1n24x5 U4117 (.a(net99),
    .b(net91),
    .c(n3145),
    .d(n3291),
    .o1(n3146));
 b15xor002an1n06x5 U4118 (.a(n3147),
    .b(n3146),
    .out0(n3150));
 b15xor002as1n06x5 U4119 (.a(net115),
    .b(net123),
    .out0(n3203));
 b15xor002an1n08x5 U4120 (.a(n3148),
    .b(n3203),
    .out0(n3149));
 b15xor002aq1n08x5 U4121 (.a(n3150),
    .b(n3149),
    .out0(n3151));
 b15xor002al1n12x5 U4122 (.a(net103),
    .b(n3151),
    .out0(n3154));
 b15xor002al1n12x5 U4123 (.a(n3152),
    .b(net46),
    .out0(n3153));
 b15qgbxo2an1n05x5 U4124 (.a(n3154),
    .b(n3153),
    .out0(n3155));
 b15qgbxo2an1n05x5 U4125 (.a(n3156),
    .b(n3155),
    .out0(n3158));
 b15xor002ah1n03x5 U4126 (.a(net126),
    .b(net121),
    .out0(n3157));
 b15xor002aq1n06x5 U4127 (.a(n3158),
    .b(n3157),
    .out0(n3175));
 b15aboi22al1n12x5 U4128 (.a(net124),
    .b(n3159),
    .c(net96),
    .d(net124),
    .out0(n3169));
 b15aboi22ar1n16x5 U4129 (.a(net107),
    .b(n3160),
    .c(net110),
    .d(net107),
    .out0(n3165));
 b15xor002as1n06x5 U4130 (.a(net101),
    .b(net119),
    .out0(n3161));
 b15xor002aq1n16x5 U4131 (.a(n3161),
    .b(net122),
    .out0(n3185));
 b15aoi022as1n08x5 U4132 (.a(net99),
    .b(net53),
    .c(n3263),
    .d(n3291),
    .o1(n3162));
 b15xor002as1n06x5 U4133 (.a(n3185),
    .b(n3162),
    .out0(n3163));
 b15xor002aq1n16x5 U4134 (.a(net102),
    .b(net120),
    .out0(n3197));
 b15xor002al1n12x5 U4135 (.a(n3163),
    .b(n3197),
    .out0(n3164));
 b15qgbxo2an1n10x5 U4136 (.a(n3165),
    .b(n3164),
    .out0(n3167));
 b15xor002al1n16x5 U4137 (.a(net117),
    .b(net49),
    .out0(n3166));
 b15qgbxo2an1n10x5 U4138 (.a(n3167),
    .b(n3166),
    .out0(n3168));
 b15xor002an1n12x5 U4139 (.a(n3169),
    .b(n3168),
    .out0(n3171));
 b15xor002ah1n03x5 U4140 (.a(net128),
    .b(net123),
    .out0(n3170));
 b15xor002aq1n08x5 U4141 (.a(n3171),
    .b(n3170),
    .out0(n3173));
 b15aoi022al1n02x5 U4142 (.a(n3176),
    .b(n3175),
    .c(n3173),
    .d(n3174),
    .o1(n3172));
 b15oai122aq1n08x5 U4143 (.a(n3172),
    .b(n3176),
    .c(n3175),
    .d(n3174),
    .e(n3173),
    .o1(n3251));
 b15aoi022an1n32x5 U4144 (.a(net43),
    .b(net50),
    .c(n3177),
    .d(n3280),
    .o1(n3181));
 b15xor002aq1n03x5 U4145 (.a(net104),
    .b(net47),
    .out0(n3179));
 b15xor002an1n06x5 U4146 (.a(net108),
    .b(net112),
    .out0(n3178));
 b15xor002an1n06x5 U4147 (.a(n3179),
    .b(n3178),
    .out0(n3180));
 b15qgbxo2an1n10x5 U4148 (.a(n3181),
    .b(n3180),
    .out0(n3183));
 b15xor002as1n03x5 U4149 (.a(net125),
    .b(net129),
    .out0(n3182));
 b15xor002as1n06x5 U4150 (.a(n3183),
    .b(n3182),
    .out0(n3190));
 b15aoi022an1n08x5 U4151 (.a(net97),
    .b(net92),
    .c(n3265),
    .d(n3372),
    .o1(n3184));
 b15xor002as1n06x5 U4152 (.a(n3185),
    .b(n3184),
    .out0(n3188));
 b15xor002ah1n03x5 U4153 (.a(net114),
    .b(n3186),
    .out0(n3187));
 b15xor002ah1n03x5 U4154 (.a(n3188),
    .b(n3187),
    .out0(n3189));
 b15xor002as1n03x5 U4155 (.a(n3190),
    .b(n3189),
    .out0(n3249));
 b15xor002ah1n08x5 U4156 (.a(net106),
    .b(net48),
    .out0(n3192));
 b15xor002as1n03x5 U4157 (.a(net113),
    .b(net111),
    .out0(n3191));
 b15xor002ar1n08x5 U4158 (.a(n3192),
    .b(n3191),
    .out0(n3202));
 b15aoi022ah1n12x5 U4159 (.a(net52),
    .b(n3193),
    .c(net51),
    .d(n3268),
    .o1(n3196));
 b15aoi022an1n16x5 U4160 (.a(net98),
    .b(net95),
    .c(n3194),
    .d(n3293),
    .o1(n3195));
 b15xor002ah1n08x5 U4161 (.a(n3196),
    .b(n3195),
    .out0(n3200));
 b15xor002an1n12x5 U4162 (.a(n3198),
    .b(n3197),
    .out0(n3199));
 b15xor002an1n16x5 U4163 (.a(n3200),
    .b(n3199),
    .out0(n3201));
 b15qgbxo2an1n05x5 U4164 (.a(n3202),
    .b(n3201),
    .out0(n3205));
 b15xor002an1n08x5 U4165 (.a(n3203),
    .b(net109),
    .out0(n3204));
 b15xor002ah1n04x5 U4166 (.a(n3205),
    .b(n3204),
    .out0(n3248));
 b15aboi22as1n04x5 U4167 (.a(net118),
    .b(net100),
    .c(net118),
    .d(n3296),
    .out0(n3206));
 b15xor002as1n04x5 U4168 (.a(net124),
    .b(n3206),
    .out0(n3207));
 b15xor002ah1n04x5 U4169 (.a(n3207),
    .b(net121),
    .out0(n3247));
 b15aoi022aq1n12x5 U4170 (.a(net66),
    .b(net814),
    .c(net63),
    .d(n4076),
    .o1(n3216));
 b15ztpn00an1n08x5 PHY_35 ();
 b15aoi022aq1n16x5 U4172 (.a(net86),
    .b(net823),
    .c(net780),
    .d(net770),
    .o1(n3212));
 b15aoi022al1n16x5 U4173 (.a(net825),
    .b(net67),
    .c(n4077),
    .d(net792),
    .o1(n3224));
 b15aoi022ah1n48x5 U4174 (.a(net62),
    .b(net70),
    .c(net810),
    .d(n4072),
    .o1(n3235));
 b15xor002ar1n12x5 U4175 (.a(n3224),
    .b(n3235),
    .out0(n3210));
 b15xor002al1n04x5 U4176 (.a(n3208),
    .b(net766),
    .out0(n3209));
 b15xor002as1n02x5 U4177 (.a(n3210),
    .b(n3209),
    .out0(n3211));
 b15xor002as1n02x5 U4178 (.a(n3212),
    .b(n3211),
    .out0(n3214));
 b15xor002as1n12x5 U4179 (.a(net73),
    .b(net83),
    .out0(n3213));
 b15xor002ah1n04x5 U4180 (.a(n3214),
    .b(n3213),
    .out0(n3215));
 b15xor002ah1n06x5 U4181 (.a(n3216),
    .b(n3215),
    .out0(n3244));
 b15aoi022an1n12x5 U4182 (.a(net828),
    .b(n4075),
    .c(net65),
    .d(net803),
    .o1(n3243));
 b15nandp2ah1n03x5 U4183 (.a(n3244),
    .b(n3243),
    .o1(n3242));
 b15aoi022ah1n06x5 U4184 (.a(net71),
    .b(net64),
    .c(n4074),
    .d(n4080),
    .o1(n3218));
 b15aoi022aq1n08x5 U4185 (.a(net88),
    .b(net832),
    .c(n4068),
    .d(n4095),
    .o1(n3217));
 b15xor002al1n08x5 U4186 (.a(n3218),
    .b(n3217),
    .out0(n3222));
 b15xor002as1n06x5 U4187 (.a(n3220),
    .b(n3219),
    .out0(n3221));
 b15xor002as1n06x5 U4188 (.a(n3222),
    .b(n3221),
    .out0(n3223));
 b15xor002an1n16x5 U4189 (.a(net72),
    .b(n3223),
    .out0(n3225));
 b15xor002aq1n06x5 U4190 (.a(n3225),
    .b(n3224),
    .out0(n3240));
 b15ztpn00an1n08x5 PHY_34 ();
 b15aoi022ah1n06x5 U4192 (.a(net826),
    .b(net827),
    .c(net800),
    .d(n4084),
    .o1(n3227));
 b15aoi022ah1n06x5 U4193 (.a(net830),
    .b(net823),
    .c(net780),
    .d(n4070),
    .o1(n3226));
 b15xor002al1n08x5 U4194 (.a(n3227),
    .b(n3226),
    .out0(n3239));
 b15aoi022as1n12x5 U4195 (.a(net65),
    .b(net831),
    .c(n4069),
    .d(n4075),
    .o1(n3229));
 b15xor002aq1n06x5 U4196 (.a(n3229),
    .b(n3228),
    .out0(n3230));
 b15qgbxo2an1n10x5 U4197 (.a(n3231),
    .b(n3230),
    .out0(n3233));
 b15xor002an1n16x5 U4198 (.a(n3233),
    .b(n3232),
    .out0(n3234));
 b15xor002ah1n16x5 U4199 (.a(net105),
    .b(n3234),
    .out0(n3236));
 b15xor002ar1n16x5 U4200 (.a(n3236),
    .b(n3235),
    .out0(n3238));
 b15nandp3an1n03x5 U4201 (.a(n3240),
    .b(n3239),
    .c(n3238),
    .o1(n3237));
 b15oai013an1n12x5 U4202 (.a(n3237),
    .b(n3240),
    .c(n3239),
    .d(n3238),
    .o1(n3241));
 b15oai112as1n16x5 U4203 (.a(n3242),
    .b(n3241),
    .c(n3244),
    .d(n3243),
    .o1(n3245));
 b15oaoi13al1n02x5 U4204 (.a(n3245),
    .b(n3247),
    .c(n3249),
    .d(n3248),
    .o1(n3246));
 b15aoai13an1n03x5 U4205 (.a(n3246),
    .b(n3247),
    .c(n3249),
    .d(n3248),
    .o1(n3250));
 b15aoi112aq1n03x5 U4206 (.a(n3251),
    .b(n3250),
    .c(n3252),
    .d(n3256),
    .o1(n3253));
 b15oai112ah1n06x5 U4207 (.a(net367),
    .b(n3253),
    .c(n3256),
    .d(n3255),
    .o1(n3257));
 b15aoi112an1n06x5 U4208 (.a(n3258),
    .b(n3257),
    .c(n3261),
    .d(n3260),
    .o1(n3259));
 b15oai012as1n16x5 U4209 (.a(n3259),
    .b(n3261),
    .c(n3260),
    .o1(n3362));
 b15aoi022ar1n08x5 U4210 (.a(net52),
    .b(net50),
    .c(net95),
    .d(n3284),
    .o1(n3262));
 b15oai122aq1n12x5 U4211 (.a(n3262),
    .b(net53),
    .c(net51),
    .d(n3263),
    .e(net50),
    .o1(n3274));
 b15aoi012ar1n04x5 U4212 (.a(net96),
    .b(n3265),
    .c(n3264),
    .o1(n3266));
 b15oaoi13an1n08x5 U4213 (.a(n3266),
    .b(net96),
    .c(net91),
    .d(net90),
    .o1(n3272));
 b15nand02an1n08x5 U4214 (.a(n3267),
    .b(net44),
    .o1(n3755));
 b15oaoi13as1n04x5 U4215 (.a(n3755),
    .b(net40),
    .c(net96),
    .d(net39),
    .o1(n3270));
 b15nand02ah1n02x5 U4216 (.a(net51),
    .b(n3268),
    .o1(n3269));
 b15oai112an1n12x5 U4217 (.a(n3270),
    .b(n3269),
    .c(n3272),
    .d(n3271),
    .o1(n3273));
 b15nor004al1n08x5 U4218 (.a(n3275),
    .b(n3362),
    .c(n3274),
    .d(n3273),
    .o1(n3283));
 b15nor004an1n06x5 U4219 (.a(net91),
    .b(net92),
    .c(net93),
    .d(net90),
    .o1(n3277));
 b15aoi022aq1n02x5 U4220 (.a(net91),
    .b(net90),
    .c(net92),
    .d(net93),
    .o1(n3276));
 b15oaoi13ar1n08x5 U4221 (.a(net40),
    .b(n3276),
    .c(n3277),
    .d(net39),
    .o1(n3278));
 b15aoi112ah1n04x5 U4222 (.a(net41),
    .b(n3278),
    .c(net90),
    .d(n3279),
    .o1(n3281));
 b15orn002ar1n08x5 U4223 (.a(net41),
    .b(n3280),
    .o(n3756));
 b15oai013ar1n12x5 U4224 (.a(n3756),
    .b(net43),
    .c(net52),
    .d(n3281),
    .o1(n3282));
 b15oai112as1n16x5 U4225 (.a(n3283),
    .b(n3282),
    .c(n3285),
    .d(n3284),
    .o1(u_reg_u_reg_if_N46));
 b15nor003as1n04x5 U4226 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .b(gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .c(n3367),
    .o1(n3366));
 b15nor002al1n02x5 U4227 (.a(n3434),
    .b(n3439),
    .o1(n3287));
 b15norp02as1n48x5 U4228 (.a(n3297),
    .b(u_reg_u_reg_if_N46),
    .o1(n3482));
 b15aoi013as1n08x5 U4229 (.a(gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q),
    .b(n3286),
    .c(net55),
    .d(n3482),
    .o1(n3363));
 b15aoi012ar1n04x5 U4230 (.a(n3363),
    .b(n3366),
    .c(n3287),
    .o1(gen_alert_tx_0__u_prim_alert_sender_alert_test_set_d));
 b15inv000aq1n24x5 U4231 (.a(n3337),
    .o1(n3294));
 b15norp02al1n32x5 U4232 (.a(n3294),
    .b(n3361),
    .o1(n3288));
 b15ztpn00an1n08x5 PHY_33 ();
 b15ztpn00an1n08x5 PHY_32 ();
 b15nor002ar1n32x5 U4235 (.a(n3442),
    .b(n3294),
    .o1(n3289));
 b15ztpn00an1n08x5 PHY_31 ();
 b15ztpn00an1n08x5 PHY_30 ();
 b15aoi022al1n32x5 U4238 (.a(reg2hw_ctrl_en_input_filter__q__27_),
    .b(net401),
    .c(reg2hw_intr_ctrl_en_lvllow__q__27_),
    .d(net395),
    .o1(n3310));
 b15norp02as1n12x5 U4239 (.a(n3299),
    .b(n3294),
    .o1(n3290));
 b15ztpn00an1n08x5 PHY_29 ();
 b15ztpn00an1n08x5 PHY_28 ();
 b15nandp2as1n48x5 U4242 (.a(n3291),
    .b(net100),
    .o1(n3371));
 b15norp02as1n48x5 U4243 (.a(n3361),
    .b(n3371),
    .o1(n3292));
 b15ztpn00an1n08x5 PHY_27 ();
 b15ztpn00an1n08x5 PHY_26 ();
 b15aoi022ah1n24x5 U4246 (.a(net567),
    .b(net388),
    .c(reg2hw_intr_ctrl_en_rising__q__27_),
    .d(net451),
    .o1(n3309));
 b15nandp2ah1n48x5 U4247 (.a(n3372),
    .b(n3293),
    .o1(n3302));
 b15nor002as1n24x5 U4248 (.a(n3294),
    .b(n3302),
    .o1(n3295));
 b15ztpn00an1n08x5 PHY_25 ();
 b15norp02as1n48x5 U4251 (.a(n3302),
    .b(n3371),
    .o1(n3982));
 b15aoi022aq1n12x5 U4252 (.a(net583),
    .b(net385),
    .c(net704),
    .d(net445),
    .o1(n3308));
 b15nandp2as1n48x5 U4253 (.a(net99),
    .b(n3296),
    .o1(n3759));
 b15norp02an1n24x5 U4254 (.a(n3299),
    .b(n3759),
    .o1(n3981));
 b15nanb02an1n04x5 U4255 (.a(u_reg_u_reg_if_N46),
    .b(n3297),
    .out0(n3298));
 b15ztpn00an1n08x5 PHY_24 ();
 b15norp02as1n48x5 U4258 (.a(n3300),
    .b(n3302),
    .o1(n3953));
 b15ztpn00an1n08x5 PHY_23 ();
 b15norp02as1n48x5 U4260 (.a(n3300),
    .b(n3299),
    .o1(n3301));
 b15ztpn00an1n08x5 PHY_22 ();
 b15nor002ah1n32x5 U4263 (.a(n3302),
    .b(n3759),
    .o1(n3303));
 b15ztpn00an1n08x5 PHY_21 ();
 b15aoi022ah1n04x5 U4266 (.a(net430),
    .b(reg2hw_intr_enable__q__27_),
    .c(net427),
    .d(net2342),
    .o1(n3304));
 b15oai012ar1n12x5 U4267 (.a(n3304),
    .b(n4123),
    .c(n3305),
    .o1(n3306));
 b15aoi112ah1n08x5 U4268 (.a(net361),
    .b(n3306),
    .c(net444),
    .d(net662),
    .o1(n3307));
 b15nand04ar1n12x5 U4269 (.a(n3310),
    .b(n3309),
    .c(n3308),
    .d(n3307),
    .o1(u_reg_u_reg_if_N41));
 b15aoi022aq1n08x5 U4270 (.a(net608),
    .b(net403),
    .c(reg2hw_intr_ctrl_en_rising__q__30_),
    .d(net451),
    .o1(n3317));
 b15ztpn00an1n08x5 PHY_20 ();
 b15aoi022aq1n08x5 U4272 (.a(reg2hw_intr_ctrl_en_lvllow__q__30_),
    .b(net397),
    .c(net442),
    .d(net651),
    .o1(n3316));
 b15ztpn00an1n08x5 PHY_19 ();
 b15aoi022an1n08x5 U4274 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__30_),
    .b(net388),
    .c(reg2hw_intr_ctrl_en_falling__q__30_),
    .d(net386),
    .o1(n3315));
 b15aoi022an1n16x5 U4275 (.a(net430),
    .b(reg2hw_intr_enable__q__30_),
    .c(net425),
    .d(net2370),
    .o1(n3311));
 b15oai012an1n24x5 U4276 (.a(n3311),
    .b(n4123),
    .c(n3312),
    .o1(n3313));
 b15aoi112as1n08x5 U4277 (.a(net363),
    .b(n3313),
    .c(net164),
    .d(net447),
    .o1(n3314));
 b15nand04as1n16x5 U4278 (.a(n3317),
    .b(n3316),
    .c(n3315),
    .d(n3314),
    .o1(u_reg_u_reg_if_N44));
 b15aoi022as1n06x5 U4279 (.a(reg2hw_ctrl_en_input_filter__q__31_),
    .b(net402),
    .c(reg2hw_intr_ctrl_en_lvllow__q__31_),
    .d(net395),
    .o1(n3324));
 b15ztpn00an1n08x5 PHY_18 ();
 b15aoi022ar1n16x5 U4281 (.a(reg2hw_intr_ctrl_en_rising__q__31_),
    .b(net451),
    .c(net426),
    .d(net2193),
    .o1(n3323));
 b15aoi022ar1n24x5 U4282 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__31_),
    .b(net388),
    .c(reg2hw_intr_ctrl_en_falling__q__31_),
    .d(net386),
    .o1(n3322));
 b15ztpn00an1n08x5 PHY_17 ();
 b15aoi022aq1n12x5 U4284 (.a(net442),
    .b(net197),
    .c(net430),
    .d(reg2hw_intr_enable__q__31_),
    .o1(n3318));
 b15oai012ah1n12x5 U4285 (.a(n3318),
    .b(n4123),
    .c(n3319),
    .o1(n3320));
 b15aoi112as1n08x5 U4286 (.a(net361),
    .b(n3320),
    .c(net698),
    .d(net446),
    .o1(n3321));
 b15nand04as1n16x5 U4287 (.a(n3324),
    .b(net2194),
    .c(n3322),
    .d(n3321),
    .o1(u_reg_u_reg_if_N45));
 b15aoi022as1n04x5 U4288 (.a(net589),
    .b(net386),
    .c(net430),
    .d(reg2hw_intr_enable__q__19_),
    .o1(n3332));
 b15ztpn00an1n08x5 PHY_16 ();
 b15aoi022ah1n08x5 U4290 (.a(reg2hw_intr_ctrl_en_rising__q__19_),
    .b(net451),
    .c(net2294),
    .d(net395),
    .o1(n3331));
 b15ztpn00an1n08x5 PHY_15 ();
 b15aoi022ah1n04x5 U4292 (.a(net628),
    .b(net402),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__19_),
    .d(net388),
    .o1(n3330));
 b15ztpn00an1n08x5 PHY_14 ();
 b15aoi022ah1n16x5 U4295 (.a(net441),
    .b(net183),
    .c(net426),
    .d(u_reg_data_in_qs[19]),
    .o1(n3326));
 b15oai012ar1n08x5 U4296 (.a(n3326),
    .b(n4123),
    .c(n3327),
    .o1(n3328));
 b15aoi112ar1n08x5 U4297 (.a(net361),
    .b(n3328),
    .c(net715),
    .d(net446),
    .o1(n3329));
 b15nand04ah1n12x5 U4298 (.a(n3332),
    .b(net2295),
    .c(n3330),
    .d(n3329),
    .o1(u_reg_u_reg_if_N33));
 b15nandp2aq1n48x5 U4299 (.a(n3482),
    .b(net451),
    .o1(n3333));
 b15ztpn00an1n08x5 PHY_13 ();
 b15ztpn00an1n08x5 PHY_12 ();
 b15nand02ar1n16x5 U4302 (.a(n3482),
    .b(n3295),
    .o1(n3334));
 b15ztpn00an1n08x5 PHY_11 ();
 b15ztpn00an1n08x5 PHY_10 ();
 b15nandp2aq1n24x5 U4305 (.a(n3482),
    .b(net403),
    .o1(n3335));
 b15ztpn00an1n08x5 PHY_9 ();
 b15nand02an1n32x5 U4308 (.a(n3482),
    .b(net394),
    .o1(n3336));
 b15ztpn00an1n08x5 PHY_8 ();
 b15ztpn00an1n08x5 PHY_7 ();
 b15inv040an1n05x5 U4311 (.a(n3442),
    .o1(n3483));
 b15nandp3ar1n08x5 U4312 (.a(n3483),
    .b(n3337),
    .c(n3482),
    .o1(n3338));
 b15ztpn00an1n08x5 PHY_6 ();
 b15ztpn00an1n08x5 PHY_5 ();
 b15ztpn00an1n08x5 PHY_4 ();
 b15ztpn00an1n08x5 PHY_3 ();
 b15nor002ar1n08x5 U4317 (.a(net779),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[25]));
 b15ztpn00an1n08x5 PHY_2 ();
 b15ztpn00an1n08x5 PHY_1 ();
 b15nor002as1n03x5 U4320 (.a(net764),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[29]));
 b15ztpn00an1n08x5 PHY_0 ();
 b15norp02aq1n04x5 U4323 (.a(net765),
    .b(n3336),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[29]));
 b15nor002ar1n08x5 U4326 (.a(net764),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[29]));
 b15nor002ah1n02x5 U4327 (.a(net764),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[29]));
 b15nor002ah1n03x5 U4328 (.a(net779),
    .b(net350),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[25]));
 b15nor002ar1n06x5 U4329 (.a(n4090),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[25]));
 b15norp02aq1n03x5 U4330 (.a(net779),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[25]));
 b15nor002ar1n06x5 U4331 (.a(net762),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[30]));
 b15norp02aq1n02x5 U4332 (.a(net776),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[26]));
 b15norp02ah1n04x5 U4333 (.a(net783),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[24]));
 b15norp02aq1n03x5 U4334 (.a(net773),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[27]));
 b15nor002ar1n04x5 U4335 (.a(net763),
    .b(net350),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[30]));
 b15norp02al1n04x5 U4336 (.a(net759),
    .b(net354),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[31]));
 b15norp02al1n04x5 U4337 (.a(net759),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[31]));
 b15nor002an1n03x5 U4338 (.a(net775),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[26]));
 b15nor002ar1n04x5 U4339 (.a(net773),
    .b(net350),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[27]));
 b15nor002an1n04x5 U4340 (.a(net776),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[26]));
 b15norp02ar1n04x5 U4341 (.a(net762),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[30]));
 b15norp02ar1n02x5 U4342 (.a(net773),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[27]));
 b15norp02as1n03x5 U4343 (.a(net772),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[27]));
 b15nor002an1n03x5 U4344 (.a(net776),
    .b(net350),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[26]));
 b15nor002ar1n08x5 U4345 (.a(net782),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[24]));
 b15nor002al1n03x5 U4346 (.a(net783),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[24]));
 b15nor002aq1n03x5 U4347 (.a(net760),
    .b(net350),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[31]));
 b15nor002an1n04x5 U4348 (.a(net783),
    .b(n3336),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[24]));
 b15nor002ah1n04x5 U4349 (.a(net763),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[30]));
 b15norp02ar1n04x5 U4350 (.a(net759),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[31]));
 b15norp02aq1n03x5 U4351 (.a(net769),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[28]));
 b15nor002as1n03x5 U4352 (.a(net769),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[28]));
 b15nor002al1n04x5 U4353 (.a(net768),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[28]));
 b15nor002aq1n04x5 U4354 (.a(net768),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[28]));
 b15norp02as1n03x5 U4356 (.a(n4077),
    .b(net355),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[11]));
 b15qgbno2an1n05x5 U4358 (.o1(u_reg_u_ctrl_en_input_filter_wr_data[4]),
    .a(net757),
    .b(net352));
 b15nor002an1n04x5 U4359 (.a(net756),
    .b(net355),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[4]));
 b15norp02an1n04x5 U4360 (.a(n4077),
    .b(net352),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[11]));
 b15qgbno2an1n10x5 U4362 (.a(n3524),
    .b(net352),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[13]));
 b15nor002aq1n03x5 U4364 (.a(n4077),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[11]));
 b15norp02an1n04x5 U4365 (.a(net756),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[4]));
 b15nor002as1n03x5 U4367 (.a(n3524),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[13]));
 b15norp02as1n03x5 U4369 (.a(n3524),
    .b(net355),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[13]));
 b15nor002aq1n03x5 U4371 (.a(n4077),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[11]));
 b15nor002as1n04x5 U4372 (.a(net756),
    .b(net350),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[4]));
 b15norp02ah1n03x5 U4374 (.a(n3524),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[13]));
 b15norp02an1n03x5 U4375 (.a(net811),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[12]));
 b15nor002aq1n04x5 U4376 (.a(n4071),
    .b(net355),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[5]));
 b15nor002ah1n04x5 U4377 (.a(n4071),
    .b(net352),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[5]));
 b15nor002ah1n04x5 U4378 (.a(net809),
    .b(net352),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[14]));
 b15nor002an1n03x5 U4379 (.a(net812),
    .b(net355),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[12]));
 b15nor002ar1n06x5 U4380 (.a(n4075),
    .b(net352),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[9]));
 b15norp02an1n04x5 U4381 (.a(net820),
    .b(n3335),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[0]));
 b15nor002aq1n03x5 U4382 (.a(n4072),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[6]));
 b15norp02an1n03x5 U4383 (.a(net814),
    .b(net352),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[7]));
 b15nor002an1n03x5 U4384 (.a(n4072),
    .b(net352),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[6]));
 b15norp02as1n03x5 U4385 (.a(net811),
    .b(net350),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[12]));
 b15norp02an1n03x5 U4386 (.a(n4072),
    .b(n3333),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[6]));
 b15nor002an1n04x5 U4387 (.a(n4075),
    .b(net355),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[9]));
 b15norp02ar1n12x5 U4388 (.a(n4078),
    .b(net352),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[12]));
 b15norp02as1n03x5 U4389 (.a(net817),
    .b(n3335),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[1]));
 b15norp02an1n04x5 U4390 (.a(net818),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[1]));
 b15norp02an1n04x5 U4391 (.a(n4075),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[9]));
 b15norp02aq1n03x5 U4392 (.a(net818),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[1]));
 b15nor002an1n03x5 U4393 (.a(n4074),
    .b(net352),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[8]));
 b15nor002as1n03x5 U4394 (.a(n4080),
    .b(net352),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[15]));
 b15norp02aq1n04x5 U4395 (.a(n4080),
    .b(net355),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[15]));
 b15nor002ar1n04x5 U4396 (.a(n4074),
    .b(net355),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[8]));
 b15nor002ah1n02x5 U4397 (.a(n4080),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[15]));
 b15norp02ar1n08x5 U4398 (.a(n4076),
    .b(net352),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[10]));
 b15nor002aq1n03x5 U4399 (.a(n4072),
    .b(net356),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[6]));
 b15norp02aq1n04x5 U4400 (.a(n4079),
    .b(net355),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[14]));
 b15norp02aq1n04x5 U4401 (.a(n4074),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[8]));
 b15nor002an1n08x5 U4402 (.a(n4069),
    .b(net352),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[2]));
 b15nor002ar1n04x5 U4403 (.a(net813),
    .b(net355),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[7]));
 b15nor002aq1n03x5 U4404 (.a(net818),
    .b(net355),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[1]));
 b15norp02an1n04x5 U4405 (.a(n4076),
    .b(net355),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[10]));
 b15norp02as1n03x5 U4406 (.a(n4076),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[10]));
 b15nor002an1n03x5 U4407 (.a(net813),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[7]));
 b15norp02aq1n03x5 U4408 (.a(net819),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[0]));
 b15nor002ah1n04x5 U4409 (.a(n4069),
    .b(net356),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[2]));
 b15nor002ar1n03x5 U4410 (.a(net809),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[14]));
 b15nor002an1n06x5 U4411 (.a(n4071),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[5]));
 b15nor002al1n03x5 U4412 (.a(n4071),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[5]));
 b15norp02aq1n03x5 U4413 (.a(n4069),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[2]));
 b15nor002ar1n06x5 U4414 (.a(net819),
    .b(net350),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[0]));
 b15nor002an1n03x5 U4415 (.a(n4073),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[7]));
 b15nor002as1n02x5 U4416 (.a(n4080),
    .b(net350),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[15]));
 b15norp02aq1n03x5 U4417 (.a(net808),
    .b(net350),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[14]));
 b15nor002ah1n04x5 U4418 (.a(net819),
    .b(net355),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[0]));
 b15norp02aq1n04x5 U4419 (.a(n4075),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[9]));
 b15norp02al1n04x5 U4420 (.a(n4076),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[10]));
 b15nor002ar1n06x5 U4421 (.a(n4074),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[8]));
 b15nor002as1n03x5 U4422 (.a(n4069),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[2]));
 b15nor002al1n04x5 U4423 (.a(n4070),
    .b(net352),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[3]));
 b15norp02an1n03x5 U4424 (.a(net816),
    .b(net355),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[3]));
 b15norp02ah1n03x5 U4425 (.a(n4070),
    .b(net357),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[3]));
 b15nor002an1n04x5 U4426 (.a(net816),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[3]));
 b15norp02al1n04x5 U4427 (.a(net784),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[23]));
 b15nor002ah1n02x5 U4428 (.a(net797),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[19]));
 b15norp02al1n04x5 U4429 (.a(net806),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[16]));
 b15norp02as1n04x5 U4430 (.a(net793),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[20]));
 b15nor002an1n08x5 U4431 (.a(net795),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[20]));
 b15nor002an1n06x5 U4432 (.a(net784),
    .b(net350),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[23]));
 b15norp02an1n04x5 U4433 (.a(n4081),
    .b(net350),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[16]));
 b15norp02al1n08x5 U4434 (.a(net806),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[16]));
 b15norp02aq1n08x5 U4435 (.a(net806),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[16]));
 b15nor002aq1n02x5 U4436 (.a(net794),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[20]));
 b15norp02al1n04x5 U4437 (.a(n4084),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[19]));
 b15nor002al1n04x5 U4438 (.a(net798),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[19]));
 b15nor002an1n03x5 U4439 (.a(net785),
    .b(net352),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[23]));
 b15norp02as1n03x5 U4440 (.a(net794),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[20]));
 b15norp02aq1n03x5 U4441 (.a(net796),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[19]));
 b15norp02aq1n04x5 U4442 (.a(net785),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[23]));
 b15nor002an1n03x5 U4443 (.a(net800),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[18]));
 b15norp02aq1n03x5 U4444 (.a(net791),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[21]));
 b15nor002as1n04x5 U4445 (.a(net788),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[22]));
 b15norp02ar1n08x5 U4446 (.a(net792),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[21]));
 b15norp02aq1n04x5 U4447 (.a(net801),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[18]));
 b15norp02as1n03x5 U4448 (.a(net804),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[17]));
 b15norp02aq1n03x5 U4449 (.a(net803),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[17]));
 b15nor002an1n03x5 U4450 (.a(net803),
    .b(net350),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[17]));
 b15norp02as1n03x5 U4451 (.a(net788),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[22]));
 b15nor002as1n04x5 U4452 (.a(net790),
    .b(net349),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[21]));
 b15nor002an1n06x5 U4453 (.a(net787),
    .b(net350),
    .o1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[22]));
 b15nor002as1n03x5 U4454 (.a(net801),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[18]));
 b15nor002ar1n04x5 U4455 (.a(net792),
    .b(net353),
    .o1(u_reg_u_intr_ctrl_en_falling_wr_data[21]));
 b15norp02aq1n04x5 U4456 (.a(net799),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[18]));
 b15nor002aq1n04x5 U4457 (.a(net804),
    .b(net351),
    .o1(u_reg_u_ctrl_en_input_filter_wr_data[17]));
 b15norp02aq1n03x5 U4458 (.a(net787),
    .b(net358),
    .o1(u_reg_u_intr_ctrl_en_rising_wr_data[22]));
 b15nand02ah1n48x5 U4459 (.a(n3482),
    .b(n3301),
    .o1(n3359));
 b15norp02as1n04x5 U4462 (.a(n3524),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[13]));
 b15norp02as1n03x5 U4465 (.a(n3538),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[4]));
 b15norp02an1n04x5 U4466 (.a(n4077),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[11]));
 b15nor002ar1n04x5 U4467 (.a(net814),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[7]));
 b15nor002aq1n03x5 U4468 (.a(n4074),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[8]));
 b15nor002as1n03x5 U4469 (.a(n4076),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[10]));
 b15norp02as1n04x5 U4470 (.a(n4078),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[12]));
 b15norp02aq1n04x5 U4471 (.a(n4080),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[15]));
 b15norp02al1n04x5 U4472 (.a(n4068),
    .b(n3359),
    .o1(u_reg_u_intr_enable_wr_data[1]));
 b15nor002al1n04x5 U4473 (.a(n4069),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[2]));
 b15nor002an1n03x5 U4474 (.a(n4075),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[9]));
 b15norp02aq1n04x5 U4475 (.a(net809),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[14]));
 b15nor002as1n04x5 U4476 (.a(n4072),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[6]));
 b15nor002aq1n03x5 U4477 (.a(net820),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[0]));
 b15norp02as1n03x5 U4478 (.a(n4071),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[5]));
 b15norp02as1n04x5 U4479 (.a(n4070),
    .b(net344),
    .o1(u_reg_u_intr_enable_wr_data[3]));
 b15norp02ah1n03x5 U4480 (.a(net795),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[20]));
 b15nor002ar1n03x5 U4481 (.a(net797),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[19]));
 b15nor002aq1n03x5 U4482 (.a(net806),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[16]));
 b15nor002ar1n08x5 U4483 (.a(net785),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[23]));
 b15norp02aq1n03x5 U4484 (.a(net804),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[17]));
 b15nor002ah1n02x5 U4485 (.a(net799),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[18]));
 b15norp02ah1n03x5 U4486 (.a(net792),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[21]));
 b15nor002an1n04x5 U4487 (.a(net788),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[22]));
 b15nor002ah1n04x5 U4490 (.a(n4090),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[25]));
 b15nor002as1n03x5 U4491 (.a(net764),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[29]));
 b15nor002aq1n03x5 U4492 (.a(net772),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[27]));
 b15norp02as1n02x5 U4493 (.a(net775),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[26]));
 b15nor002ar1n06x5 U4494 (.a(net782),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[24]));
 b15nor002aq1n02x5 U4495 (.a(net762),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[30]));
 b15nor002aq1n04x5 U4496 (.a(net759),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[31]));
 b15norp02al1n04x5 U4497 (.a(net768),
    .b(net345),
    .o1(u_reg_u_intr_enable_wr_data[28]));
 b15nandp2as1n48x5 U4498 (.a(n3482),
    .b(net444),
    .o1(n3443));
 b15norp02ar1n48x5 U4500 (.a(n3361),
    .b(n3759),
    .o1(n3870));
 b15nand02ar1n24x5 U4501 (.a(n3482),
    .b(net418),
    .o1(n3389));
 b15nand02as1n06x5 U4502 (.a(net341),
    .b(net330),
    .o1(N55));
 b15ao0012ah1n04x5 U4503 (.a(net2446),
    .b(net44),
    .c(n3362),
    .o(n1439));
 b15orn002an1n03x5 U4504 (.a(net2318),
    .b(n1439),
    .o(gen_alert_tx_0__u_prim_alert_sender_alert_req_trigger));
 b15nonb02al1n06x5 U4505 (.a(n3363),
    .b(gen_alert_tx_0__u_prim_alert_sender_alert_req_trigger),
    .out0(n3433));
 b15nor003al1n08x5 U4506 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .b(n3364),
    .c(gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .o1(n3437));
 b15aoi022ar1n02x5 U4507 (.a(n3433),
    .b(n3437),
    .c(n3365),
    .d(gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .o1(n3370));
 b15orn002ar1n02x5 U4508 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .b(gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .o(n3368));
 b15aoi112al1n03x5 U4509 (.a(n3366),
    .b(n3435),
    .c(n3368),
    .d(n3367),
    .o1(n3369));
 b15aoi112an1n03x5 U4510 (.a(n3369),
    .b(n3439),
    .c(n3370),
    .d(n3435),
    .o1(gen_alert_tx_0__u_prim_alert_sender_state_d[1]));
 b15norp02ar1n48x5 U4511 (.a(n3371),
    .b(net98),
    .o1(n3871));
 b15and002as1n24x5 U4512 (.a(net417),
    .b(n3482),
    .o(N113));
 b15nor002ah1n16x5 U4513 (.a(n3442),
    .b(n3371),
    .o1(n3877));
 b15nand02al1n24x5 U4514 (.a(n3482),
    .b(net410),
    .o1(n3431));
 b15nand02aq1n32x5 U4515 (.a(N113),
    .b(n3372),
    .o1(n3400));
 b15nand02an1n03x5 U4517 (.a(n3431),
    .b(n3400),
    .o1(N130));
 b15norp02as1n24x5 U4518 (.a(n4096),
    .b(n4080),
    .o1(n3466));
 b15aoi012aq1n16x5 U4519 (.a(n3466),
    .b(net648),
    .c(net758),
    .o1(n3373));
 b15oai022an1n32x5 U4521 (.a(n3373),
    .b(net332),
    .c(net760),
    .d(net338),
    .o1(N71));
 b15aoi012as1n24x5 U4522 (.a(n3450),
    .b(net668),
    .c(net778),
    .o1(n3374));
 b15oai022as1n16x5 U4523 (.a(n3374),
    .b(net333),
    .c(net779),
    .d(net335),
    .o1(N65));
 b15norp02as1n24x5 U4524 (.a(net815),
    .b(net796),
    .o1(n3476));
 b15aoi012ar1n08x5 U4525 (.a(n3476),
    .b(net183),
    .c(net796),
    .o1(n3375));
 b15oai022aq1n08x5 U4526 (.a(n3375),
    .b(net331),
    .c(net796),
    .d(net342),
    .o1(N59));
 b15nor002as1n06x5 U4527 (.a(n4088),
    .b(net814),
    .o1(n3473));
 b15aoi012ah1n06x5 U4528 (.a(n3473),
    .b(net673),
    .c(n4088),
    .o1(n3376));
 b15oai022aq1n16x5 U4529 (.a(n3376),
    .b(net333),
    .c(n4088),
    .d(net343),
    .o1(N63));
 b15aoi012ah1n32x5 U4530 (.a(n3460),
    .b(net656),
    .c(n4094),
    .o1(n3377));
 b15oai022as1n16x5 U4531 (.a(n3377),
    .b(net332),
    .c(net766),
    .d(net340),
    .o1(N69));
 b15norp02as1n24x5 U4532 (.a(n4067),
    .b(net806),
    .o1(n3456));
 b15aoi012as1n02x5 U4533 (.a(n3456),
    .b(net685),
    .c(net807),
    .o1(n3378));
 b15oai022an1n02x5 U4534 (.a(n3378),
    .b(net329),
    .c(net807),
    .d(net339),
    .o1(N56));
 b15aoi012an1n24x5 U4535 (.a(net736),
    .b(net185),
    .c(net793),
    .o1(n3379));
 b15oai022ar1n32x5 U4536 (.a(n3379),
    .b(net332),
    .c(net793),
    .d(net337),
    .o1(N60));
 b15norp02al1n16x5 U4537 (.a(net771),
    .b(n4077),
    .o1(n3448));
 b15aoi012aq1n16x5 U4538 (.a(net735),
    .b(net661),
    .c(net772),
    .o1(n3380));
 b15oai022as1n32x5 U4539 (.a(n3380),
    .b(net330),
    .c(net772),
    .d(net341),
    .o1(N67));
 b15nor002ar1n08x5 U4540 (.a(net786),
    .b(n4072),
    .o1(n3471));
 b15aoi012ar1n08x5 U4541 (.a(n3471),
    .b(net678),
    .c(net786),
    .o1(n3381));
 b15oai022aq1n16x5 U4542 (.a(n3381),
    .b(net333),
    .c(net786),
    .d(net336),
    .o1(N62));
 b15norp02as1n32x5 U4543 (.a(net805),
    .b(net817),
    .o1(n3452));
 b15aoi012al1n04x5 U4544 (.a(n3452),
    .b(net2313),
    .c(net802),
    .o1(n3382));
 b15oai022ah1n04x5 U4545 (.a(n3382),
    .b(net329),
    .c(net802),
    .d(net339),
    .o1(N57));
 b15norp02al1n48x5 U4546 (.a(n4071),
    .b(net792),
    .o1(n3446));
 b15aoi012al1n04x5 U4547 (.a(n3446),
    .b(net186),
    .c(net790),
    .o1(n3383));
 b15oai022as1n02x5 U4548 (.a(n3383),
    .b(net334),
    .c(net790),
    .d(net337),
    .o1(N61));
 b15norp02ar1n48x5 U4549 (.a(net763),
    .b(net808),
    .o1(n3458));
 b15aoi012aq1n12x5 U4550 (.a(n3458),
    .b(net651),
    .c(net762),
    .o1(n3384));
 b15oai022aq1n12x5 U4551 (.a(n3384),
    .b(net332),
    .c(net763),
    .d(net338),
    .o1(N70));
 b15nor002ah1n16x5 U4552 (.a(net801),
    .b(n4069),
    .o1(n3468));
 b15aoi012an1n16x5 U4553 (.a(n3468),
    .b(net680),
    .c(net801),
    .o1(n3385));
 b15oai022ah1n04x5 U4554 (.a(n3385),
    .b(net331),
    .c(net799),
    .d(net342),
    .o1(N58));
 b15nor002ah1n16x5 U4555 (.a(net774),
    .b(n4076),
    .o1(n3464));
 b15aoi012ah1n12x5 U4556 (.a(net734),
    .b(net664),
    .c(net775),
    .o1(n3386));
 b15oai022as1n32x5 U4557 (.a(n3386),
    .b(net330),
    .c(net775),
    .d(net341),
    .o1(N66));
 b15nor002aq1n04x5 U4558 (.a(n4074),
    .b(net783),
    .o1(n3444));
 b15aoi012an1n16x5 U4559 (.a(net733),
    .b(net670),
    .c(net783),
    .o1(n3387));
 b15oai022al1n16x5 U4560 (.a(n3387),
    .b(net329),
    .c(net781),
    .d(net340),
    .o1(N64));
 b15norp02an1n04x5 U4561 (.a(net812),
    .b(net770),
    .o1(n3454));
 b15aoi012as1n02x5 U4562 (.a(net732),
    .b(net659),
    .c(net768),
    .o1(n3390));
 b15oai022ah1n02x5 U4563 (.a(n3390),
    .b(net331),
    .c(net768),
    .d(net342),
    .o1(N68));
 b15aoi022ar1n24x5 U4564 (.a(net73),
    .b(net55),
    .c(net723),
    .d(net807),
    .o1(n3392));
 b15oai022aq1n08x5 U4566 (.a(n3392),
    .b(net325),
    .c(net807),
    .d(n3400),
    .o1(N131));
 b15nor002aq1n04x5 U4569 (.a(net779),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[25]));
 b15nor002aq1n03x5 U4570 (.a(net764),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[29]));
 b15nor002aq1n03x5 U4571 (.a(net759),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[31]));
 b15norp02as1n03x5 U4572 (.a(net782),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[24]));
 b15nor002an1n04x5 U4573 (.a(net772),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[27]));
 b15norp02as1n03x5 U4574 (.a(net775),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[26]));
 b15norp02as1n03x5 U4575 (.a(net762),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[30]));
 b15nor002aq1n03x5 U4576 (.a(net769),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[28]));
 b15nor002as1n04x5 U4578 (.a(n3524),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[13]));
 b15nor002as1n03x5 U4580 (.a(net756),
    .b(net348),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[4]));
 b15nor002as1n03x5 U4581 (.a(n4077),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[11]));
 b15nor002aq1n03x5 U4582 (.a(net813),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[7]));
 b15nor002as1n03x5 U4583 (.a(n4071),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[5]));
 b15nor002an1n03x5 U4584 (.a(n4080),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[15]));
 b15norp02as1n03x5 U4585 (.a(n4075),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[9]));
 b15norp02as1n03x5 U4586 (.a(net810),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[14]));
 b15nor002aq1n04x5 U4587 (.a(n4076),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[10]));
 b15norp02as1n03x5 U4588 (.a(net812),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[12]));
 b15norp02as1n03x5 U4589 (.a(n4069),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[2]));
 b15nor002al1n04x5 U4590 (.a(n4074),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[8]));
 b15norp02aq1n04x5 U4591 (.a(n4072),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[6]));
 b15norp02al1n08x5 U4592 (.a(net818),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[1]));
 b15norp02ah1n04x5 U4593 (.a(net819),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[0]));
 b15norp02as1n03x5 U4594 (.a(net816),
    .b(net346),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[3]));
 b15norp02aq1n04x5 U4595 (.a(net794),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[20]));
 b15norp02an1n03x5 U4596 (.a(net796),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[19]));
 b15nor002an1n03x5 U4597 (.a(net784),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[23]));
 b15norp02as1n03x5 U4598 (.a(net806),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[16]));
 b15norp02as1n03x5 U4599 (.a(net791),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[21]));
 b15norp02aq1n03x5 U4600 (.a(net804),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[17]));
 b15nor002aq1n03x5 U4601 (.a(net787),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[22]));
 b15nor002ar1n03x5 U4602 (.a(net799),
    .b(net347),
    .o1(u_reg_u_intr_ctrl_en_lvllow_wr_data[18]));
 b15aoi012aq1n08x5 U4603 (.a(n3462),
    .b(net696),
    .c(net795),
    .o1(n3397));
 b15nandp2as1n48x5 U4604 (.a(net97),
    .b(N113),
    .o1(n3414));
 b15oai022aq1n24x5 U4605 (.a(n3397),
    .b(n3414),
    .c(net757),
    .d(net311),
    .o1(N118));
 b15aoi012as1n02x5 U4606 (.a(n3460),
    .b(net145),
    .c(n4094),
    .o1(n3398));
 b15oai022an1n08x5 U4607 (.a(n3398),
    .b(n3414),
    .c(n3524),
    .d(net309),
    .o1(N127));
 b15aoi022ah1n06x5 U4608 (.a(net85),
    .b(net67),
    .c(net143),
    .d(net771),
    .o1(n3399));
 b15oai022al1n08x5 U4609 (.a(n3399),
    .b(n3414),
    .c(n4077),
    .d(net309),
    .o1(N125));
 b15aoi022ar1n24x5 U4610 (.a(net73),
    .b(net55),
    .c(net141),
    .d(net807),
    .o1(n3401));
 b15oai022al1n12x5 U4612 (.a(n3401),
    .b(n3414),
    .c(net820),
    .d(net311),
    .o1(N114));
 b15aoi022ar1n32x5 U4613 (.a(net88),
    .b(net70),
    .c(net727),
    .d(net761),
    .o1(n3402));
 b15oai022aq1n24x5 U4614 (.a(n3402),
    .b(n3414),
    .c(net810),
    .d(net309),
    .o1(N128));
 b15aoi022as1n02x5 U4615 (.a(net80),
    .b(net63),
    .c(net170),
    .d(n4088),
    .o1(n3403));
 b15oai022al1n02x5 U4616 (.a(n3403),
    .b(n3414),
    .c(n4073),
    .d(net313),
    .o1(N121));
 b15aoi012ah1n24x5 U4617 (.a(n3450),
    .b(net694),
    .c(net778),
    .o1(n3404));
 b15oai022aq1n06x5 U4618 (.a(n3404),
    .b(n3414),
    .c(n4075),
    .d(net313),
    .o1(N123));
 b15aoi022aq1n08x5 U4619 (.a(net79),
    .b(net62),
    .c(net169),
    .d(net786),
    .o1(n3405));
 b15oai022ah1n08x5 U4620 (.a(n3405),
    .b(n3414),
    .c(n4072),
    .d(net313),
    .o1(N120));
 b15aoi022ar1n04x5 U4621 (.a(net823),
    .b(net64),
    .c(net171),
    .d(n4089),
    .o1(n3406));
 b15oai022an1n02x5 U4622 (.a(n3406),
    .b(n3414),
    .c(n4074),
    .d(net313),
    .o1(N122));
 b15aoi022aq1n32x5 U4623 (.a(net74),
    .b(net56),
    .c(net152),
    .d(net802),
    .o1(n3407));
 b15oai022al1n24x5 U4624 (.a(n3407),
    .b(n3414),
    .c(net817),
    .d(net311),
    .o1(N115));
 b15aoi022aq1n02x5 U4625 (.a(net821),
    .b(net68),
    .c(net144),
    .d(net770),
    .o1(n3408));
 b15oai022as1n06x5 U4626 (.a(n3408),
    .b(n3414),
    .c(n4078),
    .d(net309),
    .o1(N126));
 b15aoi022as1n24x5 U4627 (.a(net89),
    .b(net71),
    .c(net725),
    .d(net758),
    .o1(n3409));
 b15oai022as1n16x5 U4628 (.a(n3409),
    .b(n3414),
    .c(n4080),
    .d(net313),
    .o1(N129));
 b15aoi022as1n32x5 U4629 (.a(net75),
    .b(net57),
    .c(net163),
    .d(net801),
    .o1(n3410));
 b15oai022ar1n32x5 U4630 (.a(n3410),
    .b(n3414),
    .c(n4069),
    .d(net308),
    .o1(N116));
 b15aoi022aq1n08x5 U4631 (.a(net84),
    .b(net66),
    .c(net142),
    .d(net774),
    .o1(n3411));
 b15oai022ah1n08x5 U4632 (.a(n3411),
    .b(n3414),
    .c(n4076),
    .d(net309),
    .o1(N124));
 b15aoi022al1n48x5 U4633 (.a(net78),
    .b(net60),
    .c(net168),
    .d(n4086),
    .o1(n3412));
 b15oai022as1n16x5 U4634 (.a(n3412),
    .b(n3414),
    .c(n4071),
    .d(net311),
    .o1(N119));
 b15aoi022ah1n48x5 U4635 (.a(net76),
    .b(net58),
    .c(net700),
    .d(net798),
    .o1(n3415));
 b15oai022ah1n24x5 U4636 (.a(n3415),
    .b(n3414),
    .c(net816),
    .d(net310),
    .o1(N117));
 b15aoi012ar1n06x5 U4637 (.a(n3450),
    .b(net708),
    .c(net779),
    .o1(n3416));
 b15oai022ah1n04x5 U4638 (.a(n3416),
    .b(net325),
    .c(net779),
    .d(net311),
    .o1(N140));
 b15aoi022as1n04x5 U4639 (.a(net80),
    .b(net63),
    .c(net2634),
    .d(n4088),
    .o1(n3417));
 b15oai022ah1n04x5 U4640 (.a(n3417),
    .b(net328),
    .c(n4088),
    .d(net313),
    .o1(N138));
 b15aoi012ar1n04x5 U4641 (.a(net736),
    .b(net153),
    .c(net793),
    .o1(n3418));
 b15oai022ah1n06x5 U4642 (.a(n3418),
    .b(net326),
    .c(net793),
    .d(net308),
    .o1(N135));
 b15aoi022an1n06x5 U4643 (.a(net826),
    .b(net830),
    .c(net716),
    .d(net798),
    .o1(n3419));
 b15oai022an1n08x5 U4644 (.a(n3419),
    .b(net326),
    .c(net798),
    .d(net308),
    .o1(N134));
 b15aoi012al1n04x5 U4645 (.a(n3460),
    .b(net162),
    .c(net765),
    .o1(n3420));
 b15oai022an1n08x5 U4646 (.a(n3420),
    .b(net327),
    .c(net765),
    .d(net310),
    .o1(N144));
 b15aoi022ar1n12x5 U4647 (.a(net84),
    .b(net66),
    .c(net159),
    .d(net774),
    .o1(n3421));
 b15oai022ar1n08x5 U4648 (.a(n3421),
    .b(net328),
    .c(net774),
    .d(net309),
    .o1(N141));
 b15aoi022an1n02x5 U4649 (.a(net85),
    .b(net67),
    .c(net160),
    .d(net771),
    .o1(n3422));
 b15oai022as1n02x5 U4650 (.a(n3422),
    .b(net328),
    .c(net771),
    .d(net309),
    .o1(N142));
 b15aoi022aq1n12x5 U4651 (.a(net828),
    .b(net56),
    .c(net149),
    .d(net802),
    .o1(n3423));
 b15oai022aq1n08x5 U4652 (.a(n3423),
    .b(net325),
    .c(net805),
    .d(net311),
    .o1(N132));
 b15aoi022ar1n02x5 U4653 (.a(net89),
    .b(net71),
    .c(net165),
    .d(net760),
    .o1(n3424));
 b15oai022ar1n02x5 U4654 (.a(n3424),
    .b(net327),
    .c(net760),
    .d(net312),
    .o1(N146));
 b15aoi022ar1n32x5 U4655 (.a(net827),
    .b(net831),
    .c(net718),
    .d(net801),
    .o1(n3425));
 b15oai022an1n24x5 U4656 (.a(n3425),
    .b(net327),
    .c(n4083),
    .d(net310),
    .o1(N133));
 b15aoi022an1n24x5 U4657 (.a(net823),
    .b(net64),
    .c(net709),
    .d(net780),
    .o1(n3426));
 b15oai022ah1n32x5 U4658 (.a(n3426),
    .b(net328),
    .c(net780),
    .d(net313),
    .o1(N139));
 b15aoi022as1n04x5 U4659 (.a(net79),
    .b(net62),
    .c(net713),
    .d(net786),
    .o1(n3427));
 b15oai022aq1n04x5 U4660 (.a(n3427),
    .b(net328),
    .c(net786),
    .d(net313),
    .o1(N137));
 b15aoi022an1n12x5 U4661 (.a(net88),
    .b(net70),
    .c(net699),
    .d(net761),
    .o1(n3428));
 b15oai022aq1n16x5 U4662 (.a(n3428),
    .b(net327),
    .c(net761),
    .d(net309),
    .o1(N145));
 b15aoi022as1n08x5 U4663 (.a(net825),
    .b(net829),
    .c(net154),
    .d(net790),
    .o1(n3429));
 b15oai022ar1n08x5 U4664 (.a(n3429),
    .b(net326),
    .c(net790),
    .d(net308),
    .o1(N136));
 b15aoi022ar1n12x5 U4665 (.a(net821),
    .b(net68),
    .c(net2232),
    .d(n4093),
    .o1(n3432));
 b15oai022ah1n04x5 U4666 (.a(n3432),
    .b(net327),
    .c(net767),
    .d(net310),
    .o1(N143));
 b15nor003ah1n04x5 U4667 (.a(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .b(gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .c(n3433),
    .o1(n3436));
 b15oaoi13as1n08x5 U4668 (.a(n3434),
    .b(n3435),
    .c(n3437),
    .d(n3436),
    .o1(n3441));
 b15norp02an1n02x5 U4669 (.a(n3441),
    .b(n3439),
    .o1(gen_alert_tx_0__u_prim_alert_sender_alert_pd));
 b15nonb02ar1n02x5 U4670 (.a(n3441),
    .b(n3439),
    .out0(gen_alert_tx_0__u_prim_alert_sender_alert_nd));
 b15inv000al1n02x5 U4671 (.a(n3438),
    .o1(n3440));
 b15aoi012aq1n02x5 U4672 (.a(n3439),
    .b(n3441),
    .c(n3440),
    .o1(gen_alert_tx_0__u_prim_alert_sender_state_d[0]));
 b15inv000ar1n20x5 U4673 (.a(n3482),
    .o1(n3481));
 b15norp03as1n24x5 U4674 (.a(n3442),
    .b(n3481),
    .c(n3759),
    .o1(n3475));
 b15nanb02ah1n16x5 U4676 (.a(net303),
    .b(net338),
    .out0(N38));
 b15aoai13as1n06x5 U4677 (.a(net302),
    .b(net733),
    .c(net203),
    .d(net781),
    .o1(n3445));
 b15oai012as1n32x5 U4678 (.a(net299),
    .b(n3443),
    .c(n4074),
    .o1(N47));
 b15aoai13as1n08x5 U4679 (.a(net305),
    .b(n3446),
    .c(net646),
    .d(net792),
    .o1(n3447));
 b15oai012an1n48x5 U4680 (.a(n3447),
    .b(net340),
    .c(n4071),
    .o1(N44));
 b15aoai13al1n04x5 U4681 (.a(net304),
    .b(n3448),
    .c(net175),
    .d(n4092),
    .o1(n3449));
 b15oai012ar1n12x5 U4682 (.a(n3449),
    .b(net338),
    .c(n4077),
    .o1(N50));
 b15aoai13as1n08x5 U4683 (.a(net302),
    .b(n3450),
    .c(net204),
    .d(net778),
    .o1(n3451));
 b15oai012ar1n48x5 U4684 (.a(n3451),
    .b(net340),
    .c(n4075),
    .o1(N48));
 b15aoai13as1n08x5 U4685 (.a(n3475),
    .b(n3452),
    .c(net184),
    .d(n4082),
    .o1(n3453));
 b15oai012ah1n24x5 U4686 (.a(n3453),
    .b(net343),
    .c(net817),
    .o1(N40));
 b15aoai13as1n02x5 U4687 (.a(net304),
    .b(net732),
    .c(net176),
    .d(n4093),
    .o1(n3455));
 b15oai012al1n04x5 U4688 (.a(n3455),
    .b(n3443),
    .c(net812),
    .o1(N51));
 b15aoai13as1n08x5 U4689 (.a(net302),
    .b(n3456),
    .c(net173),
    .d(net807),
    .o1(n3457));
 b15oai012an1n32x5 U4690 (.a(n3457),
    .b(net339),
    .c(n4067),
    .o1(N39));
 b15aoai13al1n08x5 U4691 (.a(net303),
    .b(n3458),
    .c(net178),
    .d(net763),
    .o1(n3459));
 b15oai012ar1n16x5 U4692 (.a(n3459),
    .b(net337),
    .c(net808),
    .o1(N53));
 b15aoai13aq1n03x5 U4693 (.a(net304),
    .b(n3460),
    .c(net177),
    .d(n4094),
    .o1(n3461));
 b15oai012ar1n03x5 U4694 (.a(n3461),
    .b(net336),
    .c(n3524),
    .o1(N52));
 b15aoai13as1n08x5 U4695 (.a(net302),
    .b(n3462),
    .c(net199),
    .d(n4085),
    .o1(n3463));
 b15oai012as1n32x5 U4696 (.a(n3463),
    .b(n3443),
    .c(net757),
    .o1(N43));
 b15aoai13al1n08x5 U4697 (.a(net304),
    .b(n3464),
    .c(net691),
    .d(net774),
    .o1(n3465));
 b15oai012an1n12x5 U4698 (.a(n3465),
    .b(net338),
    .c(n4076),
    .o1(N49));
 b15aoai13as1n08x5 U4699 (.a(net303),
    .b(n3466),
    .c(net686),
    .d(net760),
    .o1(n3467));
 b15oai012ar1n24x5 U4700 (.a(n3467),
    .b(net337),
    .c(n4080),
    .o1(N54));
 b15aoai13as1n08x5 U4701 (.a(net303),
    .b(n3468),
    .c(net655),
    .d(net801),
    .o1(n3469));
 b15oai012ah1n12x5 U4702 (.a(n3469),
    .b(net337),
    .c(n4069),
    .o1(N41));
 b15aoai13ar1n03x5 U4703 (.a(net304),
    .b(n3471),
    .c(net201),
    .d(net786),
    .o1(n3472));
 b15oai012ar1n02x5 U4704 (.a(n3472),
    .b(net336),
    .c(n4072),
    .o1(N45));
 b15aoai13aq1n03x5 U4705 (.a(net304),
    .b(n3473),
    .c(net202),
    .d(n4088),
    .o1(n3474));
 b15oai012al1n03x5 U4706 (.a(n3474),
    .b(net336),
    .c(net814),
    .o1(N46));
 b15aoai13as1n08x5 U4707 (.a(net303),
    .b(n3476),
    .c(net652),
    .d(net798),
    .o1(n3477));
 b15oai012al1n32x5 U4708 (.a(n3477),
    .b(net337),
    .c(net816),
    .o1(N42));
 b15inv000ah1n02x5 U4709 (.a(gen_filter_11__u_filter_filter_synced),
    .o1(n3480));
 b15nand02ar1n04x5 U4710 (.a(net638),
    .b(gen_filter_11__u_filter_stored_value_q),
    .o1(n3479));
 b15oai012ar1n08x5 U4711 (.a(n3479),
    .b(net638),
    .c(n3480),
    .o1(u_reg_u_data_in_wr_data[11]));
 b15norp02ar1n48x5 U4712 (.a(n3481),
    .b(n4123),
    .o1(n3497));
 b15nonb02aq1n03x5 U4713 (.a(reg2hw_intr_ctrl_en_rising__q__11_),
    .b(data_in_q[11]),
    .out0(n3488));
 b15aoi012al1n02x5 U4714 (.a(reg2hw_intr_ctrl_en_lvllow__q__11_),
    .b(data_in_q[11]),
    .c(reg2hw_intr_ctrl_en_falling__q__11_),
    .o1(n3486));
 b15nandp3an1n24x5 U4715 (.a(n3484),
    .b(n3483),
    .c(n3482),
    .o1(n3498));
 b15oai022ah1n04x5 U4717 (.a(n3486),
    .b(net380),
    .c(n4077),
    .d(net323),
    .o1(n3487));
 b15oaoi13as1n08x5 U4718 (.a(n3487),
    .b(net380),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__11_),
    .d(n3488),
    .o1(n3726));
 b15aboi22ar1n08x5 U4719 (.a(reg2hw_intr_state__q__11_),
    .b(n3726),
    .c(net67),
    .d(n3497),
    .out0(u_reg_u_intr_state_wr_data[11]));
 b15nand02an1n08x5 U4720 (.a(reg2hw_ctrl_en_input_filter__q__25_),
    .b(net2314),
    .o1(n3489));
 b15oai012as1n24x5 U4721 (.a(n3489),
    .b(reg2hw_ctrl_en_input_filter__q__25_),
    .c(n3490),
    .o1(u_reg_u_data_in_wr_data[25]));
 b15nonb02ar1n04x5 U4722 (.a(net549),
    .b(data_in_q[25]),
    .out0(n3494));
 b15aoi012ah1n02x5 U4723 (.a(net555),
    .b(data_in_q[25]),
    .c(reg2hw_intr_ctrl_en_falling__q__25_),
    .o1(n3492));
 b15oai022ah1n06x5 U4724 (.a(n3492),
    .b(u_reg_u_data_in_wr_data[25]),
    .c(net779),
    .d(net321),
    .o1(n3493));
 b15oaoi13as1n08x5 U4725 (.a(n3493),
    .b(u_reg_u_data_in_wr_data[25]),
    .c(net568),
    .d(n3494),
    .o1(n3727));
 b15aoi022ah1n12x5 U4726 (.a(net822),
    .b(n3497),
    .c(n3727),
    .d(n3947),
    .o1(u_reg_u_intr_state_wr_data[25]));
 b15inv040aq1n05x5 U4727 (.a(gen_filter_9__u_filter_filter_synced),
    .o1(n3496));
 b15nand02an1n12x5 U4728 (.a(net595),
    .b(net2567),
    .o1(n3495));
 b15oai012as1n32x5 U4729 (.a(n3495),
    .b(net595),
    .c(n3496),
    .o1(u_reg_u_data_in_wr_data[9]));
 b15inv000al1n02x5 U4733 (.a(data_in_q[9]),
    .o1(n3499));
 b15aoai13as1n04x5 U4734 (.a(u_reg_u_data_in_wr_data[9]),
    .b(net561),
    .c(reg2hw_intr_ctrl_en_rising__q__9_),
    .d(n3499),
    .o1(n3502));
 b15inv000al1n02x5 U4735 (.a(u_reg_u_data_in_wr_data[9]),
    .o1(n3500));
 b15aoai13ah1n04x5 U4736 (.a(n3500),
    .b(net552),
    .c(net580),
    .d(net2539),
    .o1(n3501));
 b15oai112as1n16x5 U4737 (.a(n3502),
    .b(n3501),
    .c(net322),
    .d(n4075),
    .o1(n3728));
 b15oa0022ah1n02x5 U4738 (.a(n4075),
    .b(net301),
    .c(n3728),
    .d(net2482),
    .o(u_reg_u_intr_state_wr_data[9]));
 b15inv040as1n06x5 U4739 (.a(gen_filter_1__u_filter_filter_synced),
    .o1(n3505));
 b15nand02ah1n12x5 U4740 (.a(net641),
    .b(gen_filter_1__u_filter_stored_value_q),
    .o1(n3504));
 b15oai012aq1n48x5 U4741 (.a(n3504),
    .b(net641),
    .c(n3505),
    .o1(u_reg_u_data_in_wr_data[1]));
 b15inv020an1n03x5 U4742 (.a(data_in_q[1]),
    .o1(n3506));
 b15aoai13as1n06x5 U4743 (.a(u_reg_u_data_in_wr_data[1]),
    .b(net576),
    .c(reg2hw_intr_ctrl_en_rising__q__1_),
    .d(n3506),
    .o1(n3509));
 b15inv040ar1n02x5 U4744 (.a(u_reg_u_data_in_wr_data[1]),
    .o1(n3507));
 b15aoai13ah1n06x5 U4745 (.a(n3507),
    .b(net558),
    .c(net592),
    .d(data_in_q[1]),
    .o1(n3508));
 b15oai112as1n16x5 U4746 (.a(n3509),
    .b(n3508),
    .c(net322),
    .d(net817),
    .o1(n3732));
 b15oa0022ar1n03x5 U4747 (.a(net817),
    .b(net301),
    .c(n3732),
    .d(net2521),
    .o(u_reg_u_intr_state_wr_data[1]));
 b15inv040an1n12x5 U4748 (.a(gen_filter_6__u_filter_filter_synced),
    .o1(n3512));
 b15nandp2al1n12x5 U4749 (.a(net600),
    .b(gen_filter_6__u_filter_stored_value_q),
    .o1(n3511));
 b15oai012aq1n48x5 U4750 (.a(n3511),
    .b(net600),
    .c(n3512),
    .o1(u_reg_u_data_in_wr_data[6]));
 b15inv000as1n02x5 U4751 (.a(data_in_q[6]),
    .o1(n3513));
 b15aoai13an1n06x5 U4752 (.a(u_reg_u_data_in_wr_data[6]),
    .b(net564),
    .c(reg2hw_intr_ctrl_en_rising__q__6_),
    .d(n3513),
    .o1(n3516));
 b15inv000al1n02x5 U4753 (.a(u_reg_u_data_in_wr_data[6]),
    .o1(n3514));
 b15aoai13al1n08x5 U4754 (.a(n3514),
    .b(reg2hw_intr_ctrl_en_lvllow__q__6_),
    .c(reg2hw_intr_ctrl_en_falling__q__6_),
    .d(data_in_q[6]),
    .o1(n3515));
 b15oai112as1n16x5 U4755 (.a(n3516),
    .b(n3515),
    .c(net323),
    .d(n4072),
    .o1(n3712));
 b15oa0022ar1n03x5 U4756 (.a(n4072),
    .b(net301),
    .c(n3712),
    .d(net2466),
    .o(u_reg_u_intr_state_wr_data[6]));
 b15inv000ah1n08x5 U4757 (.a(gen_filter_13__u_filter_filter_synced),
    .o1(n3519));
 b15nand02aq1n16x5 U4758 (.a(reg2hw_ctrl_en_input_filter__q__13_),
    .b(gen_filter_13__u_filter_stored_value_q),
    .o1(n3518));
 b15oai012as1n48x5 U4759 (.a(n3518),
    .b(net635),
    .c(n3519),
    .o1(u_reg_u_data_in_wr_data[13]));
 b15inv000aq1n02x5 U4760 (.a(data_in_q[13]),
    .o1(n3520));
 b15aoai13ah1n04x5 U4761 (.a(u_reg_u_data_in_wr_data[13]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__13_),
    .c(reg2hw_intr_ctrl_en_rising__q__13_),
    .d(n3520),
    .o1(n3523));
 b15inv000al1n02x5 U4762 (.a(u_reg_u_data_in_wr_data[13]),
    .o1(n3521));
 b15aoai13as1n06x5 U4763 (.a(n3521),
    .b(reg2hw_intr_ctrl_en_lvllow__q__13_),
    .c(reg2hw_intr_ctrl_en_falling__q__13_),
    .d(data_in_q[13]),
    .o1(n3522));
 b15oai112as1n16x5 U4764 (.a(n3523),
    .b(n3522),
    .c(net323),
    .d(n3524),
    .o1(n3737));
 b15oa0022ah1n03x5 U4765 (.a(n3524),
    .b(net301),
    .c(n3737),
    .d(reg2hw_intr_state__q__13_),
    .o(u_reg_u_intr_state_wr_data[13]));
 b15inv040ar1n02x5 U4766 (.a(net744),
    .o1(n3526));
 b15nandp2aq1n03x5 U4767 (.a(net611),
    .b(gen_filter_3__u_filter_stored_value_q),
    .o1(n3525));
 b15oai012ar1n08x5 U4768 (.a(n3525),
    .b(net611),
    .c(n3526),
    .o1(u_reg_u_data_in_wr_data[3]));
 b15inv000al1n02x5 U4769 (.a(data_in_q[3]),
    .o1(n3527));
 b15aoai13as1n04x5 U4770 (.a(net379),
    .b(net566),
    .c(net546),
    .d(n3527),
    .o1(n3530));
 b15inv000al1n02x5 U4771 (.a(net379),
    .o1(n3528));
 b15aoai13as1n06x5 U4772 (.a(n3528),
    .b(reg2hw_intr_ctrl_en_lvllow__q__3_),
    .c(reg2hw_intr_ctrl_en_falling__q__3_),
    .d(data_in_q[3]),
    .o1(n3529));
 b15oai112ah1n16x5 U4773 (.a(n3530),
    .b(n3529),
    .c(net323),
    .d(net815),
    .o1(n3721));
 b15oa0022ar1n06x5 U4774 (.a(net816),
    .b(net301),
    .c(n3721),
    .d(net520),
    .o(u_reg_u_intr_state_wr_data[3]));
 b15inv040ah1n06x5 U4775 (.a(net743),
    .o1(n3533));
 b15nandp2al1n12x5 U4776 (.a(net604),
    .b(gen_filter_4__u_filter_stored_value_q),
    .o1(n3532));
 b15oai012aq1n48x5 U4777 (.a(n3532),
    .b(net604),
    .c(n3533),
    .o1(u_reg_u_data_in_wr_data[4]));
 b15inv000al1n02x5 U4778 (.a(data_in_q[4]),
    .o1(n3534));
 b15aoai13an1n06x5 U4779 (.a(u_reg_u_data_in_wr_data[4]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__4_),
    .c(reg2hw_intr_ctrl_en_rising__q__4_),
    .d(n3534),
    .o1(n3537));
 b15inv000al1n02x5 U4780 (.a(u_reg_u_data_in_wr_data[4]),
    .o1(n3535));
 b15aoai13ah1n04x5 U4781 (.a(n3535),
    .b(reg2hw_intr_ctrl_en_lvllow__q__4_),
    .c(reg2hw_intr_ctrl_en_falling__q__4_),
    .d(data_in_q[4]),
    .o1(n3536));
 b15oai112as1n16x5 U4782 (.a(n3537),
    .b(n3536),
    .c(net323),
    .d(net756),
    .o1(n3750));
 b15oa0022an1n02x5 U4783 (.a(net756),
    .b(net300),
    .c(n3750),
    .d(net2563),
    .o(u_reg_u_intr_state_wr_data[4]));
 b15nand02ar1n03x5 U4784 (.a(net631),
    .b(gen_filter_15__u_filter_stored_value_q),
    .o1(n3539));
 b15oai012al1n06x5 U4785 (.a(n3539),
    .b(net631),
    .c(n3540),
    .o1(u_reg_u_data_in_wr_data[15]));
 b15inv000ah1n02x5 U4787 (.a(data_in_q[15]),
    .o1(n3541));
 b15aoai13aq1n06x5 U4788 (.a(net378),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__15_),
    .c(reg2hw_intr_ctrl_en_rising__q__15_),
    .d(n3541),
    .o1(n3544));
 b15inv000al1n02x5 U4789 (.a(net378),
    .o1(n3542));
 b15aoai13as1n06x5 U4790 (.a(n3542),
    .b(reg2hw_intr_ctrl_en_lvllow__q__15_),
    .c(reg2hw_intr_ctrl_en_falling__q__15_),
    .d(data_in_q[15]),
    .o1(n3543));
 b15oai112as1n16x5 U4791 (.a(n3544),
    .b(n3543),
    .c(net323),
    .d(n4080),
    .o1(n3738));
 b15oa0022as1n03x5 U4792 (.a(n4080),
    .b(net301),
    .c(n3738),
    .d(reg2hw_intr_state__q__15_),
    .o(u_reg_u_intr_state_wr_data[15]));
 b15inv040aq1n05x5 U4793 (.a(net742),
    .o1(n3547));
 b15nand02an1n12x5 U4794 (.a(net602),
    .b(net2354),
    .o1(n3546));
 b15oai012as1n32x5 U4795 (.a(n3546),
    .b(net602),
    .c(n3547),
    .o1(u_reg_u_data_in_wr_data[5]));
 b15inv000al1n02x5 U4796 (.a(data_in_q[5]),
    .o1(n3548));
 b15aoai13aq1n04x5 U4797 (.a(u_reg_u_data_in_wr_data[5]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__5_),
    .c(reg2hw_intr_ctrl_en_rising__q__5_),
    .d(n3548),
    .o1(n3551));
 b15inv000al1n02x5 U4798 (.a(u_reg_u_data_in_wr_data[5]),
    .o1(n3549));
 b15aoai13ah1n04x5 U4799 (.a(n3549),
    .b(reg2hw_intr_ctrl_en_lvllow__q__5_),
    .c(reg2hw_intr_ctrl_en_falling__q__5_),
    .d(data_in_q[5]),
    .o1(n3550));
 b15oai112aq1n16x5 U4800 (.a(n3551),
    .b(n3550),
    .c(net323),
    .d(n4071),
    .o1(n3734));
 b15oa0022ar1n04x5 U4801 (.a(n4071),
    .b(net301),
    .c(n3734),
    .d(net2559),
    .o(u_reg_u_intr_state_wr_data[5]));
 b15inv000al1n02x5 U4802 (.a(gen_filter_12__u_filter_filter_synced),
    .o1(n3554));
 b15nand02ah1n03x5 U4803 (.a(reg2hw_ctrl_en_input_filter__q__12_),
    .b(gen_filter_12__u_filter_stored_value_q),
    .o1(n3553));
 b15oai012al1n08x5 U4804 (.a(n3553),
    .b(reg2hw_ctrl_en_input_filter__q__12_),
    .c(n3554),
    .o1(u_reg_u_data_in_wr_data[12]));
 b15inv020aq1n03x5 U4805 (.a(data_in_q[12]),
    .o1(n3555));
 b15aoai13as1n06x5 U4806 (.a(net377),
    .b(net572),
    .c(reg2hw_intr_ctrl_en_rising__q__12_),
    .d(n3555),
    .o1(n3558));
 b15inv040as1n02x5 U4807 (.a(net377),
    .o1(n3556));
 b15aoai13as1n08x5 U4808 (.a(n3556),
    .b(reg2hw_intr_ctrl_en_lvllow__q__12_),
    .c(reg2hw_intr_ctrl_en_falling__q__12_),
    .d(data_in_q[12]),
    .o1(n3557));
 b15oai112as1n16x5 U4809 (.a(n3558),
    .b(n3557),
    .c(net323),
    .d(net811),
    .o1(n3714));
 b15oa0022ah1n03x5 U4810 (.a(net811),
    .b(net301),
    .c(n3714),
    .d(reg2hw_intr_state__q__12_),
    .o(u_reg_u_intr_state_wr_data[12]));
 b15inv000ah1n05x5 U4811 (.a(net740),
    .o1(n3561));
 b15nand02aq1n08x5 U4812 (.a(net597),
    .b(gen_filter_8__u_filter_stored_value_q),
    .o1(n3560));
 b15oai012ar1n32x5 U4813 (.a(n3560),
    .b(net597),
    .c(n3561),
    .o1(u_reg_u_data_in_wr_data[8]));
 b15inv040ah1n03x5 U4814 (.a(data_in_q[8]),
    .o1(n3562));
 b15aoai13ah1n08x5 U4815 (.a(u_reg_u_data_in_wr_data[8]),
    .b(net562),
    .c(reg2hw_intr_ctrl_en_rising__q__8_),
    .d(n3562),
    .o1(n3565));
 b15inv000al1n02x5 U4816 (.a(u_reg_u_data_in_wr_data[8]),
    .o1(n3563));
 b15aoai13as1n08x5 U4817 (.a(n3563),
    .b(net553),
    .c(reg2hw_intr_ctrl_en_falling__q__8_),
    .d(net2560),
    .o1(n3564));
 b15oai112as1n16x5 U4818 (.a(n3565),
    .b(n3564),
    .c(net322),
    .d(n4074),
    .o1(n3722));
 b15oa0022al1n02x5 U4819 (.a(n4074),
    .b(net301),
    .c(n3722),
    .d(reg2hw_intr_state__q__8_),
    .o(u_reg_u_intr_state_wr_data[8]));
 b15inv020as1n06x5 U4820 (.a(net755),
    .o1(n3568));
 b15nandp2ah1n05x5 U4821 (.a(reg2hw_ctrl_en_input_filter__q__0_),
    .b(gen_filter_0__u_filter_stored_value_q),
    .o1(n3567));
 b15oai012as1n24x5 U4822 (.a(n3567),
    .b(reg2hw_ctrl_en_input_filter__q__0_),
    .c(n3568),
    .o1(u_reg_u_data_in_wr_data[0]));
 b15inv000an1n03x5 U4823 (.a(data_in_q[0]),
    .o1(n3569));
 b15aoai13al1n08x5 U4824 (.a(u_reg_u_data_in_wr_data[0]),
    .b(net579),
    .c(reg2hw_intr_ctrl_en_rising__q__0_),
    .d(n3569),
    .o1(n3572));
 b15inv040al1n02x5 U4825 (.a(u_reg_u_data_in_wr_data[0]),
    .o1(n3570));
 b15aoai13ar1n08x5 U4826 (.a(n3570),
    .b(net560),
    .c(net594),
    .d(data_in_q[0]),
    .o1(n3571));
 b15oai112as1n16x5 U4827 (.a(n3572),
    .b(n3571),
    .c(net319),
    .d(net819),
    .o1(n3730));
 b15oa0022an1n02x5 U4828 (.a(net819),
    .b(net301),
    .c(n3730),
    .d(reg2hw_intr_state__q__0_),
    .o(u_reg_u_intr_state_wr_data[0]));
 b15inv040an1n04x5 U4829 (.a(net751),
    .o1(n3575));
 b15nand02ar1n24x5 U4830 (.a(net620),
    .b(gen_filter_23__u_filter_stored_value_q),
    .o1(n3574));
 b15oai012as1n24x5 U4831 (.a(n3574),
    .b(net619),
    .c(n3575),
    .o1(u_reg_u_data_in_wr_data[23]));
 b15inv040ah1n02x5 U4832 (.a(data_in_q[23]),
    .o1(n3576));
 b15aoai13as1n08x5 U4833 (.a(u_reg_u_data_in_wr_data[23]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__23_),
    .c(reg2hw_intr_ctrl_en_rising__q__23_),
    .d(n3576),
    .o1(n3579));
 b15inv000al1n02x5 U4834 (.a(u_reg_u_data_in_wr_data[23]),
    .o1(n3577));
 b15aoai13aq1n08x5 U4835 (.a(n3577),
    .b(reg2hw_intr_ctrl_en_lvllow__q__23_),
    .c(reg2hw_intr_ctrl_en_falling__q__23_),
    .d(data_in_q[23]),
    .o1(n3578));
 b15oai112as1n16x5 U4836 (.a(n3579),
    .b(n3578),
    .c(net320),
    .d(net784),
    .o1(n3736));
 b15oa0022al1n04x5 U4837 (.a(net784),
    .b(net300),
    .c(n3736),
    .d(reg2hw_intr_state__q__23_),
    .o(u_reg_u_intr_state_wr_data[23]));
 b15inv000as1n08x5 U4838 (.a(gen_filter_7__u_filter_filter_synced),
    .o1(n3582));
 b15nand02al1n16x5 U4839 (.a(net598),
    .b(gen_filter_7__u_filter_stored_value_q),
    .o1(n3581));
 b15oai012aq1n48x5 U4840 (.a(n3581),
    .b(net598),
    .c(n3582),
    .o1(u_reg_u_data_in_wr_data[7]));
 b15inv020as1n04x5 U4841 (.a(data_in_q[7]),
    .o1(n3583));
 b15aoai13as1n08x5 U4842 (.a(u_reg_u_data_in_wr_data[7]),
    .b(net563),
    .c(reg2hw_intr_ctrl_en_rising__q__7_),
    .d(n3583),
    .o1(n3586));
 b15inv040ar1n03x5 U4843 (.a(u_reg_u_data_in_wr_data[7]),
    .o1(n3584));
 b15aoai13as1n08x5 U4844 (.a(n3584),
    .b(reg2hw_intr_ctrl_en_lvllow__q__7_),
    .c(reg2hw_intr_ctrl_en_falling__q__7_),
    .d(data_in_q[7]),
    .o1(n3585));
 b15oai112as1n16x5 U4845 (.a(n3586),
    .b(n3585),
    .c(net323),
    .d(net813),
    .o1(n3731));
 b15oa0022an1n02x5 U4846 (.a(n4073),
    .b(net301),
    .c(n3731),
    .d(reg2hw_intr_state__q__7_),
    .o(u_reg_u_intr_state_wr_data[7]));
 b15inv040as1n04x5 U4847 (.a(gen_filter_14__u_filter_filter_synced),
    .o1(n3589));
 b15nand02al1n08x5 U4848 (.a(net632),
    .b(net2414),
    .o1(n3588));
 b15oai012ah1n24x5 U4849 (.a(n3588),
    .b(net632),
    .c(n3589),
    .o1(u_reg_u_data_in_wr_data[14]));
 b15inv020ah1n03x5 U4850 (.a(data_in_q[14]),
    .o1(n3590));
 b15aoai13al1n08x5 U4851 (.a(u_reg_u_data_in_wr_data[14]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__14_),
    .c(reg2hw_intr_ctrl_en_rising__q__14_),
    .d(n3590),
    .o1(n3593));
 b15inv000al1n02x5 U4852 (.a(u_reg_u_data_in_wr_data[14]),
    .o1(n3591));
 b15aoai13as1n06x5 U4853 (.a(n3591),
    .b(reg2hw_intr_ctrl_en_lvllow__q__14_),
    .c(reg2hw_intr_ctrl_en_falling__q__14_),
    .d(data_in_q[14]),
    .o1(n3592));
 b15oai112as1n16x5 U4854 (.a(n3593),
    .b(n3592),
    .c(net323),
    .d(net808),
    .o1(n3743));
 b15oa0022al1n04x5 U4855 (.a(net808),
    .b(net301),
    .c(n3743),
    .d(reg2hw_intr_state__q__14_),
    .o(u_reg_u_intr_state_wr_data[14]));
 b15inv000al1n12x5 U4856 (.a(gen_filter_2__u_filter_filter_synced),
    .o1(n3596));
 b15nand02aq1n16x5 U4857 (.a(reg2hw_ctrl_en_input_filter__q__2_),
    .b(net2465),
    .o1(n3595));
 b15oai012ah1n48x5 U4858 (.a(n3595),
    .b(net613),
    .c(n3596),
    .o1(u_reg_u_data_in_wr_data[2]));
 b15inv040aq1n02x5 U4859 (.a(data_in_q[2]),
    .o1(n3597));
 b15aoai13al1n08x5 U4860 (.a(u_reg_u_data_in_wr_data[2]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__2_),
    .c(net548),
    .d(n3597),
    .o1(n3600));
 b15inv040al1n02x5 U4861 (.a(u_reg_u_data_in_wr_data[2]),
    .o1(n3598));
 b15aoai13aq1n08x5 U4862 (.a(n3598),
    .b(reg2hw_intr_ctrl_en_lvllow__q__2_),
    .c(reg2hw_intr_ctrl_en_falling__q__2_),
    .d(data_in_q[2]),
    .o1(n3599));
 b15oai112as1n16x5 U4863 (.a(n3600),
    .b(n3599),
    .c(net324),
    .d(n4069),
    .o1(n3723));
 b15oa0022ar1n06x5 U4864 (.a(n4069),
    .b(net301),
    .c(n3723),
    .d(net521),
    .o(u_reg_u_intr_state_wr_data[2]));
 b15inv000an1n08x5 U4865 (.a(gen_filter_10__u_filter_filter_synced),
    .o1(n3603));
 b15nand02al1n16x5 U4866 (.a(net640),
    .b(net2568),
    .o1(n3602));
 b15oai012aq1n48x5 U4867 (.a(n3602),
    .b(net640),
    .c(n3603),
    .o1(u_reg_u_data_in_wr_data[10]));
 b15inv000al1n02x5 U4868 (.a(data_in_q[10]),
    .o1(n3604));
 b15aoai13ah1n03x5 U4869 (.a(u_reg_u_data_in_wr_data[10]),
    .b(net574),
    .c(reg2hw_intr_ctrl_en_rising__q__10_),
    .d(n3604),
    .o1(n3607));
 b15inv000al1n02x5 U4870 (.a(u_reg_u_data_in_wr_data[10]),
    .o1(n3605));
 b15aoai13aq1n06x5 U4871 (.a(n3605),
    .b(reg2hw_intr_ctrl_en_lvllow__q__10_),
    .c(reg2hw_intr_ctrl_en_falling__q__10_),
    .d(data_in_q[10]),
    .o1(n3606));
 b15oai112as1n12x5 U4872 (.a(n3607),
    .b(n3606),
    .c(net323),
    .d(n4076),
    .o1(n3739));
 b15oa0022ar1n06x5 U4873 (.a(n4076),
    .b(net301),
    .c(n3739),
    .d(reg2hw_intr_state__q__10_),
    .o(u_reg_u_intr_state_wr_data[10]));
 b15inv020ah1n05x5 U4874 (.a(net747),
    .o1(n3611));
 b15nandp2ah1n05x5 U4875 (.a(net615),
    .b(gen_filter_29__u_filter_stored_value_q),
    .o1(n3610));
 b15oai012as1n24x5 U4876 (.a(n3610),
    .b(net615),
    .c(n3611),
    .o1(u_reg_u_data_in_wr_data[29]));
 b15inv020an1n04x5 U4878 (.a(net2337),
    .o1(n3613));
 b15aoai13al1n08x5 U4879 (.a(u_reg_u_data_in_wr_data[29]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__29_),
    .c(reg2hw_intr_ctrl_en_rising__q__29_),
    .d(n3613),
    .o1(n3616));
 b15inv000al1n02x5 U4880 (.a(u_reg_u_data_in_wr_data[29]),
    .o1(n3614));
 b15aoai13an1n06x5 U4881 (.a(n3614),
    .b(reg2hw_intr_ctrl_en_lvllow__q__29_),
    .c(reg2hw_intr_ctrl_en_falling__q__29_),
    .d(net2337),
    .o1(n3615));
 b15oai112as1n16x5 U4882 (.a(n3616),
    .b(n3615),
    .c(net320),
    .d(net764),
    .o1(n3717));
 b15oa0022as1n02x5 U4883 (.a(net764),
    .b(net300),
    .c(n3717),
    .d(reg2hw_intr_state__q__29_),
    .o(u_reg_u_intr_state_wr_data[29]));
 b15nandp2al1n08x5 U4884 (.a(net624),
    .b(gen_filter_21__u_filter_stored_value_q),
    .o1(n3618));
 b15oai012an1n32x5 U4885 (.a(n3618),
    .b(net624),
    .c(n3619),
    .o1(u_reg_u_data_in_wr_data[21]));
 b15inv040al1n02x5 U4886 (.a(data_in_q[21]),
    .o1(n3620));
 b15aoai13as1n06x5 U4887 (.a(u_reg_u_data_in_wr_data[21]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__21_),
    .c(reg2hw_intr_ctrl_en_rising__q__21_),
    .d(n3620),
    .o1(n3623));
 b15inv040ar1n02x5 U4888 (.a(u_reg_u_data_in_wr_data[21]),
    .o1(n3621));
 b15aoai13al1n08x5 U4889 (.a(n3621),
    .b(reg2hw_intr_ctrl_en_lvllow__q__21_),
    .c(reg2hw_intr_ctrl_en_falling__q__21_),
    .d(data_in_q[21]),
    .o1(n3622));
 b15oai112as1n16x5 U4890 (.a(n3623),
    .b(n3622),
    .c(net320),
    .d(net791),
    .o1(n3720));
 b15oa0022al1n04x5 U4891 (.a(net791),
    .b(net300),
    .c(n3720),
    .d(reg2hw_intr_state__q__21_),
    .o(u_reg_u_intr_state_wr_data[21]));
 b15inv000ah1n04x5 U4892 (.a(gen_filter_26__u_filter_filter_synced),
    .o1(n3626));
 b15nand02al1n08x5 U4893 (.a(reg2hw_ctrl_en_input_filter__q__26_),
    .b(gen_filter_26__u_filter_stored_value_q),
    .o1(n3625));
 b15oai012ar1n24x5 U4894 (.a(n3625),
    .b(reg2hw_ctrl_en_input_filter__q__26_),
    .c(n3626),
    .o1(u_reg_u_data_in_wr_data[26]));
 b15inv000aq1n02x5 U4895 (.a(data_in_q[26]),
    .o1(n3627));
 b15aoai13as1n06x5 U4896 (.a(u_reg_u_data_in_wr_data[26]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__26_),
    .c(reg2hw_intr_ctrl_en_rising__q__26_),
    .d(n3627),
    .o1(n3630));
 b15inv000al1n02x5 U4897 (.a(u_reg_u_data_in_wr_data[26]),
    .o1(n3628));
 b15aoai13as1n06x5 U4898 (.a(n3628),
    .b(reg2hw_intr_ctrl_en_lvllow__q__26_),
    .c(net586),
    .d(data_in_q[26]),
    .o1(n3629));
 b15oai112as1n16x5 U4899 (.a(n3630),
    .b(n3629),
    .c(net320),
    .d(net775),
    .o1(n3740));
 b15oa0022ar1n02x5 U4900 (.a(net776),
    .b(net300),
    .c(n3740),
    .d(reg2hw_intr_state__q__26_),
    .o(u_reg_u_intr_state_wr_data[26]));
 b15inv040as1n04x5 U4901 (.a(gen_filter_24__u_filter_filter_synced),
    .o1(n3633));
 b15nandp2as1n05x5 U4902 (.a(reg2hw_ctrl_en_input_filter__q__24_),
    .b(net2457),
    .o1(n3632));
 b15oai012ar1n32x5 U4903 (.a(n3632),
    .b(reg2hw_ctrl_en_input_filter__q__24_),
    .c(n3633),
    .o1(u_reg_u_data_in_wr_data[24]));
 b15inv000al1n02x5 U4904 (.a(data_in_q[24]),
    .o1(n3634));
 b15aoai13as1n04x5 U4905 (.a(u_reg_u_data_in_wr_data[24]),
    .b(net569),
    .c(reg2hw_intr_ctrl_en_rising__q__24_),
    .d(n3634),
    .o1(n3637));
 b15inv000an1n02x5 U4906 (.a(u_reg_u_data_in_wr_data[24]),
    .o1(n3635));
 b15aoai13aq1n06x5 U4907 (.a(n3635),
    .b(net556),
    .c(reg2hw_intr_ctrl_en_falling__q__24_),
    .d(data_in_q[24]),
    .o1(n3636));
 b15oai112as1n16x5 U4908 (.a(n3637),
    .b(n3636),
    .c(net321),
    .d(net781),
    .o1(n3716));
 b15oa0022an1n04x5 U4909 (.a(net782),
    .b(net300),
    .c(n3716),
    .d(net2557),
    .o(u_reg_u_intr_state_wr_data[24]));
 b15qgbin1an1n05x5 U4910 (.a(gen_filter_19__u_filter_filter_synced),
    .o1(n3640));
 b15nand02as1n06x5 U4911 (.a(net627),
    .b(net2349),
    .o1(n3639));
 b15oai012an1n24x5 U4912 (.a(n3639),
    .b(net627),
    .c(n3640),
    .o1(u_reg_u_data_in_wr_data[19]));
 b15inv040an1n02x5 U4913 (.a(data_in_q[19]),
    .o1(n3641));
 b15aoai13ar1n08x5 U4914 (.a(u_reg_u_data_in_wr_data[19]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__19_),
    .c(reg2hw_intr_ctrl_en_rising__q__19_),
    .d(n3641),
    .o1(n3644));
 b15inv000as1n02x5 U4915 (.a(u_reg_u_data_in_wr_data[19]),
    .o1(n3642));
 b15aoai13as1n06x5 U4916 (.a(n3642),
    .b(reg2hw_intr_ctrl_en_lvllow__q__19_),
    .c(net589),
    .d(data_in_q[19]),
    .o1(n3643));
 b15oai112as1n16x5 U4917 (.a(n3644),
    .b(n3643),
    .c(net321),
    .d(net796),
    .o1(n3741));
 b15oa0022aq1n03x5 U4918 (.a(net797),
    .b(net300),
    .c(n3741),
    .d(reg2hw_intr_state__q__19_),
    .o(u_reg_u_intr_state_wr_data[19]));
 b15inv040as1n04x5 U4919 (.a(gen_filter_30__u_filter_filter_synced),
    .o1(n3647));
 b15nand02an1n12x5 U4920 (.a(net607),
    .b(net2347),
    .o1(n3646));
 b15oai012as1n32x5 U4921 (.a(n3646),
    .b(net607),
    .c(n3647),
    .o1(u_reg_u_data_in_wr_data[30]));
 b15inv020ar1n04x5 U4922 (.a(data_in_q[30]),
    .o1(n3648));
 b15aoai13ar1n08x5 U4923 (.a(u_reg_u_data_in_wr_data[30]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__30_),
    .c(reg2hw_intr_ctrl_en_rising__q__30_),
    .d(n3648),
    .o1(n3651));
 b15inv000al1n02x5 U4924 (.a(u_reg_u_data_in_wr_data[30]),
    .o1(n3649));
 b15aoai13as1n04x5 U4925 (.a(n3649),
    .b(reg2hw_intr_ctrl_en_lvllow__q__30_),
    .c(reg2hw_intr_ctrl_en_falling__q__30_),
    .d(data_in_q[30]),
    .o1(n3650));
 b15oai112as1n16x5 U4926 (.a(n3651),
    .b(n3650),
    .c(net320),
    .d(net762),
    .o1(n3733));
 b15oa0022ar1n06x5 U4927 (.a(net763),
    .b(net300),
    .c(n3733),
    .d(reg2hw_intr_state__q__30_),
    .o(u_reg_u_intr_state_wr_data[30]));
 b15inv020ah1n05x5 U4928 (.a(gen_filter_18__u_filter_filter_synced),
    .o1(n3654));
 b15nandp2ar1n08x5 U4929 (.a(net629),
    .b(gen_filter_18__u_filter_stored_value_q),
    .o1(n3653));
 b15oai012al1n24x5 U4930 (.a(n3653),
    .b(net629),
    .c(n3654),
    .o1(u_reg_u_data_in_wr_data[18]));
 b15inv020an1n03x5 U4931 (.a(data_in_q[18]),
    .o1(n3655));
 b15aoai13ar1n08x5 U4932 (.a(u_reg_u_data_in_wr_data[18]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__18_),
    .c(reg2hw_intr_ctrl_en_rising__q__18_),
    .d(n3655),
    .o1(n3658));
 b15inv000al1n02x5 U4933 (.a(u_reg_u_data_in_wr_data[18]),
    .o1(n3656));
 b15aoai13ar1n08x5 U4934 (.a(n3656),
    .b(reg2hw_intr_ctrl_en_lvllow__q__18_),
    .c(net590),
    .d(data_in_q[18]),
    .o1(n3657));
 b15oai112as1n16x5 U4935 (.a(n3658),
    .b(n3657),
    .c(net321),
    .d(net799),
    .o1(n3713));
 b15oa0022ah1n02x5 U4936 (.a(net800),
    .b(net300),
    .c(n3713),
    .d(reg2hw_intr_state__q__18_),
    .o(u_reg_u_intr_state_wr_data[18]));
 b15inv020an1n04x5 U4937 (.a(net754),
    .o1(n3661));
 b15nand02aq1n04x5 U4938 (.a(net626),
    .b(gen_filter_20__u_filter_stored_value_q),
    .o1(n3660));
 b15oai012al1n06x5 U4939 (.a(n3660),
    .b(net626),
    .c(n3661),
    .o1(u_reg_u_data_in_wr_data[20]));
 b15inv020ah1n03x5 U4940 (.a(data_in_q[20]),
    .o1(n3662));
 b15aoai13as1n08x5 U4941 (.a(net376),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__20_),
    .c(reg2hw_intr_ctrl_en_rising__q__20_),
    .d(n3662),
    .o1(n3665));
 b15inv000al1n02x5 U4942 (.a(net376),
    .o1(n3663));
 b15aoai13al1n08x5 U4943 (.a(n3663),
    .b(reg2hw_intr_ctrl_en_lvllow__q__20_),
    .c(reg2hw_intr_ctrl_en_falling__q__20_),
    .d(data_in_q[20]),
    .o1(n3664));
 b15oai112aq1n16x5 U4944 (.a(n3665),
    .b(n3664),
    .c(net320),
    .d(net793),
    .o1(n3742));
 b15oa0022ah1n03x5 U4945 (.a(net794),
    .b(net300),
    .c(n3742),
    .d(reg2hw_intr_state__q__20_),
    .o(u_reg_u_intr_state_wr_data[20]));
 b15inv000aq1n08x5 U4946 (.a(gen_filter_28__u_filter_filter_synced),
    .o1(n3668));
 b15nand02ah1n12x5 U4947 (.a(net616),
    .b(net2540),
    .o1(n3667));
 b15oai012aq1n48x5 U4948 (.a(n3667),
    .b(net616),
    .c(n3668),
    .o1(u_reg_u_data_in_wr_data[28]));
 b15inv020ah1n03x5 U4949 (.a(data_in_q[28]),
    .o1(n3669));
 b15aoai13al1n08x5 U4950 (.a(u_reg_u_data_in_wr_data[28]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__28_),
    .c(reg2hw_intr_ctrl_en_rising__q__28_),
    .d(n3669),
    .o1(n3672));
 b15inv000al1n02x5 U4951 (.a(u_reg_u_data_in_wr_data[28]),
    .o1(n3670));
 b15aoai13ar1n08x5 U4952 (.a(n3670),
    .b(reg2hw_intr_ctrl_en_lvllow__q__28_),
    .c(reg2hw_intr_ctrl_en_falling__q__28_),
    .d(net2428),
    .o1(n3671));
 b15oai112as1n16x5 U4953 (.a(n3672),
    .b(n3671),
    .c(net320),
    .d(net769),
    .o1(n3729));
 b15oa0022ah1n02x5 U4954 (.a(net769),
    .b(net300),
    .c(net2429),
    .d(reg2hw_intr_state__q__28_),
    .o(u_reg_u_intr_state_wr_data[28]));
 b15inv000as1n03x5 U4955 (.a(gen_filter_27__u_filter_filter_synced),
    .o1(n3675));
 b15nandp2ah1n04x5 U4956 (.a(net618),
    .b(net2256),
    .o1(n3674));
 b15oai012ah1n16x5 U4957 (.a(n3674),
    .b(net618),
    .c(n3675),
    .o1(u_reg_u_data_in_wr_data[27]));
 b15inv000al1n02x5 U4958 (.a(data_in_q[27]),
    .o1(n3676));
 b15aoai13as1n04x5 U4959 (.a(u_reg_u_data_in_wr_data[27]),
    .b(net567),
    .c(reg2hw_intr_ctrl_en_rising__q__27_),
    .d(n3676),
    .o1(n3679));
 b15inv000al1n02x5 U4960 (.a(u_reg_u_data_in_wr_data[27]),
    .o1(n3677));
 b15aoai13as1n04x5 U4961 (.a(n3677),
    .b(reg2hw_intr_ctrl_en_lvllow__q__27_),
    .c(net584),
    .d(net2470),
    .o1(n3678));
 b15oai112as1n16x5 U4962 (.a(n3679),
    .b(n3678),
    .c(net321),
    .d(net772),
    .o1(n3718));
 b15oa0022an1n03x5 U4963 (.a(net773),
    .b(net300),
    .c(n3718),
    .d(reg2hw_intr_state__q__27_),
    .o(u_reg_u_intr_state_wr_data[27]));
 b15inv000an1n05x5 U4964 (.a(gen_filter_16__u_filter_filter_synced),
    .o1(n3682));
 b15nandp2an1n05x5 U4965 (.a(reg2hw_ctrl_en_input_filter__q__16_),
    .b(gen_filter_16__u_filter_stored_value_q),
    .o1(n3681));
 b15oai012an1n24x5 U4966 (.a(n3681),
    .b(reg2hw_ctrl_en_input_filter__q__16_),
    .c(n3682),
    .o1(u_reg_u_data_in_wr_data[16]));
 b15inv000aq1n02x5 U4967 (.a(data_in_q[16]),
    .o1(n3683));
 b15aoai13an1n06x5 U4968 (.a(u_reg_u_data_in_wr_data[16]),
    .b(net571),
    .c(net551),
    .d(n3683),
    .o1(n3686));
 b15inv000al1n02x5 U4969 (.a(u_reg_u_data_in_wr_data[16]),
    .o1(n3684));
 b15aoai13as1n04x5 U4970 (.a(n3684),
    .b(reg2hw_intr_ctrl_en_lvllow__q__16_),
    .c(reg2hw_intr_ctrl_en_falling__q__16_),
    .d(net2505),
    .o1(n3685));
 b15oai112as1n16x5 U4971 (.a(n3686),
    .b(n3685),
    .c(net321),
    .d(net806),
    .o1(n3715));
 b15oa0022ah1n02x5 U4972 (.a(net806),
    .b(net300),
    .c(n3715),
    .d(reg2hw_intr_state__q__16_),
    .o(u_reg_u_intr_state_wr_data[16]));
 b15inv000ar1n12x5 U4973 (.a(net746),
    .o1(n3689));
 b15nandp2ah1n08x5 U4974 (.a(reg2hw_ctrl_en_input_filter__q__31_),
    .b(net2333),
    .o1(n3688));
 b15oai012an1n48x5 U4975 (.a(n3688),
    .b(net606),
    .c(n3689),
    .o1(u_reg_u_data_in_wr_data[31]));
 b15inv020an1n04x5 U4976 (.a(data_in_q[31]),
    .o1(n3690));
 b15aoai13al1n08x5 U4977 (.a(u_reg_u_data_in_wr_data[31]),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__31_),
    .c(reg2hw_intr_ctrl_en_rising__q__31_),
    .d(n3690),
    .o1(n3693));
 b15inv020ah1n03x5 U4978 (.a(u_reg_u_data_in_wr_data[31]),
    .o1(n3691));
 b15aoai13al1n08x5 U4979 (.a(n3691),
    .b(reg2hw_intr_ctrl_en_lvllow__q__31_),
    .c(reg2hw_intr_ctrl_en_falling__q__31_),
    .d(data_in_q[31]),
    .o1(n3692));
 b15oai112as1n16x5 U4980 (.a(n3693),
    .b(n3692),
    .c(net320),
    .d(net759),
    .o1(n3751));
 b15oa0022ar1n06x5 U4981 (.a(net759),
    .b(net300),
    .c(n3751),
    .d(reg2hw_intr_state__q__31_),
    .o(u_reg_u_intr_state_wr_data[31]));
 b15inv000ah1n05x5 U4982 (.a(net753),
    .o1(n3697));
 b15nandp2ar1n03x5 U4983 (.a(net622),
    .b(gen_filter_22__u_filter_stored_value_q),
    .o1(n3696));
 b15oai012ar1n08x5 U4984 (.a(n3696),
    .b(net622),
    .c(n3697),
    .o1(u_reg_u_data_in_wr_data[22]));
 b15inv000ar1n03x5 U4985 (.a(data_in_q[22]),
    .o1(n3698));
 b15aoai13as1n04x5 U4986 (.a(net375),
    .b(reg2hw_intr_ctrl_en_lvlhigh__q__22_),
    .c(reg2hw_intr_ctrl_en_rising__q__22_),
    .d(n3698),
    .o1(n3701));
 b15inv020ar1n04x5 U4987 (.a(net375),
    .o1(n3699));
 b15aoai13ar1n08x5 U4988 (.a(n3699),
    .b(reg2hw_intr_ctrl_en_lvllow__q__22_),
    .c(reg2hw_intr_ctrl_en_falling__q__22_),
    .d(data_in_q[22]),
    .o1(n3700));
 b15oai112as1n16x5 U4989 (.a(n3701),
    .b(n3700),
    .c(net320),
    .d(net787),
    .o1(n3735));
 b15oa0022al1n04x5 U4990 (.a(net787),
    .b(net300),
    .c(n3735),
    .d(net2569),
    .o(u_reg_u_intr_state_wr_data[22]));
 b15inv020as1n05x5 U4991 (.a(gen_filter_17__u_filter_filter_synced),
    .o1(n3704));
 b15nand02ar1n12x5 U4992 (.a(reg2hw_ctrl_en_input_filter__q__17_),
    .b(gen_filter_17__u_filter_stored_value_q),
    .o1(n3703));
 b15oai012ah1n24x5 U4993 (.a(n3703),
    .b(reg2hw_ctrl_en_input_filter__q__17_),
    .c(n3704),
    .o1(u_reg_u_data_in_wr_data[17]));
 b15inv000ar1n04x5 U4994 (.a(data_in_q[17]),
    .o1(n3705));
 b15aoai13ar1n08x5 U4995 (.a(u_reg_u_data_in_wr_data[17]),
    .b(net570),
    .c(net550),
    .d(n3705),
    .o1(n3708));
 b15inv000al1n02x5 U4996 (.a(u_reg_u_data_in_wr_data[17]),
    .o1(n3706));
 b15aoai13as1n04x5 U4997 (.a(n3706),
    .b(reg2hw_intr_ctrl_en_lvllow__q__17_),
    .c(reg2hw_intr_ctrl_en_falling__q__17_),
    .d(net2502),
    .o1(n3707));
 b15oai112as1n16x5 U4998 (.a(n3708),
    .b(n3707),
    .c(net804),
    .d(net322),
    .o1(n3719));
 b15oa0022ah1n02x5 U4999 (.a(net804),
    .b(net300),
    .c(n3719),
    .d(reg2hw_intr_state__q__17_),
    .o(u_reg_u_intr_state_wr_data[17]));
 b15nor004ah1n04x5 U5000 (.a(n3715),
    .b(n3714),
    .c(n3713),
    .d(n3712),
    .o1(n3754));
 b15nor004as1n12x5 U5001 (.a(n3719),
    .b(n3718),
    .c(n3717),
    .d(n3716),
    .o1(n3753));
 b15nor004ar1n08x5 U5002 (.a(n3723),
    .b(n3722),
    .c(n3721),
    .d(n3720),
    .o1(n3725));
 b15nand04ah1n08x5 U5003 (.a(n3727),
    .b(n3726),
    .c(n3725),
    .d(net301),
    .o1(n3749));
 b15nor004aq1n08x5 U5004 (.a(n3731),
    .b(n3730),
    .c(n3729),
    .d(n3728),
    .o1(n3747));
 b15nor004ah1n04x5 U5005 (.a(n3735),
    .b(n3734),
    .c(n3733),
    .d(n3732),
    .o1(n3746));
 b15nor004an1n12x5 U5006 (.a(n3739),
    .b(n3738),
    .c(n3737),
    .d(n3736),
    .o1(n3745));
 b15nor004as1n12x5 U5007 (.a(n3743),
    .b(n3742),
    .c(n3741),
    .d(n3740),
    .o1(n3744));
 b15nand04al1n12x5 U5008 (.a(n3747),
    .b(n3746),
    .c(n3745),
    .d(n3744),
    .o1(n3748));
 b15nor004al1n12x5 U5009 (.a(n3751),
    .b(n3750),
    .c(n3749),
    .d(n3748),
    .o1(n3752));
 b15nand03as1n12x5 U5010 (.a(n3754),
    .b(n3753),
    .c(n3752),
    .o1(u_reg_u_intr_state_n1));
 b15norp03ah1n08x5 U5011 (.a(net2019),
    .b(n3756),
    .c(n3755),
    .o1(u_reg_u_reg_if_rd_req));
 b15aoi022as1n12x5 U5013 (.a(reg2hw_intr_ctrl_en_rising__q__0_),
    .b(net455),
    .c(net594),
    .d(net387),
    .o1(n3764));
 b15aoi022ar1n32x5 U5014 (.a(n3877),
    .b(net148),
    .c(net431),
    .d(net542),
    .o1(n3763));
 b15aoi022an1n08x5 U5016 (.a(reg2hw_ctrl_en_input_filter__q__0_),
    .b(net400),
    .c(net429),
    .d(net2345),
    .o1(n3762));
 b15nor002an1n24x5 U5017 (.a(n3760),
    .b(n3759),
    .o1(n3872));
 b15aoi022ah1n48x5 U5018 (.a(net577),
    .b(net394),
    .c(net173),
    .d(net373),
    .o1(n3761));
 b15nand04as1n16x5 U5019 (.a(n3764),
    .b(n3763),
    .c(n3762),
    .d(n3761),
    .o1(n3767));
 b15aoi022as1n48x5 U5020 (.a(net439),
    .b(net525),
    .c(n3871),
    .d(net141),
    .o1(n3766));
 b15aoi022al1n32x5 U5021 (.a(net559),
    .b(n3289),
    .c(net422),
    .d(net685),
    .o1(n3765));
 b15nona23as1n32x5 U5022 (.a(net362),
    .b(n3767),
    .c(n3766),
    .d(n3765),
    .out0(u_reg_u_reg_if_N14));
 b15aoi022ah1n24x5 U5023 (.a(reg2hw_intr_ctrl_en_rising__q__1_),
    .b(n3292),
    .c(net558),
    .d(net399),
    .o1(n3773));
 b15aoi022an1n16x5 U5024 (.a(net575),
    .b(net394),
    .c(net410),
    .d(net149),
    .o1(n3772));
 b15aoi022ah1n06x5 U5026 (.a(net642),
    .b(net405),
    .c(net592),
    .d(net381),
    .o1(n3771));
 b15aoi022as1n48x5 U5028 (.a(net184),
    .b(net373),
    .c(n3301),
    .d(net539),
    .o1(n3770));
 b15nand04ah1n12x5 U5029 (.a(n3773),
    .b(n3772),
    .c(n3771),
    .d(n3770),
    .o1(n3776));
 b15aoi022as1n48x5 U5030 (.a(net414),
    .b(net731),
    .c(net422),
    .d(net682),
    .o1(n3775));
 b15aoi022ar1n32x5 U5031 (.a(net435),
    .b(net524),
    .c(net429),
    .d(u_reg_data_in_qs[1]),
    .o1(n3774));
 b15nona23as1n32x5 U5032 (.a(net365),
    .b(n3776),
    .c(n3775),
    .d(n3774),
    .out0(u_reg_u_reg_if_N15));
 b15aoi022as1n12x5 U5033 (.a(net554),
    .b(net395),
    .c(net416),
    .d(net163),
    .o1(n3780));
 b15aoi022ar1n02x5 U5034 (.a(net420),
    .b(net680),
    .c(net430),
    .d(net529),
    .o1(n3779));
 b15aoi022ar1n02x5 U5035 (.a(net612),
    .b(net401),
    .c(reg2hw_intr_ctrl_en_falling__q__2_),
    .d(net383),
    .o1(n3778));
 b15aoi022ah1n12x5 U5036 (.a(net411),
    .b(net150),
    .c(net654),
    .d(net371),
    .o1(n3777));
 b15nand04aq1n04x5 U5037 (.a(n3780),
    .b(n3779),
    .c(n3778),
    .d(n3777),
    .o1(n3783));
 b15aoi022ah1n12x5 U5038 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__2_),
    .b(net392),
    .c(net423),
    .d(net2306),
    .o1(n3782));
 b15aoi022an1n12x5 U5039 (.a(net548),
    .b(net453),
    .c(net437),
    .d(net521),
    .o1(n3781));
 b15nona23aq1n12x5 U5040 (.a(net360),
    .b(n3783),
    .c(n3782),
    .d(n3781),
    .out0(u_reg_u_reg_if_N16));
 b15aoi022as1n48x5 U5041 (.a(net609),
    .b(net402),
    .c(net419),
    .d(net183),
    .o1(n3787));
 b15aoi022al1n48x5 U5042 (.a(net547),
    .b(n3292),
    .c(net428),
    .d(u_reg_data_in_qs[3]),
    .o1(n3786));
 b15aoi022ar1n48x5 U5043 (.a(net412),
    .b(net714),
    .c(net432),
    .d(net527),
    .o1(n3785));
 b15aoi022ah1n08x5 U5044 (.a(net437),
    .b(net520),
    .c(net653),
    .d(net371),
    .o1(n3784));
 b15nand04as1n16x5 U5045 (.a(n3787),
    .b(n3786),
    .c(n3785),
    .d(n3784),
    .o1(n3790));
 b15aoi022aq1n32x5 U5046 (.a(reg2hw_intr_ctrl_en_lvllow__q__3_),
    .b(net399),
    .c(reg2hw_intr_ctrl_en_falling__q__3_),
    .d(net383),
    .o1(n3789));
 b15aoi022al1n48x5 U5047 (.a(net565),
    .b(net390),
    .c(net416),
    .d(net166),
    .o1(n3788));
 b15nona23aq1n12x5 U5048 (.a(net361),
    .b(n3790),
    .c(n3789),
    .d(n3788),
    .out0(u_reg_u_reg_if_N17));
 b15aoi022aq1n16x5 U5049 (.a(net417),
    .b(net696),
    .c(net434),
    .d(reg2hw_intr_enable__q__4_),
    .o1(n3794));
 b15aoi022al1n12x5 U5050 (.a(net545),
    .b(net455),
    .c(net428),
    .d(net2315),
    .o1(n3793));
 b15aoi022ah1n24x5 U5051 (.a(reg2hw_intr_ctrl_en_lvllow__q__4_),
    .b(net395),
    .c(reg2hw_intr_ctrl_en_falling__q__4_),
    .d(net383),
    .o1(n3792));
 b15aoi022as1n48x5 U5052 (.a(n3953),
    .b(net518),
    .c(net199),
    .d(net373),
    .o1(n3791));
 b15nand04as1n16x5 U5053 (.a(n3794),
    .b(n3793),
    .c(n3792),
    .d(n3791),
    .o1(n3797));
 b15aoi022ah1n12x5 U5054 (.a(net603),
    .b(net406),
    .c(net420),
    .d(net185),
    .o1(n3796));
 b15aoi022an1n12x5 U5055 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__4_),
    .b(net392),
    .c(net411),
    .d(net153),
    .o1(n3795));
 b15nona23as1n12x5 U5056 (.a(net364),
    .b(n3797),
    .c(n3796),
    .d(n3795),
    .out0(u_reg_u_reg_if_N18));
 b15aoi022an1n12x5 U5057 (.a(reg2hw_intr_ctrl_en_rising__q__5_),
    .b(net453),
    .c(reg2hw_intr_ctrl_en_lvllow__q__5_),
    .d(net395),
    .o1(n3801));
 b15aoi022an1n16x5 U5058 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__5_),
    .b(net392),
    .c(net411),
    .d(net154),
    .o1(n3800));
 b15aoi022an1n48x5 U5059 (.a(net601),
    .b(net405),
    .c(net428),
    .d(u_reg_data_in_qs[5]),
    .o1(n3799));
 b15aoi022aq1n16x5 U5060 (.a(net645),
    .b(net371),
    .c(net420),
    .d(net186),
    .o1(n3798));
 b15nand04as1n16x5 U5061 (.a(n3801),
    .b(n3800),
    .c(n3799),
    .d(n3798),
    .o1(n3804));
 b15aoi022an1n16x5 U5062 (.a(net581),
    .b(net387),
    .c(net430),
    .d(reg2hw_intr_enable__q__5_),
    .o1(n3803));
 b15aoi022as1n48x5 U5063 (.a(n3953),
    .b(net515),
    .c(net414),
    .d(net695),
    .o1(n3802));
 b15nona23ah1n32x5 U5064 (.a(net366),
    .b(n3804),
    .c(n3803),
    .d(n3802),
    .out0(u_reg_u_reg_if_N19));
 b15aoi022aq1n08x5 U5065 (.a(net599),
    .b(net404),
    .c(net428),
    .d(u_reg_data_in_qs[6]),
    .o1(n3808));
 b15aoi022an1n08x5 U5066 (.a(reg2hw_intr_ctrl_en_falling__q__6_),
    .b(net387),
    .c(net417),
    .d(net169),
    .o1(n3807));
 b15aoi022aq1n24x5 U5067 (.a(reg2hw_intr_ctrl_en_rising__q__6_),
    .b(net454),
    .c(reg2hw_intr_ctrl_en_lvllow__q__6_),
    .d(net398),
    .o1(n3806));
 b15aoi022al1n24x5 U5068 (.a(net436),
    .b(net513),
    .c(net201),
    .d(net374),
    .o1(n3805));
 b15nand04as1n12x5 U5069 (.a(n3808),
    .b(n3807),
    .c(n3806),
    .d(n3805),
    .o1(n3811));
 b15aoi022al1n24x5 U5070 (.a(net413),
    .b(net155),
    .c(net434),
    .d(reg2hw_intr_enable__q__6_),
    .o1(n3810));
 b15aoi022al1n16x5 U5071 (.a(net564),
    .b(net391),
    .c(net421),
    .d(net676),
    .o1(n3809));
 b15nona23as1n24x5 U5072 (.a(net365),
    .b(n3811),
    .c(n3810),
    .d(n3809),
    .out0(u_reg_u_reg_if_N20));
 b15aoi022ar1n12x5 U5073 (.a(net421),
    .b(net674),
    .c(net434),
    .d(reg2hw_intr_enable__q__7_),
    .o1(n3815));
 b15aoi022ah1n06x5 U5074 (.a(net544),
    .b(net455),
    .c(net428),
    .d(u_reg_data_in_qs[7]),
    .o1(n3814));
 b15aoi022aq1n08x5 U5075 (.a(reg2hw_ctrl_en_input_filter__q__7_),
    .b(net404),
    .c(net417),
    .d(net170),
    .o1(n3813));
 b15aoi022ar1n32x5 U5076 (.a(net436),
    .b(net512),
    .c(net202),
    .d(net374),
    .o1(n3812));
 b15nand04as1n16x5 U5077 (.a(n3815),
    .b(n3814),
    .c(n3813),
    .d(n3812),
    .o1(n3818));
 b15aoi022ar1n16x5 U5078 (.a(net563),
    .b(net391),
    .c(net413),
    .d(net712),
    .o1(n3817));
 b15aoi022as1n16x5 U5079 (.a(reg2hw_intr_ctrl_en_lvllow__q__7_),
    .b(net398),
    .c(reg2hw_intr_ctrl_en_falling__q__7_),
    .d(net382),
    .o1(n3816));
 b15nona23aq1n24x5 U5080 (.a(net365),
    .b(n3818),
    .c(n3817),
    .d(n3816),
    .out0(u_reg_u_reg_if_N21));
 b15aoi022an1n12x5 U5081 (.a(net417),
    .b(net171),
    .c(net428),
    .d(u_reg_data_in_qs[8]),
    .o1(n3822));
 b15aoi022aq1n32x5 U5082 (.a(net543),
    .b(net455),
    .c(net413),
    .d(net710),
    .o1(n3821));
 b15aoi022as1n08x5 U5083 (.a(net553),
    .b(net399),
    .c(net438),
    .d(reg2hw_intr_state__q__8_),
    .o1(n3820));
 b15aoi022as1n48x5 U5084 (.a(net644),
    .b(net373),
    .c(n3870),
    .d(net671),
    .o1(n3819));
 b15nand04an1n16x5 U5085 (.a(n3822),
    .b(n3821),
    .c(n3820),
    .d(n3819),
    .o1(n3825));
 b15aoi022aq1n12x5 U5086 (.a(net562),
    .b(net389),
    .c(net433),
    .d(reg2hw_intr_enable__q__8_),
    .o1(n3824));
 b15aoi022aq1n12x5 U5087 (.a(net596),
    .b(net404),
    .c(reg2hw_intr_ctrl_en_falling__q__8_),
    .d(net387),
    .o1(n3823));
 b15nona23ar1n32x5 U5088 (.a(net365),
    .b(n3825),
    .c(n3824),
    .d(n3823),
    .out0(u_reg_u_reg_if_N22));
 b15aoi022aq1n12x5 U5089 (.a(net561),
    .b(net393),
    .c(net433),
    .d(reg2hw_intr_enable__q__9_),
    .o1(n3829));
 b15aoi022as1n48x5 U5090 (.a(net414),
    .b(net692),
    .c(net422),
    .d(net667),
    .o1(n3828));
 b15aoi022as1n06x5 U5091 (.a(net580),
    .b(net387),
    .c(net438),
    .d(reg2hw_intr_state__q__9_),
    .o1(n3827));
 b15aoi022as1n32x5 U5092 (.a(net410),
    .b(net708),
    .c(net643),
    .d(n3872),
    .o1(n3826));
 b15nand04al1n04x5 U5093 (.a(n3829),
    .b(n3828),
    .c(n3827),
    .d(n3826),
    .o1(n3832));
 b15aoi022an1n04x5 U5094 (.a(reg2hw_ctrl_en_input_filter__q__9_),
    .b(net405),
    .c(net552),
    .d(net399),
    .o1(n3831));
 b15aoi022an1n12x5 U5095 (.a(reg2hw_intr_ctrl_en_rising__q__9_),
    .b(net455),
    .c(net428),
    .d(u_reg_data_in_qs[9]),
    .o1(n3830));
 b15nona23aq1n08x5 U5096 (.a(net365),
    .b(n3832),
    .c(n3831),
    .d(n3830),
    .out0(u_reg_u_reg_if_N23));
 b15aoi022an1n04x5 U5097 (.a(reg2hw_intr_ctrl_en_lvllow__q__10_),
    .b(net395),
    .c(net425),
    .d(net2203),
    .o1(n3836));
 b15aoi022an1n06x5 U5098 (.a(reg2hw_intr_ctrl_en_rising__q__10_),
    .b(net454),
    .c(net437),
    .d(reg2hw_intr_state__q__10_),
    .o1(n3835));
 b15aoi022ah1n32x5 U5099 (.a(net573),
    .b(net388),
    .c(net419),
    .d(net666),
    .o1(n3834));
 b15aoi022ar1n48x5 U5100 (.a(net415),
    .b(net729),
    .c(net690),
    .d(net372),
    .o1(n3833));
 b15nand04ah1n08x5 U5101 (.a(net2204),
    .b(n3835),
    .c(n3834),
    .d(n3833),
    .o1(n3839));
 b15aoi022aq1n48x5 U5102 (.a(net591),
    .b(net382),
    .c(net412),
    .d(net159),
    .o1(n3838));
 b15aoi022al1n48x5 U5103 (.a(net639),
    .b(net404),
    .c(net433),
    .d(net538),
    .o1(n3837));
 b15nona23ah1n32x5 U5104 (.a(net364),
    .b(n3839),
    .c(n3838),
    .d(n3837),
    .out0(u_reg_u_reg_if_N24));
 b15aoi022as1n48x5 U5105 (.a(net435),
    .b(net522),
    .c(net419),
    .d(net663),
    .o1(n3843));
 b15aoi022aq1n12x5 U5106 (.a(reg2hw_intr_ctrl_en_falling__q__11_),
    .b(net382),
    .c(net415),
    .d(net143),
    .o1(n3842));
 b15aoi022an1n12x5 U5107 (.a(net638),
    .b(net404),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__11_),
    .d(net391),
    .o1(n3841));
 b15aoi022al1n16x5 U5108 (.a(net412),
    .b(net160),
    .c(net175),
    .d(net372),
    .o1(n3840));
 b15nand04as1n16x5 U5109 (.a(n3843),
    .b(n3842),
    .c(n3841),
    .d(n3840),
    .o1(n3847));
 b15aoi022an1n12x5 U5110 (.a(reg2hw_intr_ctrl_en_lvllow__q__11_),
    .b(net395),
    .c(net424),
    .d(u_reg_data_in_qs[11]),
    .o1(n3846));
 b15aoi022ah1n24x5 U5111 (.a(reg2hw_intr_ctrl_en_rising__q__11_),
    .b(net453),
    .c(net430),
    .d(net537),
    .o1(n3845));
 b15nona23ah1n24x5 U5112 (.a(net363),
    .b(n3847),
    .c(n3846),
    .d(net2340),
    .out0(u_reg_u_reg_if_N25));
 b15aoi022ah1n12x5 U5113 (.a(net430),
    .b(reg2hw_intr_enable__q__12_),
    .c(net425),
    .d(u_reg_data_in_qs[12]),
    .o1(n3852));
 b15aoi022as1n24x5 U5114 (.a(reg2hw_intr_ctrl_en_lvllow__q__12_),
    .b(net398),
    .c(net412),
    .d(net703),
    .o1(n3851));
 b15aoi022ah1n08x5 U5115 (.a(reg2hw_intr_ctrl_en_falling__q__12_),
    .b(net382),
    .c(net415),
    .d(net144),
    .o1(n3850));
 b15aoi022as1n12x5 U5116 (.a(reg2hw_intr_ctrl_en_rising__q__12_),
    .b(net454),
    .c(net689),
    .d(net372),
    .o1(n3849));
 b15nand04as1n16x5 U5117 (.a(n3852),
    .b(n3851),
    .c(n3850),
    .d(n3849),
    .o1(n3855));
 b15aoi022as1n16x5 U5118 (.a(net572),
    .b(net393),
    .c(net437),
    .d(reg2hw_intr_state__q__12_),
    .o1(n3854));
 b15aoi022ar1n48x5 U5119 (.a(net636),
    .b(net403),
    .c(net419),
    .d(net193),
    .o1(n3853));
 b15nona23an1n32x5 U5120 (.a(net360),
    .b(n3855),
    .c(n3854),
    .d(n3853),
    .out0(u_reg_u_reg_if_N26));
 b15aoi022ar1n16x5 U5121 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__13_),
    .b(net389),
    .c(net433),
    .d(reg2hw_intr_enable__q__13_),
    .o1(n3859));
 b15aoi022ar1n24x5 U5122 (.a(reg2hw_intr_ctrl_en_rising__q__13_),
    .b(net454),
    .c(reg2hw_intr_ctrl_en_falling__q__13_),
    .d(net382),
    .o1(n3858));
 b15aoi022ar1n24x5 U5123 (.a(net557),
    .b(net398),
    .c(net413),
    .d(net701),
    .o1(n3857));
 b15aoi022as1n08x5 U5124 (.a(net438),
    .b(reg2hw_intr_state__q__13_),
    .c(net177),
    .d(net372),
    .o1(n3856));
 b15nand04as1n16x5 U5125 (.a(n3859),
    .b(n3858),
    .c(n3857),
    .d(n3856),
    .o1(n3862));
 b15aoi022aq1n48x5 U5126 (.a(net634),
    .b(net404),
    .c(net415),
    .d(net728),
    .o1(n3861));
 b15aoi022an1n32x5 U5127 (.a(net420),
    .b(net194),
    .c(net429),
    .d(net738),
    .o1(n3860));
 b15nona23as1n32x5 U5128 (.a(net364),
    .b(n3862),
    .c(n3861),
    .d(n3860),
    .out0(u_reg_u_reg_if_N27));
 b15aoi022as1n16x5 U5129 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__14_),
    .b(net393),
    .c(net415),
    .d(net726),
    .o1(n3866));
 b15aoi022as1n32x5 U5130 (.a(net420),
    .b(net196),
    .c(net426),
    .d(net739),
    .o1(n3865));
 b15aoi022as1n08x5 U5131 (.a(reg2hw_intr_ctrl_en_rising__q__14_),
    .b(net453),
    .c(reg2hw_intr_ctrl_en_lvllow__q__14_),
    .d(net395),
    .o1(n3864));
 b15aoi022ah1n04x5 U5132 (.a(net437),
    .b(reg2hw_intr_state__q__14_),
    .c(net688),
    .d(net371),
    .o1(n3863));
 b15nand04as1n06x5 U5133 (.a(n3866),
    .b(n3865),
    .c(n3864),
    .d(n3863),
    .o1(n3869));
 b15aoi022aq1n32x5 U5134 (.a(reg2hw_intr_ctrl_en_falling__q__14_),
    .b(net382),
    .c(net412),
    .d(net164),
    .o1(n3868));
 b15aoi022ar1n24x5 U5135 (.a(net633),
    .b(net405),
    .c(net432),
    .d(net536),
    .o1(n3867));
 b15nona23aq1n32x5 U5136 (.a(net364),
    .b(n3869),
    .c(n3868),
    .d(n3867),
    .out0(u_reg_u_reg_if_N28));
 b15aoi022an1n24x5 U5137 (.a(net438),
    .b(reg2hw_intr_state__q__15_),
    .c(net421),
    .d(net649),
    .o1(n3876));
 b15aoi022ar1n32x5 U5138 (.a(reg2hw_intr_ctrl_en_lvllow__q__15_),
    .b(net398),
    .c(net415),
    .d(net724),
    .o1(n3875));
 b15aoi022ah1n08x5 U5139 (.a(net630),
    .b(net406),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__15_),
    .d(net393),
    .o1(n3874));
 b15aoi022ar1n16x5 U5140 (.a(net687),
    .b(net371),
    .c(net430),
    .d(reg2hw_intr_enable__q__15_),
    .o1(n3873));
 b15nand04ah1n08x5 U5141 (.a(n3876),
    .b(n3875),
    .c(n3874),
    .d(n3873),
    .o1(n3880));
 b15aoi022ah1n12x5 U5142 (.a(reg2hw_intr_ctrl_en_rising__q__15_),
    .b(net453),
    .c(reg2hw_intr_ctrl_en_falling__q__15_),
    .d(net382),
    .o1(n3879));
 b15aoi022ar1n24x5 U5143 (.a(net411),
    .b(net165),
    .c(net425),
    .d(u_reg_data_in_qs[15]),
    .o1(n3878));
 b15nona23as1n32x5 U5144 (.a(net363),
    .b(n3880),
    .c(n3879),
    .d(n3878),
    .out0(u_reg_u_reg_if_N29));
 b15aoi022ar1n12x5 U5145 (.a(reg2hw_ctrl_en_input_filter__q__16_),
    .b(net400),
    .c(net571),
    .d(net394),
    .o1(n3887));
 b15aoi022ah1n16x5 U5146 (.a(net440),
    .b(net685),
    .c(net427),
    .d(net2240),
    .o1(n3886));
 b15aoi022al1n12x5 U5147 (.a(reg2hw_intr_ctrl_en_lvllow__q__16_),
    .b(net396),
    .c(net431),
    .d(reg2hw_intr_enable__q__16_),
    .o1(n3885));
 b15aoi022as1n12x5 U5148 (.a(reg2hw_intr_ctrl_en_falling__q__16_),
    .b(net384),
    .c(net723),
    .d(n3982),
    .o1(n3881));
 b15oai012ah1n04x5 U5149 (.a(n3881),
    .b(n4123),
    .c(n3882),
    .o1(n3883));
 b15aoi112ah1n06x5 U5150 (.a(net362),
    .b(n3883),
    .c(net551),
    .d(net449),
    .o1(n3884));
 b15nand04as1n16x5 U5151 (.a(n3887),
    .b(net2241),
    .c(n3885),
    .d(n3884),
    .o1(u_reg_u_reg_if_N30));
 b15aoi022ar1n12x5 U5152 (.a(net570),
    .b(net394),
    .c(net427),
    .d(net2279),
    .o1(n3895));
 b15aoi022ah1n06x5 U5153 (.a(reg2hw_ctrl_en_input_filter__q__17_),
    .b(net400),
    .c(net550),
    .d(net449),
    .o1(n3894));
 b15aoi022as1n06x5 U5154 (.a(reg2hw_intr_ctrl_en_falling__q__17_),
    .b(net384),
    .c(net431),
    .d(reg2hw_intr_enable__q__17_),
    .o1(n3893));
 b15aoi022al1n48x5 U5155 (.a(net721),
    .b(n3982),
    .c(net440),
    .d(net683),
    .o1(n3889));
 b15oai012an1n04x5 U5156 (.a(n3889),
    .b(n4123),
    .c(n3890),
    .o1(n3891));
 b15aoi112an1n06x5 U5157 (.a(net359),
    .b(n3891),
    .c(reg2hw_intr_ctrl_en_lvllow__q__17_),
    .d(net396),
    .o1(n3892));
 b15nand04as1n16x5 U5158 (.a(net2280),
    .b(n3894),
    .c(n3893),
    .d(n3892),
    .o1(u_reg_u_reg_if_N31));
 b15aoi022al1n08x5 U5159 (.a(net590),
    .b(net386),
    .c(net430),
    .d(net535),
    .o1(n3902));
 b15aoi022al1n12x5 U5160 (.a(reg2hw_intr_ctrl_en_lvllow__q__18_),
    .b(net395),
    .c(net441),
    .d(net681),
    .o1(n3901));
 b15aoi022aq1n08x5 U5161 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__18_),
    .b(net388),
    .c(net717),
    .d(net446),
    .o1(n3900));
 b15aoi022ar1n02x5 U5162 (.a(reg2hw_intr_ctrl_en_rising__q__18_),
    .b(net451),
    .c(net426),
    .d(net2236),
    .o1(n3896));
 b15oai012ah1n03x5 U5163 (.a(net2237),
    .b(n4123),
    .c(n3897),
    .o1(n3898));
 b15aoi112an1n06x5 U5164 (.a(net361),
    .b(n3898),
    .c(net629),
    .d(net402),
    .o1(n3899));
 b15nand04ah1n12x5 U5165 (.a(n3902),
    .b(n3901),
    .c(n3900),
    .d(net2238),
    .o1(u_reg_u_reg_if_N32));
 b15aoi022aq1n08x5 U5166 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__20_),
    .b(net390),
    .c(net153),
    .d(net446),
    .o1(n3909));
 b15aoi022ah1n16x5 U5167 (.a(reg2hw_intr_ctrl_en_rising__q__20_),
    .b(net453),
    .c(net442),
    .d(net185),
    .o1(n3908));
 b15aoi022as1n16x5 U5168 (.a(net2518),
    .b(net395),
    .c(reg2hw_intr_ctrl_en_falling__q__20_),
    .d(net383),
    .o1(n3907));
 b15aoi022aq1n04x5 U5169 (.a(net430),
    .b(net534),
    .c(net424),
    .d(u_reg_data_in_qs[20]),
    .o1(n3903));
 b15oai012ar1n12x5 U5170 (.a(n3903),
    .b(n4123),
    .c(n3904),
    .o1(n3905));
 b15aoi112aq1n06x5 U5171 (.a(net360),
    .b(n3905),
    .c(net625),
    .d(net401),
    .o1(n3906));
 b15nand04aq1n16x5 U5172 (.a(n3909),
    .b(n3908),
    .c(n3907),
    .d(n3906),
    .o1(u_reg_u_reg_if_N34));
 b15aoi022ah1n12x5 U5173 (.a(net2321),
    .b(net450),
    .c(reg2hw_intr_ctrl_en_falling__q__21_),
    .d(net383),
    .o1(n3918));
 b15aoi022an1n16x5 U5174 (.a(net442),
    .b(net186),
    .c(net424),
    .d(u_reg_data_in_qs[21]),
    .o1(n3917));
 b15aoi022as1n12x5 U5175 (.a(net154),
    .b(net446),
    .c(net432),
    .d(net533),
    .o1(n3916));
 b15aoi022as1n04x5 U5176 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__21_),
    .b(net390),
    .c(reg2hw_intr_ctrl_en_lvllow__q__21_),
    .d(net395),
    .o1(n3911));
 b15oai012an1n06x5 U5177 (.a(n3911),
    .b(n4123),
    .c(n3912),
    .o1(n3913));
 b15aoi112aq1n08x5 U5178 (.a(net360),
    .b(n3913),
    .c(net623),
    .d(net401),
    .o1(n3915));
 b15nand04as1n16x5 U5179 (.a(n3918),
    .b(n3917),
    .c(n3916),
    .d(n3915),
    .o1(u_reg_u_reg_if_N35));
 b15aoi022an1n12x5 U5180 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__22_),
    .b(net390),
    .c(reg2hw_intr_ctrl_en_falling__q__22_),
    .d(net383),
    .o1(n3927));
 b15aoi022ah1n06x5 U5181 (.a(reg2hw_intr_ctrl_en_lvllow__q__22_),
    .b(net395),
    .c(net430),
    .d(net532),
    .o1(n3926));
 b15aoi022as1n08x5 U5182 (.a(net621),
    .b(net401),
    .c(net424),
    .d(u_reg_data_in_qs[22]),
    .o1(n3925));
 b15aoi022al1n48x5 U5184 (.a(net713),
    .b(net448),
    .c(net443),
    .d(net677),
    .o1(n3920));
 b15oai012as1n03x5 U5185 (.a(net370),
    .b(n4123),
    .c(n3921),
    .o1(n3922));
 b15aoi112as1n06x5 U5186 (.a(net360),
    .b(n3922),
    .c(net2287),
    .d(net450),
    .o1(n3924));
 b15nand04as1n16x5 U5187 (.a(n3927),
    .b(n3926),
    .c(n3925),
    .d(net2288),
    .o1(u_reg_u_reg_if_N36));
 b15aoi022as1n06x5 U5188 (.a(net619),
    .b(net401),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__23_),
    .d(net390),
    .o1(n3938));
 b15aoi022ar1n12x5 U5189 (.a(reg2hw_intr_ctrl_en_lvllow__q__23_),
    .b(net395),
    .c(net430),
    .d(reg2hw_intr_enable__q__23_),
    .o1(n3937));
 b15aoi022as1n08x5 U5190 (.a(reg2hw_intr_ctrl_en_rising__q__23_),
    .b(net450),
    .c(net423),
    .d(net2282),
    .o1(n3936));
 b15aoi022as1n48x5 U5192 (.a(net711),
    .b(net448),
    .c(net443),
    .d(net672),
    .o1(n3931));
 b15oai012al1n08x5 U5193 (.a(n3931),
    .b(n4123),
    .c(n3932),
    .o1(n3933));
 b15aoi112aq1n06x5 U5194 (.a(net360),
    .b(n3933),
    .c(reg2hw_intr_ctrl_en_falling__q__23_),
    .d(net383),
    .o1(n3935));
 b15nand04as1n16x5 U5195 (.a(n3938),
    .b(n3937),
    .c(net2283),
    .d(n3935),
    .o1(u_reg_u_reg_if_N37));
 b15aoi022ar1n12x5 U5196 (.a(net569),
    .b(net394),
    .c(net556),
    .d(net396),
    .o1(n3945));
 b15aoi022aq1n08x5 U5197 (.a(n3981),
    .b(net189),
    .c(net434),
    .d(reg2hw_intr_enable__q__24_),
    .o1(n3944));
 b15aoi022as1n08x5 U5198 (.a(reg2hw_ctrl_en_input_filter__q__24_),
    .b(net405),
    .c(reg2hw_intr_ctrl_en_rising__q__24_),
    .d(net449),
    .o1(n3943));
 b15aoi022an1n02x5 U5199 (.a(net157),
    .b(n3982),
    .c(net429),
    .d(net2402),
    .o1(n3939));
 b15oai012aq1n06x5 U5200 (.a(n3939),
    .b(n4123),
    .c(n3940),
    .o1(n3941));
 b15aoi112an1n06x5 U5201 (.a(net365),
    .b(n3941),
    .c(reg2hw_intr_ctrl_en_falling__q__24_),
    .d(n3295),
    .o1(n3942));
 b15nand04as1n16x5 U5202 (.a(n3945),
    .b(n3944),
    .c(n3943),
    .d(n3942),
    .o1(u_reg_u_reg_if_N38));
 b15aoi022an1n08x5 U5203 (.a(reg2hw_ctrl_en_input_filter__q__25_),
    .b(net403),
    .c(net427),
    .d(net2188),
    .o1(n3952));
 b15aoi022al1n24x5 U5204 (.a(net568),
    .b(net394),
    .c(net549),
    .d(net449),
    .o1(n3951));
 b15aoi022ah1n48x5 U5205 (.a(net587),
    .b(net385),
    .c(net706),
    .d(net445),
    .o1(n3950));
 b15aoi022as1n16x5 U5206 (.a(net440),
    .b(net190),
    .c(net431),
    .d(net530),
    .o1(n3946));
 b15oai012aq1n12x5 U5207 (.a(n3946),
    .b(n4123),
    .c(n3947),
    .o1(n3948));
 b15aoi112ah1n06x5 U5208 (.a(net359),
    .b(n3948),
    .c(net555),
    .d(net396),
    .o1(n3949));
 b15nand04as1n16x5 U5209 (.a(net2189),
    .b(n3951),
    .c(n3950),
    .d(n3949),
    .o1(u_reg_u_reg_if_N39));
 b15aoi022aq1n12x5 U5210 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__26_),
    .b(net388),
    .c(net435),
    .d(reg2hw_intr_state__q__26_),
    .o1(n3961));
 b15aoi022an1n08x5 U5211 (.a(reg2hw_ctrl_en_input_filter__q__26_),
    .b(net402),
    .c(net430),
    .d(reg2hw_intr_enable__q__26_),
    .o1(n3960));
 b15aoi022as1n08x5 U5212 (.a(reg2hw_intr_ctrl_en_lvllow__q__26_),
    .b(net397),
    .c(net427),
    .d(net2211),
    .o1(n3959));
 b15aoi022aq1n12x5 U5213 (.a(net585),
    .b(net382),
    .c(net159),
    .d(net447),
    .o1(n3954));
 b15aob012ar1n12x5 U5214 (.a(net368),
    .b(net444),
    .c(net665),
    .out0(n3955));
 b15aoi112ah1n08x5 U5215 (.a(net360),
    .b(n3955),
    .c(reg2hw_intr_ctrl_en_rising__q__26_),
    .d(net451),
    .o1(n3958));
 b15nand04as1n16x5 U5216 (.a(n3961),
    .b(n3960),
    .c(net2212),
    .d(n3958),
    .o1(u_reg_u_reg_if_N40));
 b15aoi022al1n24x5 U5217 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__28_),
    .b(net388),
    .c(reg2hw_intr_ctrl_en_lvllow__q__28_),
    .d(net395),
    .o1(n3973));
 b15aoi022al1n16x5 U5218 (.a(reg2hw_intr_ctrl_en_rising__q__28_),
    .b(net450),
    .c(net441),
    .d(net659),
    .o1(n3972));
 b15aoi022aq1n12x5 U5219 (.a(net430),
    .b(reg2hw_intr_enable__q__28_),
    .c(net426),
    .d(net2244),
    .o1(n3971));
 b15aoi022an1n16x5 U5221 (.a(net582),
    .b(net386),
    .c(net702),
    .d(net446),
    .o1(n3966));
 b15oai012an1n24x5 U5222 (.a(n3966),
    .b(n4123),
    .c(n3967),
    .o1(n3968));
 b15aoi112aq1n08x5 U5223 (.a(net361),
    .b(n3968),
    .c(net617),
    .d(net402),
    .o1(n3970));
 b15nand04as1n16x5 U5224 (.a(n3973),
    .b(n3972),
    .c(net2245),
    .d(n3970),
    .o1(u_reg_u_reg_if_N42));
 b15aoi022aq1n08x5 U5225 (.a(reg2hw_intr_ctrl_en_lvllow__q__29_),
    .b(net395),
    .c(reg2hw_intr_ctrl_en_falling__q__29_),
    .d(net386),
    .o1(n3992));
 b15aoi022aq1n08x5 U5226 (.a(reg2hw_intr_ctrl_en_rising__q__29_),
    .b(net450),
    .c(net423),
    .d(net2159),
    .o1(n3991));
 b15aoi022al1n12x5 U5227 (.a(net614),
    .b(net401),
    .c(net430),
    .d(reg2hw_intr_enable__q__29_),
    .o1(n3990));
 b15aoi022ah1n06x5 U5229 (.a(net701),
    .b(net447),
    .c(net443),
    .d(net656),
    .o1(n3983));
 b15oai012aq1n08x5 U5230 (.a(net369),
    .b(n4123),
    .c(n3984),
    .o1(n3986));
 b15aoi112ar1n08x5 U5231 (.a(net360),
    .b(n3986),
    .c(reg2hw_intr_ctrl_en_lvlhigh__q__29_),
    .d(net388),
    .o1(n3989));
 b15nand04as1n16x5 U5232 (.a(n3992),
    .b(net2160),
    .c(n3990),
    .d(n3989),
    .o1(u_reg_u_reg_if_N43));
 b15nano23ah1n16x5 U5234 (.a(gen_filter_4__u_filter_diff_ctr_d[1]),
    .b(gen_filter_4__u_filter_diff_ctr_d[0]),
    .c(n3994),
    .d(n3993),
    .out0(eq_x_161_n25));
 b15nano23al1n05x5 U5235 (.a(gen_filter_25__u_filter_diff_ctr_q[3]),
    .b(gen_filter_25__u_filter_diff_ctr_d[0]),
    .c(n3996),
    .d(n3995),
    .out0(eq_x_56_n25));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_0__cio_gpio_en_q_reg_1_ (.rb(net862),
    .clk(clknet_1_1__leaf_net2050),
    .d1(N114),
    .d2(N115),
    .o1(net141),
    .o2(net152),
    .si1(net871),
    .si2(net872),
    .ssb(net1610));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_10__cio_gpio_en_q_reg_11_ (.rb(net846),
    .clk(clknet_1_0__leaf_net2050),
    .d1(N124),
    .d2(N125),
    .o1(net142),
    .o2(net143),
    .si1(net873),
    .si2(net874),
    .ssb(net1611));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_12__cio_gpio_en_q_reg_13_ (.rb(net846),
    .clk(clknet_1_0__leaf_net2050),
    .d1(N126),
    .d2(N127),
    .o1(net144),
    .o2(net145),
    .si1(net875),
    .si2(net876),
    .ssb(net1612));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_14__cio_gpio_en_q_reg_15_ (.rb(net860),
    .clk(clknet_1_1__leaf_net2050),
    .d1(N128),
    .d2(N129),
    .o1(net146),
    .o2(net147),
    .si1(net877),
    .si2(net878),
    .ssb(net1613));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_16__cio_gpio_en_q_reg_17_ (.rb(net859),
    .clk(clknet_1_1__leaf_net2045),
    .d1(N131),
    .d2(N132),
    .o1(net148),
    .o2(net149),
    .si1(net879),
    .si2(net880),
    .ssb(net1614));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_18__cio_gpio_en_q_reg_19_ (.rb(net840),
    .clk(clknet_1_0__leaf_net2045),
    .d1(N133),
    .d2(N134),
    .o1(net150),
    .o2(net151),
    .si1(net881),
    .si2(net882),
    .ssb(net1615));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_20__cio_gpio_en_q_reg_21_ (.rb(net840),
    .clk(clknet_1_0__leaf_net2045),
    .d1(N135),
    .d2(N136),
    .o1(net153),
    .o2(net154),
    .si1(net883),
    .si2(net884),
    .ssb(net1616));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_22__cio_gpio_en_q_reg_23_ (.rb(net860),
    .clk(clknet_1_1__leaf_net2045),
    .d1(N137),
    .d2(N138),
    .o1(net155),
    .o2(net156),
    .si1(net885),
    .si2(net886),
    .ssb(net1617));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_24__cio_gpio_en_q_reg_25_ (.rb(net859),
    .clk(clknet_1_1__leaf_net2045),
    .d1(N139),
    .d2(N140),
    .o1(net157),
    .o2(net158),
    .si1(net887),
    .si2(net888),
    .ssb(net1618));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_26__cio_gpio_en_q_reg_27_ (.rb(net846),
    .clk(clknet_1_1__leaf_net2045),
    .d1(N141),
    .d2(N142),
    .o1(net159),
    .o2(net160),
    .si1(net889),
    .si2(net890),
    .ssb(net1619));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_28__cio_gpio_en_q_reg_29_ (.rb(net841),
    .clk(clknet_1_0__leaf_net2045),
    .d1(N143),
    .d2(N144),
    .o1(net161),
    .o2(net162),
    .si1(net891),
    .si2(net892),
    .ssb(net1620));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_2__cio_gpio_en_q_reg_3_ (.rb(net840),
    .clk(clknet_1_0__leaf_net2050),
    .d1(N116),
    .d2(N117),
    .o1(net163),
    .o2(net166),
    .si1(net893),
    .si2(net894),
    .ssb(net1621));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_30__cio_gpio_en_q_reg_31_ (.rb(net841),
    .clk(clknet_1_0__leaf_net2045),
    .d1(N145),
    .d2(N146),
    .o1(net164),
    .o2(net165),
    .si1(net895),
    .si2(net896),
    .ssb(net1622));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_4__cio_gpio_en_q_reg_5_ (.rb(net862),
    .clk(clknet_1_1__leaf_net2050),
    .d1(N118),
    .d2(N119),
    .o1(net167),
    .o2(net168),
    .si1(net897),
    .si2(net898),
    .ssb(net1623));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_6__cio_gpio_en_q_reg_7_ (.rb(net846),
    .clk(clknet_1_0__leaf_net2050),
    .d1(N120),
    .d2(N121),
    .o1(net169),
    .o2(net170),
    .si1(net899),
    .si2(net900),
    .ssb(net1624));
 b15fqy203ar1n02x5 cio_gpio_en_q_reg_8__cio_gpio_en_q_reg_9_ (.rb(net860),
    .clk(clknet_1_1__leaf_net2050),
    .d1(N122),
    .d2(N123),
    .o1(net171),
    .o2(net172),
    .si1(net901),
    .si2(net902),
    .ssb(net1625));
 b15fqy203ar1n02x5 cio_gpio_q_reg_0__cio_gpio_q_reg_1_ (.rb(net856),
    .clk(clknet_1_1__leaf_net2040),
    .d1(N39),
    .d2(N40),
    .o1(net173),
    .o2(net184),
    .si1(net903),
    .si2(net904),
    .ssb(net1626));
 b15fqy203ar1n02x5 cio_gpio_q_reg_10__cio_gpio_q_reg_11_ (.rb(net846),
    .clk(clknet_1_0__leaf_net2040),
    .d1(N49),
    .d2(N50),
    .o1(net174),
    .o2(net175),
    .si1(net905),
    .si2(net906),
    .ssb(net1627));
 b15fqy203ar1n02x5 cio_gpio_q_reg_12__cio_gpio_q_reg_13_ (.rb(net846),
    .clk(clknet_1_0__leaf_net2040),
    .d1(N51),
    .d2(N52),
    .o1(net176),
    .o2(net177),
    .si1(net907),
    .si2(net908),
    .ssb(net1628));
 b15fqy203ar1n02x5 cio_gpio_q_reg_14__cio_gpio_q_reg_15_ (.rb(net844),
    .clk(clknet_1_0__leaf_net2040),
    .d1(N53),
    .d2(N54),
    .o1(net178),
    .o2(net179),
    .si1(net909),
    .si2(net910),
    .ssb(net1629));
 b15fqy203ar1n02x5 cio_gpio_q_reg_16__cio_gpio_q_reg_17_ (.rb(net856),
    .clk(clknet_1_1__leaf_net2034),
    .d1(N56),
    .d2(N57),
    .o1(net180),
    .o2(net181),
    .si1(net911),
    .si2(net912),
    .ssb(net1630));
 b15fqy203ar1n02x5 cio_gpio_q_reg_18__cio_gpio_q_reg_19_ (.rb(net833),
    .clk(clknet_1_0__leaf_net2034),
    .d1(N58),
    .d2(N59),
    .o1(net182),
    .o2(net183),
    .si1(net913),
    .si2(net914),
    .ssb(net1631));
 b15fqy203ar1n02x5 cio_gpio_q_reg_20__cio_gpio_q_reg_21_ (.rb(net840),
    .clk(clknet_1_0__leaf_net2034),
    .d1(N60),
    .d2(N61),
    .o1(net185),
    .o2(net186),
    .si1(net915),
    .si2(net916),
    .ssb(net1632));
 b15fqy203ar1n02x5 cio_gpio_q_reg_22__cio_gpio_q_reg_23_ (.rb(net851),
    .clk(clknet_1_1__leaf_net2034),
    .d1(net306),
    .d2(net307),
    .o1(net187),
    .o2(net188),
    .si1(net917),
    .si2(net918),
    .ssb(net1633));
 b15fqy203ar1n02x5 cio_gpio_q_reg_24__cio_gpio_q_reg_25_ (.rb(net856),
    .clk(clknet_1_1__leaf_net2034),
    .d1(N64),
    .d2(N65),
    .o1(net189),
    .o2(net190),
    .si1(net919),
    .si2(net920),
    .ssb(net1634));
 b15fqy203ar1n02x5 cio_gpio_q_reg_26__cio_gpio_q_reg_27_ (.rb(net844),
    .clk(clknet_1_0__leaf_net2034),
    .d1(N66),
    .d2(N67),
    .o1(net191),
    .o2(net192),
    .si1(net921),
    .si2(net922),
    .ssb(net1635));
 b15fqy203ar1n02x5 cio_gpio_q_reg_28__cio_gpio_q_reg_29_ (.rb(net839),
    .clk(clknet_1_1__leaf_net2034),
    .d1(N68),
    .d2(N69),
    .o1(net193),
    .o2(net194),
    .si1(net923),
    .si2(net924),
    .ssb(net1636));
 b15fqy203ar1n02x5 cio_gpio_q_reg_2__cio_gpio_q_reg_3_ (.rb(net846),
    .clk(clknet_1_0__leaf_net2040),
    .d1(N41),
    .d2(N42),
    .o1(net195),
    .o2(net198),
    .si1(net925),
    .si2(net926),
    .ssb(net1637));
 b15fqy203ar1n02x5 cio_gpio_q_reg_30__cio_gpio_q_reg_31_ (.rb(net839),
    .clk(clknet_1_0__leaf_net2034),
    .d1(N70),
    .d2(N71),
    .o1(net196),
    .o2(net197),
    .si1(net927),
    .si2(net928),
    .ssb(net1638));
 b15fqy203ar1n02x5 cio_gpio_q_reg_4__cio_gpio_q_reg_5_ (.rb(net862),
    .clk(clknet_1_1__leaf_net2040),
    .d1(N43),
    .d2(N44),
    .o1(net199),
    .o2(net200),
    .si1(net929),
    .si2(net930),
    .ssb(net1639));
 b15fqy203ar1n02x5 cio_gpio_q_reg_6__cio_gpio_q_reg_7_ (.rb(net860),
    .clk(clknet_1_1__leaf_net2040),
    .d1(N45),
    .d2(N46),
    .o1(net201),
    .o2(net202),
    .si1(net931),
    .si2(net932),
    .ssb(net1640));
 b15fqy203ar1n02x5 cio_gpio_q_reg_8__cio_gpio_q_reg_9_ (.rb(net856),
    .clk(clknet_1_1__leaf_net2040),
    .d1(N47),
    .d2(N48),
    .o1(net203),
    .o2(net204),
    .si1(net933),
    .si2(net934),
    .ssb(net1641));
 b15cilb05ah1n02x3 clk_gate_cio_gpio_en_q_reg_0_latch (.clk(clknet_leaf_7_clk_i),
    .clkout(net2050),
    .en(N113),
    .te(net935));
 b15cilb05ah1n02x3 clk_gate_cio_gpio_en_q_reg_latch (.clk(clknet_leaf_7_clk_i),
    .clkout(net2045),
    .en(N130),
    .te(net936));
 b15cilb05ah1n02x3 clk_gate_cio_gpio_q_reg_0_latch (.clk(clknet_leaf_8_clk_i),
    .clkout(net2040),
    .en(N38),
    .te(net937));
 b15cilb05ah1n02x3 clk_gate_cio_gpio_q_reg_latch (.clk(clknet_leaf_9_clk_i),
    .clkout(net2034),
    .en(net314),
    .te(net938));
 b15fpy200ar1n02x5 data_in_q_reg_0__data_in_q_reg_1_ (.clk(clknet_leaf_4_clk_i),
    .d1(u_reg_u_data_in_wr_data[0]),
    .d2(u_reg_u_data_in_wr_data[1]),
    .o1(data_in_q[0]),
    .o2(data_in_q[1]),
    .si1(net939),
    .si2(net940),
    .ssb(net1642));
 b15fpy200ar1n02x5 data_in_q_reg_10__data_in_q_reg_11_ (.clk(clknet_leaf_9_clk_i),
    .d1(u_reg_u_data_in_wr_data[10]),
    .d2(net380),
    .o1(data_in_q[10]),
    .o2(data_in_q[11]),
    .si1(net941),
    .si2(net942),
    .ssb(net1643));
 b15fpy200ar1n02x5 data_in_q_reg_12__data_in_q_reg_13_ (.clk(clknet_leaf_8_clk_i),
    .d1(net377),
    .d2(u_reg_u_data_in_wr_data[13]),
    .o1(data_in_q[12]),
    .o2(data_in_q[13]),
    .si1(net943),
    .si2(net944),
    .ssb(net1644));
 b15fpy200ar1n02x5 data_in_q_reg_14__data_in_q_reg_15_ (.clk(clknet_leaf_9_clk_i),
    .d1(u_reg_u_data_in_wr_data[14]),
    .d2(net378),
    .o1(data_in_q[14]),
    .o2(data_in_q[15]),
    .si1(net945),
    .si2(net946),
    .ssb(net1645));
 b15fpy200ar1n02x5 data_in_q_reg_16__data_in_q_reg_17_ (.clk(clknet_leaf_4_clk_i),
    .d1(u_reg_u_data_in_wr_data[16]),
    .d2(u_reg_u_data_in_wr_data[17]),
    .o1(data_in_q[16]),
    .o2(data_in_q[17]),
    .si1(net947),
    .si2(net948),
    .ssb(net1646));
 b15fpy200ar1n02x5 data_in_q_reg_18__data_in_q_reg_19_ (.clk(clknet_leaf_11_clk_i),
    .d1(u_reg_u_data_in_wr_data[18]),
    .d2(u_reg_u_data_in_wr_data[19]),
    .o1(data_in_q[18]),
    .o2(data_in_q[19]),
    .si1(net949),
    .si2(net950),
    .ssb(net1647));
 b15fpy200ar1n02x5 data_in_q_reg_20__data_in_q_reg_21_ (.clk(clknet_leaf_10_clk_i),
    .d1(net376),
    .d2(u_reg_u_data_in_wr_data[21]),
    .o1(data_in_q[20]),
    .o2(data_in_q[21]),
    .si1(net951),
    .si2(net952),
    .ssb(net1648));
 b15fpy200ar1n02x5 data_in_q_reg_22__data_in_q_reg_23_ (.clk(clknet_leaf_9_clk_i),
    .d1(net375),
    .d2(u_reg_u_data_in_wr_data[23]),
    .o1(data_in_q[22]),
    .o2(data_in_q[23]),
    .si1(net953),
    .si2(net954),
    .ssb(net1649));
 b15fpy200ar1n02x5 data_in_q_reg_24__data_in_q_reg_25_ (.clk(clknet_leaf_1_clk_i),
    .d1(u_reg_u_data_in_wr_data[24]),
    .d2(u_reg_u_data_in_wr_data[25]),
    .o1(data_in_q[24]),
    .o2(data_in_q[25]),
    .si1(net955),
    .si2(net956),
    .ssb(net1650));
 b15fpy200ar1n02x5 data_in_q_reg_26__data_in_q_reg_27_ (.clk(clknet_leaf_1_clk_i),
    .d1(u_reg_u_data_in_wr_data[26]),
    .d2(u_reg_u_data_in_wr_data[27]),
    .o1(data_in_q[26]),
    .o2(data_in_q[27]),
    .si1(net957),
    .si2(net958),
    .ssb(net1651));
 b15fpy200ar1n02x5 data_in_q_reg_28__data_in_q_reg_29_ (.clk(clknet_leaf_10_clk_i),
    .d1(u_reg_u_data_in_wr_data[28]),
    .d2(u_reg_u_data_in_wr_data[29]),
    .o1(data_in_q[28]),
    .o2(data_in_q[29]),
    .si1(net959),
    .si2(net960),
    .ssb(net1652));
 b15fpy200ar1n02x5 data_in_q_reg_2__data_in_q_reg_3_ (.clk(clknet_leaf_9_clk_i),
    .d1(u_reg_u_data_in_wr_data[2]),
    .d2(net379),
    .o1(data_in_q[2]),
    .o2(data_in_q[3]),
    .si1(net961),
    .si2(net962),
    .ssb(net1653));
 b15fpy200ar1n02x5 data_in_q_reg_30__data_in_q_reg_31_ (.clk(clknet_leaf_1_clk_i),
    .d1(u_reg_u_data_in_wr_data[30]),
    .d2(u_reg_u_data_in_wr_data[31]),
    .o1(data_in_q[30]),
    .o2(data_in_q[31]),
    .si1(net963),
    .si2(net964),
    .ssb(net1654));
 b15fpy200ar1n02x5 data_in_q_reg_4__data_in_q_reg_5_ (.clk(clknet_leaf_9_clk_i),
    .d1(u_reg_u_data_in_wr_data[4]),
    .d2(net2355),
    .o1(data_in_q[4]),
    .o2(data_in_q[5]),
    .si1(net965),
    .si2(net966),
    .ssb(net1655));
 b15fpy200ar1n02x5 data_in_q_reg_6__data_in_q_reg_7_ (.clk(clknet_leaf_8_clk_i),
    .d1(u_reg_u_data_in_wr_data[6]),
    .d2(u_reg_u_data_in_wr_data[7]),
    .o1(data_in_q[6]),
    .o2(data_in_q[7]),
    .si1(net967),
    .si2(net968),
    .ssb(net1656));
 b15fpy200ar1n02x5 data_in_q_reg_8__data_in_q_reg_9_ (.clk(clknet_leaf_7_clk_i),
    .d1(u_reg_u_data_in_wr_data[8]),
    .d2(u_reg_u_data_in_wr_data[9]),
    .o1(data_in_q[8]),
    .o2(data_in_q[9]),
    .si1(net969),
    .si2(net970),
    .ssb(net1657));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_alert_set_q_reg_gen_filter_5__u_filter_filter_q_reg (.rb(net856),
    .clk(clknet_leaf_3_clk_i),
    .d1(gen_alert_tx_0__u_prim_alert_sender_alert_req_trigger),
    .d2(net741),
    .o1(gen_alert_tx_0__u_prim_alert_sender_n1),
    .o2(gen_filter_5__u_filter_filter_q),
    .si1(net971),
    .si2(net972),
    .ssb(net1658));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_0_ (.rb(net854),
    .clk(clknet_leaf_3_clk_i),
    .d1(gen_alert_tx_0__u_prim_alert_sender_alert_test_set_d),
    .d2(gen_alert_tx_0__u_prim_alert_sender_state_d[0]),
    .o1(gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q),
    .o2(gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .si1(net973),
    .si2(net974),
    .ssb(net1659));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_ping_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_1_ (.rb(net854),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2444),
    .d2(gen_alert_tx_0__u_prim_alert_sender_state_d[1]),
    .o1(gen_alert_tx_0__u_prim_alert_sender_ping_set_q),
    .o2(gen_alert_tx_0__u_prim_alert_sender_state_q[1]),
    .si1(net975),
    .si2(net976),
    .ssb(net1660));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_state_q_reg_2__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq_reg (.rb(net854),
    .clk(clknet_leaf_3_clk_i),
    .d1(gen_alert_tx_0__u_prim_alert_sender_state_d[2]),
    .d2(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .o1(gen_alert_tx_0__u_prim_alert_sender_state_q[2]),
    .o2(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq),
    .si1(net977),
    .si2(net978),
    .ssb(net1661));
 b15fqy00car1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq_reg (.clk(clknet_leaf_3_clk_i),
    .d(net2374),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq),
    .psb(net854),
    .si(net979),
    .ssb(net1662));
 b15fqy00car1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.clk(clknet_leaf_3_clk_i),
    .d(net1),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_intq_0_),
    .psb(net855),
    .si(net980),
    .ssb(net1663));
 b15fqy00car1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.clk(clknet_leaf_3_clk_i),
    .d(net2309),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nd),
    .psb(net855),
    .si(net981),
    .ssb(net1664));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net855),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2),
    .d2(net2266),
    .o1(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_intq_0_),
    .o2(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pd),
    .si1(net982),
    .si2(net983),
    .ssb(net1665));
 b15fqy043ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_0_ (.clk(clknet_leaf_3_clk_i),
    .d(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[0]),
    .den(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[0]),
    .rb(net855),
    .si(net984),
    .ssb(net1666));
 b15fqy043ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_1_ (.clk(clknet_leaf_2_clk_i),
    .d(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_d[1]),
    .den(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_N39),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[1]),
    .rb(net855),
    .si(net985),
    .ssb(net1667));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q_reg_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq_reg (.rb(net855),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2439),
    .d2(net2516),
    .o1(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q),
    .o2(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq),
    .si1(net986),
    .si2(net987),
    .ssb(net1668));
 b15fqy00car1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq_reg (.clk(clknet_leaf_2_clk_i),
    .d(net2533),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq),
    .psb(net854),
    .si(net988),
    .ssb(net1669));
 b15fqy00car1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.clk(clknet_leaf_2_clk_i),
    .d(net3),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_intq_0_),
    .psb(net854),
    .si(net989),
    .ssb(net1670));
 b15fqy00car1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.clk(clknet_leaf_2_clk_i),
    .d(net2230),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd),
    .psb(net854),
    .si(net990),
    .ssb(net1671));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net855),
    .clk(clknet_leaf_2_clk_i),
    .d1(net4),
    .d2(net2265),
    .o1(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_intq_0_),
    .o2(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd),
    .si1(net991),
    .si2(net992),
    .ssb(net1672));
 b15fqy043ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_0_ (.clk(clknet_leaf_2_clk_i),
    .d(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[0]),
    .den(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[0]),
    .rb(net854),
    .si(net993),
    .ssb(net1673));
 b15fqy043ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_1_ (.clk(clknet_leaf_2_clk_i),
    .d(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_d[1]),
    .den(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_N39),
    .o(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .rb(net854),
    .si(net994),
    .ssb(net1674));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q_reg_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net854),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_n3),
    .d2(net5),
    .o1(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q),
    .o2(gen_filter_0__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net995),
    .si2(net996),
    .ssb(net1675));
 b15fqy203ar1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_0__u_filter_diff_ctr_q_reg_0_ (.rb(net854),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_alert_tx_0__u_prim_alert_sender_alert_pd),
    .d2(net2387),
    .o1(net140),
    .o2(gen_filter_0__u_filter_diff_ctr_q[0]),
    .si1(net997),
    .si2(net998),
    .ssb(net1676));
 b15fqy00car1n02x5 gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_1_ (.clk(clknet_leaf_2_clk_i),
    .d(gen_alert_tx_0__u_prim_alert_sender_alert_nd),
    .o(net139),
    .psb(net854),
    .si(net999),
    .ssb(net1677));
 b15fqy203ar1n02x5 gen_filter_0__u_filter_diff_ctr_q_reg_1__gen_filter_0__u_filter_diff_ctr_q_reg_2_ (.rb(net854),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_filter_0__u_filter_diff_ctr_d[1]),
    .d2(net2508),
    .o1(gen_filter_0__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_0__u_filter_diff_ctr_q[2]),
    .si1(net1000),
    .si2(net1001),
    .ssb(net1678));
 b15fqy203ar1n02x5 gen_filter_0__u_filter_diff_ctr_q_reg_3__gen_filter_0__u_filter_filter_q_reg (.rb(net851),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_filter_0__u_filter_diff_ctr_d[3]),
    .d2(net2547),
    .o1(gen_filter_0__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_0__u_filter_filter_q),
    .si1(net1002),
    .si2(net1003),
    .ssb(net1679));
 b15fqy203ar1n02x5 gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_16__u_filter_diff_ctr_q_reg_0_ (.rb(net851),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2385),
    .d2(gen_filter_16__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_0__u_filter_filter_synced),
    .o2(gen_filter_16__u_filter_diff_ctr_q[0]),
    .si1(net1004),
    .si2(net1005),
    .ssb(net1680));
 b15fqy043ar1n02x5 gen_filter_0__u_filter_stored_value_q_reg (.clk(clknet_leaf_3_clk_i),
    .d(net755),
    .den(eq_x_181_n25),
    .o(gen_filter_0__u_filter_stored_value_q),
    .rb(net854),
    .si(net1006),
    .ssb(net1681));
 b15fqy203ar1n02x5 gen_filter_10__u_filter_diff_ctr_q_reg_0__gen_filter_10__u_filter_diff_ctr_q_reg_3_ (.rb(net862),
    .clk(clknet_leaf_5_clk_i),
    .d1(gen_filter_10__u_filter_diff_ctr_d[0]),
    .d2(gen_filter_10__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_10__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_10__u_filter_diff_ctr_q[3]),
    .si1(net1007),
    .si2(net1008),
    .ssb(net1682));
 b15fqy203ar1n02x5 gen_filter_10__u_filter_diff_ctr_q_reg_1__gen_filter_10__u_filter_diff_ctr_q_reg_2_ (.rb(net862),
    .clk(clknet_leaf_5_clk_i),
    .d1(gen_filter_10__u_filter_diff_ctr_d[1]),
    .d2(gen_filter_10__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_10__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_10__u_filter_diff_ctr_q[2]),
    .si1(net1009),
    .si2(net1010),
    .ssb(net1683));
 b15fqy203ar1n02x5 gen_filter_10__u_filter_filter_q_reg_gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net860),
    .clk(clknet_leaf_6_clk_i),
    .d1(gen_filter_10__u_filter_filter_synced),
    .d2(net2395),
    .o1(gen_filter_10__u_filter_filter_q),
    .o2(gen_filter_10__u_filter_filter_synced),
    .si1(net1011),
    .si2(net1012),
    .ssb(net1684));
 b15fqy043ar1n02x5 gen_filter_10__u_filter_stored_value_q_reg (.clk(clknet_leaf_4_clk_i),
    .d(gen_filter_10__u_filter_filter_synced),
    .den(eq_x_131_n25),
    .o(gen_filter_10__u_filter_stored_value_q),
    .rb(net862),
    .si(net1013),
    .ssb(net1685));
 b15fqy203ar1n02x5 gen_filter_11__u_filter_diff_ctr_q_reg_0__gen_filter_11__u_filter_diff_ctr_q_reg_1_ (.rb(net861),
    .clk(clknet_leaf_6_clk_i),
    .d1(gen_filter_11__u_filter_diff_ctr_d[0]),
    .d2(gen_filter_11__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_11__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_11__u_filter_diff_ctr_q[1]),
    .si1(net1014),
    .si2(net1015),
    .ssb(net1686));
 b15fqy203ar1n02x5 gen_filter_11__u_filter_diff_ctr_q_reg_3__gen_filter_11__u_filter_filter_q_reg (.rb(net861),
    .clk(clknet_leaf_6_clk_i),
    .d1(net2373),
    .d2(net2555),
    .o1(gen_filter_11__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_11__u_filter_filter_q),
    .si1(net1016),
    .si2(net1017),
    .ssb(net1687));
 b15fqy203ar1n02x5 gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net861),
    .clk(clknet_leaf_6_clk_i),
    .d1(net7),
    .d2(net2270),
    .o1(gen_filter_11__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_11__u_filter_filter_synced),
    .si1(net1018),
    .si2(net1019),
    .ssb(net1688));
 b15fqy043ar1n02x5 gen_filter_11__u_filter_stored_value_q_reg (.clk(clknet_leaf_6_clk_i),
    .d(gen_filter_11__u_filter_filter_synced),
    .den(eq_x_126_n25),
    .o(gen_filter_11__u_filter_stored_value_q),
    .rb(net861),
    .si(net1020),
    .ssb(net1689));
 b15fqy203ar1n02x5 gen_filter_12__u_filter_diff_ctr_q_reg_0__gen_filter_12__u_filter_diff_ctr_q_reg_1_ (.rb(net862),
    .clk(clknet_leaf_4_clk_i),
    .d1(gen_filter_12__u_filter_diff_ctr_d[0]),
    .d2(gen_filter_12__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_12__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_12__u_filter_diff_ctr_q[1]),
    .si1(net1021),
    .si2(net1022),
    .ssb(net1690));
 b15fqy203ar1n02x5 gen_filter_12__u_filter_diff_ctr_q_reg_2__gen_filter_12__u_filter_diff_ctr_q_reg_3_ (.rb(net859),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2328),
    .d2(gen_filter_12__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_12__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_12__u_filter_diff_ctr_q[3]),
    .si1(net1023),
    .si2(net1024),
    .ssb(net1691));
 b15fqy203ar1n02x5 gen_filter_12__u_filter_filter_q_reg_gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net861),
    .clk(clknet_leaf_7_clk_i),
    .d1(gen_filter_12__u_filter_filter_synced),
    .d2(net824),
    .o1(gen_filter_12__u_filter_filter_q),
    .o2(gen_filter_12__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1025),
    .si2(net1026),
    .ssb(net1692));
 b15fqy203ar1n02x5 gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_13__u_filter_diff_ctr_q_reg_0_ (.rb(net859),
    .clk(clknet_leaf_7_clk_i),
    .d1(net2310),
    .d2(gen_filter_13__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_12__u_filter_filter_synced),
    .o2(gen_filter_13__u_filter_diff_ctr_q[0]),
    .si1(net1027),
    .si2(net1028),
    .ssb(net1693));
 b15fqy043ar1n02x5 gen_filter_12__u_filter_stored_value_q_reg (.clk(clknet_leaf_4_clk_i),
    .d(gen_filter_12__u_filter_filter_synced),
    .den(eq_x_121_n25),
    .o(gen_filter_12__u_filter_stored_value_q),
    .rb(net859),
    .si(net1029),
    .ssb(net1694));
 b15fqy203ar1n02x5 gen_filter_13__u_filter_diff_ctr_q_reg_1__gen_filter_13__u_filter_diff_ctr_q_reg_2_ (.rb(net862),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2330),
    .d2(net2364),
    .o1(gen_filter_13__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_13__u_filter_diff_ctr_q[2]),
    .si1(net1030),
    .si2(net1031),
    .ssb(net1695));
 b15fqy203ar1n02x5 gen_filter_13__u_filter_diff_ctr_q_reg_3__gen_filter_13__u_filter_filter_q_reg (.rb(net863),
    .clk(clknet_leaf_6_clk_i),
    .d1(gen_filter_13__u_filter_diff_ctr_d[3]),
    .d2(gen_filter_13__u_filter_filter_synced),
    .o1(gen_filter_13__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_13__u_filter_filter_q),
    .si1(net1032),
    .si2(net1033),
    .ssb(net1696));
 b15fqy203ar1n02x5 gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net861),
    .clk(clknet_leaf_6_clk_i),
    .d1(net9),
    .d2(net2268),
    .o1(gen_filter_13__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_13__u_filter_filter_synced),
    .si1(net1034),
    .si2(net1035),
    .ssb(net1697));
 b15fqy043ar1n02x5 gen_filter_13__u_filter_stored_value_q_reg (.clk(clknet_leaf_6_clk_i),
    .d(gen_filter_13__u_filter_filter_synced),
    .den(eq_x_116_n25),
    .o(gen_filter_13__u_filter_stored_value_q),
    .rb(net861),
    .si(net1036),
    .ssb(net1698));
 b15fqy203ar1n02x5 gen_filter_14__u_filter_diff_ctr_q_reg_0__gen_filter_14__u_filter_diff_ctr_q_reg_1_ (.rb(net841),
    .clk(clknet_leaf_8_clk_i),
    .d1(net2464),
    .d2(gen_filter_14__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_14__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_14__u_filter_diff_ctr_q[1]),
    .si1(net1037),
    .si2(net1038),
    .ssb(net1699));
 b15fqy203ar1n02x5 gen_filter_14__u_filter_diff_ctr_q_reg_2__gen_filter_14__u_filter_diff_ctr_q_reg_3_ (.rb(net841),
    .clk(clknet_leaf_8_clk_i),
    .d1(gen_filter_14__u_filter_diff_ctr_d[2]),
    .d2(gen_filter_14__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_14__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_14__u_filter_diff_ctr_q[3]),
    .si1(net1039),
    .si2(net1040),
    .ssb(net1700));
 b15fqy203ar1n02x5 gen_filter_14__u_filter_filter_q_reg_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net840),
    .clk(clknet_leaf_9_clk_i),
    .d1(gen_filter_14__u_filter_filter_synced),
    .d2(net10),
    .o1(gen_filter_14__u_filter_filter_q),
    .o2(gen_filter_14__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1041),
    .si2(net1042),
    .ssb(net1701));
 b15fqy203ar1n02x5 gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net840),
    .clk(clknet_leaf_9_clk_i),
    .d1(net2301),
    .d2(net15),
    .o1(gen_filter_14__u_filter_filter_synced),
    .o2(gen_filter_19__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1043),
    .si2(net1044),
    .ssb(net1702));
 b15fqy043ar1n02x5 gen_filter_14__u_filter_stored_value_q_reg (.clk(clknet_leaf_9_clk_i),
    .d(gen_filter_14__u_filter_filter_synced),
    .den(eq_x_111_n25),
    .o(gen_filter_14__u_filter_stored_value_q),
    .rb(net841),
    .si(net1045),
    .ssb(net1703));
 b15fqy203ar1n02x5 gen_filter_15__u_filter_diff_ctr_q_reg_1__gen_filter_15__u_filter_diff_ctr_q_reg_2_ (.rb(net864),
    .clk(clknet_leaf_5_clk_i),
    .d1(gen_filter_15__u_filter_diff_ctr_d[1]),
    .d2(gen_filter_15__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_15__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_15__u_filter_diff_ctr_q[2]),
    .si1(net1046),
    .si2(net1047),
    .ssb(net1704));
 b15fqy203ar1n02x5 gen_filter_15__u_filter_diff_ctr_q_reg_3__gen_filter_15__u_filter_filter_q_reg (.rb(net864),
    .clk(clknet_leaf_5_clk_i),
    .d1(gen_filter_15__u_filter_diff_ctr_d[3]),
    .d2(gen_filter_15__u_filter_filter_synced),
    .o1(gen_filter_15__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_15__u_filter_filter_q),
    .si1(net1048),
    .si2(net1049),
    .ssb(net1705));
 b15fqy203ar1n02x5 gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net863),
    .clk(clknet_leaf_5_clk_i),
    .d1(net11),
    .d2(net2260),
    .o1(gen_filter_15__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_15__u_filter_filter_synced),
    .si1(net1050),
    .si2(net1051),
    .ssb(net1706));
 b15fqy043ar1n02x5 gen_filter_15__u_filter_stored_value_q_reg (.clk(clknet_leaf_5_clk_i),
    .d(gen_filter_15__u_filter_filter_synced),
    .den(eq_x_106_n25),
    .o(gen_filter_15__u_filter_stored_value_q),
    .rb(net862),
    .si(net1052),
    .ssb(net1707));
 b15fqy203ar1n02x5 gen_filter_16__u_filter_diff_ctr_q_reg_1__gen_filter_16__u_filter_diff_ctr_q_reg_2_ (.rb(net851),
    .clk(clknet_leaf_2_clk_i),
    .d1(net2461),
    .d2(net2369),
    .o1(gen_filter_16__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_16__u_filter_diff_ctr_q[2]),
    .si1(net1053),
    .si2(net1054),
    .ssb(net1708));
 b15fqy203ar1n02x5 gen_filter_16__u_filter_diff_ctr_q_reg_3__gen_filter_16__u_filter_filter_q_reg (.rb(net851),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_filter_16__u_filter_diff_ctr_d[3]),
    .d2(gen_filter_16__u_filter_filter_synced),
    .o1(gen_filter_16__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_16__u_filter_filter_q),
    .si1(net1055),
    .si2(net1056),
    .ssb(net1709));
 b15fqy203ar1n02x5 gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_diff_ctr_q_reg_0_ (.rb(net851),
    .clk(clknet_leaf_2_clk_i),
    .d1(net12),
    .d2(gen_filter_17__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_16__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_17__u_filter_diff_ctr_q[0]),
    .si1(net1057),
    .si2(net1058),
    .ssb(net1710));
 b15fqy203ar1n02x5 gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_30__u_filter_diff_ctr_q_reg_0_ (.rb(net837),
    .clk(clknet_leaf_1_clk_i),
    .d1(net2299),
    .d2(net2366),
    .o1(gen_filter_16__u_filter_filter_synced),
    .o2(gen_filter_30__u_filter_diff_ctr_q[0]),
    .si1(net1059),
    .si2(net1060),
    .ssb(net1711));
 b15fqy043ar1n02x5 gen_filter_16__u_filter_stored_value_q_reg (.clk(clknet_leaf_1_clk_i),
    .d(gen_filter_16__u_filter_filter_synced),
    .den(eq_x_101_n25),
    .o(gen_filter_16__u_filter_stored_value_q),
    .rb(net851),
    .si(net1061),
    .ssb(net1712));
 b15fqy203ar1n02x5 gen_filter_17__u_filter_diff_ctr_q_reg_1__gen_filter_17__u_filter_diff_ctr_q_reg_2_ (.rb(net851),
    .clk(clknet_leaf_1_clk_i),
    .d1(net2352),
    .d2(net2361),
    .o1(gen_filter_17__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_17__u_filter_diff_ctr_q[2]),
    .si1(net1062),
    .si2(net1063),
    .ssb(net1713));
 b15fqy203ar1n02x5 gen_filter_17__u_filter_diff_ctr_q_reg_3__gen_filter_17__u_filter_filter_q_reg (.rb(net851),
    .clk(clknet_leaf_1_clk_i),
    .d1(gen_filter_17__u_filter_diff_ctr_d[3]),
    .d2(net2545),
    .o1(gen_filter_17__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_17__u_filter_filter_q),
    .si1(net1064),
    .si2(net1065),
    .ssb(net1714));
 b15fqy203ar1n02x5 gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net851),
    .clk(clknet_leaf_2_clk_i),
    .d1(net13),
    .d2(net2267),
    .o1(gen_filter_17__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_17__u_filter_filter_synced),
    .si1(net1066),
    .si2(net1067),
    .ssb(net1715));
 b15fqy043ar1n02x5 gen_filter_17__u_filter_stored_value_q_reg (.clk(clknet_leaf_1_clk_i),
    .d(gen_filter_17__u_filter_filter_synced),
    .den(eq_x_96_n25),
    .o(gen_filter_17__u_filter_stored_value_q),
    .rb(net851),
    .si(net1068),
    .ssb(net1716));
 b15fqy203ar1n02x5 gen_filter_18__u_filter_diff_ctr_q_reg_0__gen_filter_18__u_filter_diff_ctr_q_reg_1_ (.rb(net833),
    .clk(clknet_leaf_0_clk_i),
    .d1(gen_filter_18__u_filter_diff_ctr_d[0]),
    .d2(gen_filter_18__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_18__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_18__u_filter_diff_ctr_q[1]),
    .si1(net1069),
    .si2(net1070),
    .ssb(net1717));
 b15fqy203ar1n02x5 gen_filter_18__u_filter_diff_ctr_q_reg_2__gen_filter_18__u_filter_diff_ctr_q_reg_3_ (.rb(net833),
    .clk(clknet_leaf_0_clk_i),
    .d1(gen_filter_18__u_filter_diff_ctr_d[2]),
    .d2(gen_filter_18__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_18__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_18__u_filter_diff_ctr_q[3]),
    .si1(net1071),
    .si2(net1072),
    .ssb(net1718));
 b15fqy203ar1n02x5 gen_filter_18__u_filter_filter_q_reg_gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net833),
    .clk(clknet_leaf_11_clk_i),
    .d1(gen_filter_18__u_filter_filter_synced),
    .d2(net14),
    .o1(gen_filter_18__u_filter_filter_q),
    .o2(gen_filter_18__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1073),
    .si2(net1074),
    .ssb(net1719));
 b15fqy203ar1n02x5 gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_diff_ctr_q_reg_0_ (.rb(net833),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2272),
    .d2(net2359),
    .o1(gen_filter_18__u_filter_filter_synced),
    .o2(gen_filter_19__u_filter_diff_ctr_q[0]),
    .si1(net1075),
    .si2(net1076),
    .ssb(net1720));
 b15fqy043ar1n02x5 gen_filter_18__u_filter_stored_value_q_reg (.clk(clknet_leaf_0_clk_i),
    .d(gen_filter_18__u_filter_filter_synced),
    .den(eq_x_91_n25),
    .o(gen_filter_18__u_filter_stored_value_q),
    .rb(net833),
    .si(net1077),
    .ssb(net1721));
 b15fqy203ar1n02x5 gen_filter_19__u_filter_diff_ctr_q_reg_1__gen_filter_19__u_filter_diff_ctr_q_reg_2_ (.rb(net833),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2475),
    .d2(gen_filter_19__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_19__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_19__u_filter_diff_ctr_q[2]),
    .si1(net1078),
    .si2(net1079),
    .ssb(net1722));
 b15fqy203ar1n02x5 gen_filter_19__u_filter_diff_ctr_q_reg_3__gen_filter_19__u_filter_filter_q_reg (.rb(net833),
    .clk(clknet_leaf_11_clk_i),
    .d1(gen_filter_19__u_filter_diff_ctr_d[3]),
    .d2(gen_filter_19__u_filter_filter_synced),
    .o1(gen_filter_19__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_19__u_filter_filter_q),
    .si1(net1080),
    .si2(net1081),
    .ssb(net1723));
 b15fqy203ar1n02x5 gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_21__u_filter_diff_ctr_q_reg_0_ (.rb(net833),
    .clk(clknet_leaf_11_clk_i),
    .d1(gen_filter_19__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .d2(gen_filter_21__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_19__u_filter_filter_synced),
    .o2(gen_filter_21__u_filter_diff_ctr_q[0]),
    .si1(net1082),
    .si2(net1083),
    .ssb(net1724));
 b15fqy043ar1n02x5 gen_filter_19__u_filter_stored_value_q_reg (.clk(clknet_leaf_11_clk_i),
    .d(gen_filter_19__u_filter_filter_synced),
    .den(eq_x_86_n25),
    .o(gen_filter_19__u_filter_stored_value_q),
    .rb(net833),
    .si(net1084),
    .ssb(net1725));
 b15fqy203ar1n02x5 gen_filter_1__u_filter_diff_ctr_q_reg_0__gen_filter_1__u_filter_diff_ctr_q_reg_1_ (.rb(net855),
    .clk(clknet_leaf_3_clk_i),
    .d1(net2500),
    .d2(net2451),
    .o1(gen_filter_1__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_1__u_filter_diff_ctr_q[1]),
    .si1(net1085),
    .si2(net1086),
    .ssb(net1726));
 b15fqy203ar1n02x5 gen_filter_1__u_filter_diff_ctr_q_reg_2__gen_filter_1__u_filter_diff_ctr_q_reg_3_ (.rb(net856),
    .clk(clknet_leaf_3_clk_i),
    .d1(net2488),
    .d2(net2425),
    .o1(gen_filter_1__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_1__u_filter_diff_ctr_q[3]),
    .si1(net1087),
    .si2(net1088),
    .ssb(net1727));
 b15fqy203ar1n02x5 gen_filter_1__u_filter_filter_q_reg_gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net856),
    .clk(clknet_leaf_3_clk_i),
    .d1(gen_filter_1__u_filter_filter_synced),
    .d2(net16),
    .o1(gen_filter_1__u_filter_filter_q),
    .o2(gen_filter_1__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1089),
    .si2(net1090),
    .ssb(net1728));
 b15fqy203ar1n02x5 gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__intr_hw_intr_o_reg_0_ (.rb(net856),
    .clk(clknet_leaf_3_clk_i),
    .d1(net2271),
    .d2(intr_hw_N32),
    .o1(gen_filter_1__u_filter_filter_synced),
    .o2(net205),
    .si1(net1091),
    .si2(net1092),
    .ssb(net1729));
 b15fqy043ar1n02x5 gen_filter_1__u_filter_stored_value_q_reg (.clk(clknet_leaf_3_clk_i),
    .d(gen_filter_1__u_filter_filter_synced),
    .den(eq_x_176_n25),
    .o(gen_filter_1__u_filter_stored_value_q),
    .rb(net856),
    .si(net1093),
    .ssb(net1730));
 b15fqy203ar1n02x5 gen_filter_20__u_filter_diff_ctr_q_reg_0__gen_filter_20__u_filter_diff_ctr_q_reg_1_ (.rb(net838),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2421),
    .d2(net2437),
    .o1(gen_filter_20__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_20__u_filter_diff_ctr_q[1]),
    .si1(net1094),
    .si2(net1095),
    .ssb(net1731));
 b15fqy203ar1n02x5 gen_filter_20__u_filter_diff_ctr_q_reg_2__gen_filter_20__u_filter_diff_ctr_q_reg_3_ (.rb(net838),
    .clk(clknet_leaf_0_clk_i),
    .d1(gen_filter_20__u_filter_diff_ctr_d[2]),
    .d2(gen_filter_20__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_20__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_20__u_filter_diff_ctr_q[3]),
    .si1(net1096),
    .si2(net1097),
    .ssb(net1732));
 b15fqy203ar1n02x5 gen_filter_20__u_filter_filter_q_reg_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net836),
    .clk(clknet_leaf_11_clk_i),
    .d1(net754),
    .d2(net870),
    .o1(gen_filter_20__u_filter_filter_q),
    .o2(gen_filter_20__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1098),
    .si2(net1099),
    .ssb(net1733));
 b15fqy203ar1n02x5 gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_diff_ctr_q_reg_0_ (.rb(net839),
    .clk(clknet_leaf_1_clk_i),
    .d1(net2390),
    .d2(gen_filter_23__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_20__u_filter_filter_synced),
    .o2(gen_filter_23__u_filter_diff_ctr_q[0]),
    .si1(net1100),
    .si2(net1101),
    .ssb(net1734));
 b15fqy043ar1n02x5 gen_filter_20__u_filter_stored_value_q_reg (.clk(clknet_leaf_0_clk_i),
    .d(gen_filter_20__u_filter_filter_synced),
    .den(eq_x_81_n25),
    .o(gen_filter_20__u_filter_stored_value_q),
    .rb(net838),
    .si(net1102),
    .ssb(net1735));
 b15fqy203ar1n02x5 gen_filter_21__u_filter_diff_ctr_q_reg_1__gen_filter_21__u_filter_diff_ctr_q_reg_2_ (.rb(net833),
    .clk(clknet_leaf_11_clk_i),
    .d1(gen_filter_21__u_filter_diff_ctr_d[1]),
    .d2(net2469),
    .o1(gen_filter_21__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_21__u_filter_diff_ctr_q[2]),
    .si1(net1103),
    .si2(net1104),
    .ssb(net1736));
 b15fqy203ar1n02x5 gen_filter_21__u_filter_diff_ctr_q_reg_3__gen_filter_21__u_filter_filter_q_reg (.rb(net833),
    .clk(clknet_leaf_11_clk_i),
    .d1(gen_filter_21__u_filter_diff_ctr_d[3]),
    .d2(net2541),
    .o1(gen_filter_21__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_21__u_filter_filter_q),
    .si1(net1105),
    .si2(net1106),
    .ssb(net1737));
 b15fqy203ar1n02x5 gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net833),
    .clk(clknet_leaf_11_clk_i),
    .d1(net18),
    .d2(net2255),
    .o1(gen_filter_21__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_21__u_filter_filter_synced),
    .si1(net1107),
    .si2(net1108),
    .ssb(net1738));
 b15fqy043ar1n02x5 gen_filter_21__u_filter_stored_value_q_reg (.clk(clknet_leaf_11_clk_i),
    .d(gen_filter_21__u_filter_filter_synced),
    .den(eq_x_76_n25),
    .o(gen_filter_21__u_filter_stored_value_q),
    .rb(net833),
    .si(net1109),
    .ssb(net1739));
 b15fqy203ar1n02x5 gen_filter_22__u_filter_diff_ctr_q_reg_0__gen_filter_22__u_filter_diff_ctr_q_reg_1_ (.rb(net852),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_filter_22__u_filter_diff_ctr_d[0]),
    .d2(gen_filter_22__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_22__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_22__u_filter_diff_ctr_q[1]),
    .si1(net1110),
    .si2(net1111),
    .ssb(net1740));
 b15fqy203ar1n02x5 gen_filter_22__u_filter_diff_ctr_q_reg_2__gen_filter_22__u_filter_diff_ctr_q_reg_3_ (.rb(net852),
    .clk(clknet_leaf_1_clk_i),
    .d1(gen_filter_22__u_filter_diff_ctr_d[2]),
    .d2(net2336),
    .o1(gen_filter_22__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_22__u_filter_diff_ctr_q[3]),
    .si1(net1112),
    .si2(net1113),
    .ssb(net1741));
 b15fqy203ar1n02x5 gen_filter_22__u_filter_filter_q_reg_gen_filter_24__u_filter_diff_ctr_q_reg_0_ (.rb(net854),
    .clk(clknet_leaf_2_clk_i),
    .d1(net752),
    .d2(gen_filter_24__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_22__u_filter_filter_q),
    .o2(gen_filter_24__u_filter_diff_ctr_q[0]),
    .si1(net1114),
    .si2(net1115),
    .ssb(net1742));
 b15fqy203ar1n02x5 gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net856),
    .clk(clknet_leaf_3_clk_i),
    .d1(net19),
    .d2(net2253),
    .o1(gen_filter_22__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_22__u_filter_filter_synced),
    .si1(net1116),
    .si2(net1117),
    .ssb(net1743));
 b15fqy043ar1n02x5 gen_filter_22__u_filter_stored_value_q_reg (.clk(clknet_leaf_4_clk_i),
    .d(net2501),
    .den(eq_x_71_n25),
    .o(gen_filter_22__u_filter_stored_value_q),
    .rb(net853),
    .si(net1118),
    .ssb(net1744));
 b15fqy203ar1n02x5 gen_filter_23__u_filter_diff_ctr_q_reg_1__gen_filter_23__u_filter_diff_ctr_q_reg_2_ (.rb(net852),
    .clk(clknet_leaf_1_clk_i),
    .d1(net2529),
    .d2(net2377),
    .o1(gen_filter_23__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_23__u_filter_diff_ctr_q[2]),
    .si1(net1119),
    .si2(net1120),
    .ssb(net1745));
 b15fqy203ar1n02x5 gen_filter_23__u_filter_diff_ctr_q_reg_3__gen_filter_23__u_filter_filter_q_reg (.rb(net853),
    .clk(clknet_leaf_1_clk_i),
    .d1(gen_filter_23__u_filter_diff_ctr_d[3]),
    .d2(net749),
    .o1(gen_filter_23__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_23__u_filter_filter_q),
    .si1(net1121),
    .si2(net1122),
    .ssb(net1746));
 b15fqy203ar1n02x5 gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net840),
    .clk(clknet_leaf_9_clk_i),
    .d1(net20),
    .d2(net2262),
    .o1(gen_filter_23__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_23__u_filter_filter_synced),
    .si1(net1123),
    .si2(net1124),
    .ssb(net1747));
 b15fqy043ar1n02x5 gen_filter_23__u_filter_stored_value_q_reg (.clk(clknet_leaf_4_clk_i),
    .d(net750),
    .den(eq_x_66_n25),
    .o(gen_filter_23__u_filter_stored_value_q),
    .rb(net853),
    .si(net1125),
    .ssb(net1748));
 b15fqy203ar1n02x5 gen_filter_24__u_filter_diff_ctr_q_reg_1__gen_filter_24__u_filter_diff_ctr_q_reg_3_ (.rb(net852),
    .clk(clknet_leaf_1_clk_i),
    .d1(net2320),
    .d2(net2324),
    .o1(gen_filter_24__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_24__u_filter_diff_ctr_q[3]),
    .si1(net1126),
    .si2(net1127),
    .ssb(net1749));
 b15fqy203ar1n02x5 gen_filter_24__u_filter_diff_ctr_q_reg_2__gen_filter_24__u_filter_filter_q_reg (.rb(net852),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_filter_24__u_filter_diff_ctr_d[2]),
    .d2(gen_filter_24__u_filter_filter_synced),
    .o1(gen_filter_24__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_24__u_filter_filter_q),
    .si1(net1128),
    .si2(net1129),
    .ssb(net1750));
 b15fqy203ar1n02x5 gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net852),
    .clk(clknet_leaf_2_clk_i),
    .d1(net21),
    .d2(net2263),
    .o1(gen_filter_24__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_24__u_filter_filter_synced),
    .si1(net1130),
    .si2(net1131),
    .ssb(net1751));
 b15fqy043ar1n02x5 gen_filter_24__u_filter_stored_value_q_reg (.clk(clknet_leaf_1_clk_i),
    .d(gen_filter_24__u_filter_filter_synced),
    .den(eq_x_61_n25),
    .o(gen_filter_24__u_filter_stored_value_q),
    .rb(net852),
    .si(net1132),
    .ssb(net1752));
 b15fqy203ar1n02x5 gen_filter_25__u_filter_diff_ctr_q_reg_0__gen_filter_25__u_filter_diff_ctr_q_reg_1_ (.rb(net856),
    .clk(clknet_leaf_3_clk_i),
    .d1(gen_filter_25__u_filter_diff_ctr_d[0]),
    .d2(gen_filter_25__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_25__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_25__u_filter_diff_ctr_q[1]),
    .si1(net1133),
    .si2(net1134),
    .ssb(net1753));
 b15fqy203ar1n02x5 gen_filter_25__u_filter_diff_ctr_q_reg_2__gen_filter_25__u_filter_diff_ctr_q_reg_3_ (.rb(net853),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2434),
    .d2(gen_filter_25__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_25__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_25__u_filter_diff_ctr_q[3]),
    .si1(net1135),
    .si2(net1136),
    .ssb(net1754));
 b15fqy003ar1n02x5 gen_filter_25__u_filter_filter_q_reg (.rb(net853),
    .clk(clknet_leaf_1_clk_i),
    .d(net748),
    .o(gen_filter_25__u_filter_filter_q),
    .si(net1137),
    .ssb(net1755));
 b15fqy203ar1n02x5 gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net862),
    .clk(clknet_leaf_5_clk_i),
    .d1(net22),
    .d2(net2261),
    .o1(gen_filter_25__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_25__u_filter_filter_synced),
    .si1(net1138),
    .si2(net1139),
    .ssb(net1756));
 b15fqy043ar1n02x5 gen_filter_25__u_filter_stored_value_q_reg (.clk(clknet_leaf_4_clk_i),
    .d(net748),
    .den(eq_x_56_n25),
    .o(gen_filter_25__u_filter_stored_value_q),
    .rb(net856),
    .si(net1140),
    .ssb(net1757));
 b15fqy203ar1n02x5 gen_filter_26__u_filter_diff_ctr_q_reg_0__gen_filter_26__u_filter_diff_ctr_q_reg_1_ (.rb(net851),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_filter_26__u_filter_diff_ctr_d[0]),
    .d2(net2524),
    .o1(gen_filter_26__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_26__u_filter_diff_ctr_q[1]),
    .si1(net1141),
    .si2(net1142),
    .ssb(net1758));
 b15fqy203ar1n02x5 gen_filter_26__u_filter_diff_ctr_q_reg_2__gen_filter_26__u_filter_diff_ctr_q_reg_3_ (.rb(net851),
    .clk(clknet_leaf_2_clk_i),
    .d1(gen_filter_26__u_filter_diff_ctr_d[2]),
    .d2(net2480),
    .o1(gen_filter_26__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_26__u_filter_diff_ctr_q[3]),
    .si1(net1143),
    .si2(net1144),
    .ssb(net1759));
 b15fqy203ar1n02x5 gen_filter_26__u_filter_filter_q_reg_gen_filter_31__u_filter_diff_ctr_q_reg_0_ (.rb(net837),
    .clk(clknet_leaf_0_clk_i),
    .d1(gen_filter_26__u_filter_filter_synced),
    .d2(gen_filter_31__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_26__u_filter_filter_q),
    .o2(gen_filter_31__u_filter_diff_ctr_q[0]),
    .si1(net1145),
    .si2(net1146),
    .ssb(net1760));
 b15fqy203ar1n02x5 gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_diff_ctr_q_reg_0_ (.rb(net838),
    .clk(clknet_leaf_0_clk_i),
    .d1(net23),
    .d2(gen_filter_28__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_26__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_28__u_filter_diff_ctr_q[0]),
    .si1(net1147),
    .si2(net1148),
    .ssb(net1761));
 b15fqy203ar1n02x5 gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_31__u_filter_diff_ctr_q_reg_1_ (.rb(net837),
    .clk(clknet_leaf_0_clk_i),
    .d1(gen_filter_26__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .d2(gen_filter_31__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_26__u_filter_filter_synced),
    .o2(gen_filter_31__u_filter_diff_ctr_q[1]),
    .si1(net1149),
    .si2(net1150),
    .ssb(net1762));
 b15fqy043ar1n02x5 gen_filter_26__u_filter_stored_value_q_reg (.clk(clknet_leaf_0_clk_i),
    .d(gen_filter_26__u_filter_filter_synced),
    .den(eq_x_51_n25),
    .o(gen_filter_26__u_filter_stored_value_q),
    .rb(net837),
    .si(net1151),
    .ssb(net1763));
 b15fqy203ar1n02x5 gen_filter_27__u_filter_diff_ctr_q_reg_0__gen_filter_27__u_filter_diff_ctr_q_reg_1_ (.rb(net838),
    .clk(clknet_leaf_0_clk_i),
    .d1(gen_filter_27__u_filter_diff_ctr_d[0]),
    .d2(net2459),
    .o1(gen_filter_27__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_27__u_filter_diff_ctr_q[1]),
    .si1(net1152),
    .si2(net1153),
    .ssb(net1764));
 b15fqy203ar1n02x5 gen_filter_27__u_filter_diff_ctr_q_reg_2__gen_filter_27__u_filter_diff_ctr_q_reg_3_ (.rb(net838),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2441),
    .d2(gen_filter_27__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_27__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_27__u_filter_diff_ctr_q[3]),
    .si1(net1154),
    .si2(net1155),
    .ssb(net1765));
 b15fqy203ar1n02x5 gen_filter_27__u_filter_filter_q_reg_gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net838),
    .clk(clknet_leaf_0_clk_i),
    .d1(gen_filter_27__u_filter_filter_synced),
    .d2(net24),
    .o1(gen_filter_27__u_filter_filter_q),
    .o2(gen_filter_27__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1156),
    .si2(net1157),
    .ssb(net1766));
 b15fqy203ar1n02x5 gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_30__u_filter_diff_ctr_q_reg_1_ (.rb(net838),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2273),
    .d2(gen_filter_30__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_27__u_filter_filter_synced),
    .o2(gen_filter_30__u_filter_diff_ctr_q[1]),
    .si1(net1158),
    .si2(net1159),
    .ssb(net1767));
 b15fqy043ar1n02x5 gen_filter_27__u_filter_stored_value_q_reg (.clk(clknet_leaf_0_clk_i),
    .d(gen_filter_27__u_filter_filter_synced),
    .den(eq_x_46_n25),
    .o(gen_filter_27__u_filter_stored_value_q),
    .rb(net838),
    .si(net1160),
    .ssb(net1768));
 b15fqy203ar1n02x5 gen_filter_28__u_filter_diff_ctr_q_reg_1__gen_filter_28__u_filter_diff_ctr_q_reg_2_ (.rb(net836),
    .clk(clknet_leaf_0_clk_i),
    .d1(gen_filter_28__u_filter_diff_ctr_d[1]),
    .d2(gen_filter_28__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_28__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_28__u_filter_diff_ctr_q[2]),
    .si1(net1161),
    .si2(net1162),
    .ssb(net1769));
 b15fqy203ar1n02x5 gen_filter_28__u_filter_diff_ctr_q_reg_3__gen_filter_28__u_filter_filter_q_reg (.rb(net833),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2455),
    .d2(gen_filter_28__u_filter_filter_synced),
    .o1(gen_filter_28__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_28__u_filter_filter_q),
    .si1(net1163),
    .si2(net1164),
    .ssb(net1770));
 b15fqy203ar1n02x5 gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net836),
    .clk(clknet_leaf_0_clk_i),
    .d1(net25),
    .d2(net2264),
    .o1(gen_filter_28__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_28__u_filter_filter_synced),
    .si1(net1165),
    .si2(net1166),
    .ssb(net1771));
 b15fqy043ar1n02x5 gen_filter_28__u_filter_stored_value_q_reg (.clk(clknet_leaf_0_clk_i),
    .d(gen_filter_28__u_filter_filter_synced),
    .den(eq_x_41_n25),
    .o(gen_filter_28__u_filter_stored_value_q),
    .rb(net836),
    .si(net1167),
    .ssb(net1772));
 b15fqy203ar1n02x5 gen_filter_29__u_filter_diff_ctr_q_reg_0__gen_filter_29__u_filter_diff_ctr_q_reg_1_ (.rb(net838),
    .clk(clknet_leaf_0_clk_i),
    .d1(net2392),
    .d2(gen_filter_29__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_29__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_29__u_filter_diff_ctr_q[1]),
    .si1(net1168),
    .si2(net1169),
    .ssb(net1773));
 b15fqy203ar1n02x5 gen_filter_29__u_filter_diff_ctr_q_reg_2__gen_filter_29__u_filter_diff_ctr_q_reg_3_ (.rb(net838),
    .clk(clknet_leaf_1_clk_i),
    .d1(net2411),
    .d2(gen_filter_29__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_29__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_29__u_filter_diff_ctr_q[3]),
    .si1(net1170),
    .si2(net1171),
    .ssb(net1774));
 b15fqy003ar1n02x5 gen_filter_29__u_filter_filter_q_reg (.rb(net838),
    .clk(clknet_leaf_1_clk_i),
    .d(net747),
    .o(gen_filter_29__u_filter_filter_q),
    .si(net1172),
    .ssb(net1775));
 b15fqy203ar1n02x5 gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net834),
    .clk(clknet_leaf_11_clk_i),
    .d1(net26),
    .d2(net2254),
    .o1(gen_filter_29__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_29__u_filter_filter_synced),
    .si1(net1173),
    .si2(net1174),
    .ssb(net1776));
 b15fqy043ar1n02x5 gen_filter_29__u_filter_stored_value_q_reg (.clk(clknet_leaf_1_clk_i),
    .d(net747),
    .den(eq_x_36_n25),
    .o(gen_filter_29__u_filter_stored_value_q),
    .rb(net838),
    .si(net1175),
    .ssb(net1777));
 b15fqy203ar1n02x5 gen_filter_2__u_filter_diff_ctr_q_reg_0__gen_filter_2__u_filter_diff_ctr_q_reg_1_ (.rb(net862),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2431),
    .d2(net2397),
    .o1(gen_filter_2__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_2__u_filter_diff_ctr_q[1]),
    .si1(net1176),
    .si2(net1177),
    .ssb(net1778));
 b15fqy203ar1n02x5 gen_filter_2__u_filter_diff_ctr_q_reg_2__gen_filter_2__u_filter_diff_ctr_q_reg_3_ (.rb(net862),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2514),
    .d2(net2405),
    .o1(gen_filter_2__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_2__u_filter_diff_ctr_q[3]),
    .si1(net1178),
    .si2(net1179),
    .ssb(net1779));
 b15fqy203ar1n02x5 gen_filter_2__u_filter_filter_q_reg_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net862),
    .clk(clknet_leaf_4_clk_i),
    .d1(gen_filter_2__u_filter_filter_synced),
    .d2(net869),
    .o1(gen_filter_2__u_filter_filter_q),
    .o2(gen_filter_2__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1180),
    .si2(net1181),
    .ssb(net1780));
 b15fqy203ar1n02x5 gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_3__u_filter_diff_ctr_q_reg_0_ (.rb(net859),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2325),
    .d2(gen_filter_3__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_2__u_filter_filter_synced),
    .o2(gen_filter_3__u_filter_diff_ctr_q[0]),
    .si1(net1182),
    .si2(net1183),
    .ssb(net1781));
 b15fqy043ar1n02x5 gen_filter_2__u_filter_stored_value_q_reg (.clk(clknet_leaf_4_clk_i),
    .d(gen_filter_2__u_filter_filter_synced),
    .den(eq_x_171_n25),
    .o(gen_filter_2__u_filter_stored_value_q),
    .rb(net859),
    .si(net1184),
    .ssb(net1782));
 b15fqy203ar1n02x5 gen_filter_30__u_filter_diff_ctr_q_reg_2__gen_filter_30__u_filter_diff_ctr_q_reg_3_ (.rb(net837),
    .clk(clknet_leaf_0_clk_i),
    .d1(gen_filter_30__u_filter_diff_ctr_d[2]),
    .d2(gen_filter_30__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_30__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_30__u_filter_diff_ctr_q[3]),
    .si1(net1185),
    .si2(net1186),
    .ssb(net1783));
 b15fqy203ar1n02x5 gen_filter_30__u_filter_filter_q_reg_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net837),
    .clk(clknet_leaf_0_clk_i),
    .d1(gen_filter_30__u_filter_filter_synced),
    .d2(net28),
    .o1(gen_filter_30__u_filter_filter_q),
    .o2(gen_filter_30__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1187),
    .si2(net1188),
    .ssb(net1784));
 b15fqy003ar1n02x5 gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net838),
    .clk(clknet_leaf_1_clk_i),
    .d(net2356),
    .o(gen_filter_30__u_filter_filter_synced),
    .si(net1189),
    .ssb(net1785));
 b15fqy043ar1n02x5 gen_filter_30__u_filter_stored_value_q_reg (.clk(clknet_leaf_0_clk_i),
    .d(gen_filter_30__u_filter_filter_synced),
    .den(eq_x_31_n25),
    .o(gen_filter_30__u_filter_stored_value_q),
    .rb(net837),
    .si(net1190),
    .ssb(net1786));
 b15fqy203ar1n02x5 gen_filter_31__u_filter_diff_ctr_q_reg_2__gen_filter_31__u_filter_diff_ctr_q_reg_3_ (.rb(net837),
    .clk(clknet_leaf_1_clk_i),
    .d1(net2536),
    .d2(net2631),
    .o1(gen_filter_31__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_31__u_filter_diff_ctr_q[3]),
    .si1(net1191),
    .si2(net1192),
    .ssb(net1787));
 b15fqy203ar1n02x5 gen_filter_31__u_filter_filter_q_reg_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net852),
    .clk(clknet_leaf_1_clk_i),
    .d1(net2348),
    .d2(net29),
    .o1(gen_filter_31__u_filter_filter_q),
    .o2(gen_filter_31__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1193),
    .si2(net1194),
    .ssb(net1788));
 b15fqy203ar1n02x5 gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_reg_err_q_reg (.rb(net854),
    .clk(clknet_leaf_3_clk_i),
    .d1(gen_filter_31__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .d2(n1439),
    .o1(gen_filter_31__u_filter_filter_synced),
    .o2(u_reg_err_q),
    .si1(net1195),
    .si2(net1196),
    .ssb(net1789));
 b15fqy043ar1n02x5 gen_filter_31__u_filter_stored_value_q_reg (.clk(clknet_leaf_1_clk_i),
    .d(net746),
    .den(eq_x_26_n25),
    .o(gen_filter_31__u_filter_stored_value_q),
    .rb(net837),
    .si(net1197),
    .ssb(net1790));
 b15fqy203ar1n02x5 gen_filter_3__u_filter_diff_ctr_q_reg_1__gen_filter_3__u_filter_diff_ctr_q_reg_2_ (.rb(net853),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2486),
    .d2(gen_filter_3__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_3__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_3__u_filter_diff_ctr_q[2]),
    .si1(net1198),
    .si2(net1199),
    .ssb(net1791));
 b15fqy203ar1n02x5 gen_filter_3__u_filter_diff_ctr_q_reg_3__gen_filter_3__u_filter_filter_q_reg (.rb(net859),
    .clk(clknet_leaf_4_clk_i),
    .d1(gen_filter_3__u_filter_diff_ctr_d[3]),
    .d2(net745),
    .o1(gen_filter_3__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_3__u_filter_filter_q),
    .si1(net1200),
    .si2(net1201),
    .ssb(net1792));
 b15fqy203ar1n02x5 gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_4__u_filter_diff_ctr_q_reg_1_ (.rb(net863),
    .clk(clknet_leaf_6_clk_i),
    .d1(net30),
    .d2(gen_filter_4__u_filter_diff_ctr_d[1]),
    .o1(gen_filter_3__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_4__u_filter_diff_ctr_q[1]),
    .si1(net1202),
    .si2(net1203),
    .ssb(net1793));
 b15fqy203ar1n02x5 gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_8__u_filter_diff_ctr_q_reg_0_ (.rb(net863),
    .clk(clknet_leaf_6_clk_i),
    .d1(net2258),
    .d2(gen_filter_8__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_3__u_filter_filter_synced),
    .o2(gen_filter_8__u_filter_diff_ctr_q[0]),
    .si1(net1204),
    .si2(net1205),
    .ssb(net1794));
 b15fqy043ar1n02x5 gen_filter_3__u_filter_stored_value_q_reg (.clk(clknet_leaf_4_clk_i),
    .d(net744),
    .den(eq_x_166_n25),
    .o(gen_filter_3__u_filter_stored_value_q),
    .rb(net853),
    .si(net1206),
    .ssb(net1795));
 b15fqy203ar1n02x5 gen_filter_4__u_filter_diff_ctr_q_reg_0__gen_filter_4__u_filter_diff_ctr_q_reg_2_ (.rb(net863),
    .clk(clknet_leaf_6_clk_i),
    .d1(net2532),
    .d2(net2504),
    .o1(gen_filter_4__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_4__u_filter_diff_ctr_q[2]),
    .si1(net1207),
    .si2(net1208),
    .ssb(net1796));
 b15fqy203ar1n02x5 gen_filter_4__u_filter_diff_ctr_q_reg_3__gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net864),
    .clk(clknet_leaf_6_clk_i),
    .d1(gen_filter_4__u_filter_diff_ctr_d[3]),
    .d2(net31),
    .o1(gen_filter_4__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_4__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1209),
    .si2(net1210),
    .ssb(net1797));
 b15fqy203ar1n02x5 gen_filter_4__u_filter_filter_q_reg_gen_filter_7__u_filter_filter_q_reg (.rb(net864),
    .clk(clknet_leaf_5_clk_i),
    .d1(gen_filter_4__u_filter_filter_synced),
    .d2(gen_filter_7__u_filter_filter_synced),
    .o1(gen_filter_4__u_filter_filter_q),
    .o2(gen_filter_7__u_filter_filter_q),
    .si1(net1211),
    .si2(net1212),
    .ssb(net1798));
 b15fqy203ar1n02x5 gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_7__u_filter_diff_ctr_q_reg_0_ (.rb(net864),
    .clk(clknet_leaf_6_clk_i),
    .d1(net2291),
    .d2(gen_filter_7__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_4__u_filter_filter_synced),
    .o2(gen_filter_7__u_filter_diff_ctr_q[0]),
    .si1(net1213),
    .si2(net1214),
    .ssb(net1799));
 b15fqy043ar1n02x5 gen_filter_4__u_filter_stored_value_q_reg (.clk(clknet_leaf_5_clk_i),
    .d(net743),
    .den(eq_x_161_n25),
    .o(gen_filter_4__u_filter_stored_value_q),
    .rb(net862),
    .si(net1215),
    .ssb(net1800));
 b15fqy203ar1n02x5 gen_filter_5__u_filter_diff_ctr_q_reg_0__gen_filter_5__u_filter_diff_ctr_q_reg_1_ (.rb(net856),
    .clk(clknet_leaf_4_clk_i),
    .d1(net2416),
    .d2(net2408),
    .o1(gen_filter_5__u_filter_diff_ctr_q[0]),
    .o2(gen_filter_5__u_filter_diff_ctr_q[1]),
    .si1(net1216),
    .si2(net1217),
    .ssb(net1801));
 b15fqy203ar1n02x5 gen_filter_5__u_filter_diff_ctr_q_reg_2__gen_filter_5__u_filter_diff_ctr_q_reg_3_ (.rb(net856),
    .clk(clknet_leaf_4_clk_i),
    .d1(gen_filter_5__u_filter_diff_ctr_d[2]),
    .d2(gen_filter_5__u_filter_diff_ctr_d[3]),
    .o1(gen_filter_5__u_filter_diff_ctr_q[2]),
    .o2(gen_filter_5__u_filter_diff_ctr_q[3]),
    .si1(net1218),
    .si2(net1219),
    .ssb(net1802));
 b15fqy203ar1n02x5 gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_diff_ctr_q_reg_0_ (.rb(net863),
    .clk(clknet_leaf_5_clk_i),
    .d1(net32),
    .d2(net2401),
    .o1(gen_filter_5__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_6__u_filter_diff_ctr_q[0]),
    .si1(net1220),
    .si2(net1221),
    .ssb(net1803));
 b15fqy203ar1n02x5 gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_filter_q_reg (.rb(net863),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2300),
    .d2(gen_filter_6__u_filter_filter_synced),
    .o1(gen_filter_5__u_filter_filter_synced),
    .o2(gen_filter_6__u_filter_filter_q),
    .si1(net1222),
    .si2(net1223),
    .ssb(net1804));
 b15fqy043ar1n02x5 gen_filter_5__u_filter_stored_value_q_reg (.clk(clknet_leaf_4_clk_i),
    .d(net742),
    .den(eq_x_156_n25),
    .o(gen_filter_5__u_filter_stored_value_q),
    .rb(net859),
    .si(net1224),
    .ssb(net1805));
 b15fqy203ar1n02x5 gen_filter_6__u_filter_diff_ctr_q_reg_1__gen_filter_6__u_filter_diff_ctr_q_reg_2_ (.rb(net863),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2399),
    .d2(net2419),
    .o1(gen_filter_6__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_6__u_filter_diff_ctr_q[2]),
    .si1(net1225),
    .si2(net1226),
    .ssb(net1806));
 b15fqy203ar1n02x5 gen_filter_6__u_filter_diff_ctr_q_reg_3__gen_filter_15__u_filter_diff_ctr_q_reg_0_ (.rb(net864),
    .clk(clknet_leaf_5_clk_i),
    .d1(gen_filter_6__u_filter_diff_ctr_d[3]),
    .d2(gen_filter_15__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_6__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_15__u_filter_diff_ctr_q[0]),
    .si1(net1227),
    .si2(net1228),
    .ssb(net1807));
 b15fqy203ar1n02x5 gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net864),
    .clk(clknet_leaf_5_clk_i),
    .d1(net33),
    .d2(net2259),
    .o1(gen_filter_6__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_6__u_filter_filter_synced),
    .si1(net1229),
    .si2(net1230),
    .ssb(net1808));
 b15fqy043ar1n02x5 gen_filter_6__u_filter_stored_value_q_reg (.clk(clknet_leaf_5_clk_i),
    .d(gen_filter_6__u_filter_filter_synced),
    .den(eq_x_151_n25),
    .o(gen_filter_6__u_filter_stored_value_q),
    .rb(net864),
    .si(net1231),
    .ssb(net1809));
 b15fqy203ar1n02x5 gen_filter_7__u_filter_diff_ctr_q_reg_1__gen_filter_7__u_filter_diff_ctr_q_reg_2_ (.rb(net864),
    .clk(clknet_leaf_5_clk_i),
    .d1(net2538),
    .d2(gen_filter_7__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_7__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_7__u_filter_diff_ctr_q[2]),
    .si1(net1232),
    .si2(net1233),
    .ssb(net1810));
 b15fqy203ar1n02x5 gen_filter_7__u_filter_diff_ctr_q_reg_3__gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net864),
    .clk(clknet_leaf_6_clk_i),
    .d1(gen_filter_7__u_filter_diff_ctr_d[3]),
    .d2(net34),
    .o1(gen_filter_7__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_7__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1234),
    .si2(net1235),
    .ssb(net1811));
 b15fqy203ar1n02x5 gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_9__u_filter_diff_ctr_q_reg_0_ (.rb(net863),
    .clk(clknet_leaf_6_clk_i),
    .d1(net2286),
    .d2(gen_filter_9__u_filter_diff_ctr_d[0]),
    .o1(gen_filter_7__u_filter_filter_synced),
    .o2(gen_filter_9__u_filter_diff_ctr_q[0]),
    .si1(net1236),
    .si2(net1237),
    .ssb(net1812));
 b15fqy043ar1n02x5 gen_filter_7__u_filter_stored_value_q_reg (.clk(clknet_leaf_6_clk_i),
    .d(gen_filter_7__u_filter_filter_synced),
    .den(eq_x_146_n25),
    .o(gen_filter_7__u_filter_stored_value_q),
    .rb(net863),
    .si(net1238),
    .ssb(net1813));
 b15fqy203ar1n02x5 gen_filter_8__u_filter_diff_ctr_q_reg_1__gen_filter_8__u_filter_diff_ctr_q_reg_2_ (.rb(net863),
    .clk(clknet_leaf_6_clk_i),
    .d1(net2494),
    .d2(gen_filter_8__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_8__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_8__u_filter_diff_ctr_q[2]),
    .si1(net1239),
    .si2(net1240),
    .ssb(net1814));
 b15fqy203ar1n02x5 gen_filter_8__u_filter_diff_ctr_q_reg_3__gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net861),
    .clk(clknet_leaf_6_clk_i),
    .d1(gen_filter_8__u_filter_diff_ctr_d[3]),
    .d2(net6),
    .o1(gen_filter_8__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_10__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1241),
    .si2(net1242),
    .ssb(net1815));
 b15fqy203ar1n02x5 gen_filter_8__u_filter_filter_q_reg_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net861),
    .clk(clknet_leaf_6_clk_i),
    .d1(net740),
    .d2(net35),
    .o1(gen_filter_8__u_filter_filter_q),
    .o2(gen_filter_8__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .si1(net1243),
    .si2(net1244),
    .ssb(net1816));
 b15fqy203ar1n02x5 gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_diff_ctr_q_reg_2_ (.rb(net863),
    .clk(clknet_leaf_6_clk_i),
    .d1(net2481),
    .d2(net2382),
    .o1(gen_filter_8__u_filter_filter_synced),
    .o2(gen_filter_11__u_filter_diff_ctr_q[2]),
    .si1(net1245),
    .si2(net1246),
    .ssb(net1817));
 b15fqy043ar1n02x5 gen_filter_8__u_filter_stored_value_q_reg (.clk(clknet_leaf_6_clk_i),
    .d(net2456),
    .den(eq_x_141_n25),
    .o(gen_filter_8__u_filter_stored_value_q),
    .rb(net863),
    .si(net1247),
    .ssb(net1818));
 b15fqy203ar1n02x5 gen_filter_9__u_filter_diff_ctr_q_reg_1__gen_filter_9__u_filter_diff_ctr_q_reg_2_ (.rb(net863),
    .clk(clknet_leaf_6_clk_i),
    .d1(gen_filter_9__u_filter_diff_ctr_d[1]),
    .d2(gen_filter_9__u_filter_diff_ctr_d[2]),
    .o1(gen_filter_9__u_filter_diff_ctr_q[1]),
    .o2(gen_filter_9__u_filter_diff_ctr_q[2]),
    .si1(net1248),
    .si2(net1249),
    .ssb(net1819));
 b15fqy203ar1n02x5 gen_filter_9__u_filter_diff_ctr_q_reg_3__gen_filter_9__u_filter_filter_q_reg (.rb(net863),
    .clk(clknet_leaf_6_clk_i),
    .d1(net2491),
    .d2(gen_filter_9__u_filter_filter_synced),
    .o1(gen_filter_9__u_filter_diff_ctr_q[3]),
    .o2(gen_filter_9__u_filter_filter_q),
    .si1(net1250),
    .si2(net1251),
    .ssb(net1820));
 b15fqy203ar1n02x5 gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0_ (.rb(net861),
    .clk(clknet_leaf_6_clk_i),
    .d1(net36),
    .d2(net2269),
    .o1(gen_filter_9__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .o2(gen_filter_9__u_filter_filter_synced),
    .si1(net1252),
    .si2(net1253),
    .ssb(net1821));
 b15fqy043ar1n02x5 gen_filter_9__u_filter_stored_value_q_reg (.clk(clknet_leaf_6_clk_i),
    .d(gen_filter_9__u_filter_filter_synced),
    .den(eq_x_136_n25),
    .o(gen_filter_9__u_filter_stored_value_q),
    .rb(net861),
    .si(net1254),
    .ssb(net1822));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_10__intr_hw_intr_o_reg_11_ (.rb(net846),
    .clk(clknet_leaf_8_clk_i),
    .d1(intr_hw_N22),
    .d2(intr_hw_N21),
    .o1(net206),
    .o2(net207),
    .si1(net1255),
    .si2(net1256),
    .ssb(net1823));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_12__intr_hw_intr_o_reg_14_ (.rb(net846),
    .clk(clknet_leaf_8_clk_i),
    .d1(intr_hw_N20),
    .d2(intr_hw_N18),
    .o1(net208),
    .o2(net210),
    .si1(net1257),
    .si2(net1258),
    .ssb(net1824));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_15__intr_hw_intr_o_reg_25_ (.rb(net846),
    .clk(clknet_leaf_8_clk_i),
    .d1(intr_hw_N17),
    .d2(intr_hw_N7),
    .o1(net211),
    .o2(net222),
    .si1(net1259),
    .si2(net1260),
    .ssb(net1825));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_16__intr_hw_intr_o_reg_17_ (.rb(net851),
    .clk(clknet_leaf_1_clk_i),
    .d1(intr_hw_N16),
    .d2(intr_hw_N15),
    .o1(net212),
    .o2(net213),
    .si1(net1261),
    .si2(net1262),
    .ssb(net1826));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_18__intr_hw_intr_o_reg_19_ (.rb(net836),
    .clk(clknet_leaf_0_clk_i),
    .d1(intr_hw_N14),
    .d2(intr_hw_N13),
    .o1(net214),
    .o2(net215),
    .si1(net1263),
    .si2(net1264),
    .ssb(net1827));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_1__intr_hw_intr_o_reg_2_ (.rb(net837),
    .clk(clknet_leaf_0_clk_i),
    .d1(intr_hw_N31),
    .d2(intr_hw_N30),
    .o1(net216),
    .o2(net227),
    .si1(net1265),
    .si2(net1266),
    .ssb(net1828));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_20__intr_hw_intr_o_reg_21_ (.rb(net840),
    .clk(clknet_leaf_9_clk_i),
    .d1(intr_hw_N12),
    .d2(intr_hw_N11),
    .o1(net217),
    .o2(net218),
    .si1(net1267),
    .si2(net1268),
    .ssb(net1829));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_22__intr_hw_intr_o_reg_23_ (.rb(net840),
    .clk(clknet_leaf_9_clk_i),
    .d1(intr_hw_N10),
    .d2(intr_hw_N9),
    .o1(net219),
    .o2(net220),
    .si1(net1269),
    .si2(net1270),
    .ssb(net1830));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_24__intr_hw_intr_o_reg_26_ (.rb(net837),
    .clk(clknet_leaf_1_clk_i),
    .d1(intr_hw_N8),
    .d2(intr_hw_N6),
    .o1(net221),
    .o2(net223),
    .si1(net1271),
    .si2(net1272),
    .ssb(net1831));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_27__intr_hw_intr_o_reg_28_ (.rb(net836),
    .clk(clknet_leaf_11_clk_i),
    .d1(intr_hw_N5),
    .d2(intr_hw_N4),
    .o1(net224),
    .o2(net225),
    .si1(net1273),
    .si2(net1274),
    .ssb(net1832));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_29__intr_hw_intr_o_reg_30_ (.rb(net840),
    .clk(clknet_leaf_9_clk_i),
    .d1(intr_hw_N3),
    .d2(intr_hw_N2),
    .o1(net226),
    .o2(net228),
    .si1(net1275),
    .si2(net1276),
    .ssb(net1833));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_31__u_reg_u_data_in_q_reg_1_ (.rb(net853),
    .clk(clknet_leaf_4_clk_i),
    .d1(intr_hw_N1),
    .d2(u_reg_u_data_in_wr_data[1]),
    .o1(net229),
    .o2(u_reg_data_in_qs[1]),
    .si1(net1277),
    .si2(net1278),
    .ssb(net1834));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_3__intr_hw_intr_o_reg_4_ (.rb(net862),
    .clk(clknet_leaf_4_clk_i),
    .d1(intr_hw_N29),
    .d2(intr_hw_N28),
    .o1(net230),
    .o2(net231),
    .si1(net1279),
    .si2(net1280),
    .ssb(net1835));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_5__intr_hw_intr_o_reg_6_ (.rb(net863),
    .clk(clknet_leaf_5_clk_i),
    .d1(intr_hw_N27),
    .d2(intr_hw_N26),
    .o1(net232),
    .o2(net233),
    .si1(net1281),
    .si2(net1282),
    .ssb(net1836));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_7__intr_hw_intr_o_reg_8_ (.rb(net861),
    .clk(clknet_leaf_6_clk_i),
    .d1(intr_hw_N25),
    .d2(intr_hw_N24),
    .o1(net234),
    .o2(net235),
    .si1(net1283),
    .si2(net1284),
    .ssb(net1837));
 b15fqy203ar1n02x5 intr_hw_intr_o_reg_9__intr_hw_intr_o_reg_13_ (.rb(net860),
    .clk(clknet_leaf_6_clk_i),
    .d1(net2483),
    .d2(intr_hw_N19),
    .o1(net236),
    .o2(net209),
    .si1(net1285),
    .si2(net1286),
    .ssb(net1838));
 b15cilb05ah1n02x3 u_reg_u_ctrl_en_input_filter_clk_gate_q_reg_0_latch (.clk(clknet_leaf_1_clk_i),
    .clkout(u_reg_u_ctrl_en_input_filter_net2073),
    .en(n4127),
    .te(net1287));
 b15cilb05ah1n02x3 u_reg_u_ctrl_en_input_filter_clk_gate_q_reg_latch (.clk(clknet_leaf_4_clk_i),
    .clkout(u_reg_u_ctrl_en_input_filter_net2067),
    .en(n4127),
    .te(net1288));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_0__u_reg_u_ctrl_en_input_filter_q_reg_1_ (.rb(net859),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2067),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[0]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[1]),
    .o1(reg2hw_ctrl_en_input_filter__q__0_),
    .o2(reg2hw_ctrl_en_input_filter__q__1_),
    .si1(net1289),
    .si2(net1290),
    .ssb(net1839));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_10__u_reg_u_ctrl_en_input_filter_q_reg_11_ (.rb(net859),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2067),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[10]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[11]),
    .o1(reg2hw_ctrl_en_input_filter__q__10_),
    .o2(reg2hw_ctrl_en_input_filter__q__11_),
    .si1(net1291),
    .si2(net1292),
    .ssb(net1840));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_12__u_reg_u_ctrl_en_input_filter_q_reg_13_ (.rb(net859),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2067),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[12]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[13]),
    .o1(reg2hw_ctrl_en_input_filter__q__12_),
    .o2(reg2hw_ctrl_en_input_filter__q__13_),
    .si1(net1293),
    .si2(net1294),
    .ssb(net1841));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_14__u_reg_u_ctrl_en_input_filter_q_reg_15_ (.rb(net867),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2067),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[14]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[15]),
    .o1(reg2hw_ctrl_en_input_filter__q__14_),
    .o2(reg2hw_ctrl_en_input_filter__q__15_),
    .si1(net1295),
    .si2(net1296),
    .ssb(net1842));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_16__u_reg_u_ctrl_en_input_filter_q_reg_17_ (.rb(net851),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2073),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[16]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[17]),
    .o1(reg2hw_ctrl_en_input_filter__q__16_),
    .o2(reg2hw_ctrl_en_input_filter__q__17_),
    .si1(net1297),
    .si2(net1298),
    .ssb(net1843));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_18__u_reg_u_ctrl_en_input_filter_q_reg_19_ (.rb(net839),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2073),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[18]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[19]),
    .o1(reg2hw_ctrl_en_input_filter__q__18_),
    .o2(reg2hw_ctrl_en_input_filter__q__19_),
    .si1(net1299),
    .si2(net1300),
    .ssb(net1844));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_20__u_reg_u_ctrl_en_input_filter_q_reg_21_ (.rb(net853),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2073),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[20]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[21]),
    .o1(reg2hw_ctrl_en_input_filter__q__20_),
    .o2(reg2hw_ctrl_en_input_filter__q__21_),
    .si1(net1301),
    .si2(net1302),
    .ssb(net1845));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_22__u_reg_u_ctrl_en_input_filter_q_reg_23_ (.rb(net853),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2073),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[22]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[23]),
    .o1(reg2hw_ctrl_en_input_filter__q__22_),
    .o2(reg2hw_ctrl_en_input_filter__q__23_),
    .si1(net1303),
    .si2(net1304),
    .ssb(net1846));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_24__u_reg_u_ctrl_en_input_filter_q_reg_25_ (.rb(net853),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2073),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[24]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[25]),
    .o1(reg2hw_ctrl_en_input_filter__q__24_),
    .o2(reg2hw_ctrl_en_input_filter__q__25_),
    .si1(net1305),
    .si2(net1306),
    .ssb(net1847));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_26__u_reg_u_ctrl_en_input_filter_q_reg_27_ (.rb(net837),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2073),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[26]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[27]),
    .o1(reg2hw_ctrl_en_input_filter__q__26_),
    .o2(reg2hw_ctrl_en_input_filter__q__27_),
    .si1(net1307),
    .si2(net1308),
    .ssb(net1848));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_28__u_reg_u_ctrl_en_input_filter_q_reg_29_ (.rb(net851),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2073),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[28]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[29]),
    .o1(reg2hw_ctrl_en_input_filter__q__28_),
    .o2(reg2hw_ctrl_en_input_filter__q__29_),
    .si1(net1309),
    .si2(net1310),
    .ssb(net1849));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_2__u_reg_u_ctrl_en_input_filter_q_reg_3_ (.rb(net867),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2067),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[2]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[3]),
    .o1(reg2hw_ctrl_en_input_filter__q__2_),
    .o2(reg2hw_ctrl_en_input_filter__q__3_),
    .si1(net1311),
    .si2(net1312),
    .ssb(net1850));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_30__u_reg_u_ctrl_en_input_filter_q_reg_31_ (.rb(net849),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2073),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[30]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[31]),
    .o1(reg2hw_ctrl_en_input_filter__q__30_),
    .o2(reg2hw_ctrl_en_input_filter__q__31_),
    .si1(net1313),
    .si2(net1314),
    .ssb(net1851));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_4__u_reg_u_ctrl_en_input_filter_q_reg_5_ (.rb(net865),
    .clk(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2067),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[4]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[5]),
    .o1(reg2hw_ctrl_en_input_filter__q__4_),
    .o2(reg2hw_ctrl_en_input_filter__q__5_),
    .si1(net1315),
    .si2(net1316),
    .ssb(net1852));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_6__u_reg_u_ctrl_en_input_filter_q_reg_7_ (.rb(net859),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2067),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[6]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[7]),
    .o1(reg2hw_ctrl_en_input_filter__q__6_),
    .o2(reg2hw_ctrl_en_input_filter__q__7_),
    .si1(net1317),
    .si2(net1318),
    .ssb(net1853));
 b15fqy203ar1n02x5 u_reg_u_ctrl_en_input_filter_q_reg_8__u_reg_u_ctrl_en_input_filter_q_reg_9_ (.rb(net866),
    .clk(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2067),
    .d1(u_reg_u_ctrl_en_input_filter_wr_data[8]),
    .d2(u_reg_u_ctrl_en_input_filter_wr_data[9]),
    .o1(reg2hw_ctrl_en_input_filter__q__8_),
    .o2(reg2hw_ctrl_en_input_filter__q__9_),
    .si1(net1319),
    .si2(net1320),
    .ssb(net1854));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_0__u_reg_u_data_in_q_reg_3_ (.rb(net859),
    .clk(clknet_leaf_7_clk_i),
    .d1(u_reg_u_data_in_wr_data[0]),
    .d2(net379),
    .o1(u_reg_data_in_qs[0]),
    .o2(u_reg_data_in_qs[3]),
    .si1(net1321),
    .si2(net1322),
    .ssb(net1855));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_10__u_reg_u_data_in_q_reg_14_ (.rb(net844),
    .clk(clknet_leaf_7_clk_i),
    .d1(u_reg_u_data_in_wr_data[10]),
    .d2(u_reg_u_data_in_wr_data[14]),
    .o1(u_reg_data_in_qs[10]),
    .o2(u_reg_data_in_qs[14]),
    .si1(net1323),
    .si2(net1324),
    .ssb(net1856));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_11__u_reg_u_data_in_q_reg_12_ (.rb(net841),
    .clk(clknet_leaf_9_clk_i),
    .d1(net380),
    .d2(net377),
    .o1(u_reg_data_in_qs[11]),
    .o2(u_reg_data_in_qs[12]),
    .si1(net1325),
    .si2(net1326),
    .ssb(net1857));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_13__u_reg_u_reg_if_rspop_reg_1_ (.rb(net856),
    .clk(clknet_leaf_4_clk_i),
    .d1(u_reg_u_data_in_wr_data[13]),
    .d2(n1429),
    .o1(u_reg_data_in_qs[13]),
    .o2(net292),
    .si1(net1327),
    .si2(net1328),
    .ssb(net1858));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_15__u_reg_u_data_in_q_reg_20_ (.rb(net841),
    .clk(clknet_leaf_9_clk_i),
    .d1(net378),
    .d2(net376),
    .o1(u_reg_data_in_qs[15]),
    .o2(u_reg_data_in_qs[20]),
    .si1(net1329),
    .si2(net1330),
    .ssb(net1859));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_16__u_reg_u_data_in_q_reg_17_ (.rb(net857),
    .clk(clknet_leaf_4_clk_i),
    .d1(u_reg_u_data_in_wr_data[16]),
    .d2(u_reg_u_data_in_wr_data[17]),
    .o1(u_reg_data_in_qs[16]),
    .o2(u_reg_data_in_qs[17]),
    .si1(net1331),
    .si2(net1332),
    .ssb(net1860));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_18__u_reg_u_data_in_q_reg_19_ (.rb(net833),
    .clk(clknet_leaf_11_clk_i),
    .d1(u_reg_u_data_in_wr_data[18]),
    .d2(u_reg_u_data_in_wr_data[19]),
    .o1(u_reg_data_in_qs[18]),
    .o2(u_reg_data_in_qs[19]),
    .si1(net1333),
    .si2(net1334),
    .ssb(net1861));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_21__u_reg_u_data_in_q_reg_22_ (.rb(net840),
    .clk(clknet_leaf_9_clk_i),
    .d1(u_reg_u_data_in_wr_data[21]),
    .d2(net375),
    .o1(u_reg_data_in_qs[21]),
    .o2(u_reg_data_in_qs[22]),
    .si1(net1335),
    .si2(net1336),
    .ssb(net1862));
 b15fqy003ar1n02x5 u_reg_u_data_in_q_reg_23_ (.rb(net840),
    .clk(clknet_leaf_9_clk_i),
    .d(u_reg_u_data_in_wr_data[23]),
    .o(u_reg_data_in_qs[23]),
    .si(net1337),
    .ssb(net1863));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_24__u_reg_u_data_in_q_reg_25_ (.rb(net853),
    .clk(clknet_leaf_4_clk_i),
    .d1(u_reg_u_data_in_wr_data[24]),
    .d2(u_reg_u_data_in_wr_data[25]),
    .o1(u_reg_data_in_qs[24]),
    .o2(u_reg_data_in_qs[25]),
    .si1(net1338),
    .si2(net1339),
    .ssb(net1864));
 b15fqy003ar1n02x5 u_reg_u_data_in_q_reg_26_ (.rb(net849),
    .clk(clknet_leaf_1_clk_i),
    .d(u_reg_u_data_in_wr_data[26]),
    .o(u_reg_data_in_qs[26]),
    .si(net1340),
    .ssb(net1865));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_27__u_reg_u_data_in_q_reg_28_ (.rb(net838),
    .clk(clknet_leaf_1_clk_i),
    .d1(u_reg_u_data_in_wr_data[27]),
    .d2(u_reg_u_data_in_wr_data[28]),
    .o1(u_reg_data_in_qs[27]),
    .o2(u_reg_data_in_qs[28]),
    .si1(net1341),
    .si2(net1342),
    .ssb(net1866));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_29__u_reg_u_data_in_q_reg_30_ (.rb(net839),
    .clk(clknet_leaf_10_clk_i),
    .d1(u_reg_u_data_in_wr_data[29]),
    .d2(u_reg_u_data_in_wr_data[30]),
    .o1(u_reg_data_in_qs[29]),
    .o2(u_reg_data_in_qs[30]),
    .si1(net1343),
    .si2(net1344),
    .ssb(net1867));
 b15fqy003ar1n02x5 u_reg_u_data_in_q_reg_2_ (.rb(net843),
    .clk(clknet_leaf_9_clk_i),
    .d(u_reg_u_data_in_wr_data[2]),
    .o(u_reg_data_in_qs[2]),
    .si(net1345),
    .ssb(net1868));
 b15fqy003ar1n02x5 u_reg_u_data_in_q_reg_31_ (.rb(net839),
    .clk(clknet_leaf_10_clk_i),
    .d(u_reg_u_data_in_wr_data[31]),
    .o(u_reg_data_in_qs[31]),
    .si(net1346),
    .ssb(net1869));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_4__u_reg_u_data_in_q_reg_5_ (.rb(net859),
    .clk(clknet_leaf_7_clk_i),
    .d1(u_reg_u_data_in_wr_data[4]),
    .d2(u_reg_u_data_in_wr_data[5]),
    .o1(u_reg_data_in_qs[4]),
    .o2(u_reg_data_in_qs[5]),
    .si1(net1347),
    .si2(net1348),
    .ssb(net1870));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_6__u_reg_u_data_in_q_reg_7_ (.rb(net860),
    .clk(clknet_leaf_6_clk_i),
    .d1(u_reg_u_data_in_wr_data[6]),
    .d2(u_reg_u_data_in_wr_data[7]),
    .o1(u_reg_data_in_qs[6]),
    .o2(u_reg_data_in_qs[7]),
    .si1(net1349),
    .si2(net1350),
    .ssb(net1871));
 b15fqy203ar1n02x5 u_reg_u_data_in_q_reg_8__u_reg_u_data_in_q_reg_9_ (.rb(net860),
    .clk(clknet_leaf_6_clk_i),
    .d1(u_reg_u_data_in_wr_data[8]),
    .d2(u_reg_u_data_in_wr_data[9]),
    .o1(u_reg_data_in_qs[8]),
    .o2(u_reg_data_in_qs[9]),
    .si1(net1351),
    .si2(net1352),
    .ssb(net1872));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_falling_clk_gate_q_reg_0_latch (.clk(clknet_leaf_1_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_falling_net2073),
    .en(n4128),
    .te(net1353));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_falling_clk_gate_q_reg_latch (.clk(clknet_leaf_8_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_falling_net2067),
    .en(n4128),
    .te(net1354));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_0__u_reg_u_intr_ctrl_en_falling_q_reg_1_ (.rb(net841),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2067),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[0]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[1]),
    .o1(reg2hw_intr_ctrl_en_falling__q__0_),
    .o2(reg2hw_intr_ctrl_en_falling__q__1_),
    .si1(net1355),
    .si2(net1356),
    .ssb(net1873));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_10__u_reg_u_intr_ctrl_en_falling_q_reg_11_ (.rb(net841),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2067),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[10]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[11]),
    .o1(reg2hw_intr_ctrl_en_falling__q__10_),
    .o2(reg2hw_intr_ctrl_en_falling__q__11_),
    .si1(net1357),
    .si2(net1358),
    .ssb(net1874));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_12__u_reg_u_intr_ctrl_en_falling_q_reg_13_ (.rb(net842),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2067),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[12]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[13]),
    .o1(reg2hw_intr_ctrl_en_falling__q__12_),
    .o2(reg2hw_intr_ctrl_en_falling__q__13_),
    .si1(net1359),
    .si2(net1360),
    .ssb(net1875));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_14__u_reg_u_intr_ctrl_en_falling_q_reg_15_ (.rb(net842),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2067),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[14]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[15]),
    .o1(reg2hw_intr_ctrl_en_falling__q__14_),
    .o2(reg2hw_intr_ctrl_en_falling__q__15_),
    .si1(net1361),
    .si2(net1362),
    .ssb(net1876));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_16__u_reg_u_intr_ctrl_en_falling_q_reg_17_ (.rb(net853),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2073),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[16]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[17]),
    .o1(reg2hw_intr_ctrl_en_falling__q__16_),
    .o2(reg2hw_intr_ctrl_en_falling__q__17_),
    .si1(net1363),
    .si2(net1364),
    .ssb(net1877));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_18__u_reg_u_intr_ctrl_en_falling_q_reg_19_ (.rb(net844),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2073),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[18]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[19]),
    .o1(reg2hw_intr_ctrl_en_falling__q__18_),
    .o2(reg2hw_intr_ctrl_en_falling__q__19_),
    .si1(net1365),
    .si2(net1366),
    .ssb(net1878));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_20__u_reg_u_intr_ctrl_en_falling_q_reg_21_ (.rb(net844),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2073),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[20]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[21]),
    .o1(reg2hw_intr_ctrl_en_falling__q__20_),
    .o2(reg2hw_intr_ctrl_en_falling__q__21_),
    .si1(net1367),
    .si2(net1368),
    .ssb(net1879));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_22__u_reg_u_intr_ctrl_en_falling_q_reg_23_ (.rb(net859),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2073),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[22]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[23]),
    .o1(reg2hw_intr_ctrl_en_falling__q__22_),
    .o2(reg2hw_intr_ctrl_en_falling__q__23_),
    .si1(net1369),
    .si2(net1370),
    .ssb(net1880));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_24__u_reg_u_intr_ctrl_en_falling_q_reg_25_ (.rb(net853),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2073),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[24]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[25]),
    .o1(reg2hw_intr_ctrl_en_falling__q__24_),
    .o2(reg2hw_intr_ctrl_en_falling__q__25_),
    .si1(net1371),
    .si2(net1372),
    .ssb(net1881));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_26__u_reg_u_intr_ctrl_en_falling_q_reg_27_ (.rb(net844),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2073),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[26]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[27]),
    .o1(reg2hw_intr_ctrl_en_falling__q__26_),
    .o2(reg2hw_intr_ctrl_en_falling__q__27_),
    .si1(net1373),
    .si2(net1374),
    .ssb(net1882));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_28__u_reg_u_intr_ctrl_en_falling_q_reg_29_ (.rb(net839),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2073),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[28]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[29]),
    .o1(reg2hw_intr_ctrl_en_falling__q__28_),
    .o2(reg2hw_intr_ctrl_en_falling__q__29_),
    .si1(net1375),
    .si2(net1376),
    .ssb(net1883));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_2__u_reg_u_intr_ctrl_en_falling_q_reg_3_ (.rb(net842),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2067),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[2]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[3]),
    .o1(reg2hw_intr_ctrl_en_falling__q__2_),
    .o2(reg2hw_intr_ctrl_en_falling__q__3_),
    .si1(net1377),
    .si2(net1378),
    .ssb(net1884));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_30__u_reg_u_intr_ctrl_en_falling_q_reg_31_ (.rb(net839),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2073),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[30]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[31]),
    .o1(reg2hw_intr_ctrl_en_falling__q__30_),
    .o2(reg2hw_intr_ctrl_en_falling__q__31_),
    .si1(net1379),
    .si2(net1380),
    .ssb(net1885));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_4__u_reg_u_intr_ctrl_en_falling_q_reg_5_ (.rb(net842),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2067),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[4]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[5]),
    .o1(reg2hw_intr_ctrl_en_falling__q__4_),
    .o2(reg2hw_intr_ctrl_en_falling__q__5_),
    .si1(net1381),
    .si2(net1382),
    .ssb(net1886));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_6__u_reg_u_intr_ctrl_en_falling_q_reg_7_ (.rb(net842),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2067),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[6]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[7]),
    .o1(reg2hw_intr_ctrl_en_falling__q__6_),
    .o2(reg2hw_intr_ctrl_en_falling__q__7_),
    .si1(net1383),
    .si2(net1384),
    .ssb(net1887));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_falling_q_reg_8__u_reg_u_intr_ctrl_en_falling_q_reg_9_ (.rb(net842),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2067),
    .d1(u_reg_u_intr_ctrl_en_falling_wr_data[8]),
    .d2(u_reg_u_intr_ctrl_en_falling_wr_data[9]),
    .o1(reg2hw_intr_ctrl_en_falling__q__8_),
    .o2(reg2hw_intr_ctrl_en_falling__q__9_),
    .si1(net1385),
    .si2(net1386),
    .ssb(net1888));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_lvlhigh_clk_gate_q_reg_0_latch (.clk(clknet_leaf_9_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_lvlhigh_net2073),
    .en(n4126),
    .te(net1387));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_lvlhigh_clk_gate_q_reg_latch (.clk(clknet_leaf_9_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_lvlhigh_net2067),
    .en(n4126),
    .te(net1388));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_0__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_1_ (.rb(net840),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[0]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[1]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__0_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__1_),
    .si1(net1389),
    .si2(net1390),
    .ssb(net1889));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_10__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_11_ (.rb(net841),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[10]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[11]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__10_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__11_),
    .si1(net1391),
    .si2(net1392),
    .ssb(net1890));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_12__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_13_ (.rb(net840),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[12]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[13]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__12_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__13_),
    .si1(net1393),
    .si2(net1394),
    .ssb(net1891));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_14__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_15_ (.rb(net840),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[14]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[15]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__14_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__15_),
    .si1(net1395),
    .si2(net1396),
    .ssb(net1892));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_16__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_17_ (.rb(net844),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[16]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[17]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__16_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__17_),
    .si1(net1397),
    .si2(net1398),
    .ssb(net1893));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_18__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_19_ (.rb(net843),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[18]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[19]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__18_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__19_),
    .si1(net1399),
    .si2(net1400),
    .ssb(net1894));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_20__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_21_ (.rb(net843),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[20]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[21]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__20_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__21_),
    .si1(net1401),
    .si2(net1402),
    .ssb(net1895));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_22__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_23_ (.rb(net843),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[22]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[23]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__22_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__23_),
    .si1(net1403),
    .si2(net1404),
    .ssb(net1896));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_24__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_25_ (.rb(net844),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[24]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[25]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__24_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__25_),
    .si1(net1405),
    .si2(net1406),
    .ssb(net1897));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_26__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_27_ (.rb(net844),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[26]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[27]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__26_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__27_),
    .si1(net1407),
    .si2(net1408),
    .ssb(net1898));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_28__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_29_ (.rb(net843),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[28]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[29]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__28_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__29_),
    .si1(net1409),
    .si2(net1410),
    .ssb(net1899));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_2__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_3_ (.rb(net841),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[2]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[3]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__2_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__3_),
    .si1(net1411),
    .si2(net1412),
    .ssb(net1900));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_30__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_31_ (.rb(net844),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[30]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[31]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__30_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__31_),
    .si1(net1413),
    .si2(net1414),
    .ssb(net1901));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_4__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_5_ (.rb(net840),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[4]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[5]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__4_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__5_),
    .si1(net1415),
    .si2(net1416),
    .ssb(net1902));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_6__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_7_ (.rb(net841),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[6]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[7]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__6_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__7_),
    .si1(net1417),
    .si2(net1418),
    .ssb(net1903));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_8__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_9_ (.rb(net841),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[8]),
    .d2(u_reg_u_intr_ctrl_en_lvlhigh_wr_data[9]),
    .o1(reg2hw_intr_ctrl_en_lvlhigh__q__8_),
    .o2(reg2hw_intr_ctrl_en_lvlhigh__q__9_),
    .si1(net1419),
    .si2(net1420),
    .ssb(net1904));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_lvllow_clk_gate_q_reg_0_latch (.clk(clknet_leaf_10_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_lvllow_net2073),
    .en(n4124),
    .te(net1421));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_lvllow_clk_gate_q_reg_latch (.clk(clknet_leaf_8_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_lvllow_net2067),
    .en(n4124),
    .te(net1422));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_0__u_reg_u_intr_ctrl_en_lvllow_q_reg_1_ (.rb(net842),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[0]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[1]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__0_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__1_),
    .si1(net1423),
    .si2(net1424),
    .ssb(net1905));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_10__u_reg_u_intr_ctrl_en_lvllow_q_reg_11_ (.rb(net842),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[10]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[11]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__10_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__11_),
    .si1(net1425),
    .si2(net1426),
    .ssb(net1906));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_12__u_reg_u_intr_ctrl_en_lvllow_q_reg_13_ (.rb(net841),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[12]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[13]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__12_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__13_),
    .si1(net1427),
    .si2(net1428),
    .ssb(net1907));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_14__u_reg_u_intr_ctrl_en_lvllow_q_reg_15_ (.rb(net841),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[14]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[15]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__14_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__15_),
    .si1(net1429),
    .si2(net1430),
    .ssb(net1908));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_16__u_reg_u_intr_ctrl_en_lvllow_q_reg_17_ (.rb(net839),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[16]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[17]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__16_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__17_),
    .si1(net1431),
    .si2(net1432),
    .ssb(net1909));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_18__u_reg_u_intr_ctrl_en_lvllow_q_reg_19_ (.rb(net834),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[18]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[19]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__18_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__19_),
    .si1(net1433),
    .si2(net1434),
    .ssb(net1910));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_20__u_reg_u_intr_ctrl_en_lvllow_q_reg_21_ (.rb(net834),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[20]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[21]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__20_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__21_),
    .si1(net1435),
    .si2(net1436),
    .ssb(net1911));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_22__u_reg_u_intr_ctrl_en_lvllow_q_reg_23_ (.rb(net834),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[22]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[23]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__22_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__23_),
    .si1(net1437),
    .si2(net1438),
    .ssb(net1912));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_24__u_reg_u_intr_ctrl_en_lvllow_q_reg_25_ (.rb(net839),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[24]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[25]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__24_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__25_),
    .si1(net1439),
    .si2(net1440),
    .ssb(net1913));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_26__u_reg_u_intr_ctrl_en_lvllow_q_reg_27_ (.rb(net839),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[26]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[27]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__26_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__27_),
    .si1(net1441),
    .si2(net1442),
    .ssb(net1914));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_28__u_reg_u_intr_ctrl_en_lvllow_q_reg_29_ (.rb(net835),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[28]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[29]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__28_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__29_),
    .si1(net1443),
    .si2(net1444),
    .ssb(net1915));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_2__u_reg_u_intr_ctrl_en_lvllow_q_reg_3_ (.rb(net841),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[2]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[3]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__2_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__3_),
    .si1(net1445),
    .si2(net1446),
    .ssb(net1916));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_30__u_reg_u_intr_ctrl_en_lvllow_q_reg_31_ (.rb(net839),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2073),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[30]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[31]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__30_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__31_),
    .si1(net1447),
    .si2(net1448),
    .ssb(net1917));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_4__u_reg_u_intr_ctrl_en_lvllow_q_reg_5_ (.rb(net842),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[4]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[5]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__4_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__5_),
    .si1(net1449),
    .si2(net1450),
    .ssb(net1918));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_6__u_reg_u_intr_ctrl_en_lvllow_q_reg_7_ (.rb(net842),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[6]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[7]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__6_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__7_),
    .si1(net1451),
    .si2(net1452),
    .ssb(net1919));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_8__u_reg_u_intr_ctrl_en_lvllow_q_reg_9_ (.rb(net842),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2067),
    .d1(u_reg_u_intr_ctrl_en_lvllow_wr_data[8]),
    .d2(u_reg_u_intr_ctrl_en_lvllow_wr_data[9]),
    .o1(reg2hw_intr_ctrl_en_lvllow__q__8_),
    .o2(reg2hw_intr_ctrl_en_lvllow__q__9_),
    .si1(net1453),
    .si2(net1454),
    .ssb(net1920));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_rising_clk_gate_q_reg_0_latch (.clk(clknet_leaf_10_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_rising_net2073),
    .en(n4129),
    .te(net1455));
 b15cilb05ah1n02x3 u_reg_u_intr_ctrl_en_rising_clk_gate_q_reg_latch (.clk(clknet_leaf_7_clk_i),
    .clkout(u_reg_u_intr_ctrl_en_rising_net2067),
    .en(n4129),
    .te(net1456));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_0__u_reg_u_intr_ctrl_en_rising_q_reg_1_ (.rb(net846),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2067),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[0]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[1]),
    .o1(reg2hw_intr_ctrl_en_rising__q__0_),
    .o2(reg2hw_intr_ctrl_en_rising__q__1_),
    .si1(net1457),
    .si2(net1458),
    .ssb(net1921));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_10__u_reg_u_intr_ctrl_en_rising_q_reg_11_ (.rb(net846),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2067),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[10]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[11]),
    .o1(reg2hw_intr_ctrl_en_rising__q__10_),
    .o2(reg2hw_intr_ctrl_en_rising__q__11_),
    .si1(net1459),
    .si2(net1460),
    .ssb(net1922));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_12__u_reg_u_intr_ctrl_en_rising_q_reg_13_ (.rb(net846),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2067),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[12]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[13]),
    .o1(reg2hw_intr_ctrl_en_rising__q__12_),
    .o2(reg2hw_intr_ctrl_en_rising__q__13_),
    .si1(net1461),
    .si2(net1462),
    .ssb(net1923));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_14__u_reg_u_intr_ctrl_en_rising_q_reg_15_ (.rb(net846),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2067),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[14]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[15]),
    .o1(reg2hw_intr_ctrl_en_rising__q__14_),
    .o2(reg2hw_intr_ctrl_en_rising__q__15_),
    .si1(net1463),
    .si2(net1464),
    .ssb(net1924));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_16__u_reg_u_intr_ctrl_en_rising_q_reg_17_ (.rb(net835),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2073),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[16]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[17]),
    .o1(reg2hw_intr_ctrl_en_rising__q__16_),
    .o2(reg2hw_intr_ctrl_en_rising__q__17_),
    .si1(net1465),
    .si2(net1466),
    .ssb(net1925));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_18__u_reg_u_intr_ctrl_en_rising_q_reg_19_ (.rb(net835),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2073),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[18]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[19]),
    .o1(reg2hw_intr_ctrl_en_rising__q__18_),
    .o2(reg2hw_intr_ctrl_en_rising__q__19_),
    .si1(net1467),
    .si2(net1468),
    .ssb(net1926));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_20__u_reg_u_intr_ctrl_en_rising_q_reg_21_ (.rb(net835),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2073),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[20]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[21]),
    .o1(reg2hw_intr_ctrl_en_rising__q__20_),
    .o2(reg2hw_intr_ctrl_en_rising__q__21_),
    .si1(net1469),
    .si2(net1470),
    .ssb(net1927));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_22__u_reg_u_intr_ctrl_en_rising_q_reg_23_ (.rb(net835),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2073),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[22]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[23]),
    .o1(reg2hw_intr_ctrl_en_rising__q__22_),
    .o2(reg2hw_intr_ctrl_en_rising__q__23_),
    .si1(net1471),
    .si2(net1472),
    .ssb(net1928));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_24__u_reg_u_intr_ctrl_en_rising_q_reg_25_ (.rb(net835),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2073),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[24]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[25]),
    .o1(reg2hw_intr_ctrl_en_rising__q__24_),
    .o2(reg2hw_intr_ctrl_en_rising__q__25_),
    .si1(net1473),
    .si2(net1474),
    .ssb(net1929));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_26__u_reg_u_intr_ctrl_en_rising_q_reg_27_ (.rb(net835),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2073),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[26]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[27]),
    .o1(reg2hw_intr_ctrl_en_rising__q__26_),
    .o2(reg2hw_intr_ctrl_en_rising__q__27_),
    .si1(net1475),
    .si2(net1476),
    .ssb(net1930));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_28__u_reg_u_intr_ctrl_en_rising_q_reg_29_ (.rb(net835),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2073),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[28]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[29]),
    .o1(reg2hw_intr_ctrl_en_rising__q__28_),
    .o2(reg2hw_intr_ctrl_en_rising__q__29_),
    .si1(net1477),
    .si2(net1478),
    .ssb(net1931));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_2__u_reg_u_intr_ctrl_en_rising_q_reg_3_ (.rb(net846),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2067),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[2]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[3]),
    .o1(reg2hw_intr_ctrl_en_rising__q__2_),
    .o2(reg2hw_intr_ctrl_en_rising__q__3_),
    .si1(net1479),
    .si2(net1480),
    .ssb(net1932));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_30__u_reg_u_intr_ctrl_en_rising_q_reg_31_ (.rb(net835),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2073),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[30]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[31]),
    .o1(reg2hw_intr_ctrl_en_rising__q__30_),
    .o2(reg2hw_intr_ctrl_en_rising__q__31_),
    .si1(net1481),
    .si2(net1482),
    .ssb(net1933));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_4__u_reg_u_intr_ctrl_en_rising_q_reg_5_ (.rb(net846),
    .clk(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2067),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[4]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[5]),
    .o1(reg2hw_intr_ctrl_en_rising__q__4_),
    .o2(reg2hw_intr_ctrl_en_rising__q__5_),
    .si1(net1483),
    .si2(net1484),
    .ssb(net1934));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_6__u_reg_u_intr_ctrl_en_rising_q_reg_7_ (.rb(net848),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2067),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[6]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[7]),
    .o1(reg2hw_intr_ctrl_en_rising__q__6_),
    .o2(reg2hw_intr_ctrl_en_rising__q__7_),
    .si1(net1485),
    .si2(net1486),
    .ssb(net1935));
 b15fqy203ar1n02x5 u_reg_u_intr_ctrl_en_rising_q_reg_8__u_reg_u_intr_ctrl_en_rising_q_reg_9_ (.rb(net848),
    .clk(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2067),
    .d1(u_reg_u_intr_ctrl_en_rising_wr_data[8]),
    .d2(u_reg_u_intr_ctrl_en_rising_wr_data[9]),
    .o1(reg2hw_intr_ctrl_en_rising__q__8_),
    .o2(reg2hw_intr_ctrl_en_rising__q__9_),
    .si1(net1487),
    .si2(net1488),
    .ssb(net1936));
 b15cilb05ah1n02x3 u_reg_u_intr_enable_clk_gate_q_reg_0_latch (.clk(clknet_leaf_1_clk_i),
    .clkout(u_reg_u_intr_enable_net2073),
    .en(n4125),
    .te(net1489));
 b15cilb05ah1n02x3 u_reg_u_intr_enable_clk_gate_q_reg_latch (.clk(clknet_leaf_7_clk_i),
    .clkout(u_reg_u_intr_enable_net2067),
    .en(n4125),
    .te(net1490));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_0__u_reg_u_intr_enable_q_reg_1_ (.rb(net860),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2067),
    .d1(u_reg_u_intr_enable_wr_data[0]),
    .d2(u_reg_u_intr_enable_wr_data[1]),
    .o1(reg2hw_intr_enable__q__0_),
    .o2(reg2hw_intr_enable__q__1_),
    .si1(net1491),
    .si2(net1492),
    .ssb(net1937));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_10__u_reg_u_intr_enable_q_reg_11_ (.rb(net860),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2067),
    .d1(u_reg_u_intr_enable_wr_data[10]),
    .d2(u_reg_u_intr_enable_wr_data[11]),
    .o1(reg2hw_intr_enable__q__10_),
    .o2(reg2hw_intr_enable__q__11_),
    .si1(net1493),
    .si2(net1494),
    .ssb(net1938));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_12__u_reg_u_intr_enable_q_reg_13_ (.rb(net860),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2067),
    .d1(u_reg_u_intr_enable_wr_data[12]),
    .d2(u_reg_u_intr_enable_wr_data[13]),
    .o1(reg2hw_intr_enable__q__12_),
    .o2(reg2hw_intr_enable__q__13_),
    .si1(net1495),
    .si2(net1496),
    .ssb(net1939));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_14__u_reg_u_intr_enable_q_reg_15_ (.rb(net860),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2067),
    .d1(u_reg_u_intr_enable_wr_data[14]),
    .d2(u_reg_u_intr_enable_wr_data[15]),
    .o1(reg2hw_intr_enable__q__14_),
    .o2(reg2hw_intr_enable__q__15_),
    .si1(net1497),
    .si2(net1498),
    .ssb(net1940));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_16__u_reg_u_intr_enable_q_reg_17_ (.rb(net853),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2073),
    .d1(u_reg_u_intr_enable_wr_data[16]),
    .d2(u_reg_u_intr_enable_wr_data[17]),
    .o1(reg2hw_intr_enable__q__16_),
    .o2(reg2hw_intr_enable__q__17_),
    .si1(net1499),
    .si2(net1500),
    .ssb(net1941));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_18__u_reg_u_intr_enable_q_reg_19_ (.rb(net839),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2073),
    .d1(u_reg_u_intr_enable_wr_data[18]),
    .d2(u_reg_u_intr_enable_wr_data[19]),
    .o1(reg2hw_intr_enable__q__18_),
    .o2(reg2hw_intr_enable__q__19_),
    .si1(net1501),
    .si2(net1502),
    .ssb(net1942));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_20__u_reg_u_intr_enable_q_reg_21_ (.rb(net839),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2073),
    .d1(u_reg_u_intr_enable_wr_data[20]),
    .d2(u_reg_u_intr_enable_wr_data[21]),
    .o1(reg2hw_intr_enable__q__20_),
    .o2(reg2hw_intr_enable__q__21_),
    .si1(net1503),
    .si2(net1504),
    .ssb(net1943));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_22__u_reg_u_intr_enable_q_reg_23_ (.rb(net839),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2073),
    .d1(u_reg_u_intr_enable_wr_data[22]),
    .d2(u_reg_u_intr_enable_wr_data[23]),
    .o1(reg2hw_intr_enable__q__22_),
    .o2(reg2hw_intr_enable__q__23_),
    .si1(net1505),
    .si2(net1506),
    .ssb(net1944));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_24__u_reg_u_intr_enable_q_reg_25_ (.rb(net853),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2073),
    .d1(u_reg_u_intr_enable_wr_data[24]),
    .d2(u_reg_u_intr_enable_wr_data[25]),
    .o1(reg2hw_intr_enable__q__24_),
    .o2(reg2hw_intr_enable__q__25_),
    .si1(net1507),
    .si2(net1508),
    .ssb(net1945));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_26__u_reg_u_intr_enable_q_reg_27_ (.rb(net839),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2073),
    .d1(u_reg_u_intr_enable_wr_data[26]),
    .d2(u_reg_u_intr_enable_wr_data[27]),
    .o1(reg2hw_intr_enable__q__26_),
    .o2(reg2hw_intr_enable__q__27_),
    .si1(net1509),
    .si2(net1510),
    .ssb(net1946));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_28__u_reg_u_intr_enable_q_reg_29_ (.rb(net849),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2073),
    .d1(u_reg_u_intr_enable_wr_data[28]),
    .d2(u_reg_u_intr_enable_wr_data[29]),
    .o1(reg2hw_intr_enable__q__28_),
    .o2(reg2hw_intr_enable__q__29_),
    .si1(net1511),
    .si2(net1512),
    .ssb(net1947));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_2__u_reg_u_intr_enable_q_reg_3_ (.rb(net860),
    .clk(clknet_1_0__leaf_u_reg_u_intr_enable_net2067),
    .d1(u_reg_u_intr_enable_wr_data[2]),
    .d2(u_reg_u_intr_enable_wr_data[3]),
    .o1(reg2hw_intr_enable__q__2_),
    .o2(reg2hw_intr_enable__q__3_),
    .si1(net1513),
    .si2(net1514),
    .ssb(net1948));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_30__u_reg_u_intr_enable_q_reg_31_ (.rb(net849),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2073),
    .d1(u_reg_u_intr_enable_wr_data[30]),
    .d2(u_reg_u_intr_enable_wr_data[31]),
    .o1(reg2hw_intr_enable__q__30_),
    .o2(reg2hw_intr_enable__q__31_),
    .si1(net1515),
    .si2(net1516),
    .ssb(net1949));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_4__u_reg_u_intr_enable_q_reg_5_ (.rb(net860),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2067),
    .d1(u_reg_u_intr_enable_wr_data[4]),
    .d2(u_reg_u_intr_enable_wr_data[5]),
    .o1(reg2hw_intr_enable__q__4_),
    .o2(reg2hw_intr_enable__q__5_),
    .si1(net1517),
    .si2(net1518),
    .ssb(net1950));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_6__u_reg_u_intr_enable_q_reg_7_ (.rb(net860),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2067),
    .d1(u_reg_u_intr_enable_wr_data[6]),
    .d2(u_reg_u_intr_enable_wr_data[7]),
    .o1(reg2hw_intr_enable__q__6_),
    .o2(reg2hw_intr_enable__q__7_),
    .si1(net1519),
    .si2(net1520),
    .ssb(net1951));
 b15fqy203ar1n02x5 u_reg_u_intr_enable_q_reg_8__u_reg_u_intr_enable_q_reg_9_ (.rb(net860),
    .clk(clknet_1_1__leaf_u_reg_u_intr_enable_net2067),
    .d1(u_reg_u_intr_enable_wr_data[8]),
    .d2(u_reg_u_intr_enable_wr_data[9]),
    .o1(reg2hw_intr_enable__q__8_),
    .o2(reg2hw_intr_enable__q__9_),
    .si1(net1521),
    .si2(net1522),
    .ssb(net1952));
 b15cilb05ah1n02x3 u_reg_u_intr_state_clk_gate_q_reg_0_latch (.clk(clknet_leaf_10_clk_i),
    .clkout(u_reg_u_intr_state_net2096),
    .en(u_reg_u_intr_state_n1),
    .te(net1523));
 b15cilb05ah1n02x3 u_reg_u_intr_state_clk_gate_q_reg_latch (.clk(clknet_leaf_7_clk_i),
    .clkout(u_reg_u_intr_state_net2090),
    .en(u_reg_u_intr_state_n1),
    .te(net1524));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_0__u_reg_u_intr_state_q_reg_1_ (.rb(net844),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2090),
    .d1(u_reg_u_intr_state_wr_data[0]),
    .d2(u_reg_u_intr_state_wr_data[1]),
    .o1(reg2hw_intr_state__q__0_),
    .o2(reg2hw_intr_state__q__1_),
    .si1(net1525),
    .si2(net1526),
    .ssb(net1953));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_10__u_reg_u_intr_state_q_reg_11_ (.rb(net844),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2090),
    .d1(u_reg_u_intr_state_wr_data[10]),
    .d2(u_reg_u_intr_state_wr_data[11]),
    .o1(reg2hw_intr_state__q__10_),
    .o2(reg2hw_intr_state__q__11_),
    .si1(net1527),
    .si2(net1528),
    .ssb(net1954));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_12__u_reg_u_intr_state_q_reg_13_ (.rb(net845),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2090),
    .d1(u_reg_u_intr_state_wr_data[12]),
    .d2(u_reg_u_intr_state_wr_data[13]),
    .o1(reg2hw_intr_state__q__12_),
    .o2(reg2hw_intr_state__q__13_),
    .si1(net1529),
    .si2(net1530),
    .ssb(net1955));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_14__u_reg_u_intr_state_q_reg_15_ (.rb(net845),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2090),
    .d1(u_reg_u_intr_state_wr_data[14]),
    .d2(u_reg_u_intr_state_wr_data[15]),
    .o1(reg2hw_intr_state__q__14_),
    .o2(reg2hw_intr_state__q__15_),
    .si1(net1531),
    .si2(net1532),
    .ssb(net1956));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_16__u_reg_u_intr_state_q_reg_17_ (.rb(net845),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2096),
    .d1(u_reg_u_intr_state_wr_data[16]),
    .d2(u_reg_u_intr_state_wr_data[17]),
    .o1(reg2hw_intr_state__q__16_),
    .o2(reg2hw_intr_state__q__17_),
    .si1(net1533),
    .si2(net1534),
    .ssb(net1957));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_18__u_reg_u_intr_state_q_reg_19_ (.rb(net844),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2096),
    .d1(u_reg_u_intr_state_wr_data[18]),
    .d2(u_reg_u_intr_state_wr_data[19]),
    .o1(reg2hw_intr_state__q__18_),
    .o2(reg2hw_intr_state__q__19_),
    .si1(net1535),
    .si2(net1536),
    .ssb(net1958));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_20__u_reg_u_intr_state_q_reg_21_ (.rb(net844),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2096),
    .d1(u_reg_u_intr_state_wr_data[20]),
    .d2(u_reg_u_intr_state_wr_data[21]),
    .o1(reg2hw_intr_state__q__20_),
    .o2(reg2hw_intr_state__q__21_),
    .si1(net1537),
    .si2(net1538),
    .ssb(net1959));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_22__u_reg_u_intr_state_q_reg_23_ (.rb(net844),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2096),
    .d1(u_reg_u_intr_state_wr_data[22]),
    .d2(u_reg_u_intr_state_wr_data[23]),
    .o1(reg2hw_intr_state__q__22_),
    .o2(reg2hw_intr_state__q__23_),
    .si1(net1539),
    .si2(net1540),
    .ssb(net1960));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_24__u_reg_u_intr_state_q_reg_25_ (.rb(net845),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2096),
    .d1(u_reg_u_intr_state_wr_data[24]),
    .d2(net2496),
    .o1(reg2hw_intr_state__q__24_),
    .o2(reg2hw_intr_state__q__25_),
    .si1(net1541),
    .si2(net1542),
    .ssb(net1961));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_26__u_reg_u_intr_state_q_reg_27_ (.rb(net845),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2096),
    .d1(u_reg_u_intr_state_wr_data[26]),
    .d2(u_reg_u_intr_state_wr_data[27]),
    .o1(reg2hw_intr_state__q__26_),
    .o2(reg2hw_intr_state__q__27_),
    .si1(net1543),
    .si2(net1544),
    .ssb(net1962));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_28__u_reg_u_intr_state_q_reg_29_ (.rb(net844),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2096),
    .d1(u_reg_u_intr_state_wr_data[28]),
    .d2(net2338),
    .o1(reg2hw_intr_state__q__28_),
    .o2(reg2hw_intr_state__q__29_),
    .si1(net1545),
    .si2(net1546),
    .ssb(net1963));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_2__u_reg_u_intr_state_q_reg_3_ (.rb(net845),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2090),
    .d1(u_reg_u_intr_state_wr_data[2]),
    .d2(u_reg_u_intr_state_wr_data[3]),
    .o1(reg2hw_intr_state__q__2_),
    .o2(reg2hw_intr_state__q__3_),
    .si1(net1547),
    .si2(net1548),
    .ssb(net1964));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_30__u_reg_u_intr_state_q_reg_31_ (.rb(net845),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2096),
    .d1(u_reg_u_intr_state_wr_data[30]),
    .d2(u_reg_u_intr_state_wr_data[31]),
    .o1(reg2hw_intr_state__q__30_),
    .o2(reg2hw_intr_state__q__31_),
    .si1(net1549),
    .si2(net1550),
    .ssb(net1965));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_4__u_reg_u_intr_state_q_reg_5_ (.rb(net845),
    .clk(clknet_1_0__leaf_u_reg_u_intr_state_net2090),
    .d1(u_reg_u_intr_state_wr_data[4]),
    .d2(u_reg_u_intr_state_wr_data[5]),
    .o1(reg2hw_intr_state__q__4_),
    .o2(reg2hw_intr_state__q__5_),
    .si1(net1551),
    .si2(net1552),
    .ssb(net1966));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_6__u_reg_u_intr_state_q_reg_7_ (.rb(net845),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2090),
    .d1(u_reg_u_intr_state_wr_data[6]),
    .d2(u_reg_u_intr_state_wr_data[7]),
    .o1(reg2hw_intr_state__q__6_),
    .o2(reg2hw_intr_state__q__7_),
    .si1(net1553),
    .si2(net1554),
    .ssb(net1967));
 b15fqy203ar1n02x5 u_reg_u_intr_state_q_reg_8__u_reg_u_intr_state_q_reg_9_ (.rb(net845),
    .clk(clknet_1_1__leaf_u_reg_u_intr_state_net2090),
    .d1(u_reg_u_intr_state_wr_data[8]),
    .d2(u_reg_u_intr_state_wr_data[9]),
    .o1(reg2hw_intr_state__q__8_),
    .o2(reg2hw_intr_state__q__9_),
    .si1(net1555),
    .si2(net1556),
    .ssb(net1968));
 b15cilb05ah1n02x3 u_reg_u_reg_if_clk_gate_rdata_reg_0_latch (.clk(clknet_leaf_1_clk_i),
    .clkout(u_reg_u_reg_if_net2124),
    .en(net408),
    .te(net1557));
 b15cilb05ah1n02x3 u_reg_u_reg_if_clk_gate_rdata_reg_latch (.clk(clknet_leaf_11_clk_i),
    .clkout(u_reg_u_reg_if_net2119),
    .en(net408),
    .te(net1558));
 b15cilb05ah1n02x3 u_reg_u_reg_if_clk_gate_reqid_reg_latch (.clk(clknet_leaf_5_clk_i),
    .clkout(u_reg_u_reg_if_net2113),
    .en(net409),
    .te(net1559));
 b15fqy043ar1n02x5 u_reg_u_reg_if_error_reg (.clk(clknet_leaf_3_clk_i),
    .d(u_reg_u_reg_if_N46),
    .den(u_reg_u_reg_if_a_ack),
    .o(net248),
    .rb(net856),
    .si(net1560),
    .ssb(net1969));
 b15fqy043ar1n02x5 u_reg_u_reg_if_outstanding_reg (.clk(clknet_leaf_3_clk_i),
    .d(u_reg_u_reg_if_a_ack),
    .den(u_reg_u_reg_if_N7),
    .o(net294),
    .rb(net858),
    .si(net1561),
    .ssb(net1970));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_0__u_reg_u_reg_if_rdata_reg_1_ (.rb(net834),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2119),
    .d1(u_reg_u_reg_if_N14),
    .d2(u_reg_u_reg_if_N15),
    .o1(net244),
    .o2(net245),
    .si1(net1562),
    .si2(net1563),
    .ssb(net1971));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_10__u_reg_u_reg_if_rdata_reg_11_ (.rb(net834),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2119),
    .d1(u_reg_u_reg_if_N24),
    .d2(net2341),
    .o1(net255),
    .o2(net256),
    .si1(net1564),
    .si2(net1565),
    .ssb(net1972));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_12__u_reg_u_reg_if_rdata_reg_13_ (.rb(net834),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2119),
    .d1(u_reg_u_reg_if_N26),
    .d2(u_reg_u_reg_if_N27),
    .o1(net257),
    .o2(net258),
    .si1(net1566),
    .si2(net1567),
    .ssb(net1973));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_14__u_reg_u_reg_if_rdata_reg_15_ (.rb(net834),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2119),
    .d1(net2423),
    .d2(u_reg_u_reg_if_N29),
    .o1(net260),
    .o2(net261),
    .si1(net1568),
    .si2(net1569),
    .ssb(net1974));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_16__u_reg_u_reg_if_rdata_reg_17_ (.rb(net837),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2124),
    .d1(net2242),
    .d2(net2281),
    .o1(net262),
    .o2(net263),
    .si1(net1570),
    .si2(net1571),
    .ssb(net1975));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_18__u_reg_u_reg_if_rdata_reg_19_ (.rb(net834),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2124),
    .d1(net2239),
    .d2(net2296),
    .o1(net264),
    .o2(net265),
    .si1(net1572),
    .si2(net1573),
    .ssb(net1976));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_20__u_reg_u_reg_if_rdata_reg_21_ (.rb(net834),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2124),
    .d1(u_reg_u_reg_if_N34),
    .d2(net2322),
    .o1(net266),
    .o2(net267),
    .si1(net1574),
    .si2(net1575),
    .ssb(net1977));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_22__u_reg_u_reg_if_rdata_reg_23_ (.rb(net834),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2124),
    .d1(net2289),
    .d2(net2284),
    .o1(net268),
    .o2(net269),
    .si1(net1576),
    .si2(net1577),
    .ssb(net1978));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_24__u_reg_u_reg_if_rdata_reg_25_ (.rb(net837),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2124),
    .d1(net2403),
    .d2(net2190),
    .o1(net271),
    .o2(net272),
    .si1(net1578),
    .si2(net1579),
    .ssb(net1979));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_26__u_reg_u_reg_if_rdata_reg_27_ (.rb(net837),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2124),
    .d1(net2213),
    .d2(net2343),
    .o1(net273),
    .o2(net274),
    .si1(net1580),
    .si2(net1581),
    .ssb(net1980));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_28__u_reg_u_reg_if_rdata_reg_29_ (.rb(net834),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2124),
    .d1(net2246),
    .d2(net2161),
    .o1(net275),
    .o2(net276),
    .si1(net1582),
    .si2(net1583),
    .ssb(net1981));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_2__u_reg_u_reg_if_rdata_reg_3_ (.rb(net834),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2119),
    .d1(net2307),
    .d2(u_reg_u_reg_if_N17),
    .o1(net246),
    .o2(net247),
    .si1(net1584),
    .si2(net1585),
    .ssb(net1982));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_30__u_reg_u_reg_if_rdata_reg_31_ (.rb(net837),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2124),
    .d1(net2371),
    .d2(net2195),
    .o1(net277),
    .o2(net278),
    .si1(net1586),
    .si2(net1587),
    .ssb(net1983));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_4__u_reg_u_reg_if_rdata_reg_5_ (.rb(net834),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2119),
    .d1(u_reg_u_reg_if_N18),
    .d2(u_reg_u_reg_if_N19),
    .o1(net249),
    .o2(net250),
    .si1(net1588),
    .si2(net1589),
    .ssb(net1984));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_6__u_reg_u_reg_if_rdata_reg_7_ (.rb(net834),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2119),
    .d1(net318),
    .d2(net317),
    .o1(net251),
    .o2(net252),
    .si1(net1590),
    .si2(net1591),
    .ssb(net1985));
 b15fqy203ar1n02x5 u_reg_u_reg_if_rdata_reg_8__u_reg_u_reg_if_rdata_reg_9_ (.rb(net834),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2119),
    .d1(net316),
    .d2(net315),
    .o1(net253),
    .o2(net254),
    .si1(net1592),
    .si2(net1593),
    .ssb(net1986));
 b15fqy203ar1n02x5 u_reg_u_reg_if_reqid_reg_0__u_reg_u_reg_if_reqid_reg_1_ (.rb(net862),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2113),
    .d1(net130),
    .d2(net131),
    .o1(net279),
    .o2(net281),
    .si1(net1594),
    .si2(net1595),
    .ssb(net1987));
 b15fqy203ar1n02x5 u_reg_u_reg_if_reqid_reg_2__u_reg_u_reg_if_reqid_reg_3_ (.rb(net866),
    .clk(clknet_1_0__leaf_u_reg_u_reg_if_net2113),
    .d1(net132),
    .d2(net133),
    .o1(net282),
    .o2(net283),
    .si1(net1596),
    .si2(net1597),
    .ssb(net1988));
 b15fqy203ar1n02x5 u_reg_u_reg_if_reqid_reg_4__u_reg_u_reg_if_reqid_reg_5_ (.rb(net866),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2113),
    .d1(net134),
    .d2(net135),
    .o1(net284),
    .o2(net285),
    .si1(net1598),
    .si2(net1599),
    .ssb(net1989));
 b15fqy203ar1n02x5 u_reg_u_reg_if_reqid_reg_6__u_reg_u_reg_if_reqid_reg_7_ (.rb(net866),
    .clk(clknet_1_1__leaf_u_reg_u_reg_if_net2113),
    .d1(net136),
    .d2(net137),
    .o1(net286),
    .o2(net287),
    .si1(net1600),
    .si2(net1601),
    .ssb(net1990));
 b15fqy043ar1n02x5 u_reg_u_reg_if_reqsz_reg_0_ (.clk(clknet_leaf_3_clk_i),
    .d(net39),
    .den(u_reg_u_reg_if_a_ack),
    .o(net288),
    .rb(net858),
    .si(net1602),
    .ssb(net1991));
 b15fqy043ar1n02x5 u_reg_u_reg_if_reqsz_reg_1_ (.clk(clknet_leaf_3_clk_i),
    .d(net40),
    .den(u_reg_u_reg_if_a_ack),
    .o(net289),
    .rb(net858),
    .si(net1603),
    .ssb(net1992));
 b15fqy043ar1n02x5 u_reg_u_reg_if_rspop_reg_0_ (.clk(clknet_leaf_5_clk_i),
    .d(u_reg_u_reg_if_rd_req),
    .den(net409),
    .o(net291),
    .rb(net867),
    .si(net1604),
    .ssb(net1993));
 b15fqy003ar1n02x5 u_reg_u_reg_if_rspop_reg_2_ (.rb(net858),
    .clk(clknet_leaf_3_clk_i),
    .d(n1432),
    .o(net293),
    .si(net1605),
    .ssb(net1994));
 b15tihi00an1n03x5 U3325_1606 (.o(net1606));
 b15cbf000an1n16x5 clkbuf_leaf_0_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_0_clk_i));
 b15ztpn00an1n08x5 PHY_98 ();
 b15ztpn00an1n08x5 PHY_99 ();
 b15ztpn00an1n08x5 PHY_100 ();
 b15ztpn00an1n08x5 PHY_101 ();
 b15ztpn00an1n08x5 PHY_102 ();
 b15ztpn00an1n08x5 PHY_103 ();
 b15ztpn00an1n08x5 PHY_104 ();
 b15ztpn00an1n08x5 PHY_105 ();
 b15ztpn00an1n08x5 PHY_106 ();
 b15ztpn00an1n08x5 PHY_107 ();
 b15ztpn00an1n08x5 PHY_108 ();
 b15ztpn00an1n08x5 PHY_109 ();
 b15ztpn00an1n08x5 PHY_110 ();
 b15ztpn00an1n08x5 PHY_111 ();
 b15ztpn00an1n08x5 PHY_112 ();
 b15ztpn00an1n08x5 PHY_113 ();
 b15ztpn00an1n08x5 PHY_114 ();
 b15ztpn00an1n08x5 PHY_115 ();
 b15ztpn00an1n08x5 PHY_116 ();
 b15ztpn00an1n08x5 PHY_117 ();
 b15ztpn00an1n08x5 PHY_118 ();
 b15ztpn00an1n08x5 PHY_119 ();
 b15ztpn00an1n08x5 PHY_120 ();
 b15ztpn00an1n08x5 PHY_121 ();
 b15ztpn00an1n08x5 PHY_122 ();
 b15ztpn00an1n08x5 PHY_123 ();
 b15ztpn00an1n08x5 PHY_124 ();
 b15ztpn00an1n08x5 PHY_125 ();
 b15ztpn00an1n08x5 PHY_126 ();
 b15ztpn00an1n08x5 PHY_127 ();
 b15ztpn00an1n08x5 PHY_128 ();
 b15ztpn00an1n08x5 PHY_129 ();
 b15ztpn00an1n08x5 PHY_130 ();
 b15ztpn00an1n08x5 PHY_131 ();
 b15ztpn00an1n08x5 PHY_132 ();
 b15ztpn00an1n08x5 PHY_133 ();
 b15ztpn00an1n08x5 PHY_134 ();
 b15ztpn00an1n08x5 PHY_135 ();
 b15ztpn00an1n08x5 PHY_136 ();
 b15ztpn00an1n08x5 PHY_137 ();
 b15ztpn00an1n08x5 PHY_138 ();
 b15ztpn00an1n08x5 PHY_139 ();
 b15ztpn00an1n08x5 PHY_140 ();
 b15ztpn00an1n08x5 PHY_141 ();
 b15ztpn00an1n08x5 PHY_142 ();
 b15ztpn00an1n08x5 PHY_143 ();
 b15ztpn00an1n08x5 PHY_144 ();
 b15ztpn00an1n08x5 PHY_145 ();
 b15ztpn00an1n08x5 PHY_146 ();
 b15ztpn00an1n08x5 PHY_147 ();
 b15ztpn00an1n08x5 PHY_148 ();
 b15ztpn00an1n08x5 PHY_149 ();
 b15ztpn00an1n08x5 PHY_150 ();
 b15ztpn00an1n08x5 PHY_151 ();
 b15ztpn00an1n08x5 PHY_152 ();
 b15ztpn00an1n08x5 PHY_153 ();
 b15ztpn00an1n08x5 PHY_154 ();
 b15ztpn00an1n08x5 PHY_155 ();
 b15ztpn00an1n08x5 PHY_156 ();
 b15ztpn00an1n08x5 PHY_157 ();
 b15ztpn00an1n08x5 PHY_158 ();
 b15ztpn00an1n08x5 PHY_159 ();
 b15ztpn00an1n08x5 PHY_160 ();
 b15ztpn00an1n08x5 PHY_161 ();
 b15ztpn00an1n08x5 PHY_162 ();
 b15ztpn00an1n08x5 PHY_163 ();
 b15ztpn00an1n08x5 PHY_164 ();
 b15ztpn00an1n08x5 PHY_165 ();
 b15ztpn00an1n08x5 PHY_166 ();
 b15ztpn00an1n08x5 PHY_167 ();
 b15ztpn00an1n08x5 PHY_168 ();
 b15ztpn00an1n08x5 PHY_169 ();
 b15ztpn00an1n08x5 PHY_170 ();
 b15ztpn00an1n08x5 PHY_171 ();
 b15ztpn00an1n08x5 PHY_172 ();
 b15ztpn00an1n08x5 PHY_173 ();
 b15ztpn00an1n08x5 PHY_174 ();
 b15ztpn00an1n08x5 PHY_175 ();
 b15ztpn00an1n08x5 PHY_176 ();
 b15ztpn00an1n08x5 PHY_177 ();
 b15ztpn00an1n08x5 PHY_178 ();
 b15ztpn00an1n08x5 PHY_179 ();
 b15ztpn00an1n08x5 PHY_180 ();
 b15ztpn00an1n08x5 PHY_181 ();
 b15ztpn00an1n08x5 PHY_182 ();
 b15ztpn00an1n08x5 PHY_183 ();
 b15ztpn00an1n08x5 PHY_184 ();
 b15ztpn00an1n08x5 PHY_185 ();
 b15ztpn00an1n08x5 PHY_186 ();
 b15ztpn00an1n08x5 PHY_187 ();
 b15ztpn00an1n08x5 PHY_188 ();
 b15ztpn00an1n08x5 PHY_189 ();
 b15ztpn00an1n08x5 PHY_190 ();
 b15ztpn00an1n08x5 PHY_191 ();
 b15ztpn00an1n08x5 PHY_192 ();
 b15ztpn00an1n08x5 PHY_193 ();
 b15ztpn00an1n08x5 PHY_194 ();
 b15ztpn00an1n08x5 PHY_195 ();
 b15ztpn00an1n08x5 PHY_196 ();
 b15ztpn00an1n08x5 PHY_197 ();
 b15ztpn00an1n08x5 PHY_198 ();
 b15ztpn00an1n08x5 PHY_199 ();
 b15ztpn00an1n08x5 PHY_200 ();
 b15ztpn00an1n08x5 PHY_201 ();
 b15ztpn00an1n08x5 PHY_202 ();
 b15ztpn00an1n08x5 PHY_203 ();
 b15ztpn00an1n08x5 PHY_204 ();
 b15ztpn00an1n08x5 PHY_205 ();
 b15ztpn00an1n08x5 PHY_206 ();
 b15ztpn00an1n08x5 PHY_207 ();
 b15ztpn00an1n08x5 PHY_208 ();
 b15ztpn00an1n08x5 PHY_209 ();
 b15ztpn00an1n08x5 PHY_210 ();
 b15ztpn00an1n08x5 PHY_211 ();
 b15ztpn00an1n08x5 PHY_212 ();
 b15ztpn00an1n08x5 PHY_213 ();
 b15ztpn00an1n08x5 PHY_214 ();
 b15ztpn00an1n08x5 PHY_215 ();
 b15ztpn00an1n08x5 PHY_216 ();
 b15ztpn00an1n08x5 PHY_217 ();
 b15ztpn00an1n08x5 PHY_218 ();
 b15ztpn00an1n08x5 PHY_219 ();
 b15ztpn00an1n08x5 PHY_220 ();
 b15ztpn00an1n08x5 PHY_221 ();
 b15ztpn00an1n08x5 PHY_222 ();
 b15ztpn00an1n08x5 PHY_223 ();
 b15ztpn00an1n08x5 PHY_224 ();
 b15ztpn00an1n08x5 PHY_225 ();
 b15ztpn00an1n08x5 PHY_226 ();
 b15ztpn00an1n08x5 PHY_227 ();
 b15ztpn00an1n08x5 PHY_228 ();
 b15ztpn00an1n08x5 PHY_229 ();
 b15ztpn00an1n08x5 PHY_230 ();
 b15ztpn00an1n08x5 PHY_231 ();
 b15ztpn00an1n08x5 PHY_232 ();
 b15ztpn00an1n08x5 PHY_233 ();
 b15ztpn00an1n08x5 PHY_234 ();
 b15ztpn00an1n08x5 PHY_235 ();
 b15ztpn00an1n08x5 PHY_236 ();
 b15ztpn00an1n08x5 PHY_237 ();
 b15ztpn00an1n08x5 PHY_238 ();
 b15ztpn00an1n08x5 PHY_239 ();
 b15ztpn00an1n08x5 PHY_240 ();
 b15ztpn00an1n08x5 PHY_241 ();
 b15ztpn00an1n08x5 PHY_242 ();
 b15ztpn00an1n08x5 PHY_243 ();
 b15ztpn00an1n08x5 PHY_244 ();
 b15ztpn00an1n08x5 PHY_245 ();
 b15ztpn00an1n08x5 PHY_246 ();
 b15ztpn00an1n08x5 PHY_247 ();
 b15ztpn00an1n08x5 PHY_248 ();
 b15ztpn00an1n08x5 PHY_249 ();
 b15ztpn00an1n08x5 PHY_250 ();
 b15ztpn00an1n08x5 PHY_251 ();
 b15ztpn00an1n08x5 PHY_252 ();
 b15ztpn00an1n08x5 PHY_253 ();
 b15ztpn00an1n08x5 PHY_254 ();
 b15ztpn00an1n08x5 PHY_255 ();
 b15ztpn00an1n08x5 PHY_256 ();
 b15ztpn00an1n08x5 PHY_257 ();
 b15ztpn00an1n08x5 PHY_258 ();
 b15ztpn00an1n08x5 PHY_259 ();
 b15ztpn00an1n08x5 PHY_260 ();
 b15ztpn00an1n08x5 PHY_261 ();
 b15ztpn00an1n08x5 PHY_262 ();
 b15ztpn00an1n08x5 PHY_263 ();
 b15ztpn00an1n08x5 PHY_264 ();
 b15ztpn00an1n08x5 PHY_265 ();
 b15ztpn00an1n08x5 PHY_266 ();
 b15ztpn00an1n08x5 PHY_267 ();
 b15ztpn00an1n08x5 PHY_268 ();
 b15ztpn00an1n08x5 PHY_269 ();
 b15ztpn00an1n08x5 PHY_270 ();
 b15ztpn00an1n08x5 PHY_271 ();
 b15ztpn00an1n08x5 PHY_272 ();
 b15ztpn00an1n08x5 PHY_273 ();
 b15ztpn00an1n08x5 PHY_274 ();
 b15ztpn00an1n08x5 PHY_275 ();
 b15ztpn00an1n08x5 PHY_276 ();
 b15ztpn00an1n08x5 PHY_277 ();
 b15ztpn00an1n08x5 PHY_278 ();
 b15ztpn00an1n08x5 PHY_279 ();
 b15ztpn00an1n08x5 PHY_280 ();
 b15ztpn00an1n08x5 PHY_281 ();
 b15ztpn00an1n08x5 PHY_282 ();
 b15ztpn00an1n08x5 PHY_283 ();
 b15ztpn00an1n08x5 PHY_284 ();
 b15ztpn00an1n08x5 PHY_285 ();
 b15ztpn00an1n08x5 PHY_286 ();
 b15ztpn00an1n08x5 PHY_287 ();
 b15ztpn00an1n08x5 PHY_288 ();
 b15ztpn00an1n08x5 PHY_289 ();
 b15ztpn00an1n08x5 PHY_290 ();
 b15ztpn00an1n08x5 PHY_291 ();
 b15ztpn00an1n08x5 PHY_292 ();
 b15ztpn00an1n08x5 PHY_293 ();
 b15ztpn00an1n08x5 PHY_294 ();
 b15ztpn00an1n08x5 PHY_295 ();
 b15ztpn00an1n08x5 PHY_296 ();
 b15ztpn00an1n08x5 PHY_297 ();
 b15ztpn00an1n08x5 PHY_298 ();
 b15ztpn00an1n08x5 PHY_299 ();
 b15ztpn00an1n08x5 PHY_300 ();
 b15ztpn00an1n08x5 PHY_301 ();
 b15ztpn00an1n08x5 PHY_302 ();
 b15ztpn00an1n08x5 PHY_303 ();
 b15ztpn00an1n08x5 PHY_304 ();
 b15ztpn00an1n08x5 PHY_305 ();
 b15ztpn00an1n08x5 PHY_306 ();
 b15ztpn00an1n08x5 PHY_307 ();
 b15ztpn00an1n08x5 PHY_308 ();
 b15ztpn00an1n08x5 PHY_309 ();
 b15ztpn00an1n08x5 PHY_310 ();
 b15ztpn00an1n08x5 PHY_311 ();
 b15ztpn00an1n08x5 PHY_312 ();
 b15ztpn00an1n08x5 PHY_313 ();
 b15ztpn00an1n08x5 PHY_314 ();
 b15ztpn00an1n08x5 PHY_315 ();
 b15ztpn00an1n08x5 PHY_316 ();
 b15ztpn00an1n08x5 PHY_317 ();
 b15ztpn00an1n08x5 PHY_318 ();
 b15ztpn00an1n08x5 PHY_319 ();
 b15ztpn00an1n08x5 PHY_320 ();
 b15ztpn00an1n08x5 PHY_321 ();
 b15ztpn00an1n08x5 PHY_322 ();
 b15ztpn00an1n08x5 PHY_323 ();
 b15ztpn00an1n08x5 PHY_324 ();
 b15ztpn00an1n08x5 PHY_325 ();
 b15ztpn00an1n08x5 PHY_326 ();
 b15ztpn00an1n08x5 PHY_327 ();
 b15ztpn00an1n08x5 PHY_328 ();
 b15ztpn00an1n08x5 PHY_329 ();
 b15ztpn00an1n08x5 PHY_330 ();
 b15ztpn00an1n08x5 PHY_331 ();
 b15ztpn00an1n08x5 PHY_332 ();
 b15ztpn00an1n08x5 PHY_333 ();
 b15ztpn00an1n08x5 PHY_334 ();
 b15ztpn00an1n08x5 PHY_335 ();
 b15ztpn00an1n08x5 PHY_336 ();
 b15ztpn00an1n08x5 PHY_337 ();
 b15ztpn00an1n08x5 PHY_338 ();
 b15ztpn00an1n08x5 PHY_339 ();
 b15ztpn00an1n08x5 PHY_340 ();
 b15ztpn00an1n08x5 PHY_341 ();
 b15ztpn00an1n08x5 PHY_342 ();
 b15ztpn00an1n08x5 PHY_343 ();
 b15ztpn00an1n08x5 PHY_344 ();
 b15ztpn00an1n08x5 PHY_345 ();
 b15ztpn00an1n08x5 PHY_346 ();
 b15ztpn00an1n08x5 PHY_347 ();
 b15ztpn00an1n08x5 PHY_348 ();
 b15ztpn00an1n08x5 PHY_349 ();
 b15ztpn00an1n08x5 PHY_350 ();
 b15ztpn00an1n08x5 PHY_351 ();
 b15ztpn00an1n08x5 PHY_352 ();
 b15ztpn00an1n08x5 PHY_353 ();
 b15ztpn00an1n08x5 PHY_354 ();
 b15ztpn00an1n08x5 PHY_355 ();
 b15ztpn00an1n08x5 PHY_356 ();
 b15ztpn00an1n08x5 PHY_357 ();
 b15ztpn00an1n08x5 PHY_358 ();
 b15ztpn00an1n08x5 PHY_359 ();
 b15ztpn00an1n08x5 PHY_360 ();
 b15ztpn00an1n08x5 PHY_361 ();
 b15ztpn00an1n08x5 PHY_362 ();
 b15ztpn00an1n08x5 PHY_363 ();
 b15ztpn00an1n08x5 PHY_364 ();
 b15ztpn00an1n08x5 PHY_365 ();
 b15ztpn00an1n08x5 PHY_366 ();
 b15ztpn00an1n08x5 PHY_367 ();
 b15ztpn00an1n08x5 PHY_368 ();
 b15ztpn00an1n08x5 PHY_369 ();
 b15ztpn00an1n08x5 PHY_370 ();
 b15ztpn00an1n08x5 PHY_371 ();
 b15ztpn00an1n08x5 PHY_372 ();
 b15ztpn00an1n08x5 PHY_373 ();
 b15ztpn00an1n08x5 PHY_374 ();
 b15ztpn00an1n08x5 PHY_375 ();
 b15ztpn00an1n08x5 PHY_376 ();
 b15ztpn00an1n08x5 PHY_377 ();
 b15ztpn00an1n08x5 PHY_378 ();
 b15ztpn00an1n08x5 PHY_379 ();
 b15ztpn00an1n08x5 PHY_380 ();
 b15ztpn00an1n08x5 PHY_381 ();
 b15ztpn00an1n08x5 PHY_382 ();
 b15ztpn00an1n08x5 PHY_383 ();
 b15ztpn00an1n08x5 PHY_384 ();
 b15ztpn00an1n08x5 PHY_385 ();
 b15ztpn00an1n08x5 PHY_386 ();
 b15ztpn00an1n08x5 PHY_387 ();
 b15ztpn00an1n08x5 PHY_388 ();
 b15ztpn00an1n08x5 PHY_389 ();
 b15ztpn00an1n08x5 TAP_390 ();
 b15ztpn00an1n08x5 TAP_391 ();
 b15ztpn00an1n08x5 TAP_392 ();
 b15ztpn00an1n08x5 TAP_393 ();
 b15ztpn00an1n08x5 TAP_394 ();
 b15ztpn00an1n08x5 TAP_395 ();
 b15ztpn00an1n08x5 TAP_396 ();
 b15ztpn00an1n08x5 TAP_397 ();
 b15ztpn00an1n08x5 TAP_398 ();
 b15ztpn00an1n08x5 TAP_399 ();
 b15ztpn00an1n08x5 TAP_400 ();
 b15ztpn00an1n08x5 TAP_401 ();
 b15ztpn00an1n08x5 TAP_402 ();
 b15ztpn00an1n08x5 TAP_403 ();
 b15ztpn00an1n08x5 TAP_404 ();
 b15ztpn00an1n08x5 TAP_405 ();
 b15ztpn00an1n08x5 TAP_406 ();
 b15ztpn00an1n08x5 TAP_407 ();
 b15ztpn00an1n08x5 TAP_408 ();
 b15ztpn00an1n08x5 TAP_409 ();
 b15ztpn00an1n08x5 TAP_410 ();
 b15ztpn00an1n08x5 TAP_411 ();
 b15ztpn00an1n08x5 TAP_412 ();
 b15ztpn00an1n08x5 TAP_413 ();
 b15ztpn00an1n08x5 TAP_414 ();
 b15ztpn00an1n08x5 TAP_415 ();
 b15ztpn00an1n08x5 TAP_416 ();
 b15ztpn00an1n08x5 TAP_417 ();
 b15ztpn00an1n08x5 TAP_418 ();
 b15ztpn00an1n08x5 TAP_419 ();
 b15ztpn00an1n08x5 TAP_420 ();
 b15ztpn00an1n08x5 TAP_421 ();
 b15ztpn00an1n08x5 TAP_422 ();
 b15ztpn00an1n08x5 TAP_423 ();
 b15ztpn00an1n08x5 TAP_424 ();
 b15ztpn00an1n08x5 TAP_425 ();
 b15ztpn00an1n08x5 TAP_426 ();
 b15ztpn00an1n08x5 TAP_427 ();
 b15ztpn00an1n08x5 TAP_428 ();
 b15ztpn00an1n08x5 TAP_429 ();
 b15ztpn00an1n08x5 TAP_430 ();
 b15ztpn00an1n08x5 TAP_431 ();
 b15ztpn00an1n08x5 TAP_432 ();
 b15ztpn00an1n08x5 TAP_433 ();
 b15ztpn00an1n08x5 TAP_434 ();
 b15ztpn00an1n08x5 TAP_435 ();
 b15ztpn00an1n08x5 TAP_436 ();
 b15ztpn00an1n08x5 TAP_437 ();
 b15ztpn00an1n08x5 TAP_438 ();
 b15ztpn00an1n08x5 TAP_439 ();
 b15ztpn00an1n08x5 TAP_440 ();
 b15ztpn00an1n08x5 TAP_441 ();
 b15ztpn00an1n08x5 TAP_442 ();
 b15ztpn00an1n08x5 TAP_443 ();
 b15ztpn00an1n08x5 TAP_444 ();
 b15ztpn00an1n08x5 TAP_445 ();
 b15ztpn00an1n08x5 TAP_446 ();
 b15ztpn00an1n08x5 TAP_447 ();
 b15ztpn00an1n08x5 TAP_448 ();
 b15ztpn00an1n08x5 TAP_449 ();
 b15ztpn00an1n08x5 TAP_450 ();
 b15ztpn00an1n08x5 TAP_451 ();
 b15ztpn00an1n08x5 TAP_452 ();
 b15ztpn00an1n08x5 TAP_453 ();
 b15ztpn00an1n08x5 TAP_454 ();
 b15ztpn00an1n08x5 TAP_455 ();
 b15ztpn00an1n08x5 TAP_456 ();
 b15ztpn00an1n08x5 TAP_457 ();
 b15ztpn00an1n08x5 TAP_458 ();
 b15ztpn00an1n08x5 TAP_459 ();
 b15ztpn00an1n08x5 TAP_460 ();
 b15ztpn00an1n08x5 TAP_461 ();
 b15ztpn00an1n08x5 TAP_462 ();
 b15ztpn00an1n08x5 TAP_463 ();
 b15ztpn00an1n08x5 TAP_464 ();
 b15ztpn00an1n08x5 TAP_465 ();
 b15ztpn00an1n08x5 TAP_466 ();
 b15ztpn00an1n08x5 TAP_467 ();
 b15ztpn00an1n08x5 TAP_468 ();
 b15ztpn00an1n08x5 TAP_469 ();
 b15ztpn00an1n08x5 TAP_470 ();
 b15ztpn00an1n08x5 TAP_471 ();
 b15ztpn00an1n08x5 TAP_472 ();
 b15ztpn00an1n08x5 TAP_473 ();
 b15ztpn00an1n08x5 TAP_474 ();
 b15ztpn00an1n08x5 TAP_475 ();
 b15ztpn00an1n08x5 TAP_476 ();
 b15ztpn00an1n08x5 TAP_477 ();
 b15ztpn00an1n08x5 TAP_478 ();
 b15ztpn00an1n08x5 TAP_479 ();
 b15ztpn00an1n08x5 TAP_480 ();
 b15ztpn00an1n08x5 TAP_481 ();
 b15ztpn00an1n08x5 TAP_482 ();
 b15ztpn00an1n08x5 TAP_483 ();
 b15ztpn00an1n08x5 TAP_484 ();
 b15ztpn00an1n08x5 TAP_485 ();
 b15ztpn00an1n08x5 TAP_486 ();
 b15ztpn00an1n08x5 TAP_487 ();
 b15ztpn00an1n08x5 TAP_488 ();
 b15ztpn00an1n08x5 TAP_489 ();
 b15ztpn00an1n08x5 TAP_490 ();
 b15ztpn00an1n08x5 TAP_491 ();
 b15ztpn00an1n08x5 TAP_492 ();
 b15ztpn00an1n08x5 TAP_493 ();
 b15ztpn00an1n08x5 TAP_494 ();
 b15ztpn00an1n08x5 TAP_495 ();
 b15ztpn00an1n08x5 TAP_496 ();
 b15ztpn00an1n08x5 TAP_497 ();
 b15ztpn00an1n08x5 TAP_498 ();
 b15ztpn00an1n08x5 TAP_499 ();
 b15ztpn00an1n08x5 TAP_500 ();
 b15ztpn00an1n08x5 TAP_501 ();
 b15ztpn00an1n08x5 TAP_502 ();
 b15ztpn00an1n08x5 TAP_503 ();
 b15ztpn00an1n08x5 TAP_504 ();
 b15ztpn00an1n08x5 TAP_505 ();
 b15ztpn00an1n08x5 TAP_506 ();
 b15ztpn00an1n08x5 TAP_507 ();
 b15ztpn00an1n08x5 TAP_508 ();
 b15ztpn00an1n08x5 TAP_509 ();
 b15ztpn00an1n08x5 TAP_510 ();
 b15ztpn00an1n08x5 TAP_511 ();
 b15ztpn00an1n08x5 TAP_512 ();
 b15ztpn00an1n08x5 TAP_513 ();
 b15ztpn00an1n08x5 TAP_514 ();
 b15ztpn00an1n08x5 TAP_515 ();
 b15ztpn00an1n08x5 TAP_516 ();
 b15ztpn00an1n08x5 TAP_517 ();
 b15ztpn00an1n08x5 TAP_518 ();
 b15ztpn00an1n08x5 TAP_519 ();
 b15ztpn00an1n08x5 TAP_520 ();
 b15ztpn00an1n08x5 TAP_521 ();
 b15ztpn00an1n08x5 TAP_522 ();
 b15ztpn00an1n08x5 TAP_523 ();
 b15ztpn00an1n08x5 TAP_524 ();
 b15ztpn00an1n08x5 TAP_525 ();
 b15ztpn00an1n08x5 TAP_526 ();
 b15ztpn00an1n08x5 TAP_527 ();
 b15ztpn00an1n08x5 TAP_528 ();
 b15ztpn00an1n08x5 TAP_529 ();
 b15ztpn00an1n08x5 TAP_530 ();
 b15ztpn00an1n08x5 TAP_531 ();
 b15ztpn00an1n08x5 TAP_532 ();
 b15ztpn00an1n08x5 TAP_533 ();
 b15ztpn00an1n08x5 TAP_534 ();
 b15ztpn00an1n08x5 TAP_535 ();
 b15ztpn00an1n08x5 TAP_536 ();
 b15ztpn00an1n08x5 TAP_537 ();
 b15ztpn00an1n08x5 TAP_538 ();
 b15ztpn00an1n08x5 TAP_539 ();
 b15ztpn00an1n08x5 TAP_540 ();
 b15ztpn00an1n08x5 TAP_541 ();
 b15ztpn00an1n08x5 TAP_542 ();
 b15ztpn00an1n08x5 TAP_543 ();
 b15ztpn00an1n08x5 TAP_544 ();
 b15ztpn00an1n08x5 TAP_545 ();
 b15ztpn00an1n08x5 TAP_546 ();
 b15ztpn00an1n08x5 TAP_547 ();
 b15ztpn00an1n08x5 TAP_548 ();
 b15ztpn00an1n08x5 TAP_549 ();
 b15ztpn00an1n08x5 TAP_550 ();
 b15ztpn00an1n08x5 TAP_551 ();
 b15ztpn00an1n08x5 TAP_552 ();
 b15ztpn00an1n08x5 TAP_553 ();
 b15ztpn00an1n08x5 TAP_554 ();
 b15ztpn00an1n08x5 TAP_555 ();
 b15ztpn00an1n08x5 TAP_556 ();
 b15ztpn00an1n08x5 TAP_557 ();
 b15ztpn00an1n08x5 TAP_558 ();
 b15ztpn00an1n08x5 TAP_559 ();
 b15ztpn00an1n08x5 TAP_560 ();
 b15ztpn00an1n08x5 TAP_561 ();
 b15ztpn00an1n08x5 TAP_562 ();
 b15ztpn00an1n08x5 TAP_563 ();
 b15ztpn00an1n08x5 TAP_564 ();
 b15ztpn00an1n08x5 TAP_565 ();
 b15ztpn00an1n08x5 TAP_566 ();
 b15ztpn00an1n08x5 TAP_567 ();
 b15ztpn00an1n08x5 TAP_568 ();
 b15ztpn00an1n08x5 TAP_569 ();
 b15ztpn00an1n08x5 TAP_570 ();
 b15ztpn00an1n08x5 TAP_571 ();
 b15ztpn00an1n08x5 TAP_572 ();
 b15ztpn00an1n08x5 TAP_573 ();
 b15ztpn00an1n08x5 TAP_574 ();
 b15ztpn00an1n08x5 TAP_575 ();
 b15ztpn00an1n08x5 TAP_576 ();
 b15ztpn00an1n08x5 TAP_577 ();
 b15ztpn00an1n08x5 TAP_578 ();
 b15ztpn00an1n08x5 TAP_579 ();
 b15ztpn00an1n08x5 TAP_580 ();
 b15ztpn00an1n08x5 TAP_581 ();
 b15ztpn00an1n08x5 TAP_582 ();
 b15ztpn00an1n08x5 TAP_583 ();
 b15ztpn00an1n08x5 TAP_584 ();
 b15ztpn00an1n08x5 TAP_585 ();
 b15ztpn00an1n08x5 TAP_586 ();
 b15ztpn00an1n08x5 TAP_587 ();
 b15ztpn00an1n08x5 TAP_588 ();
 b15ztpn00an1n08x5 TAP_589 ();
 b15ztpn00an1n08x5 TAP_590 ();
 b15ztpn00an1n08x5 TAP_591 ();
 b15ztpn00an1n08x5 TAP_592 ();
 b15ztpn00an1n08x5 TAP_593 ();
 b15ztpn00an1n08x5 TAP_594 ();
 b15ztpn00an1n08x5 TAP_595 ();
 b15ztpn00an1n08x5 TAP_596 ();
 b15ztpn00an1n08x5 TAP_597 ();
 b15ztpn00an1n08x5 TAP_598 ();
 b15ztpn00an1n08x5 TAP_599 ();
 b15ztpn00an1n08x5 TAP_600 ();
 b15ztpn00an1n08x5 TAP_601 ();
 b15ztpn00an1n08x5 TAP_602 ();
 b15ztpn00an1n08x5 TAP_603 ();
 b15ztpn00an1n08x5 TAP_604 ();
 b15ztpn00an1n08x5 TAP_605 ();
 b15ztpn00an1n08x5 TAP_606 ();
 b15ztpn00an1n08x5 TAP_607 ();
 b15ztpn00an1n08x5 TAP_608 ();
 b15ztpn00an1n08x5 TAP_609 ();
 b15ztpn00an1n08x5 TAP_610 ();
 b15ztpn00an1n08x5 TAP_611 ();
 b15ztpn00an1n08x5 TAP_612 ();
 b15ztpn00an1n08x5 TAP_613 ();
 b15ztpn00an1n08x5 TAP_614 ();
 b15ztpn00an1n08x5 TAP_615 ();
 b15ztpn00an1n08x5 TAP_616 ();
 b15ztpn00an1n08x5 TAP_617 ();
 b15ztpn00an1n08x5 TAP_618 ();
 b15ztpn00an1n08x5 TAP_619 ();
 b15ztpn00an1n08x5 TAP_620 ();
 b15ztpn00an1n08x5 TAP_621 ();
 b15ztpn00an1n08x5 TAP_622 ();
 b15ztpn00an1n08x5 TAP_623 ();
 b15ztpn00an1n08x5 TAP_624 ();
 b15ztpn00an1n08x5 TAP_625 ();
 b15ztpn00an1n08x5 TAP_626 ();
 b15ztpn00an1n08x5 TAP_627 ();
 b15ztpn00an1n08x5 TAP_628 ();
 b15ztpn00an1n08x5 TAP_629 ();
 b15ztpn00an1n08x5 TAP_630 ();
 b15ztpn00an1n08x5 TAP_631 ();
 b15ztpn00an1n08x5 TAP_632 ();
 b15ztpn00an1n08x5 TAP_633 ();
 b15ztpn00an1n08x5 TAP_634 ();
 b15ztpn00an1n08x5 TAP_635 ();
 b15ztpn00an1n08x5 TAP_636 ();
 b15ztpn00an1n08x5 TAP_637 ();
 b15ztpn00an1n08x5 TAP_638 ();
 b15ztpn00an1n08x5 TAP_639 ();
 b15ztpn00an1n08x5 TAP_640 ();
 b15ztpn00an1n08x5 TAP_641 ();
 b15ztpn00an1n08x5 TAP_642 ();
 b15ztpn00an1n08x5 TAP_643 ();
 b15ztpn00an1n08x5 TAP_644 ();
 b15ztpn00an1n08x5 TAP_645 ();
 b15ztpn00an1n08x5 TAP_646 ();
 b15ztpn00an1n08x5 TAP_647 ();
 b15ztpn00an1n08x5 TAP_648 ();
 b15ztpn00an1n08x5 TAP_649 ();
 b15ztpn00an1n08x5 TAP_650 ();
 b15ztpn00an1n08x5 TAP_651 ();
 b15ztpn00an1n08x5 TAP_652 ();
 b15ztpn00an1n08x5 TAP_653 ();
 b15ztpn00an1n08x5 TAP_654 ();
 b15ztpn00an1n08x5 TAP_655 ();
 b15ztpn00an1n08x5 TAP_656 ();
 b15ztpn00an1n08x5 TAP_657 ();
 b15ztpn00an1n08x5 TAP_658 ();
 b15ztpn00an1n08x5 TAP_659 ();
 b15ztpn00an1n08x5 TAP_660 ();
 b15ztpn00an1n08x5 TAP_661 ();
 b15ztpn00an1n08x5 TAP_662 ();
 b15ztpn00an1n08x5 TAP_663 ();
 b15ztpn00an1n08x5 TAP_664 ();
 b15ztpn00an1n08x5 TAP_665 ();
 b15ztpn00an1n08x5 TAP_666 ();
 b15ztpn00an1n08x5 TAP_667 ();
 b15ztpn00an1n08x5 TAP_668 ();
 b15ztpn00an1n08x5 TAP_669 ();
 b15ztpn00an1n08x5 TAP_670 ();
 b15ztpn00an1n08x5 TAP_671 ();
 b15ztpn00an1n08x5 TAP_672 ();
 b15ztpn00an1n08x5 TAP_673 ();
 b15ztpn00an1n08x5 TAP_674 ();
 b15ztpn00an1n08x5 TAP_675 ();
 b15ztpn00an1n08x5 TAP_676 ();
 b15ztpn00an1n08x5 TAP_677 ();
 b15ztpn00an1n08x5 TAP_678 ();
 b15ztpn00an1n08x5 TAP_679 ();
 b15ztpn00an1n08x5 TAP_680 ();
 b15ztpn00an1n08x5 TAP_681 ();
 b15ztpn00an1n08x5 TAP_682 ();
 b15ztpn00an1n08x5 TAP_683 ();
 b15ztpn00an1n08x5 TAP_684 ();
 b15ztpn00an1n08x5 TAP_685 ();
 b15ztpn00an1n08x5 TAP_686 ();
 b15ztpn00an1n08x5 TAP_687 ();
 b15ztpn00an1n08x5 TAP_688 ();
 b15ztpn00an1n08x5 TAP_689 ();
 b15ztpn00an1n08x5 TAP_690 ();
 b15ztpn00an1n08x5 TAP_691 ();
 b15ztpn00an1n08x5 TAP_692 ();
 b15ztpn00an1n08x5 TAP_693 ();
 b15ztpn00an1n08x5 TAP_694 ();
 b15ztpn00an1n08x5 TAP_695 ();
 b15ztpn00an1n08x5 TAP_696 ();
 b15ztpn00an1n08x5 TAP_697 ();
 b15ztpn00an1n08x5 TAP_698 ();
 b15ztpn00an1n08x5 TAP_699 ();
 b15ztpn00an1n08x5 TAP_700 ();
 b15ztpn00an1n08x5 TAP_701 ();
 b15ztpn00an1n08x5 TAP_702 ();
 b15ztpn00an1n08x5 TAP_703 ();
 b15ztpn00an1n08x5 TAP_704 ();
 b15ztpn00an1n08x5 TAP_705 ();
 b15ztpn00an1n08x5 TAP_706 ();
 b15ztpn00an1n08x5 TAP_707 ();
 b15ztpn00an1n08x5 TAP_708 ();
 b15ztpn00an1n08x5 TAP_709 ();
 b15ztpn00an1n08x5 TAP_710 ();
 b15ztpn00an1n08x5 TAP_711 ();
 b15ztpn00an1n08x5 TAP_712 ();
 b15ztpn00an1n08x5 TAP_713 ();
 b15ztpn00an1n08x5 TAP_714 ();
 b15ztpn00an1n08x5 TAP_715 ();
 b15ztpn00an1n08x5 TAP_716 ();
 b15ztpn00an1n08x5 TAP_717 ();
 b15ztpn00an1n08x5 TAP_718 ();
 b15ztpn00an1n08x5 TAP_719 ();
 b15ztpn00an1n08x5 TAP_720 ();
 b15ztpn00an1n08x5 TAP_721 ();
 b15ztpn00an1n08x5 TAP_722 ();
 b15ztpn00an1n08x5 TAP_723 ();
 b15ztpn00an1n08x5 TAP_724 ();
 b15ztpn00an1n08x5 TAP_725 ();
 b15ztpn00an1n08x5 TAP_726 ();
 b15ztpn00an1n08x5 TAP_727 ();
 b15ztpn00an1n08x5 TAP_728 ();
 b15ztpn00an1n08x5 TAP_729 ();
 b15ztpn00an1n08x5 TAP_730 ();
 b15ztpn00an1n08x5 TAP_731 ();
 b15ztpn00an1n08x5 TAP_732 ();
 b15ztpn00an1n08x5 TAP_733 ();
 b15ztpn00an1n08x5 TAP_734 ();
 b15ztpn00an1n08x5 TAP_735 ();
 b15ztpn00an1n08x5 TAP_736 ();
 b15ztpn00an1n08x5 TAP_737 ();
 b15ztpn00an1n08x5 TAP_738 ();
 b15ztpn00an1n08x5 TAP_739 ();
 b15ztpn00an1n08x5 TAP_740 ();
 b15ztpn00an1n08x5 TAP_741 ();
 b15ztpn00an1n08x5 TAP_742 ();
 b15ztpn00an1n08x5 TAP_743 ();
 b15ztpn00an1n08x5 TAP_744 ();
 b15ztpn00an1n08x5 TAP_745 ();
 b15ztpn00an1n08x5 TAP_746 ();
 b15ztpn00an1n08x5 TAP_747 ();
 b15ztpn00an1n08x5 TAP_748 ();
 b15ztpn00an1n08x5 TAP_749 ();
 b15ztpn00an1n08x5 TAP_750 ();
 b15ztpn00an1n08x5 TAP_751 ();
 b15ztpn00an1n08x5 TAP_752 ();
 b15ztpn00an1n08x5 TAP_753 ();
 b15ztpn00an1n08x5 TAP_754 ();
 b15ztpn00an1n08x5 TAP_755 ();
 b15ztpn00an1n08x5 TAP_756 ();
 b15ztpn00an1n08x5 TAP_757 ();
 b15ztpn00an1n08x5 TAP_758 ();
 b15ztpn00an1n08x5 TAP_759 ();
 b15ztpn00an1n08x5 TAP_760 ();
 b15ztpn00an1n08x5 TAP_761 ();
 b15ztpn00an1n08x5 TAP_762 ();
 b15ztpn00an1n08x5 TAP_763 ();
 b15ztpn00an1n08x5 TAP_764 ();
 b15ztpn00an1n08x5 TAP_765 ();
 b15ztpn00an1n08x5 TAP_766 ();
 b15ztpn00an1n08x5 TAP_767 ();
 b15ztpn00an1n08x5 TAP_768 ();
 b15ztpn00an1n08x5 TAP_769 ();
 b15ztpn00an1n08x5 TAP_770 ();
 b15ztpn00an1n08x5 TAP_771 ();
 b15ztpn00an1n08x5 TAP_772 ();
 b15ztpn00an1n08x5 TAP_773 ();
 b15ztpn00an1n08x5 TAP_774 ();
 b15ztpn00an1n08x5 TAP_775 ();
 b15ztpn00an1n08x5 TAP_776 ();
 b15ztpn00an1n08x5 TAP_777 ();
 b15ztpn00an1n08x5 TAP_778 ();
 b15ztpn00an1n08x5 TAP_779 ();
 b15ztpn00an1n08x5 TAP_780 ();
 b15bfn000ah1n02x5 input1 (.a(alert_rx_i[0]),
    .o(net1));
 b15bfn000ah1n04x5 input2 (.a(alert_rx_i[1]),
    .o(net2));
 b15bfn000ah1n04x5 input3 (.a(alert_rx_i[2]),
    .o(net3));
 b15bfn000ah1n03x5 input4 (.a(alert_rx_i[3]),
    .o(net4));
 b15qgbbf1an1n05x5 input5 (.a(cio_gpio_i[0]),
    .o(net5));
 b15bfn001ah1n08x5 input6 (.a(cio_gpio_i[10]),
    .o(net6));
 b15bfn001as1n08x5 input7 (.a(cio_gpio_i[11]),
    .o(net7));
 b15bfn001as1n12x5 input8 (.a(cio_gpio_i[12]),
    .o(net8));
 b15bfn001ah1n16x5 input9 (.a(cio_gpio_i[13]),
    .o(net9));
 b15bfn000ar1n02x5 input10 (.a(cio_gpio_i[14]),
    .o(net10));
 b15bfn001ah1n08x5 input11 (.a(cio_gpio_i[15]),
    .o(net11));
 b15bfn000as1n03x5 input12 (.a(cio_gpio_i[16]),
    .o(net12));
 b15bfn001aq1n06x5 input13 (.a(cio_gpio_i[17]),
    .o(net13));
 b15bfn001aq1n06x5 input14 (.a(cio_gpio_i[18]),
    .o(net14));
 b15bfn000as1n02x5 input15 (.a(cio_gpio_i[19]),
    .o(net15));
 b15bfn000as1n04x5 input16 (.a(cio_gpio_i[1]),
    .o(net16));
 b15bfn001as1n12x5 input17 (.a(cio_gpio_i[20]),
    .o(net17));
 b15bfn001as1n08x5 input18 (.a(cio_gpio_i[21]),
    .o(net18));
 b15bfn001as1n06x5 input19 (.a(cio_gpio_i[22]),
    .o(net19));
 b15bfn000as1n03x5 input20 (.a(cio_gpio_i[23]),
    .o(net20));
 b15bfn000ah1n03x5 input21 (.a(cio_gpio_i[24]),
    .o(net21));
 b15bfn001aq1n06x5 input22 (.a(cio_gpio_i[25]),
    .o(net22));
 b15bfn000as1n03x5 input23 (.a(cio_gpio_i[26]),
    .o(net23));
 b15bfm201as1n04x5 input24 (.a(cio_gpio_i[27]),
    .o(net24));
 b15bfn000ah1n04x5 input25 (.a(cio_gpio_i[28]),
    .o(net25));
 b15bfn000as1n03x5 input26 (.a(cio_gpio_i[29]),
    .o(net26));
 b15bfn001as1n16x5 input27 (.a(cio_gpio_i[2]),
    .o(net27));
 b15bfn001ah1n08x5 input28 (.a(cio_gpio_i[30]),
    .o(net28));
 b15bfn001ah1n08x5 input29 (.a(cio_gpio_i[31]),
    .o(net29));
 b15bfn001as1n06x5 input30 (.a(cio_gpio_i[3]),
    .o(net30));
 b15bfn001ah1n08x5 input31 (.a(cio_gpio_i[4]),
    .o(net31));
 b15bfn000ah1n06x5 input32 (.a(cio_gpio_i[5]),
    .o(net32));
 b15bfn000as1n03x5 input33 (.a(cio_gpio_i[6]),
    .o(net33));
 b15bfn001ah1n06x5 input34 (.a(cio_gpio_i[7]),
    .o(net34));
 b15bfn001as1n06x5 input35 (.a(cio_gpio_i[8]),
    .o(net35));
 b15bfn001as1n08x5 input36 (.a(cio_gpio_i[9]),
    .o(net36));
 b15bfn001as1n32x5 input37 (.a(net2305),
    .o(net37));
 b15bfn000al1n02x5 input38 (.a(tl_i[0]),
    .o(net38));
 b15bfn001as1n08x5 input39 (.a(tl_i[100]),
    .o(net39));
 b15bfn001ah1n08x5 input40 (.a(tl_i[101]),
    .o(net40));
 b15bfn001as1n08x5 input41 (.a(tl_i[105]),
    .o(net41));
 b15bfn000ah1n06x5 input42 (.a(tl_i[106]),
    .o(net42));
 b15bfn001as1n16x5 input43 (.a(tl_i[107]),
    .o(net43));
 b15bfn001ah1n12x5 input44 (.a(tl_i[108]),
    .o(net44));
 b15qgbbf1an1n05x5 input45 (.a(tl_i[10]),
    .o(net45));
 b15bfn001aq1n06x5 input46 (.a(tl_i[11]),
    .o(net46));
 b15bfn000as1n03x5 input47 (.a(tl_i[12]),
    .o(net47));
 b15bfn000as1n03x5 input48 (.a(tl_i[13]),
    .o(net48));
 b15bfn000ah1n06x5 input49 (.a(tl_i[14]),
    .o(net49));
 b15bfn001as1n16x5 input50 (.a(tl_i[15]),
    .o(net50));
 b15bfn001ah1n16x5 input51 (.a(tl_i[16]),
    .o(net51));
 b15bfn001ah1n16x5 input52 (.a(tl_i[17]),
    .o(net52));
 b15bfn001as1n12x5 input53 (.a(tl_i[18]),
    .o(net53));
 b15bfn001as1n08x5 input54 (.a(tl_i[1]),
    .o(net54));
 b15bfn001ah1n64x5 input55 (.a(tl_i[24]),
    .o(net55));
 b15bfn001as1n48x5 input56 (.a(tl_i[25]),
    .o(net56));
 b15bfn001as1n48x5 input57 (.a(tl_i[26]),
    .o(net57));
 b15bfn001as1n32x5 input58 (.a(tl_i[27]),
    .o(net58));
 b15bfn001ah1n24x5 input59 (.a(tl_i[28]),
    .o(net59));
 b15bfn001ah1n64x5 input60 (.a(tl_i[29]),
    .o(net60));
 b15bfn001ah1n16x5 input61 (.a(tl_i[2]),
    .o(net61));
 b15bfn001ah1n48x5 input62 (.a(tl_i[30]),
    .o(net62));
 b15bfn001ah1n48x5 input63 (.a(tl_i[31]),
    .o(net63));
 b15bfn001as1n32x5 input64 (.a(tl_i[32]),
    .o(net64));
 b15bfn001ah1n32x5 input65 (.a(tl_i[33]),
    .o(net65));
 b15bfn000as1n32x5 input66 (.a(tl_i[34]),
    .o(net66));
 b15bfn001as1n32x5 input67 (.a(tl_i[35]),
    .o(net67));
 b15bfn001as1n32x5 input68 (.a(tl_i[36]),
    .o(net68));
 b15bfn001as1n16x5 input69 (.a(tl_i[37]),
    .o(net69));
 b15bfn001as1n32x5 input70 (.a(tl_i[38]),
    .o(net70));
 b15bfn001ah1n48x5 input71 (.a(tl_i[39]),
    .o(net71));
 b15bfn001as1n08x5 input72 (.a(tl_i[3]),
    .o(net72));
 b15bfn001as1n48x5 input73 (.a(tl_i[40]),
    .o(net73));
 b15bfn001as1n24x5 input74 (.a(tl_i[41]),
    .o(net74));
 b15bfn001ah1n48x5 input75 (.a(net2549),
    .o(net75));
 b15bfn001as1n48x5 input76 (.a(tl_i[43]),
    .o(net76));
 b15bfn001ah1n32x5 input77 (.a(tl_i[44]),
    .o(net77));
 b15bfn001as1n48x5 input78 (.a(tl_i[45]),
    .o(net78));
 b15bfn001ah1n24x5 input79 (.a(tl_i[46]),
    .o(net79));
 b15bfn001as1n32x5 input80 (.a(tl_i[47]),
    .o(net80));
 b15bfn001as1n24x5 input81 (.a(tl_i[48]),
    .o(net81));
 b15bfn001as1n16x5 input82 (.a(tl_i[49]),
    .o(net82));
 b15bfn001as1n12x5 input83 (.a(tl_i[4]),
    .o(net83));
 b15bfn001ah1n24x5 input84 (.a(tl_i[50]),
    .o(net84));
 b15bfn000ah1n24x5 input85 (.a(tl_i[51]),
    .o(net85));
 b15bfn001as1n24x5 input86 (.a(tl_i[52]),
    .o(net86));
 b15bfn001ah1n16x5 input87 (.a(tl_i[53]),
    .o(net87));
 b15bfn000as1n32x5 input88 (.a(tl_i[54]),
    .o(net88));
 b15bfn001as1n32x5 input89 (.a(tl_i[55]),
    .o(net89));
 b15bfn001ah1n24x5 input90 (.a(tl_i[56]),
    .o(net90));
 b15bfn001ah1n24x5 input91 (.a(tl_i[57]),
    .o(net91));
 b15bfn001ah1n16x5 input92 (.a(tl_i[58]),
    .o(net92));
 b15bfn001as1n16x5 input93 (.a(tl_i[59]),
    .o(net93));
 b15bfn001as1n08x5 input94 (.a(tl_i[5]),
    .o(net94));
 b15bfn001ah1n16x5 input95 (.a(tl_i[60]),
    .o(net95));
 b15bfn001as1n16x5 input96 (.a(tl_i[61]),
    .o(net96));
 b15bfn001ah1n48x5 input97 (.a(tl_i[62]),
    .o(net97));
 b15bfn001as1n32x5 input98 (.a(tl_i[63]),
    .o(net98));
 b15bfn001as1n24x5 input99 (.a(tl_i[64]),
    .o(net99));
 b15bfn001ah1n24x5 input100 (.a(tl_i[65]),
    .o(net100));
 b15bfn001ah1n08x5 input101 (.a(tl_i[66]),
    .o(net101));
 b15bfn001as1n08x5 input102 (.a(tl_i[67]),
    .o(net102));
 b15bfn001as1n12x5 input103 (.a(tl_i[68]),
    .o(net103));
 b15bfn001as1n06x5 input104 (.a(tl_i[69]),
    .o(net104));
 b15bfn001ah1n08x5 input105 (.a(tl_i[6]),
    .o(net105));
 b15bfn001ah1n08x5 input106 (.a(tl_i[70]),
    .o(net106));
 b15bfn001as1n12x5 input107 (.a(tl_i[71]),
    .o(net107));
 b15bfn001ah1n08x5 input108 (.a(tl_i[72]),
    .o(net108));
 b15bfn001ah1n08x5 input109 (.a(tl_i[73]),
    .o(net109));
 b15bfn001ah1n12x5 input110 (.a(tl_i[74]),
    .o(net110));
 b15bfn001as1n12x5 input111 (.a(tl_i[75]),
    .o(net111));
 b15bfn001as1n08x5 input112 (.a(tl_i[76]),
    .o(net112));
 b15bfn001as1n06x5 input113 (.a(tl_i[77]),
    .o(net113));
 b15bfn001ah1n16x5 input114 (.a(tl_i[78]),
    .o(net114));
 b15bfn001as1n06x5 input115 (.a(tl_i[79]),
    .o(net115));
 b15bfn001aq1n06x5 input116 (.a(tl_i[7]),
    .o(net116));
 b15bfn001ah1n08x5 input117 (.a(tl_i[80]),
    .o(net117));
 b15bfn001as1n08x5 input118 (.a(tl_i[81]),
    .o(net118));
 b15bfn001ah1n08x5 input119 (.a(tl_i[82]),
    .o(net119));
 b15bfn000as1n12x5 input120 (.a(tl_i[83]),
    .o(net120));
 b15bfn001ah1n08x5 input121 (.a(tl_i[84]),
    .o(net121));
 b15bfn000as1n12x5 input122 (.a(tl_i[85]),
    .o(net122));
 b15bfn000ah1n06x5 input123 (.a(tl_i[86]),
    .o(net123));
 b15bfn001as1n12x5 input124 (.a(tl_i[87]),
    .o(net124));
 b15bfn001as1n08x5 input125 (.a(tl_i[88]),
    .o(net125));
 b15bfn001as1n08x5 input126 (.a(tl_i[89]),
    .o(net126));
 b15bfn000as1n04x5 input127 (.a(tl_i[8]),
    .o(net127));
 b15bfn001ah1n08x5 input128 (.a(tl_i[90]),
    .o(net128));
 b15bfn001as1n12x5 input129 (.a(tl_i[91]),
    .o(net129));
 b15bfn000ah1n03x5 input130 (.a(tl_i[92]),
    .o(net130));
 b15bfn000ah1n03x5 input131 (.a(tl_i[93]),
    .o(net131));
 b15bfn000ah1n04x5 input132 (.a(tl_i[94]),
    .o(net132));
 b15bfn000ah1n04x5 input133 (.a(tl_i[95]),
    .o(net133));
 b15bfn000ah1n03x5 input134 (.a(tl_i[96]),
    .o(net134));
 b15bfn000ah1n03x5 input135 (.a(tl_i[97]),
    .o(net135));
 b15bfn000as1n02x5 input136 (.a(tl_i[98]),
    .o(net136));
 b15bfn000as1n02x5 input137 (.a(tl_i[99]),
    .o(net137));
 b15bfn001as1n06x5 input138 (.a(tl_i[9]),
    .o(net138));
 b15bfn000ah1n03x5 output139 (.a(net2585),
    .o(net2029));
 b15bfn000ah1n03x5 output140 (.a(net2583),
    .o(net2038));
 b15bfn000ah1n03x5 output141 (.a(net2247),
    .o(cio_gpio_en_o[0]));
 b15bfn000ah1n03x5 output142 (.a(net2174),
    .o(cio_gpio_en_o[10]));
 b15bfn000ah1n03x5 output143 (.a(net2243),
    .o(cio_gpio_en_o[11]));
 b15bfn000ah1n03x5 output144 (.a(net2252),
    .o(cio_gpio_en_o[12]));
 b15bfn000ah1n03x5 output145 (.a(net2152),
    .o(net2153));
 b15bfn000ah1n03x5 output146 (.a(net2225),
    .o(cio_gpio_en_o[14]));
 b15bfn000ah1n03x5 output147 (.a(net2235),
    .o(cio_gpio_en_o[15]));
 b15bfn000ah1n03x5 output148 (.a(net722),
    .o(cio_gpio_en_o[16]));
 b15bfn000ah1n03x5 output149 (.a(net720),
    .o(cio_gpio_en_o[17]));
 b15bfn000ah1n03x5 output150 (.a(net717),
    .o(cio_gpio_en_o[18]));
 b15bfn000ah1n03x5 output151 (.a(net715),
    .o(cio_gpio_en_o[19]));
 b15bfn000ah1n03x5 output152 (.a(net2162),
    .o(net2163));
 b15bfn000ah1n03x5 output153 (.a(net2290),
    .o(cio_gpio_en_o[20]));
 b15bfn000ah1n03x5 output154 (.a(net2186),
    .o(net2187));
 b15bfn000ah1n03x5 output155 (.a(net713),
    .o(cio_gpio_en_o[22]));
 b15bfn000ah1n03x5 output156 (.a(net2196),
    .o(net2197));
 b15bfn000ah1n03x5 output157 (.a(net709),
    .o(cio_gpio_en_o[24]));
 b15bfn000ah1n03x5 output158 (.a(net2227),
    .o(cio_gpio_en_o[25]));
 b15bfn000ah1n03x5 output159 (.a(net2478),
    .o(cio_gpio_en_o[26]));
 b15bfn000ah1n03x5 output160 (.a(net704),
    .o(cio_gpio_en_o[27]));
 b15bfn000ah1n03x5 output161 (.a(net702),
    .o(cio_gpio_en_o[28]));
 b15bfn000ah1n03x5 output162 (.a(net701),
    .o(cio_gpio_en_o[29]));
 b15bfn000ah1n03x5 output163 (.a(net2219),
    .o(cio_gpio_en_o[2]));
 b15bfn000ah1n03x5 output164 (.a(net699),
    .o(cio_gpio_en_o[30]));
 b15bfn000ah1n03x5 output165 (.a(net697),
    .o(cio_gpio_en_o[31]));
 b15bfn000ah1n03x5 output166 (.a(net700),
    .o(cio_gpio_en_o[3]));
 b15bfn000ah1n03x5 output167 (.a(net2169),
    .o(net2170));
 b15bfn000ah1n03x5 output168 (.a(net695),
    .o(cio_gpio_en_o[5]));
 b15bfn000ah1n03x5 output169 (.a(net2222),
    .o(net2223));
 b15bfn000ah1n03x5 output170 (.a(net2198),
    .o(net2199));
 b15bfn000ah1n03x5 output171 (.a(net2171),
    .o(net2172));
 b15bfn000ah1n03x5 output172 (.a(net693),
    .o(cio_gpio_en_o[9]));
 b15bfn000ah1n03x5 output173 (.a(net173),
    .o(cio_gpio_o[0]));
 b15bfn000ah1n03x5 output174 (.a(net2530),
    .o(cio_gpio_o[10]));
 b15bfn000ah1n03x5 output175 (.a(net175),
    .o(cio_gpio_o[11]));
 b15bfn000ah1n03x5 output176 (.a(net176),
    .o(cio_gpio_o[12]));
 b15bfn000ah1n03x5 output177 (.a(net177),
    .o(cio_gpio_o[13]));
 b15bfn000ah1n03x5 output178 (.a(net688),
    .o(cio_gpio_o[14]));
 b15bfn000ah1n03x5 output179 (.a(net686),
    .o(cio_gpio_o[15]));
 b15bfn000ah1n03x5 output180 (.a(net684),
    .o(cio_gpio_o[16]));
 b15bfn000ah1n03x5 output181 (.a(net682),
    .o(cio_gpio_o[17]));
 b15bfn000ah1n03x5 output182 (.a(net182),
    .o(cio_gpio_o[18]));
 b15bfn000ah1n03x5 output183 (.a(net183),
    .o(cio_gpio_o[19]));
 b15bfn000ah1n03x5 output184 (.a(net184),
    .o(cio_gpio_o[1]));
 b15bfn000ah1n03x5 output185 (.a(net185),
    .o(cio_gpio_o[20]));
 b15bfn000ah1n03x5 output186 (.a(net186),
    .o(cio_gpio_o[21]));
 b15bfn000ah1n03x5 output187 (.a(net677),
    .o(cio_gpio_o[22]));
 b15bfn000ah1n03x5 output188 (.a(net673),
    .o(cio_gpio_o[23]));
 b15bfn000ah1n03x5 output189 (.a(net669),
    .o(cio_gpio_o[24]));
 b15bfn000ah1n03x5 output190 (.a(net667),
    .o(cio_gpio_o[25]));
 b15bfn000ah1n03x5 output191 (.a(net664),
    .o(cio_gpio_o[26]));
 b15bfn000ah1n03x5 output192 (.a(net660),
    .o(cio_gpio_o[27]));
 b15bfn000ah1n03x5 output193 (.a(net658),
    .o(cio_gpio_o[28]));
 b15bfn000ah1n03x5 output194 (.a(net656),
    .o(cio_gpio_o[29]));
 b15bfn000ah1n03x5 output195 (.a(net654),
    .o(cio_gpio_o[2]));
 b15bfn000ah1n03x5 output196 (.a(net650),
    .o(cio_gpio_o[30]));
 b15bfn000ah1n03x5 output197 (.a(net648),
    .o(cio_gpio_o[31]));
 b15bfn000ah1n03x5 output198 (.a(net652),
    .o(cio_gpio_o[3]));
 b15bfn000ah1n03x5 output199 (.a(net199),
    .o(cio_gpio_o[4]));
 b15bfn000ah1n03x5 output200 (.a(net2346),
    .o(cio_gpio_o[5]));
 b15bfn000ah1n03x5 output201 (.a(net201),
    .o(cio_gpio_o[6]));
 b15bfn000ah1n03x5 output202 (.a(net202),
    .o(cio_gpio_o[7]));
 b15bfn000ah1n03x5 output203 (.a(net203),
    .o(cio_gpio_o[8]));
 b15bfn000ah1n03x5 output204 (.a(net204),
    .o(cio_gpio_o[9]));
 b15bfn000ah1n03x5 output205 (.a(net2571),
    .o(net2004));
 b15bfn000ah1n03x5 output206 (.a(net2579),
    .o(net2022));
 b15bfn000ah1n03x5 output207 (.a(net2577),
    .o(net2016));
 b15bfn000ah1n03x5 output208 (.a(net2090),
    .o(net2091));
 b15bfn000ah1n03x5 output209 (.a(net2067),
    .o(net2068));
 b15bfn000ah1n03x5 output210 (.a(net2084),
    .o(net2085));
 b15bfn000ah1n03x5 output211 (.a(net2575),
    .o(net2010));
 b15bfn000ah1n03x5 output212 (.a(net2096),
    .o(net2097));
 b15bfn000ah1n03x5 output213 (.a(net2106),
    .o(net2107));
 b15bfn000ah1n03x5 output214 (.a(net2063),
    .o(net2064));
 b15bfn000ah1n03x5 output215 (.a(net2086),
    .o(net2087));
 b15bfn000ah1n03x5 output216 (.a(net2581),
    .o(net2018));
 b15bfn000ah1n03x5 output217 (.a(net2035),
    .o(net2036));
 b15bfn000ah1n03x5 output218 (.a(net2032),
    .o(net2033));
 b15bfn000ah1n03x5 output219 (.a(net2052),
    .o(net2053));
 b15bfn000ah1n03x5 output220 (.a(net2049),
    .o(net2051));
 b15bfn000ah1n03x5 output221 (.a(net2112),
    .o(net2113));
 b15bfn000ah1n03x5 output222 (.a(net2573),
    .o(net2006));
 b15bfn000ah1n03x5 output223 (.a(net2125),
    .o(net2126));
 b15bfn000ah1n03x5 output224 (.a(net2591),
    .o(net2048));
 b15bfn000ah1n03x5 output225 (.a(net2589),
    .o(net2046));
 b15bfn000ah1n03x5 output226 (.a(net2110),
    .o(net2111));
 b15bfn000ah1n03x5 output227 (.a(net2587),
    .o(net2024));
 b15bfn000ah1n03x5 output228 (.a(net2108),
    .o(net2109));
 b15bfn000ah1n03x5 output229 (.a(net2123),
    .o(net2124));
 b15bfn000ah1n03x5 output230 (.a(net2597),
    .o(net2066));
 b15bfn000ah1n03x5 output231 (.a(net2595),
    .o(net2062));
 b15bfn000ah1n03x5 output232 (.a(net2071),
    .o(net2072));
 b15bfn000ah1n03x5 output233 (.a(net2069),
    .o(net2070));
 b15bfn000ah1n03x5 output234 (.a(net2073),
    .o(net2074));
 b15bfn000ah1n03x5 output235 (.a(net2059),
    .o(net2060));
 b15bfn000ah1n03x5 output236 (.a(net2078),
    .o(net2079));
 b15bfn000ah1n03x5 output237 (.a(net2083),
    .o(tl_o[0]));
 b15bfn000ah1n03x5 output238 (.a(net2077),
    .o(tl_o[10]));
 b15bfn000ah1n03x5 output239 (.a(net2013),
    .o(net2014));
 b15bfn000ah1n03x5 output240 (.a(net2042),
    .o(net2043));
 b15bfn000ah1n03x5 output241 (.a(net2027),
    .o(tl_o[13]));
 b15bfn000ah1n03x5 output242 (.a(net242),
    .o(tl_o[14]));
 b15bfn000ah1n03x5 output243 (.a(net243),
    .o(tl_o[15]));
 b15bfn000ah1n03x5 output244 (.a(net509),
    .o(tl_o[16]));
 b15bfn000ah1n03x5 output245 (.a(net507),
    .o(tl_o[17]));
 b15bfn000ah1n03x5 output246 (.a(net2157),
    .o(net2158));
 b15bfn000ah1n03x5 output247 (.a(net2115),
    .o(net2116));
 b15bfn000ah1n03x5 output248 (.a(net2012),
    .o(net2000));
 b15bfn000ah1n03x5 output249 (.a(net468),
    .o(tl_o[20]));
 b15bfn000ah1n03x5 output250 (.a(net465),
    .o(tl_o[21]));
 b15bfn000ah1n03x5 output251 (.a(net2127),
    .o(net2128));
 b15bfn000ah1n03x5 output252 (.a(net2167),
    .o(net2168));
 b15bfn000ah1n03x5 output253 (.a(net2180),
    .o(net2181));
 b15bfn000ah1n03x5 output254 (.a(net459),
    .o(tl_o[25]));
 b15bfn000ah1n03x5 output255 (.a(net2145),
    .o(tl_o[26]));
 b15bfn000ah1n03x5 output256 (.a(net2139),
    .o(net2140));
 b15bfn000ah1n03x5 output257 (.a(net2146),
    .o(net2147));
 b15bfn000ah1n03x5 output258 (.a(net2141),
    .o(net2142));
 b15bfn000ah1n03x5 output259 (.a(net2293),
    .o(tl_o[2]));
 b15bfn000ah1n03x5 output260 (.a(net2129),
    .o(net2130));
 b15bfn000ah1n03x5 output261 (.a(net2134),
    .o(net2135));
 b15bfn000ah1n03x5 output262 (.a(net2205),
    .o(net2206));
 b15bfn000ah1n03x5 output263 (.a(net2292),
    .o(tl_o[33]));
 b15bfn000ah1n03x5 output264 (.a(net2182),
    .o(net2183));
 b15bfn000ah1n03x5 output265 (.a(net2257),
    .o(tl_o[35]));
 b15bfn000ah1n03x5 output266 (.a(net2308),
    .o(tl_o[36]));
 b15bfn000ah1n03x5 output267 (.a(net2131),
    .o(net2132));
 b15bfn000ah1n03x5 output268 (.a(net2278),
    .o(tl_o[38]));
 b15bfn000ah1n03x5 output269 (.a(net2136),
    .o(tl_o[39]));
 b15bfn000ah1n03x5 output270 (.a(net2179),
    .o(tl_o[3]));
 b15bfn000ah1n03x5 output271 (.a(net2148),
    .o(net2149));
 b15bfn000ah1n03x5 output272 (.a(net488),
    .o(tl_o[41]));
 b15bfn000ah1n03x5 output273 (.a(net486),
    .o(tl_o[42]));
 b15bfn000ah1n03x5 output274 (.a(net2191),
    .o(net2192));
 b15bfn000ah1n03x5 output275 (.a(net2175),
    .o(net2176));
 b15bfn000ah1n03x5 output276 (.a(net2150),
    .o(net2151));
 b15bfn000ah1n03x5 output277 (.a(net2276),
    .o(tl_o[46]));
 b15bfn000ah1n03x5 output278 (.a(net2220),
    .o(tl_o[47]));
 b15bfn000ah1n03x5 output279 (.a(net2102),
    .o(net2103));
 b15bfn000ah1n03x5 output280 (.a(net2277),
    .o(tl_o[4]));
 b15bfn000ah1n03x5 output281 (.a(net2100),
    .o(net2101));
 b15bfn000ah1n03x5 output282 (.a(net2117),
    .o(net2118));
 b15bfn000ah1n03x5 output283 (.a(net2119),
    .o(net2120));
 b15bfn000ah1n03x5 output284 (.a(net2098),
    .o(net2099));
 b15bfn000ah1n03x5 output285 (.a(net2104),
    .o(net2105));
 b15bfn000ah1n03x5 output286 (.a(net2094),
    .o(net2095));
 b15bfn000ah1n03x5 output287 (.a(net2092),
    .o(net2093));
 b15bfn000ah1n03x5 output288 (.a(net2076),
    .o(net2031));
 b15bfn000ah1n03x5 output289 (.a(net2026),
    .o(net2002));
 b15bfn000ah1n03x5 output290 (.a(net2202),
    .o(tl_o[5]));
 b15bfn000ah1n03x5 output291 (.a(net2088),
    .o(net2089));
 b15bfn000ah1n03x5 output292 (.a(net2055),
    .o(tl_o[63]));
 b15bfn000ah1n03x5 output293 (.a(net2041),
    .o(net2008));
 b15bfn000ah1n03x5 output294 (.a(net2082),
    .o(net2020));
 b15bfn000ah1n03x5 output295 (.a(net2138),
    .o(tl_o[6]));
 b15bfn000ah1n03x5 output296 (.a(net2185),
    .o(tl_o[7]));
 b15bfn000ah1n03x5 output297 (.a(net2217),
    .o(tl_o[8]));
 b15bfn000ah1n03x5 output298 (.a(net2058),
    .o(tl_o[9]));
 b15bfn000as1n24x5 wire299 (.a(n3445),
    .o(net299));
 b15bfn001as1n16x5 fanout300 (.a(n4130),
    .o(net300));
 b15bfn001ah1n24x5 fanout301 (.a(n4130),
    .o(net301));
 b15bfn001as1n64x5 fanout302 (.a(n3475),
    .o(net302));
 b15bfn001ah1n32x5 wire303 (.a(net305),
    .o(net303));
 b15bfn001as1n24x5 wire304 (.a(net305),
    .o(net304));
 b15bfn001as1n24x5 max_length305 (.a(net302),
    .o(net305));
 b15bfn001as1n16x5 wire306 (.a(N62),
    .o(net306));
 b15bfn001as1n16x5 wire307 (.a(N63),
    .o(net307));
 b15bfn001as1n48x5 fanout308 (.a(net312),
    .o(net308));
 b15bfn001ah1n32x5 max_length309 (.a(net310),
    .o(net309));
 b15bfn001as1n32x5 max_length310 (.a(net308),
    .o(net310));
 b15bfn001as1n64x5 fanout311 (.a(n3400),
    .o(net311));
 b15bfn001as1n32x5 max_length312 (.a(net313),
    .o(net312));
 b15bfn001as1n32x5 wire313 (.a(net311),
    .o(net313));
 b15bfn001as1n16x5 wire314 (.a(N55),
    .o(net314));
 b15bfn001as1n16x5 wire315 (.a(u_reg_u_reg_if_N23),
    .o(net315));
 b15bfn001ah1n24x5 wire316 (.a(u_reg_u_reg_if_N22),
    .o(net316));
 b15bfn001as1n24x5 wire317 (.a(u_reg_u_reg_if_N21),
    .o(net317));
 b15bfn001as1n24x5 wire318 (.a(u_reg_u_reg_if_N20),
    .o(net318));
 b15bfn001as1n48x5 fanout319 (.a(net322),
    .o(net319));
 b15bfn001as1n48x5 max_length320 (.a(net321),
    .o(net320));
 b15bfn001as1n32x5 wire321 (.a(net319),
    .o(net321));
 b15bfn001as1n64x5 fanout322 (.a(n3498),
    .o(net322));
 b15bfn001ah1n48x5 wire323 (.a(net322),
    .o(net323));
 b15bfn001ah1n24x5 wire324 (.a(n3498),
    .o(net324));
 b15bfn001as1n48x5 fanout325 (.a(n3431),
    .o(net325));
 b15bfn001ah1n24x5 wire326 (.a(net325),
    .o(net326));
 b15bfn001ah1n32x5 wire327 (.a(net328),
    .o(net327));
 b15bfn001as1n32x5 wire328 (.a(net325),
    .o(net328));
 b15bfn001as1n48x5 fanout329 (.a(n3389),
    .o(net329));
 b15bfn001as1n32x5 max_length330 (.a(net331),
    .o(net330));
 b15bfn001as1n24x5 wire331 (.a(net332),
    .o(net331));
 b15bfn001as1n32x5 wire332 (.a(net333),
    .o(net332));
 b15bfn001ah1n32x5 max_length333 (.a(net329),
    .o(net333));
 b15bfn001as1n16x5 wire334 (.a(n3389),
    .o(net334));
 b15bfn001as1n48x5 fanout335 (.a(net340),
    .o(net335));
 b15bfn000as1n24x5 wire336 (.a(net335),
    .o(net336));
 b15bfn001ah1n48x5 wire337 (.a(net338),
    .o(net337));
 b15bfn001ah1n48x5 wire338 (.a(net335),
    .o(net338));
 b15bfn001as1n64x5 fanout339 (.a(n3443),
    .o(net339));
 b15bfn001as1n48x5 max_length340 (.a(net343),
    .o(net340));
 b15bfn001as1n32x5 max_length341 (.a(net342),
    .o(net341));
 b15bfn001as1n24x5 wire342 (.a(net339),
    .o(net342));
 b15bfn001as1n32x5 max_length343 (.a(net339),
    .o(net343));
 b15bfn001ah1n32x5 fanout344 (.a(n3359),
    .o(net344));
 b15bfn000as1n24x5 fanout345 (.a(n3359),
    .o(net345));
 b15bfn001ah1n32x5 fanout346 (.a(net348),
    .o(net346));
 b15bfn001ah1n24x5 fanout347 (.a(net348),
    .o(net347));
 b15bfn001ah1n32x5 wire348 (.a(n3338),
    .o(net348));
 b15bfn000as1n24x5 fanout349 (.a(net350),
    .o(net349));
 b15bfn001ah1n32x5 fanout350 (.a(n3336),
    .o(net350));
 b15bfn001ah1n32x5 fanout351 (.a(net352),
    .o(net351));
 b15bfn001as1n32x5 fanout352 (.a(n3335),
    .o(net352));
 b15bfn001as1n32x5 fanout353 (.a(net354),
    .o(net353));
 b15bfn001as1n24x5 fanout354 (.a(n3334),
    .o(net354));
 b15bfn001as1n32x5 wire355 (.a(net354),
    .o(net355));
 b15bfn001ah1n24x5 wire356 (.a(n3334),
    .o(net356));
 b15bfn001ah1n32x5 fanout357 (.a(n3333),
    .o(net357));
 b15bfn001as1n24x5 fanout358 (.a(n3333),
    .o(net358));
 b15bfn001as1n32x5 fanout359 (.a(net362),
    .o(net359));
 b15bfn001ah1n48x5 max_length360 (.a(net361),
    .o(net360));
 b15bfn001aq1n48x5 wire361 (.a(net359),
    .o(net361));
 b15bfn001as1n48x5 fanout362 (.a(net366),
    .o(net362));
 b15bfn001as1n24x5 max_length363 (.a(net364),
    .o(net363));
 b15bfn001as1n32x5 max_length364 (.a(net365),
    .o(net364));
 b15bfn000as1n32x5 wire365 (.a(net362),
    .o(net365));
 b15bfn001as1n24x5 wire366 (.a(n3298),
    .o(net366));
 b15bfn001ah1n24x5 wire367 (.a(n3254),
    .o(net367));
 b15bfn001ah1n24x5 wire368 (.a(n3954),
    .o(net368));
 b15bfn001as1n16x5 wire369 (.a(n3983),
    .o(net369));
 b15bfn001as1n24x5 wire370 (.a(n3920),
    .o(net370));
 b15bfn001ah1n32x5 wire371 (.a(net372),
    .o(net371));
 b15bfn001as1n32x5 load_slew372 (.a(net374),
    .o(net372));
 b15bfn001ah1n48x5 load_slew373 (.a(n3872),
    .o(net373));
 b15bfn001as1n32x5 max_length374 (.a(n3872),
    .o(net374));
 b15bfn001ah1n24x5 wire375 (.a(u_reg_u_data_in_wr_data[22]),
    .o(net375));
 b15bfn001as1n24x5 wire376 (.a(u_reg_u_data_in_wr_data[20]),
    .o(net376));
 b15bfn001ah1n32x5 wire377 (.a(u_reg_u_data_in_wr_data[12]),
    .o(net377));
 b15bfn001as1n24x5 wire378 (.a(u_reg_u_data_in_wr_data[15]),
    .o(net378));
 b15bfn001ah1n24x5 wire379 (.a(u_reg_u_data_in_wr_data[3]),
    .o(net379));
 b15bfn001ah1n24x5 wire380 (.a(u_reg_u_data_in_wr_data[11]),
    .o(net380));
 b15bfn001as1n48x5 fanout381 (.a(net384),
    .o(net381));
 b15bfn001ah1n48x5 load_slew382 (.a(net383),
    .o(net382));
 b15bfn001ah1n48x5 wire383 (.a(net381),
    .o(net383));
 b15bfn001as1n64x5 fanout384 (.a(n3295),
    .o(net384));
 b15bfn001as1n32x5 wire385 (.a(net384),
    .o(net385));
 b15bfn001as1n32x5 wire386 (.a(net384),
    .o(net386));
 b15bfn001as1n24x5 wire387 (.a(net384),
    .o(net387));
 b15bfn001as1n64x5 fanout388 (.a(net394),
    .o(net388));
 b15bfn001ah1n24x5 wire389 (.a(net388),
    .o(net389));
 b15bfn001as1n32x5 max_length390 (.a(net388),
    .o(net390));
 b15bfn001as1n48x5 fanout391 (.a(net394),
    .o(net391));
 b15bfn001ah1n32x5 max_length392 (.a(net393),
    .o(net392));
 b15bfn001as1n32x5 max_length393 (.a(net391),
    .o(net393));
 b15bfn001ah1n80x5 fanout394 (.a(n3290),
    .o(net394));
 b15bfn001as1n80x5 fanout395 (.a(net397),
    .o(net395));
 b15bfn001as1n64x5 fanout396 (.a(n3289),
    .o(net396));
 b15bfn001ah1n32x5 max_length397 (.a(net396),
    .o(net397));
 b15bfn001aq1n48x5 wire398 (.a(net399),
    .o(net398));
 b15bfn001as1n32x5 wire399 (.a(net396),
    .o(net399));
 b15bfn001as1n64x5 fanout400 (.a(net403),
    .o(net400));
 b15bfn001ah1n48x5 max_length401 (.a(net402),
    .o(net401));
 b15bfn001ah1n48x5 wire402 (.a(net400),
    .o(net402));
 b15bfn001as1n64x5 fanout403 (.a(n3288),
    .o(net403));
 b15bfn001ah1n48x5 max_length404 (.a(net405),
    .o(net404));
 b15bfn001as1n32x5 wire405 (.a(net403),
    .o(net405));
 b15bfn001as1n32x5 wire406 (.a(n3288),
    .o(net406));
 b15bfn001ah1n24x5 wire407 (.a(n3017),
    .o(net407));
 b15bfn001ah1n32x5 wire408 (.a(u_reg_u_reg_if_a_ack),
    .o(net408));
 b15bfn001as1n24x5 max_length409 (.a(u_reg_u_reg_if_a_ack),
    .o(net409));
 b15bfn001as1n64x5 fanout410 (.a(n3877),
    .o(net410));
 b15bfn001as1n32x5 max_length411 (.a(net412),
    .o(net411));
 b15bfn001ah1n48x5 load_slew412 (.a(net413),
    .o(net412));
 b15bfn001ah1n48x5 wire413 (.a(net410),
    .o(net413));
 b15bfn001as1n64x5 fanout414 (.a(n3871),
    .o(net414));
 b15bfn001ah1n48x5 max_length415 (.a(net417),
    .o(net415));
 b15bfn001ah1n48x5 max_length416 (.a(net417),
    .o(net416));
 b15bfn001ah1n48x5 wire417 (.a(net414),
    .o(net417));
 b15bfn001as1n64x5 fanout418 (.a(n3870),
    .o(net418));
 b15bfn001ah1n48x5 wire419 (.a(net420),
    .o(net419));
 b15bfn001ah1n48x5 wire420 (.a(net418),
    .o(net420));
 b15bfn001as1n24x5 wire421 (.a(net418),
    .o(net421));
 b15bfn001ah1n48x5 load_slew422 (.a(net418),
    .o(net422));
 b15bfn001as1n64x5 fanout423 (.a(n3303),
    .o(net423));
 b15bfn001as1n24x5 max_length424 (.a(net423),
    .o(net424));
 b15bfn001ah1n32x5 max_length425 (.a(net423),
    .o(net425));
 b15bfn001ah1n48x5 max_length426 (.a(net423),
    .o(net426));
 b15bfn001as1n64x5 fanout427 (.a(n3303),
    .o(net427));
 b15bfn001ah1n48x5 wire428 (.a(net429),
    .o(net428));
 b15bfn001ah1n32x5 max_length429 (.a(net427),
    .o(net429));
 b15bfn001ah1n80x5 fanout430 (.a(net432),
    .o(net430));
 b15bfn001as1n64x5 fanout431 (.a(n3301),
    .o(net431));
 b15bfn001ah1n48x5 wire432 (.a(net431),
    .o(net432));
 b15bfn001as1n24x5 max_length433 (.a(net434),
    .o(net433));
 b15bfn001as1n24x5 max_length434 (.a(net431),
    .o(net434));
 b15bfn001as1n64x5 fanout435 (.a(n3953),
    .o(net435));
 b15bfn001as1n16x5 max_length436 (.a(net438),
    .o(net436));
 b15bfn001as1n32x5 max_length437 (.a(net438),
    .o(net437));
 b15bfn001as1n32x5 wire438 (.a(net435),
    .o(net438));
 b15bfn001as1n48x5 max_length439 (.a(net435),
    .o(net439));
 b15bfn001as1n64x5 fanout440 (.a(n3981),
    .o(net440));
 b15bfn001ah1n32x5 max_length441 (.a(net444),
    .o(net441));
 b15bfn001ah1n32x5 max_length442 (.a(net444),
    .o(net442));
 b15bfn001ah1n48x5 wire443 (.a(net444),
    .o(net443));
 b15bfn001ah1n48x5 wire444 (.a(net440),
    .o(net444));
 b15bfn000as1n32x5 wire445 (.a(n3982),
    .o(net445));
 b15bfn001ah1n48x5 wire446 (.a(n3982),
    .o(net446));
 b15bfn001as1n32x5 max_length447 (.a(net448),
    .o(net447));
 b15bfn001as1n32x5 wire448 (.a(n3982),
    .o(net448));
 b15bfn001as1n48x5 fanout449 (.a(net452),
    .o(net449));
 b15bfn001as1n32x5 max_length450 (.a(net451),
    .o(net450));
 b15bfn001ah1n48x5 max_length451 (.a(net449),
    .o(net451));
 b15bfn001as1n48x5 fanout452 (.a(n3292),
    .o(net452));
 b15bfn001ah1n48x5 max_length453 (.a(net454),
    .o(net453));
 b15bfn001ah1n48x5 max_length454 (.a(net455),
    .o(net454));
 b15bfn001as1n32x5 wire455 (.a(net452),
    .o(net455));
 b15bfn000as1n32x5 wire456 (.a(n3007),
    .o(net456));
 b15bfn001ah1n32x5 wire457 (.a(n3029),
    .o(net457));
 b15bfn001ah1n32x5 wire458 (.a(n3000),
    .o(net458));
 b15bfn001as1n08x5 load_slew459 (.a(net460),
    .o(net459));
 b15bfn001as1n24x5 wire460 (.a(net2155),
    .o(net460));
 b15bfn001as1n12x5 wire461 (.a(net2154),
    .o(net461));
 b15bfn001as1n12x5 max_cap462 (.a(net463),
    .o(net462));
 b15bfn001ah1n12x5 load_slew463 (.a(net2166),
    .o(net463));
 b15bfn001ah1n16x5 wire464 (.a(net2127),
    .o(net464));
 b15bfn001ah1n12x5 wire465 (.a(net466),
    .o(net465));
 b15bfn001as1n24x5 wire466 (.a(net2165),
    .o(net466));
 b15bfn001as1n12x5 wire467 (.a(net2164),
    .o(net467));
 b15bfn001as1n12x5 wire468 (.a(net469),
    .o(net468));
 b15bfn001as1n24x5 wire469 (.a(net470),
    .o(net469));
 b15bfn001as1n12x5 wire470 (.a(net2177),
    .o(net470));
 b15bfn001ah1n12x5 wire471 (.a(net472),
    .o(net471));
 b15bfn001as1n16x5 wire472 (.a(net278),
    .o(net472));
 b15bfn001as1n08x5 load_slew473 (.a(net2115),
    .o(net473));
 b15bfn001as1n12x5 max_cap474 (.a(net475),
    .o(net474));
 b15bfn001ah1n12x5 wire475 (.a(net2114),
    .o(net475));
 b15bfn001ah1n12x5 load_slew476 (.a(net477),
    .o(net476));
 b15bfn001as1n12x5 max_cap477 (.a(net2156),
    .o(net477));
 b15bfn001as1n24x5 wire478 (.a(net479),
    .o(net478));
 b15bfn001as1n12x5 wire479 (.a(net276),
    .o(net479));
 b15bfn001ah1n24x5 wire480 (.a(net481),
    .o(net480));
 b15bfn001ah1n12x5 load_slew481 (.a(net482),
    .o(net481));
 b15bfn001ah1n12x5 load_slew482 (.a(net2175),
    .o(net482));
 b15bfn001ah1n12x5 load_slew483 (.a(net484),
    .o(net483));
 b15bfn001ah1n16x5 wire484 (.a(net274),
    .o(net484));
 b15bfn001ah1n24x5 wire485 (.a(net273),
    .o(net485));
 b15bfn001ah1n12x5 wire486 (.a(net487),
    .o(net486));
 b15bfn001ah1n16x5 max_cap487 (.a(net2312),
    .o(net487));
 b15bfn001ah1n12x5 load_slew488 (.a(net489),
    .o(net488));
 b15bfn001ah1n12x5 load_slew489 (.a(net2218),
    .o(net489));
 b15bfn001as1n12x5 wire490 (.a(net491),
    .o(net490));
 b15bfn001as1n12x5 wire491 (.a(net2148),
    .o(net491));
 b15bfn001as1n24x5 wire492 (.a(net493),
    .o(net492));
 b15bfn001as1n12x5 wire493 (.a(net494),
    .o(net493));
 b15bfn001ah1n12x5 wire494 (.a(net2131),
    .o(net494));
 b15bfn001ah1n16x5 max_cap495 (.a(net264),
    .o(net495));
 b15bfn001as1n12x5 max_cap496 (.a(net262),
    .o(net496));
 b15bfn001as1n12x5 max_cap497 (.a(net2133),
    .o(net497));
 b15bfn001ah1n12x5 load_slew498 (.a(net2129),
    .o(net498));
 b15bfn001as1n16x5 wire499 (.a(net500),
    .o(net499));
 b15bfn001as1n08x5 load_slew500 (.a(net2141),
    .o(net500));
 b15bfn001as1n12x5 max_cap501 (.a(net258),
    .o(net501));
 b15bfn001ah1n12x5 wire502 (.a(net2146),
    .o(net502));
 b15bfn001ah1n12x5 load_slew503 (.a(net257),
    .o(net503));
 b15bfn001as1n16x5 wire504 (.a(net2139),
    .o(net504));
 b15bfn001ah1n16x5 max_cap505 (.a(net2144),
    .o(net505));
 b15bfn001ah1n12x5 load_slew506 (.a(net2143),
    .o(net506));
 b15bfn001ah1n32x5 wire507 (.a(net508),
    .o(net507));
 b15bfn001ah1n16x5 wire508 (.a(net2214),
    .o(net508));
 b15bfn001ah1n12x5 load_slew509 (.a(net510),
    .o(net509));
 b15bfn001ah1n12x5 wire510 (.a(net2275),
    .o(net510));
 b15bfn001ah1n24x5 wire511 (.a(net2274),
    .o(net511));
 b15bfn001as1n16x5 wire512 (.a(reg2hw_intr_state__q__7_),
    .o(net512));
 b15bfn001ah1n12x5 wire513 (.a(net514),
    .o(net513));
 b15bfn001as1n08x5 load_slew514 (.a(net2466),
    .o(net514));
 b15bfn001ah1n24x5 wire515 (.a(net516),
    .o(net515));
 b15bfn001ah1n12x5 load_slew516 (.a(net517),
    .o(net516));
 b15bfn001ah1n12x5 load_slew517 (.a(net2638),
    .o(net517));
 b15bfn001ah1n16x5 wire518 (.a(net519),
    .o(net518));
 b15bfn001ah1n16x5 wire519 (.a(reg2hw_intr_state__q__4_),
    .o(net519));
 b15bfn001ah1n12x5 wire520 (.a(reg2hw_intr_state__q__3_),
    .o(net520));
 b15bfn001ah1n12x5 wire521 (.a(reg2hw_intr_state__q__2_),
    .o(net521));
 b15bfn001as1n16x5 wire522 (.a(net523),
    .o(net522));
 b15bfn001ah1n08x5 load_slew523 (.a(reg2hw_intr_state__q__11_),
    .o(net523));
 b15bfn001as1n12x5 wire524 (.a(reg2hw_intr_state__q__1_),
    .o(net524));
 b15bfn001as1n16x5 wire525 (.a(net526),
    .o(net525));
 b15bfn001as1n16x5 wire526 (.a(reg2hw_intr_state__q__0_),
    .o(net526));
 b15bfn001as1n16x5 wire527 (.a(net528),
    .o(net527));
 b15bfn001as1n06x5 load_slew528 (.a(reg2hw_intr_enable__q__3_),
    .o(net528));
 b15bfn001ah1n12x5 wire529 (.a(reg2hw_intr_enable__q__2_),
    .o(net529));
 b15bfn001ah1n16x5 wire530 (.a(reg2hw_intr_enable__q__25_),
    .o(net530));
 b15bfn001ah1n08x5 load_slew531 (.a(reg2hw_intr_enable__q__25_),
    .o(net531));
 b15bfn001ah1n16x5 wire532 (.a(reg2hw_intr_enable__q__22_),
    .o(net532));
 b15bfn001ah1n24x5 wire533 (.a(reg2hw_intr_enable__q__21_),
    .o(net533));
 b15bfn001as1n16x5 wire534 (.a(reg2hw_intr_enable__q__20_),
    .o(net534));
 b15bfn001ah1n16x5 wire535 (.a(reg2hw_intr_enable__q__18_),
    .o(net535));
 b15bfn001ah1n16x5 wire536 (.a(net2520),
    .o(net536));
 b15bfn001as1n16x5 wire537 (.a(net2339),
    .o(net537));
 b15bfn001ah1n12x5 load_slew538 (.a(reg2hw_intr_enable__q__10_),
    .o(net538));
 b15bfn001ah1n24x5 wire539 (.a(net540),
    .o(net539));
 b15bfn001ah1n12x5 load_slew540 (.a(net541),
    .o(net540));
 b15bfn001as1n12x5 wire541 (.a(net2562),
    .o(net541));
 b15bfn001as1n16x5 wire542 (.a(reg2hw_intr_enable__q__0_),
    .o(net542));
 b15bfn001as1n12x5 wire543 (.a(reg2hw_intr_ctrl_en_rising__q__8_),
    .o(net543));
 b15bfn001ah1n16x5 max_cap544 (.a(reg2hw_intr_ctrl_en_rising__q__7_),
    .o(net544));
 b15bfn001ah1n16x5 max_cap545 (.a(reg2hw_intr_ctrl_en_rising__q__4_),
    .o(net545));
 b15bfn001as1n12x5 max_cap546 (.a(net547),
    .o(net546));
 b15bfn001as1n12x5 wire547 (.a(net2542),
    .o(net547));
 b15bfn001as1n16x5 wire548 (.a(reg2hw_intr_ctrl_en_rising__q__2_),
    .o(net548));
 b15bfn001ah1n16x5 wire549 (.a(reg2hw_intr_ctrl_en_rising__q__25_),
    .o(net549));
 b15bfn001as1n16x5 wire550 (.a(reg2hw_intr_ctrl_en_rising__q__17_),
    .o(net550));
 b15bfn001ah1n16x5 wire551 (.a(reg2hw_intr_ctrl_en_rising__q__16_),
    .o(net551));
 b15bfn001as1n16x5 wire552 (.a(reg2hw_intr_ctrl_en_lvllow__q__9_),
    .o(net552));
 b15bfn001ah1n16x5 wire553 (.a(reg2hw_intr_ctrl_en_lvllow__q__8_),
    .o(net553));
 b15bfn001as1n08x5 load_slew554 (.a(reg2hw_intr_ctrl_en_lvllow__q__2_),
    .o(net554));
 b15bfn001ah1n16x5 wire555 (.a(reg2hw_intr_ctrl_en_lvllow__q__25_),
    .o(net555));
 b15bfn001ah1n16x5 wire556 (.a(reg2hw_intr_ctrl_en_lvllow__q__24_),
    .o(net556));
 b15bfn001ah1n12x5 load_slew557 (.a(reg2hw_intr_ctrl_en_lvllow__q__13_),
    .o(net557));
 b15bfn001ah1n24x5 wire558 (.a(reg2hw_intr_ctrl_en_lvllow__q__1_),
    .o(net558));
 b15bfn001ah1n16x5 wire559 (.a(net560),
    .o(net559));
 b15bfn001ah1n24x5 wire560 (.a(reg2hw_intr_ctrl_en_lvllow__q__0_),
    .o(net560));
 b15bfn001ah1n16x5 wire561 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__9_),
    .o(net561));
 b15bfn001ah1n16x5 wire562 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__8_),
    .o(net562));
 b15bfn001as1n16x5 wire563 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__7_),
    .o(net563));
 b15bfn001as1n16x5 wire564 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__6_),
    .o(net564));
 b15bfn001ah1n16x5 wire565 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__3_),
    .o(net565));
 b15bfn001as1n08x5 load_slew566 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__3_),
    .o(net566));
 b15bfn001ah1n16x5 wire567 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__27_),
    .o(net567));
 b15bfn001as1n16x5 wire568 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__25_),
    .o(net568));
 b15bfn001ah1n16x5 wire569 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__24_),
    .o(net569));
 b15bfn001as1n16x5 wire570 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__17_),
    .o(net570));
 b15bfn001as1n16x5 wire571 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__16_),
    .o(net571));
 b15bfn001ah1n16x5 wire572 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__12_),
    .o(net572));
 b15bfn001as1n16x5 wire573 (.a(net574),
    .o(net573));
 b15bfn001ah1n12x5 wire574 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__10_),
    .o(net574));
 b15bfn001ah1n12x5 wire575 (.a(net576),
    .o(net575));
 b15bfn001as1n16x5 wire576 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__1_),
    .o(net576));
 b15bfn001as1n24x5 wire577 (.a(net578),
    .o(net577));
 b15bfn001as1n12x5 wire578 (.a(net579),
    .o(net578));
 b15bfn001as1n16x5 wire579 (.a(reg2hw_intr_ctrl_en_lvlhigh__q__0_),
    .o(net579));
 b15bfn001ah1n16x5 wire580 (.a(reg2hw_intr_ctrl_en_falling__q__9_),
    .o(net580));
 b15bfn001as1n08x5 load_slew581 (.a(reg2hw_intr_ctrl_en_falling__q__5_),
    .o(net581));
 b15bfn001ah1n08x5 load_slew582 (.a(reg2hw_intr_ctrl_en_falling__q__28_),
    .o(net582));
 b15bfn001ah1n12x5 wire583 (.a(net584),
    .o(net583));
 b15bfn001ah1n12x5 wire584 (.a(reg2hw_intr_ctrl_en_falling__q__27_),
    .o(net584));
 b15bfn001ah1n16x5 wire585 (.a(reg2hw_intr_ctrl_en_falling__q__26_),
    .o(net585));
 b15bfn001ah1n12x5 load_slew586 (.a(reg2hw_intr_ctrl_en_falling__q__26_),
    .o(net586));
 b15bfn001as1n24x5 wire587 (.a(net588),
    .o(net587));
 b15bfn001as1n12x5 wire588 (.a(reg2hw_intr_ctrl_en_falling__q__25_),
    .o(net588));
 b15bfn001as1n16x5 wire589 (.a(reg2hw_intr_ctrl_en_falling__q__19_),
    .o(net589));
 b15bfn001as1n16x5 wire590 (.a(reg2hw_intr_ctrl_en_falling__q__18_),
    .o(net590));
 b15bfn001ah1n12x5 wire591 (.a(reg2hw_intr_ctrl_en_falling__q__10_),
    .o(net591));
 b15bfn001ah1n24x5 wire592 (.a(net593),
    .o(net592));
 b15bfn001ah1n12x5 wire593 (.a(reg2hw_intr_ctrl_en_falling__q__1_),
    .o(net593));
 b15bfn001as1n16x5 wire594 (.a(reg2hw_intr_ctrl_en_falling__q__0_),
    .o(net594));
 b15bfn001as1n12x5 wire595 (.a(reg2hw_ctrl_en_input_filter__q__9_),
    .o(net595));
 b15bfn001as1n08x5 load_slew596 (.a(net597),
    .o(net596));
 b15bfn001as1n12x5 wire597 (.a(net2498),
    .o(net597));
 b15bfn001as1n12x5 wire598 (.a(reg2hw_ctrl_en_input_filter__q__7_),
    .o(net598));
 b15bfn001as1n12x5 max_cap599 (.a(net600),
    .o(net599));
 b15bfn001ah1n16x5 wire600 (.a(net2565),
    .o(net600));
 b15bfn001ah1n12x5 wire601 (.a(reg2hw_ctrl_en_input_filter__q__5_),
    .o(net601));
 b15bfn001ah1n12x5 load_slew602 (.a(reg2hw_ctrl_en_input_filter__q__5_),
    .o(net602));
 b15bfn001ah1n24x5 wire603 (.a(net605),
    .o(net603));
 b15bfn001ah1n16x5 wire604 (.a(reg2hw_ctrl_en_input_filter__q__4_),
    .o(net604));
 b15bfn001ah1n12x5 load_slew605 (.a(reg2hw_ctrl_en_input_filter__q__4_),
    .o(net605));
 b15bfn001as1n08x5 load_slew606 (.a(reg2hw_ctrl_en_input_filter__q__31_),
    .o(net606));
 b15bfn001ah1n16x5 wire607 (.a(reg2hw_ctrl_en_input_filter__q__30_),
    .o(net607));
 b15bfn001as1n08x5 load_slew608 (.a(reg2hw_ctrl_en_input_filter__q__30_),
    .o(net608));
 b15bfn000as1n32x5 wire609 (.a(net610),
    .o(net609));
 b15bfn001as1n16x5 wire610 (.a(net611),
    .o(net610));
 b15bfn001ah1n12x5 wire611 (.a(reg2hw_ctrl_en_input_filter__q__3_),
    .o(net611));
 b15bfn001ah1n16x5 wire612 (.a(reg2hw_ctrl_en_input_filter__q__2_),
    .o(net612));
 b15bfn001ah1n12x5 load_slew613 (.a(reg2hw_ctrl_en_input_filter__q__2_),
    .o(net613));
 b15bfn001ah1n12x5 load_slew614 (.a(net615),
    .o(net614));
 b15bfn001ah1n16x5 wire615 (.a(reg2hw_ctrl_en_input_filter__q__29_),
    .o(net615));
 b15bfn001ah1n16x5 wire616 (.a(net617),
    .o(net616));
 b15bfn001as1n12x5 wire617 (.a(reg2hw_ctrl_en_input_filter__q__28_),
    .o(net617));
 b15bfn001as1n08x5 load_slew618 (.a(reg2hw_ctrl_en_input_filter__q__27_),
    .o(net618));
 b15bfn001as1n12x5 wire619 (.a(net620),
    .o(net619));
 b15bfn001as1n12x5 wire620 (.a(reg2hw_ctrl_en_input_filter__q__23_),
    .o(net620));
 b15bfn001as1n16x5 wire621 (.a(net622),
    .o(net621));
 b15bfn001ah1n12x5 wire622 (.a(reg2hw_ctrl_en_input_filter__q__22_),
    .o(net622));
 b15bfn001ah1n12x5 load_slew623 (.a(net624),
    .o(net623));
 b15bfn001as1n16x5 wire624 (.a(reg2hw_ctrl_en_input_filter__q__21_),
    .o(net624));
 b15bfn001ah1n12x5 wire625 (.a(net626),
    .o(net625));
 b15bfn001ah1n12x5 wire626 (.a(reg2hw_ctrl_en_input_filter__q__20_),
    .o(net626));
 b15bfn001as1n08x5 load_slew627 (.a(net628),
    .o(net627));
 b15bfn001ah1n12x5 wire628 (.a(reg2hw_ctrl_en_input_filter__q__19_),
    .o(net628));
 b15bfn001as1n16x5 wire629 (.a(reg2hw_ctrl_en_input_filter__q__18_),
    .o(net629));
 b15bfn001ah1n16x5 wire630 (.a(reg2hw_ctrl_en_input_filter__q__15_),
    .o(net630));
 b15bfn001ah1n12x5 load_slew631 (.a(reg2hw_ctrl_en_input_filter__q__15_),
    .o(net631));
 b15bfn001as1n12x5 wire632 (.a(net633),
    .o(net632));
 b15bfn001ah1n16x5 wire633 (.a(reg2hw_ctrl_en_input_filter__q__14_),
    .o(net633));
 b15bfn001as1n12x5 wire634 (.a(net635),
    .o(net634));
 b15bfn001ah1n12x5 wire635 (.a(reg2hw_ctrl_en_input_filter__q__13_),
    .o(net635));
 b15bfn001ah1n24x5 wire636 (.a(net637),
    .o(net636));
 b15bfn001ah1n12x5 load_slew637 (.a(reg2hw_ctrl_en_input_filter__q__12_),
    .o(net637));
 b15bfn001ah1n16x5 wire638 (.a(reg2hw_ctrl_en_input_filter__q__11_),
    .o(net638));
 b15bfn001as1n12x5 wire639 (.a(reg2hw_ctrl_en_input_filter__q__10_),
    .o(net639));
 b15bfn001as1n12x5 wire640 (.a(reg2hw_ctrl_en_input_filter__q__10_),
    .o(net640));
 b15bfn001as1n16x5 wire641 (.a(net642),
    .o(net641));
 b15bfn001ah1n12x5 wire642 (.a(reg2hw_ctrl_en_input_filter__q__1_),
    .o(net642));
 b15bfn001ah1n12x5 load_slew643 (.a(net204),
    .o(net643));
 b15bfn001as1n12x5 max_cap644 (.a(net203),
    .o(net644));
 b15bfn001ah1n16x5 wire645 (.a(net646),
    .o(net645));
 b15bfn001ah1n24x5 wire646 (.a(net647),
    .o(net646));
 b15bfn001as1n08x5 wire647 (.a(net200),
    .o(net647));
 b15bfn001as1n08x5 load_slew648 (.a(net649),
    .o(net648));
 b15bfn001ah1n16x5 wire649 (.a(net197),
    .o(net649));
 b15bfn001as1n12x5 wire650 (.a(net651),
    .o(net650));
 b15bfn001as1n08x5 load_slew651 (.a(net196),
    .o(net651));
 b15bfn001ah1n12x5 wire652 (.a(net653),
    .o(net652));
 b15bfn001as1n12x5 wire653 (.a(net198),
    .o(net653));
 b15bfn001ah1n12x5 wire654 (.a(net655),
    .o(net654));
 b15bfn001as1n12x5 wire655 (.a(net195),
    .o(net655));
 b15bfn001as1n24x5 wire656 (.a(net657),
    .o(net656));
 b15bfn001as1n12x5 wire657 (.a(net194),
    .o(net657));
 b15bfn001as1n08x5 wire658 (.a(net659),
    .o(net658));
 b15bfn001ah1n12x5 load_slew659 (.a(net193),
    .o(net659));
 b15bfn001as1n12x5 max_cap660 (.a(net661),
    .o(net660));
 b15bfn001ah1n12x5 load_slew661 (.a(net662),
    .o(net661));
 b15bfn001as1n12x5 max_cap662 (.a(net663),
    .o(net662));
 b15bfn001as1n16x5 wire663 (.a(net192),
    .o(net663));
 b15bfn001ah1n12x5 wire664 (.a(net665),
    .o(net664));
 b15bfn001ah1n12x5 load_slew665 (.a(net666),
    .o(net665));
 b15bfn001ah1n16x5 wire666 (.a(net191),
    .o(net666));
 b15bfn001as1n12x5 load_slew667 (.a(net668),
    .o(net667));
 b15bfn001ah1n12x5 wire668 (.a(net190),
    .o(net668));
 b15bfn001ah1n12x5 wire669 (.a(net670),
    .o(net669));
 b15bfn001ah1n12x5 load_slew670 (.a(net189),
    .o(net670));
 b15bfn001ah1n16x5 max_cap671 (.a(net189),
    .o(net671));
 b15bfn001ah1n12x5 wire672 (.a(net673),
    .o(net672));
 b15bfn001ah1n08x5 load_slew673 (.a(net674),
    .o(net673));
 b15bfn001as1n24x5 wire674 (.a(net675),
    .o(net674));
 b15bfn001as1n12x5 wire675 (.a(net188),
    .o(net675));
 b15bfn001as1n08x5 wire676 (.a(net678),
    .o(net676));
 b15bfn001as1n12x5 wire677 (.a(net678),
    .o(net677));
 b15bfn001as1n24x5 wire678 (.a(net679),
    .o(net678));
 b15bfn001as1n12x5 wire679 (.a(net187),
    .o(net679));
 b15bfn001as1n12x5 wire680 (.a(net681),
    .o(net680));
 b15bfn001as1n08x5 wire681 (.a(net182),
    .o(net681));
 b15bfn001ah1n16x5 wire682 (.a(net683),
    .o(net682));
 b15bfn001ah1n12x5 wire683 (.a(net181),
    .o(net683));
 b15bfn001as1n12x5 wire684 (.a(net685),
    .o(net684));
 b15bfn001ah1n12x5 wire685 (.a(net2302),
    .o(net685));
 b15bfn001as1n16x5 wire686 (.a(net687),
    .o(net686));
 b15bfn001ah1n12x5 wire687 (.a(net179),
    .o(net687));
 b15bfn001ah1n12x5 load_slew688 (.a(net178),
    .o(net688));
 b15bfn001ah1n08x5 load_slew689 (.a(net176),
    .o(net689));
 b15bfn001as1n08x5 load_slew690 (.a(net691),
    .o(net690));
 b15bfn001as1n08x5 load_slew691 (.a(net174),
    .o(net691));
 b15bfn001ah1n12x5 load_slew692 (.a(net693),
    .o(net692));
 b15bfn001ah1n12x5 wire693 (.a(net2249),
    .o(net693));
 b15bfn001as1n16x5 wire694 (.a(net2248),
    .o(net694));
 b15bfn001ah1n16x5 max_cap695 (.a(net2221),
    .o(net695));
 b15bfn001as1n16x5 wire696 (.a(net167),
    .o(net696));
 b15bfn001ah1n08x5 load_slew697 (.a(net698),
    .o(net697));
 b15bfn001ah1n16x5 wire698 (.a(net2316),
    .o(net698));
 b15bfn001as1n08x5 wire699 (.a(net2250),
    .o(net699));
 b15bfn001as1n12x5 max_cap700 (.a(net2251),
    .o(net700));
 b15bfn001as1n16x5 wire701 (.a(net2304),
    .o(net701));
 b15bfn001as1n16x5 wire702 (.a(net2233),
    .o(net702));
 b15bfn001ah1n12x5 load_slew703 (.a(net2232),
    .o(net703));
 b15bfn001ah1n32x5 wire704 (.a(net705),
    .o(net704));
 b15bfn001as1n16x5 wire705 (.a(net2548),
    .o(net705));
 b15bfn001as1n12x5 wire706 (.a(net707),
    .o(net706));
 b15bfn001as1n16x5 wire707 (.a(net2226),
    .o(net707));
 b15bfn001as1n12x5 wire708 (.a(net158),
    .o(net708));
 b15bfn001as1n16x5 wire709 (.a(net2208),
    .o(net709));
 b15bfn001ah1n12x5 load_slew710 (.a(net2207),
    .o(net710));
 b15bfn001ah1n12x5 load_slew711 (.a(net712),
    .o(net711));
 b15bfn001ah1n12x5 load_slew712 (.a(net156),
    .o(net712));
 b15bfn000as1n12x5 wire713 (.a(net2231),
    .o(net713));
 b15bfn001ah1n16x5 wire714 (.a(net151),
    .o(net714));
 b15bfn001as1n16x5 wire715 (.a(net2210),
    .o(net715));
 b15bfn001ah1n12x5 load_slew716 (.a(net2209),
    .o(net716));
 b15bfn001as1n16x5 wire717 (.a(net719),
    .o(net717));
 b15bfn001ah1n12x5 load_slew718 (.a(net150),
    .o(net718));
 b15bfn001as1n08x5 load_slew719 (.a(net2228),
    .o(net719));
 b15bfn001ah1n12x5 load_slew720 (.a(net721),
    .o(net720));
 b15bfn001ah1n12x5 wire721 (.a(net2297),
    .o(net721));
 b15bfn001as1n12x5 wire722 (.a(net723),
    .o(net722));
 b15bfn001ah1n12x5 load_slew723 (.a(net2311),
    .o(net723));
 b15bfn001as1n08x5 load_slew724 (.a(net725),
    .o(net724));
 b15bfn001ah1n24x5 wire725 (.a(net2234),
    .o(net725));
 b15bfn001ah1n12x5 load_slew726 (.a(net727),
    .o(net726));
 b15bfn001ah1n24x5 wire727 (.a(net2224),
    .o(net727));
 b15bfn001as1n12x5 max_cap728 (.a(net145),
    .o(net728));
 b15bfn001as1n08x5 load_slew729 (.a(net730),
    .o(net729));
 b15bfn001as1n08x5 wire730 (.a(net2173),
    .o(net730));
 b15bfn001ah1n12x5 load_slew731 (.a(net152),
    .o(net731));
 b15bfn001ah1n24x5 wire732 (.a(n3454),
    .o(net732));
 b15bfn001ah1n32x5 wire733 (.a(n3444),
    .o(net733));
 b15bfn001ah1n24x5 wire734 (.a(n3464),
    .o(net734));
 b15bfn001ah1n24x5 wire735 (.a(n3448),
    .o(net735));
 b15bfn001ah1n24x5 wire736 (.a(n3462),
    .o(net736));
 b15bfn001ah1n12x5 load_slew737 (.a(net2054),
    .o(net737));
 b15bfn001ah1n16x5 wire738 (.a(net2445),
    .o(net738));
 b15bfn001ah1n16x5 wire739 (.a(net2422),
    .o(net739));
 b15bfn001as1n12x5 wire740 (.a(net2456),
    .o(net740));
 b15bfn001ah1n16x5 wire741 (.a(gen_filter_5__u_filter_filter_synced),
    .o(net741));
 b15bfn001as1n08x5 wire742 (.a(gen_filter_5__u_filter_filter_synced),
    .o(net742));
 b15bfn001ah1n12x5 load_slew743 (.a(gen_filter_4__u_filter_filter_synced),
    .o(net743));
 b15bfn001as1n08x5 load_slew744 (.a(net745),
    .o(net744));
 b15bfn001as1n12x5 wire745 (.a(gen_filter_3__u_filter_filter_synced),
    .o(net745));
 b15bfn001as1n12x5 wire746 (.a(gen_filter_31__u_filter_filter_synced),
    .o(net746));
 b15bfn001as1n16x5 wire747 (.a(net2362),
    .o(net747));
 b15bfn001as1n16x5 wire748 (.a(gen_filter_25__u_filter_filter_synced),
    .o(net748));
 b15bfn001as1n08x5 load_slew749 (.a(net750),
    .o(net749));
 b15bfn001ah1n12x5 wire750 (.a(net751),
    .o(net750));
 b15bfn001ah1n16x5 wire751 (.a(gen_filter_23__u_filter_filter_synced),
    .o(net751));
 b15bfn001ah1n12x5 load_slew752 (.a(net753),
    .o(net752));
 b15bfn001ah1n06x5 load_slew753 (.a(net2501),
    .o(net753));
 b15bfn001ah1n12x5 load_slew754 (.a(gen_filter_20__u_filter_filter_synced),
    .o(net754));
 b15bfn000as1n12x5 wire755 (.a(gen_filter_0__u_filter_filter_synced),
    .o(net755));
 b15bfn001as1n24x5 wire756 (.a(net757),
    .o(net756));
 b15bfn001ah1n48x5 load_slew757 (.a(n3538),
    .o(net757));
 b15bfn001as1n64x5 fanout758 (.a(n4096),
    .o(net758));
 b15bfn001as1n24x5 wire759 (.a(net760),
    .o(net759));
 b15bfn001aq1n48x5 wire760 (.a(net758),
    .o(net760));
 b15bfn001as1n64x5 fanout761 (.a(n4095),
    .o(net761));
 b15bfn001as1n24x5 max_length762 (.a(net763),
    .o(net762));
 b15bfn001ah1n48x5 wire763 (.a(net761),
    .o(net763));
 b15bfn001as1n24x5 wire764 (.a(net766),
    .o(net764));
 b15bfn001ah1n32x5 wire765 (.a(n4094),
    .o(net765));
 b15bfn001ah1n24x5 max_length766 (.a(n4094),
    .o(net766));
 b15bfn001as1n48x5 fanout767 (.a(n4093),
    .o(net767));
 b15bfn001ah1n24x5 max_length768 (.a(net769),
    .o(net768));
 b15bfn001as1n32x5 wire769 (.a(net767),
    .o(net769));
 b15bfn001as1n24x5 wire770 (.a(net767),
    .o(net770));
 b15bfn001as1n64x5 fanout771 (.a(n4092),
    .o(net771));
 b15bfn000as1n32x5 max_length772 (.a(net773),
    .o(net772));
 b15bfn000as1n32x5 wire773 (.a(net771),
    .o(net773));
 b15bfn001as1n64x5 fanout774 (.a(n4091),
    .o(net774));
 b15bfn001ah1n32x5 max_length775 (.a(net776),
    .o(net775));
 b15bfn001as1n32x5 wire776 (.a(net774),
    .o(net776));
 b15bfn001as1n32x5 max_length777 (.a(net779),
    .o(net777));
 b15bfn001as1n32x5 wire778 (.a(net779),
    .o(net778));
 b15bfn001as1n32x5 wire779 (.a(n4090),
    .o(net779));
 b15bfn001as1n64x5 fanout780 (.a(n4089),
    .o(net780));
 b15bfn001ah1n32x5 max_length781 (.a(net783),
    .o(net781));
 b15bfn001as1n24x5 max_length782 (.a(net783),
    .o(net782));
 b15bfn001as1n32x5 wire783 (.a(net780),
    .o(net783));
 b15bfn001as1n24x5 wire784 (.a(net785),
    .o(net784));
 b15bfn001as1n24x5 wire785 (.a(n4088),
    .o(net785));
 b15bfn001as1n64x5 fanout786 (.a(n4087),
    .o(net786));
 b15bfn001as1n24x5 wire787 (.a(net788),
    .o(net787));
 b15bfn001ah1n32x5 wire788 (.a(net786),
    .o(net788));
 b15bfn001as1n48x5 fanout789 (.a(n4086),
    .o(net789));
 b15bfn001ah1n24x5 max_length790 (.a(net791),
    .o(net790));
 b15bfn001as1n24x5 max_length791 (.a(net792),
    .o(net791));
 b15bfn001as1n32x5 wire792 (.a(net789),
    .o(net792));
 b15bfn001as1n32x5 max_length793 (.a(net794),
    .o(net793));
 b15bfn000as1n24x5 wire794 (.a(net795),
    .o(net794));
 b15bfn001aq1n48x5 wire795 (.a(n4085),
    .o(net795));
 b15bfn001ah1n32x5 wire796 (.a(net798),
    .o(net796));
 b15bfn001as1n48x5 max_length797 (.a(n4084),
    .o(net797));
 b15bfn001ah1n48x5 max_length798 (.a(n4084),
    .o(net798));
 b15bfn001as1n64x5 fanout799 (.a(n4083),
    .o(net799));
 b15bfn001ah1n24x5 wire800 (.a(net799),
    .o(net800));
 b15bfn001ah1n48x5 wire801 (.a(net799),
    .o(net801));
 b15bfn001as1n64x5 fanout802 (.a(n4082),
    .o(net802));
 b15bfn001as1n16x5 max_length803 (.a(net805),
    .o(net803));
 b15bfn001ah1n32x5 wire804 (.a(net802),
    .o(net804));
 b15bfn001ah1n48x5 max_length805 (.a(net802),
    .o(net805));
 b15bfn001ah1n32x5 wire806 (.a(n4081),
    .o(net806));
 b15bfn001ah1n32x5 wire807 (.a(n4081),
    .o(net807));
 b15bfn001ah1n32x5 max_length808 (.a(net809),
    .o(net808));
 b15bfn001ah1n24x5 max_length809 (.a(n4079),
    .o(net809));
 b15bfn001ah1n32x5 max_length810 (.a(n4079),
    .o(net810));
 b15bfn001ah1n32x5 max_length811 (.a(net812),
    .o(net811));
 b15bfn001ah1n32x5 max_length812 (.a(n4078),
    .o(net812));
 b15bfn001ah1n24x5 max_length813 (.a(n4073),
    .o(net813));
 b15bfn001as1n32x5 max_length814 (.a(n4073),
    .o(net814));
 b15bfn001as1n32x5 max_length815 (.a(net816),
    .o(net815));
 b15bfn001as1n32x5 wire816 (.a(n4070),
    .o(net816));
 b15bfn001as1n32x5 wire817 (.a(n4068),
    .o(net817));
 b15bfn001as1n24x5 wire818 (.a(n4068),
    .o(net818));
 b15bfn001ah1n32x5 wire819 (.a(net820),
    .o(net819));
 b15bfn001as1n32x5 wire820 (.a(n4067),
    .o(net820));
 b15bfn001ah1n32x5 max_length821 (.a(net86),
    .o(net821));
 b15bfn001ah1n48x5 wire822 (.a(net82),
    .o(net822));
 b15bfn001ah1n48x5 wire823 (.a(net81),
    .o(net823));
 b15bfn001as1n16x5 wire824 (.a(net8),
    .o(net824));
 b15bfn000ah1n48x5 wire825 (.a(net78),
    .o(net825));
 b15bfn001ah1n48x5 wire826 (.a(net76),
    .o(net826));
 b15bfn001as1n24x5 wire827 (.a(net75),
    .o(net827));
 b15bfn001as1n32x5 wire828 (.a(net74),
    .o(net828));
 b15bfn001ah1n48x5 load_slew829 (.a(net60),
    .o(net829));
 b15bfn001as1n32x5 wire830 (.a(net58),
    .o(net830));
 b15bfn001ah1n48x5 wire831 (.a(net57),
    .o(net831));
 b15bfn001as1n32x5 wire832 (.a(net56),
    .o(net832));
 b15bfn001as1n48x5 fanout833 (.a(net836),
    .o(net833));
 b15bfn001as1n48x5 fanout834 (.a(net836),
    .o(net834));
 b15bfn001as1n24x5 fanout835 (.a(net836),
    .o(net835));
 b15bfn001as1n48x5 fanout836 (.a(net847),
    .o(net836));
 b15bfn001as1n48x5 fanout837 (.a(net838),
    .o(net837));
 b15bfn001as1n48x5 fanout838 (.a(net847),
    .o(net838));
 b15bfn001ah1n64x5 fanout839 (.a(net849),
    .o(net839));
 b15bfn001as1n48x5 fanout840 (.a(net843),
    .o(net840));
 b15bfn001ah1n64x5 fanout841 (.a(net843),
    .o(net841));
 b15bfn000as1n32x5 fanout842 (.a(net843),
    .o(net842));
 b15bfn001ah1n48x5 fanout843 (.a(net850),
    .o(net843));
 b15bfn001ah1n64x5 fanout844 (.a(net848),
    .o(net844));
 b15bfn001ah1n32x5 fanout845 (.a(net848),
    .o(net845));
 b15bfn001ah1n64x5 fanout846 (.a(net848),
    .o(net846));
 b15bfn001as1n64x5 fanout847 (.a(net37),
    .o(net847));
 b15bfn001ah1n48x5 wire848 (.a(net849),
    .o(net848));
 b15bfn001as1n32x5 wire849 (.a(net847),
    .o(net849));
 b15bfn001ah1n32x5 max_length850 (.a(net847),
    .o(net850));
 b15bfn001as1n48x5 fanout851 (.a(net857),
    .o(net851));
 b15bfn001ah1n32x5 fanout852 (.a(net857),
    .o(net852));
 b15bfn001ah1n64x5 fanout853 (.a(net857),
    .o(net853));
 b15bfn001ah1n48x5 fanout854 (.a(net858),
    .o(net854));
 b15bfn001ah1n24x5 fanout855 (.a(net858),
    .o(net855));
 b15bfn001ah1n64x5 fanout856 (.a(net858),
    .o(net856));
 b15bfn001as1n48x5 fanout857 (.a(net868),
    .o(net857));
 b15bfn001as1n32x5 wire858 (.a(net857),
    .o(net858));
 b15bfn001ah1n64x5 fanout859 (.a(net865),
    .o(net859));
 b15bfn001ah1n64x5 fanout860 (.a(net867),
    .o(net860));
 b15bfn001ah1n48x5 fanout861 (.a(net866),
    .o(net861));
 b15bfn001ah1n64x5 fanout862 (.a(net867),
    .o(net862));
 b15bfn001as1n48x5 fanout863 (.a(net866),
    .o(net863));
 b15bfn001as1n32x5 fanout864 (.a(net866),
    .o(net864));
 b15bfn001as1n64x5 fanout865 (.a(net868),
    .o(net865));
 b15bfn001ah1n48x5 max_length866 (.a(net867),
    .o(net866));
 b15bfn001ah1n48x5 load_slew867 (.a(net865),
    .o(net867));
 b15bfn001as1n32x5 wire868 (.a(net37),
    .o(net868));
 b15bfn001as1n32x5 wire869 (.a(net27),
    .o(net869));
 b15bfn001as1n16x5 wire870 (.a(net17),
    .o(net870));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_0__cio_gpio_en_q_reg_1__871 (.o(net871));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_0__cio_gpio_en_q_reg_1__872 (.o(net872));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_10__cio_gpio_en_q_reg_11__873 (.o(net873));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_10__cio_gpio_en_q_reg_11__874 (.o(net874));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_12__cio_gpio_en_q_reg_13__875 (.o(net875));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_12__cio_gpio_en_q_reg_13__876 (.o(net876));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_14__cio_gpio_en_q_reg_15__877 (.o(net877));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_14__cio_gpio_en_q_reg_15__878 (.o(net878));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_16__cio_gpio_en_q_reg_17__879 (.o(net879));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_16__cio_gpio_en_q_reg_17__880 (.o(net880));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_18__cio_gpio_en_q_reg_19__881 (.o(net881));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_18__cio_gpio_en_q_reg_19__882 (.o(net882));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_20__cio_gpio_en_q_reg_21__883 (.o(net883));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_20__cio_gpio_en_q_reg_21__884 (.o(net884));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_22__cio_gpio_en_q_reg_23__885 (.o(net885));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_22__cio_gpio_en_q_reg_23__886 (.o(net886));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_24__cio_gpio_en_q_reg_25__887 (.o(net887));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_24__cio_gpio_en_q_reg_25__888 (.o(net888));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_26__cio_gpio_en_q_reg_27__889 (.o(net889));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_26__cio_gpio_en_q_reg_27__890 (.o(net890));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_28__cio_gpio_en_q_reg_29__891 (.o(net891));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_28__cio_gpio_en_q_reg_29__892 (.o(net892));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_2__cio_gpio_en_q_reg_3__893 (.o(net893));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_2__cio_gpio_en_q_reg_3__894 (.o(net894));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_30__cio_gpio_en_q_reg_31__895 (.o(net895));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_30__cio_gpio_en_q_reg_31__896 (.o(net896));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_4__cio_gpio_en_q_reg_5__897 (.o(net897));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_4__cio_gpio_en_q_reg_5__898 (.o(net898));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_6__cio_gpio_en_q_reg_7__899 (.o(net899));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_6__cio_gpio_en_q_reg_7__900 (.o(net900));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_8__cio_gpio_en_q_reg_9__901 (.o(net901));
 b15tilo00an1n03x5 cio_gpio_en_q_reg_8__cio_gpio_en_q_reg_9__902 (.o(net902));
 b15tilo00an1n03x5 cio_gpio_q_reg_0__cio_gpio_q_reg_1__903 (.o(net903));
 b15tilo00an1n03x5 cio_gpio_q_reg_0__cio_gpio_q_reg_1__904 (.o(net904));
 b15tilo00an1n03x5 cio_gpio_q_reg_10__cio_gpio_q_reg_11__905 (.o(net905));
 b15tilo00an1n03x5 cio_gpio_q_reg_10__cio_gpio_q_reg_11__906 (.o(net906));
 b15tilo00an1n03x5 cio_gpio_q_reg_12__cio_gpio_q_reg_13__907 (.o(net907));
 b15tilo00an1n03x5 cio_gpio_q_reg_12__cio_gpio_q_reg_13__908 (.o(net908));
 b15tilo00an1n03x5 cio_gpio_q_reg_14__cio_gpio_q_reg_15__909 (.o(net909));
 b15tilo00an1n03x5 cio_gpio_q_reg_14__cio_gpio_q_reg_15__910 (.o(net910));
 b15tilo00an1n03x5 cio_gpio_q_reg_16__cio_gpio_q_reg_17__911 (.o(net911));
 b15tilo00an1n03x5 cio_gpio_q_reg_16__cio_gpio_q_reg_17__912 (.o(net912));
 b15tilo00an1n03x5 cio_gpio_q_reg_18__cio_gpio_q_reg_19__913 (.o(net913));
 b15tilo00an1n03x5 cio_gpio_q_reg_18__cio_gpio_q_reg_19__914 (.o(net914));
 b15tilo00an1n03x5 cio_gpio_q_reg_20__cio_gpio_q_reg_21__915 (.o(net915));
 b15tilo00an1n03x5 cio_gpio_q_reg_20__cio_gpio_q_reg_21__916 (.o(net916));
 b15tilo00an1n03x5 cio_gpio_q_reg_22__cio_gpio_q_reg_23__917 (.o(net917));
 b15tilo00an1n03x5 cio_gpio_q_reg_22__cio_gpio_q_reg_23__918 (.o(net918));
 b15tilo00an1n03x5 cio_gpio_q_reg_24__cio_gpio_q_reg_25__919 (.o(net919));
 b15tilo00an1n03x5 cio_gpio_q_reg_24__cio_gpio_q_reg_25__920 (.o(net920));
 b15tilo00an1n03x5 cio_gpio_q_reg_26__cio_gpio_q_reg_27__921 (.o(net921));
 b15tilo00an1n03x5 cio_gpio_q_reg_26__cio_gpio_q_reg_27__922 (.o(net922));
 b15tilo00an1n03x5 cio_gpio_q_reg_28__cio_gpio_q_reg_29__923 (.o(net923));
 b15tilo00an1n03x5 cio_gpio_q_reg_28__cio_gpio_q_reg_29__924 (.o(net924));
 b15tilo00an1n03x5 cio_gpio_q_reg_2__cio_gpio_q_reg_3__925 (.o(net925));
 b15tilo00an1n03x5 cio_gpio_q_reg_2__cio_gpio_q_reg_3__926 (.o(net926));
 b15tilo00an1n03x5 cio_gpio_q_reg_30__cio_gpio_q_reg_31__927 (.o(net927));
 b15tilo00an1n03x5 cio_gpio_q_reg_30__cio_gpio_q_reg_31__928 (.o(net928));
 b15tilo00an1n03x5 cio_gpio_q_reg_4__cio_gpio_q_reg_5__929 (.o(net929));
 b15tilo00an1n03x5 cio_gpio_q_reg_4__cio_gpio_q_reg_5__930 (.o(net930));
 b15tilo00an1n03x5 cio_gpio_q_reg_6__cio_gpio_q_reg_7__931 (.o(net931));
 b15tilo00an1n03x5 cio_gpio_q_reg_6__cio_gpio_q_reg_7__932 (.o(net932));
 b15tilo00an1n03x5 cio_gpio_q_reg_8__cio_gpio_q_reg_9__933 (.o(net933));
 b15tilo00an1n03x5 cio_gpio_q_reg_8__cio_gpio_q_reg_9__934 (.o(net934));
 b15tilo00an1n03x5 clk_gate_cio_gpio_en_q_reg_0_latch_935 (.o(net935));
 b15tilo00an1n03x5 clk_gate_cio_gpio_en_q_reg_latch_936 (.o(net936));
 b15tilo00an1n03x5 clk_gate_cio_gpio_q_reg_0_latch_937 (.o(net937));
 b15tilo00an1n03x5 clk_gate_cio_gpio_q_reg_latch_938 (.o(net938));
 b15tilo00an1n03x5 data_in_q_reg_0__data_in_q_reg_1__939 (.o(net939));
 b15tilo00an1n03x5 data_in_q_reg_0__data_in_q_reg_1__940 (.o(net940));
 b15tilo00an1n03x5 data_in_q_reg_10__data_in_q_reg_11__941 (.o(net941));
 b15tilo00an1n03x5 data_in_q_reg_10__data_in_q_reg_11__942 (.o(net942));
 b15tilo00an1n03x5 data_in_q_reg_12__data_in_q_reg_13__943 (.o(net943));
 b15tilo00an1n03x5 data_in_q_reg_12__data_in_q_reg_13__944 (.o(net944));
 b15tilo00an1n03x5 data_in_q_reg_14__data_in_q_reg_15__945 (.o(net945));
 b15tilo00an1n03x5 data_in_q_reg_14__data_in_q_reg_15__946 (.o(net946));
 b15tilo00an1n03x5 data_in_q_reg_16__data_in_q_reg_17__947 (.o(net947));
 b15tilo00an1n03x5 data_in_q_reg_16__data_in_q_reg_17__948 (.o(net948));
 b15tilo00an1n03x5 data_in_q_reg_18__data_in_q_reg_19__949 (.o(net949));
 b15tilo00an1n03x5 data_in_q_reg_18__data_in_q_reg_19__950 (.o(net950));
 b15tilo00an1n03x5 data_in_q_reg_20__data_in_q_reg_21__951 (.o(net951));
 b15tilo00an1n03x5 data_in_q_reg_20__data_in_q_reg_21__952 (.o(net952));
 b15tilo00an1n03x5 data_in_q_reg_22__data_in_q_reg_23__953 (.o(net953));
 b15tilo00an1n03x5 data_in_q_reg_22__data_in_q_reg_23__954 (.o(net954));
 b15tilo00an1n03x5 data_in_q_reg_24__data_in_q_reg_25__955 (.o(net955));
 b15tilo00an1n03x5 data_in_q_reg_24__data_in_q_reg_25__956 (.o(net956));
 b15tilo00an1n03x5 data_in_q_reg_26__data_in_q_reg_27__957 (.o(net957));
 b15tilo00an1n03x5 data_in_q_reg_26__data_in_q_reg_27__958 (.o(net958));
 b15tilo00an1n03x5 data_in_q_reg_28__data_in_q_reg_29__959 (.o(net959));
 b15tilo00an1n03x5 data_in_q_reg_28__data_in_q_reg_29__960 (.o(net960));
 b15tilo00an1n03x5 data_in_q_reg_2__data_in_q_reg_3__961 (.o(net961));
 b15tilo00an1n03x5 data_in_q_reg_2__data_in_q_reg_3__962 (.o(net962));
 b15tilo00an1n03x5 data_in_q_reg_30__data_in_q_reg_31__963 (.o(net963));
 b15tilo00an1n03x5 data_in_q_reg_30__data_in_q_reg_31__964 (.o(net964));
 b15tilo00an1n03x5 data_in_q_reg_4__data_in_q_reg_5__965 (.o(net965));
 b15tilo00an1n03x5 data_in_q_reg_4__data_in_q_reg_5__966 (.o(net966));
 b15tilo00an1n03x5 data_in_q_reg_6__data_in_q_reg_7__967 (.o(net967));
 b15tilo00an1n03x5 data_in_q_reg_6__data_in_q_reg_7__968 (.o(net968));
 b15tilo00an1n03x5 data_in_q_reg_8__data_in_q_reg_9__969 (.o(net969));
 b15tilo00an1n03x5 data_in_q_reg_8__data_in_q_reg_9__970 (.o(net970));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_alert_set_q_reg_gen_filter_5__u_filter_filter_q_reg_971 (.o(net971));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_alert_set_q_reg_gen_filter_5__u_filter_filter_q_reg_972 (.o(net972));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_0__973 (.o(net973));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_0__974 (.o(net974));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_ping_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_1__975 (.o(net975));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_ping_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_1__976 (.o(net976));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_state_q_reg_2__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq_reg_977 (.o(net977));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_state_q_reg_2__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq_reg_978 (.o(net978));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq_reg_979 (.o(net979));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__980 (.o(net980));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__981 (.o(net981));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__982 (.o(net982));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__983 (.o(net983));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_0__984 (.o(net984));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_1__985 (.o(net985));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q_reg_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq_reg_986 (.o(net986));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q_reg_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq_reg_987 (.o(net987));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq_reg_988 (.o(net988));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__989 (.o(net989));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__990 (.o(net990));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__991 (.o(net991));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__992 (.o(net992));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_0__993 (.o(net993));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_1__994 (.o(net994));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q_reg_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__995 (.o(net995));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q_reg_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__996 (.o(net996));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_0__u_filter_diff_ctr_q_reg_0__997 (.o(net997));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_0__u_filter_diff_ctr_q_reg_0__998 (.o(net998));
 b15tilo00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_1__999 (.o(net999));
 b15tilo00an1n03x5 gen_filter_0__u_filter_diff_ctr_q_reg_1__gen_filter_0__u_filter_diff_ctr_q_reg_2__1000 (.o(net1000));
 b15tilo00an1n03x5 gen_filter_0__u_filter_diff_ctr_q_reg_1__gen_filter_0__u_filter_diff_ctr_q_reg_2__1001 (.o(net1001));
 b15tilo00an1n03x5 gen_filter_0__u_filter_diff_ctr_q_reg_3__gen_filter_0__u_filter_filter_q_reg_1002 (.o(net1002));
 b15tilo00an1n03x5 gen_filter_0__u_filter_diff_ctr_q_reg_3__gen_filter_0__u_filter_filter_q_reg_1003 (.o(net1003));
 b15tilo00an1n03x5 gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_16__u_filter_diff_ctr_q_reg_0__1004 (.o(net1004));
 b15tilo00an1n03x5 gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_16__u_filter_diff_ctr_q_reg_0__1005 (.o(net1005));
 b15tilo00an1n03x5 gen_filter_0__u_filter_stored_value_q_reg_1006 (.o(net1006));
 b15tilo00an1n03x5 gen_filter_10__u_filter_diff_ctr_q_reg_0__gen_filter_10__u_filter_diff_ctr_q_reg_3__1007 (.o(net1007));
 b15tilo00an1n03x5 gen_filter_10__u_filter_diff_ctr_q_reg_0__gen_filter_10__u_filter_diff_ctr_q_reg_3__1008 (.o(net1008));
 b15tilo00an1n03x5 gen_filter_10__u_filter_diff_ctr_q_reg_1__gen_filter_10__u_filter_diff_ctr_q_reg_2__1009 (.o(net1009));
 b15tilo00an1n03x5 gen_filter_10__u_filter_diff_ctr_q_reg_1__gen_filter_10__u_filter_diff_ctr_q_reg_2__1010 (.o(net1010));
 b15tilo00an1n03x5 gen_filter_10__u_filter_filter_q_reg_gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1011 (.o(net1011));
 b15tilo00an1n03x5 gen_filter_10__u_filter_filter_q_reg_gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1012 (.o(net1012));
 b15tilo00an1n03x5 gen_filter_10__u_filter_stored_value_q_reg_1013 (.o(net1013));
 b15tilo00an1n03x5 gen_filter_11__u_filter_diff_ctr_q_reg_0__gen_filter_11__u_filter_diff_ctr_q_reg_1__1014 (.o(net1014));
 b15tilo00an1n03x5 gen_filter_11__u_filter_diff_ctr_q_reg_0__gen_filter_11__u_filter_diff_ctr_q_reg_1__1015 (.o(net1015));
 b15tilo00an1n03x5 gen_filter_11__u_filter_diff_ctr_q_reg_3__gen_filter_11__u_filter_filter_q_reg_1016 (.o(net1016));
 b15tilo00an1n03x5 gen_filter_11__u_filter_diff_ctr_q_reg_3__gen_filter_11__u_filter_filter_q_reg_1017 (.o(net1017));
 b15tilo00an1n03x5 gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1018 (.o(net1018));
 b15tilo00an1n03x5 gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1019 (.o(net1019));
 b15tilo00an1n03x5 gen_filter_11__u_filter_stored_value_q_reg_1020 (.o(net1020));
 b15tilo00an1n03x5 gen_filter_12__u_filter_diff_ctr_q_reg_0__gen_filter_12__u_filter_diff_ctr_q_reg_1__1021 (.o(net1021));
 b15tilo00an1n03x5 gen_filter_12__u_filter_diff_ctr_q_reg_0__gen_filter_12__u_filter_diff_ctr_q_reg_1__1022 (.o(net1022));
 b15tilo00an1n03x5 gen_filter_12__u_filter_diff_ctr_q_reg_2__gen_filter_12__u_filter_diff_ctr_q_reg_3__1023 (.o(net1023));
 b15tilo00an1n03x5 gen_filter_12__u_filter_diff_ctr_q_reg_2__gen_filter_12__u_filter_diff_ctr_q_reg_3__1024 (.o(net1024));
 b15tilo00an1n03x5 gen_filter_12__u_filter_filter_q_reg_gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1025 (.o(net1025));
 b15tilo00an1n03x5 gen_filter_12__u_filter_filter_q_reg_gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1026 (.o(net1026));
 b15tilo00an1n03x5 gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_13__u_filter_diff_ctr_q_reg_0__1027 (.o(net1027));
 b15tilo00an1n03x5 gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_13__u_filter_diff_ctr_q_reg_0__1028 (.o(net1028));
 b15tilo00an1n03x5 gen_filter_12__u_filter_stored_value_q_reg_1029 (.o(net1029));
 b15tilo00an1n03x5 gen_filter_13__u_filter_diff_ctr_q_reg_1__gen_filter_13__u_filter_diff_ctr_q_reg_2__1030 (.o(net1030));
 b15tilo00an1n03x5 gen_filter_13__u_filter_diff_ctr_q_reg_1__gen_filter_13__u_filter_diff_ctr_q_reg_2__1031 (.o(net1031));
 b15tilo00an1n03x5 gen_filter_13__u_filter_diff_ctr_q_reg_3__gen_filter_13__u_filter_filter_q_reg_1032 (.o(net1032));
 b15tilo00an1n03x5 gen_filter_13__u_filter_diff_ctr_q_reg_3__gen_filter_13__u_filter_filter_q_reg_1033 (.o(net1033));
 b15tilo00an1n03x5 gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1034 (.o(net1034));
 b15tilo00an1n03x5 gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1035 (.o(net1035));
 b15tilo00an1n03x5 gen_filter_13__u_filter_stored_value_q_reg_1036 (.o(net1036));
 b15tilo00an1n03x5 gen_filter_14__u_filter_diff_ctr_q_reg_0__gen_filter_14__u_filter_diff_ctr_q_reg_1__1037 (.o(net1037));
 b15tilo00an1n03x5 gen_filter_14__u_filter_diff_ctr_q_reg_0__gen_filter_14__u_filter_diff_ctr_q_reg_1__1038 (.o(net1038));
 b15tilo00an1n03x5 gen_filter_14__u_filter_diff_ctr_q_reg_2__gen_filter_14__u_filter_diff_ctr_q_reg_3__1039 (.o(net1039));
 b15tilo00an1n03x5 gen_filter_14__u_filter_diff_ctr_q_reg_2__gen_filter_14__u_filter_diff_ctr_q_reg_3__1040 (.o(net1040));
 b15tilo00an1n03x5 gen_filter_14__u_filter_filter_q_reg_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1041 (.o(net1041));
 b15tilo00an1n03x5 gen_filter_14__u_filter_filter_q_reg_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1042 (.o(net1042));
 b15tilo00an1n03x5 gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1043 (.o(net1043));
 b15tilo00an1n03x5 gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1044 (.o(net1044));
 b15tilo00an1n03x5 gen_filter_14__u_filter_stored_value_q_reg_1045 (.o(net1045));
 b15tilo00an1n03x5 gen_filter_15__u_filter_diff_ctr_q_reg_1__gen_filter_15__u_filter_diff_ctr_q_reg_2__1046 (.o(net1046));
 b15tilo00an1n03x5 gen_filter_15__u_filter_diff_ctr_q_reg_1__gen_filter_15__u_filter_diff_ctr_q_reg_2__1047 (.o(net1047));
 b15tilo00an1n03x5 gen_filter_15__u_filter_diff_ctr_q_reg_3__gen_filter_15__u_filter_filter_q_reg_1048 (.o(net1048));
 b15tilo00an1n03x5 gen_filter_15__u_filter_diff_ctr_q_reg_3__gen_filter_15__u_filter_filter_q_reg_1049 (.o(net1049));
 b15tilo00an1n03x5 gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1050 (.o(net1050));
 b15tilo00an1n03x5 gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1051 (.o(net1051));
 b15tilo00an1n03x5 gen_filter_15__u_filter_stored_value_q_reg_1052 (.o(net1052));
 b15tilo00an1n03x5 gen_filter_16__u_filter_diff_ctr_q_reg_1__gen_filter_16__u_filter_diff_ctr_q_reg_2__1053 (.o(net1053));
 b15tilo00an1n03x5 gen_filter_16__u_filter_diff_ctr_q_reg_1__gen_filter_16__u_filter_diff_ctr_q_reg_2__1054 (.o(net1054));
 b15tilo00an1n03x5 gen_filter_16__u_filter_diff_ctr_q_reg_3__gen_filter_16__u_filter_filter_q_reg_1055 (.o(net1055));
 b15tilo00an1n03x5 gen_filter_16__u_filter_diff_ctr_q_reg_3__gen_filter_16__u_filter_filter_q_reg_1056 (.o(net1056));
 b15tilo00an1n03x5 gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_diff_ctr_q_reg_0__1057 (.o(net1057));
 b15tilo00an1n03x5 gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_diff_ctr_q_reg_0__1058 (.o(net1058));
 b15tilo00an1n03x5 gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_30__u_filter_diff_ctr_q_reg_0__1059 (.o(net1059));
 b15tilo00an1n03x5 gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_30__u_filter_diff_ctr_q_reg_0__1060 (.o(net1060));
 b15tilo00an1n03x5 gen_filter_16__u_filter_stored_value_q_reg_1061 (.o(net1061));
 b15tilo00an1n03x5 gen_filter_17__u_filter_diff_ctr_q_reg_1__gen_filter_17__u_filter_diff_ctr_q_reg_2__1062 (.o(net1062));
 b15tilo00an1n03x5 gen_filter_17__u_filter_diff_ctr_q_reg_1__gen_filter_17__u_filter_diff_ctr_q_reg_2__1063 (.o(net1063));
 b15tilo00an1n03x5 gen_filter_17__u_filter_diff_ctr_q_reg_3__gen_filter_17__u_filter_filter_q_reg_1064 (.o(net1064));
 b15tilo00an1n03x5 gen_filter_17__u_filter_diff_ctr_q_reg_3__gen_filter_17__u_filter_filter_q_reg_1065 (.o(net1065));
 b15tilo00an1n03x5 gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1066 (.o(net1066));
 b15tilo00an1n03x5 gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1067 (.o(net1067));
 b15tilo00an1n03x5 gen_filter_17__u_filter_stored_value_q_reg_1068 (.o(net1068));
 b15tilo00an1n03x5 gen_filter_18__u_filter_diff_ctr_q_reg_0__gen_filter_18__u_filter_diff_ctr_q_reg_1__1069 (.o(net1069));
 b15tilo00an1n03x5 gen_filter_18__u_filter_diff_ctr_q_reg_0__gen_filter_18__u_filter_diff_ctr_q_reg_1__1070 (.o(net1070));
 b15tilo00an1n03x5 gen_filter_18__u_filter_diff_ctr_q_reg_2__gen_filter_18__u_filter_diff_ctr_q_reg_3__1071 (.o(net1071));
 b15tilo00an1n03x5 gen_filter_18__u_filter_diff_ctr_q_reg_2__gen_filter_18__u_filter_diff_ctr_q_reg_3__1072 (.o(net1072));
 b15tilo00an1n03x5 gen_filter_18__u_filter_filter_q_reg_gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1073 (.o(net1073));
 b15tilo00an1n03x5 gen_filter_18__u_filter_filter_q_reg_gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1074 (.o(net1074));
 b15tilo00an1n03x5 gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_diff_ctr_q_reg_0__1075 (.o(net1075));
 b15tilo00an1n03x5 gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_diff_ctr_q_reg_0__1076 (.o(net1076));
 b15tilo00an1n03x5 gen_filter_18__u_filter_stored_value_q_reg_1077 (.o(net1077));
 b15tilo00an1n03x5 gen_filter_19__u_filter_diff_ctr_q_reg_1__gen_filter_19__u_filter_diff_ctr_q_reg_2__1078 (.o(net1078));
 b15tilo00an1n03x5 gen_filter_19__u_filter_diff_ctr_q_reg_1__gen_filter_19__u_filter_diff_ctr_q_reg_2__1079 (.o(net1079));
 b15tilo00an1n03x5 gen_filter_19__u_filter_diff_ctr_q_reg_3__gen_filter_19__u_filter_filter_q_reg_1080 (.o(net1080));
 b15tilo00an1n03x5 gen_filter_19__u_filter_diff_ctr_q_reg_3__gen_filter_19__u_filter_filter_q_reg_1081 (.o(net1081));
 b15tilo00an1n03x5 gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_21__u_filter_diff_ctr_q_reg_0__1082 (.o(net1082));
 b15tilo00an1n03x5 gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_21__u_filter_diff_ctr_q_reg_0__1083 (.o(net1083));
 b15tilo00an1n03x5 gen_filter_19__u_filter_stored_value_q_reg_1084 (.o(net1084));
 b15tilo00an1n03x5 gen_filter_1__u_filter_diff_ctr_q_reg_0__gen_filter_1__u_filter_diff_ctr_q_reg_1__1085 (.o(net1085));
 b15tilo00an1n03x5 gen_filter_1__u_filter_diff_ctr_q_reg_0__gen_filter_1__u_filter_diff_ctr_q_reg_1__1086 (.o(net1086));
 b15tilo00an1n03x5 gen_filter_1__u_filter_diff_ctr_q_reg_2__gen_filter_1__u_filter_diff_ctr_q_reg_3__1087 (.o(net1087));
 b15tilo00an1n03x5 gen_filter_1__u_filter_diff_ctr_q_reg_2__gen_filter_1__u_filter_diff_ctr_q_reg_3__1088 (.o(net1088));
 b15tilo00an1n03x5 gen_filter_1__u_filter_filter_q_reg_gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1089 (.o(net1089));
 b15tilo00an1n03x5 gen_filter_1__u_filter_filter_q_reg_gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1090 (.o(net1090));
 b15tilo00an1n03x5 gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__intr_hw_intr_o_reg_0__1091 (.o(net1091));
 b15tilo00an1n03x5 gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__intr_hw_intr_o_reg_0__1092 (.o(net1092));
 b15tilo00an1n03x5 gen_filter_1__u_filter_stored_value_q_reg_1093 (.o(net1093));
 b15tilo00an1n03x5 gen_filter_20__u_filter_diff_ctr_q_reg_0__gen_filter_20__u_filter_diff_ctr_q_reg_1__1094 (.o(net1094));
 b15tilo00an1n03x5 gen_filter_20__u_filter_diff_ctr_q_reg_0__gen_filter_20__u_filter_diff_ctr_q_reg_1__1095 (.o(net1095));
 b15tilo00an1n03x5 gen_filter_20__u_filter_diff_ctr_q_reg_2__gen_filter_20__u_filter_diff_ctr_q_reg_3__1096 (.o(net1096));
 b15tilo00an1n03x5 gen_filter_20__u_filter_diff_ctr_q_reg_2__gen_filter_20__u_filter_diff_ctr_q_reg_3__1097 (.o(net1097));
 b15tilo00an1n03x5 gen_filter_20__u_filter_filter_q_reg_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1098 (.o(net1098));
 b15tilo00an1n03x5 gen_filter_20__u_filter_filter_q_reg_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1099 (.o(net1099));
 b15tilo00an1n03x5 gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_diff_ctr_q_reg_0__1100 (.o(net1100));
 b15tilo00an1n03x5 gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_diff_ctr_q_reg_0__1101 (.o(net1101));
 b15tilo00an1n03x5 gen_filter_20__u_filter_stored_value_q_reg_1102 (.o(net1102));
 b15tilo00an1n03x5 gen_filter_21__u_filter_diff_ctr_q_reg_1__gen_filter_21__u_filter_diff_ctr_q_reg_2__1103 (.o(net1103));
 b15tilo00an1n03x5 gen_filter_21__u_filter_diff_ctr_q_reg_1__gen_filter_21__u_filter_diff_ctr_q_reg_2__1104 (.o(net1104));
 b15tilo00an1n03x5 gen_filter_21__u_filter_diff_ctr_q_reg_3__gen_filter_21__u_filter_filter_q_reg_1105 (.o(net1105));
 b15tilo00an1n03x5 gen_filter_21__u_filter_diff_ctr_q_reg_3__gen_filter_21__u_filter_filter_q_reg_1106 (.o(net1106));
 b15tilo00an1n03x5 gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1107 (.o(net1107));
 b15tilo00an1n03x5 gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1108 (.o(net1108));
 b15tilo00an1n03x5 gen_filter_21__u_filter_stored_value_q_reg_1109 (.o(net1109));
 b15tilo00an1n03x5 gen_filter_22__u_filter_diff_ctr_q_reg_0__gen_filter_22__u_filter_diff_ctr_q_reg_1__1110 (.o(net1110));
 b15tilo00an1n03x5 gen_filter_22__u_filter_diff_ctr_q_reg_0__gen_filter_22__u_filter_diff_ctr_q_reg_1__1111 (.o(net1111));
 b15tilo00an1n03x5 gen_filter_22__u_filter_diff_ctr_q_reg_2__gen_filter_22__u_filter_diff_ctr_q_reg_3__1112 (.o(net1112));
 b15tilo00an1n03x5 gen_filter_22__u_filter_diff_ctr_q_reg_2__gen_filter_22__u_filter_diff_ctr_q_reg_3__1113 (.o(net1113));
 b15tilo00an1n03x5 gen_filter_22__u_filter_filter_q_reg_gen_filter_24__u_filter_diff_ctr_q_reg_0__1114 (.o(net1114));
 b15tilo00an1n03x5 gen_filter_22__u_filter_filter_q_reg_gen_filter_24__u_filter_diff_ctr_q_reg_0__1115 (.o(net1115));
 b15tilo00an1n03x5 gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1116 (.o(net1116));
 b15tilo00an1n03x5 gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1117 (.o(net1117));
 b15tilo00an1n03x5 gen_filter_22__u_filter_stored_value_q_reg_1118 (.o(net1118));
 b15tilo00an1n03x5 gen_filter_23__u_filter_diff_ctr_q_reg_1__gen_filter_23__u_filter_diff_ctr_q_reg_2__1119 (.o(net1119));
 b15tilo00an1n03x5 gen_filter_23__u_filter_diff_ctr_q_reg_1__gen_filter_23__u_filter_diff_ctr_q_reg_2__1120 (.o(net1120));
 b15tilo00an1n03x5 gen_filter_23__u_filter_diff_ctr_q_reg_3__gen_filter_23__u_filter_filter_q_reg_1121 (.o(net1121));
 b15tilo00an1n03x5 gen_filter_23__u_filter_diff_ctr_q_reg_3__gen_filter_23__u_filter_filter_q_reg_1122 (.o(net1122));
 b15tilo00an1n03x5 gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1123 (.o(net1123));
 b15tilo00an1n03x5 gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1124 (.o(net1124));
 b15tilo00an1n03x5 gen_filter_23__u_filter_stored_value_q_reg_1125 (.o(net1125));
 b15tilo00an1n03x5 gen_filter_24__u_filter_diff_ctr_q_reg_1__gen_filter_24__u_filter_diff_ctr_q_reg_3__1126 (.o(net1126));
 b15tilo00an1n03x5 gen_filter_24__u_filter_diff_ctr_q_reg_1__gen_filter_24__u_filter_diff_ctr_q_reg_3__1127 (.o(net1127));
 b15tilo00an1n03x5 gen_filter_24__u_filter_diff_ctr_q_reg_2__gen_filter_24__u_filter_filter_q_reg_1128 (.o(net1128));
 b15tilo00an1n03x5 gen_filter_24__u_filter_diff_ctr_q_reg_2__gen_filter_24__u_filter_filter_q_reg_1129 (.o(net1129));
 b15tilo00an1n03x5 gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1130 (.o(net1130));
 b15tilo00an1n03x5 gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1131 (.o(net1131));
 b15tilo00an1n03x5 gen_filter_24__u_filter_stored_value_q_reg_1132 (.o(net1132));
 b15tilo00an1n03x5 gen_filter_25__u_filter_diff_ctr_q_reg_0__gen_filter_25__u_filter_diff_ctr_q_reg_1__1133 (.o(net1133));
 b15tilo00an1n03x5 gen_filter_25__u_filter_diff_ctr_q_reg_0__gen_filter_25__u_filter_diff_ctr_q_reg_1__1134 (.o(net1134));
 b15tilo00an1n03x5 gen_filter_25__u_filter_diff_ctr_q_reg_2__gen_filter_25__u_filter_diff_ctr_q_reg_3__1135 (.o(net1135));
 b15tilo00an1n03x5 gen_filter_25__u_filter_diff_ctr_q_reg_2__gen_filter_25__u_filter_diff_ctr_q_reg_3__1136 (.o(net1136));
 b15tilo00an1n03x5 gen_filter_25__u_filter_filter_q_reg_1137 (.o(net1137));
 b15tilo00an1n03x5 gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1138 (.o(net1138));
 b15tilo00an1n03x5 gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1139 (.o(net1139));
 b15tilo00an1n03x5 gen_filter_25__u_filter_stored_value_q_reg_1140 (.o(net1140));
 b15tilo00an1n03x5 gen_filter_26__u_filter_diff_ctr_q_reg_0__gen_filter_26__u_filter_diff_ctr_q_reg_1__1141 (.o(net1141));
 b15tilo00an1n03x5 gen_filter_26__u_filter_diff_ctr_q_reg_0__gen_filter_26__u_filter_diff_ctr_q_reg_1__1142 (.o(net1142));
 b15tilo00an1n03x5 gen_filter_26__u_filter_diff_ctr_q_reg_2__gen_filter_26__u_filter_diff_ctr_q_reg_3__1143 (.o(net1143));
 b15tilo00an1n03x5 gen_filter_26__u_filter_diff_ctr_q_reg_2__gen_filter_26__u_filter_diff_ctr_q_reg_3__1144 (.o(net1144));
 b15tilo00an1n03x5 gen_filter_26__u_filter_filter_q_reg_gen_filter_31__u_filter_diff_ctr_q_reg_0__1145 (.o(net1145));
 b15tilo00an1n03x5 gen_filter_26__u_filter_filter_q_reg_gen_filter_31__u_filter_diff_ctr_q_reg_0__1146 (.o(net1146));
 b15tilo00an1n03x5 gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_diff_ctr_q_reg_0__1147 (.o(net1147));
 b15tilo00an1n03x5 gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_diff_ctr_q_reg_0__1148 (.o(net1148));
 b15tilo00an1n03x5 gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_31__u_filter_diff_ctr_q_reg_1__1149 (.o(net1149));
 b15tilo00an1n03x5 gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_31__u_filter_diff_ctr_q_reg_1__1150 (.o(net1150));
 b15tilo00an1n03x5 gen_filter_26__u_filter_stored_value_q_reg_1151 (.o(net1151));
 b15tilo00an1n03x5 gen_filter_27__u_filter_diff_ctr_q_reg_0__gen_filter_27__u_filter_diff_ctr_q_reg_1__1152 (.o(net1152));
 b15tilo00an1n03x5 gen_filter_27__u_filter_diff_ctr_q_reg_0__gen_filter_27__u_filter_diff_ctr_q_reg_1__1153 (.o(net1153));
 b15tilo00an1n03x5 gen_filter_27__u_filter_diff_ctr_q_reg_2__gen_filter_27__u_filter_diff_ctr_q_reg_3__1154 (.o(net1154));
 b15tilo00an1n03x5 gen_filter_27__u_filter_diff_ctr_q_reg_2__gen_filter_27__u_filter_diff_ctr_q_reg_3__1155 (.o(net1155));
 b15tilo00an1n03x5 gen_filter_27__u_filter_filter_q_reg_gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1156 (.o(net1156));
 b15tilo00an1n03x5 gen_filter_27__u_filter_filter_q_reg_gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1157 (.o(net1157));
 b15tilo00an1n03x5 gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_30__u_filter_diff_ctr_q_reg_1__1158 (.o(net1158));
 b15tilo00an1n03x5 gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_30__u_filter_diff_ctr_q_reg_1__1159 (.o(net1159));
 b15tilo00an1n03x5 gen_filter_27__u_filter_stored_value_q_reg_1160 (.o(net1160));
 b15tilo00an1n03x5 gen_filter_28__u_filter_diff_ctr_q_reg_1__gen_filter_28__u_filter_diff_ctr_q_reg_2__1161 (.o(net1161));
 b15tilo00an1n03x5 gen_filter_28__u_filter_diff_ctr_q_reg_1__gen_filter_28__u_filter_diff_ctr_q_reg_2__1162 (.o(net1162));
 b15tilo00an1n03x5 gen_filter_28__u_filter_diff_ctr_q_reg_3__gen_filter_28__u_filter_filter_q_reg_1163 (.o(net1163));
 b15tilo00an1n03x5 gen_filter_28__u_filter_diff_ctr_q_reg_3__gen_filter_28__u_filter_filter_q_reg_1164 (.o(net1164));
 b15tilo00an1n03x5 gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1165 (.o(net1165));
 b15tilo00an1n03x5 gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1166 (.o(net1166));
 b15tilo00an1n03x5 gen_filter_28__u_filter_stored_value_q_reg_1167 (.o(net1167));
 b15tilo00an1n03x5 gen_filter_29__u_filter_diff_ctr_q_reg_0__gen_filter_29__u_filter_diff_ctr_q_reg_1__1168 (.o(net1168));
 b15tilo00an1n03x5 gen_filter_29__u_filter_diff_ctr_q_reg_0__gen_filter_29__u_filter_diff_ctr_q_reg_1__1169 (.o(net1169));
 b15tilo00an1n03x5 gen_filter_29__u_filter_diff_ctr_q_reg_2__gen_filter_29__u_filter_diff_ctr_q_reg_3__1170 (.o(net1170));
 b15tilo00an1n03x5 gen_filter_29__u_filter_diff_ctr_q_reg_2__gen_filter_29__u_filter_diff_ctr_q_reg_3__1171 (.o(net1171));
 b15tilo00an1n03x5 gen_filter_29__u_filter_filter_q_reg_1172 (.o(net1172));
 b15tilo00an1n03x5 gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1173 (.o(net1173));
 b15tilo00an1n03x5 gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1174 (.o(net1174));
 b15tilo00an1n03x5 gen_filter_29__u_filter_stored_value_q_reg_1175 (.o(net1175));
 b15tilo00an1n03x5 gen_filter_2__u_filter_diff_ctr_q_reg_0__gen_filter_2__u_filter_diff_ctr_q_reg_1__1176 (.o(net1176));
 b15tilo00an1n03x5 gen_filter_2__u_filter_diff_ctr_q_reg_0__gen_filter_2__u_filter_diff_ctr_q_reg_1__1177 (.o(net1177));
 b15tilo00an1n03x5 gen_filter_2__u_filter_diff_ctr_q_reg_2__gen_filter_2__u_filter_diff_ctr_q_reg_3__1178 (.o(net1178));
 b15tilo00an1n03x5 gen_filter_2__u_filter_diff_ctr_q_reg_2__gen_filter_2__u_filter_diff_ctr_q_reg_3__1179 (.o(net1179));
 b15tilo00an1n03x5 gen_filter_2__u_filter_filter_q_reg_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1180 (.o(net1180));
 b15tilo00an1n03x5 gen_filter_2__u_filter_filter_q_reg_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1181 (.o(net1181));
 b15tilo00an1n03x5 gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_3__u_filter_diff_ctr_q_reg_0__1182 (.o(net1182));
 b15tilo00an1n03x5 gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_3__u_filter_diff_ctr_q_reg_0__1183 (.o(net1183));
 b15tilo00an1n03x5 gen_filter_2__u_filter_stored_value_q_reg_1184 (.o(net1184));
 b15tilo00an1n03x5 gen_filter_30__u_filter_diff_ctr_q_reg_2__gen_filter_30__u_filter_diff_ctr_q_reg_3__1185 (.o(net1185));
 b15tilo00an1n03x5 gen_filter_30__u_filter_diff_ctr_q_reg_2__gen_filter_30__u_filter_diff_ctr_q_reg_3__1186 (.o(net1186));
 b15tilo00an1n03x5 gen_filter_30__u_filter_filter_q_reg_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1187 (.o(net1187));
 b15tilo00an1n03x5 gen_filter_30__u_filter_filter_q_reg_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1188 (.o(net1188));
 b15tilo00an1n03x5 gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1189 (.o(net1189));
 b15tilo00an1n03x5 gen_filter_30__u_filter_stored_value_q_reg_1190 (.o(net1190));
 b15tilo00an1n03x5 gen_filter_31__u_filter_diff_ctr_q_reg_2__gen_filter_31__u_filter_diff_ctr_q_reg_3__1191 (.o(net1191));
 b15tilo00an1n03x5 gen_filter_31__u_filter_diff_ctr_q_reg_2__gen_filter_31__u_filter_diff_ctr_q_reg_3__1192 (.o(net1192));
 b15tilo00an1n03x5 gen_filter_31__u_filter_filter_q_reg_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1193 (.o(net1193));
 b15tilo00an1n03x5 gen_filter_31__u_filter_filter_q_reg_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1194 (.o(net1194));
 b15tilo00an1n03x5 gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_reg_err_q_reg_1195 (.o(net1195));
 b15tilo00an1n03x5 gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_reg_err_q_reg_1196 (.o(net1196));
 b15tilo00an1n03x5 gen_filter_31__u_filter_stored_value_q_reg_1197 (.o(net1197));
 b15tilo00an1n03x5 gen_filter_3__u_filter_diff_ctr_q_reg_1__gen_filter_3__u_filter_diff_ctr_q_reg_2__1198 (.o(net1198));
 b15tilo00an1n03x5 gen_filter_3__u_filter_diff_ctr_q_reg_1__gen_filter_3__u_filter_diff_ctr_q_reg_2__1199 (.o(net1199));
 b15tilo00an1n03x5 gen_filter_3__u_filter_diff_ctr_q_reg_3__gen_filter_3__u_filter_filter_q_reg_1200 (.o(net1200));
 b15tilo00an1n03x5 gen_filter_3__u_filter_diff_ctr_q_reg_3__gen_filter_3__u_filter_filter_q_reg_1201 (.o(net1201));
 b15tilo00an1n03x5 gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_4__u_filter_diff_ctr_q_reg_1__1202 (.o(net1202));
 b15tilo00an1n03x5 gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_4__u_filter_diff_ctr_q_reg_1__1203 (.o(net1203));
 b15tilo00an1n03x5 gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_8__u_filter_diff_ctr_q_reg_0__1204 (.o(net1204));
 b15tilo00an1n03x5 gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_8__u_filter_diff_ctr_q_reg_0__1205 (.o(net1205));
 b15tilo00an1n03x5 gen_filter_3__u_filter_stored_value_q_reg_1206 (.o(net1206));
 b15tilo00an1n03x5 gen_filter_4__u_filter_diff_ctr_q_reg_0__gen_filter_4__u_filter_diff_ctr_q_reg_2__1207 (.o(net1207));
 b15tilo00an1n03x5 gen_filter_4__u_filter_diff_ctr_q_reg_0__gen_filter_4__u_filter_diff_ctr_q_reg_2__1208 (.o(net1208));
 b15tilo00an1n03x5 gen_filter_4__u_filter_diff_ctr_q_reg_3__gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1209 (.o(net1209));
 b15tilo00an1n03x5 gen_filter_4__u_filter_diff_ctr_q_reg_3__gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1210 (.o(net1210));
 b15tilo00an1n03x5 gen_filter_4__u_filter_filter_q_reg_gen_filter_7__u_filter_filter_q_reg_1211 (.o(net1211));
 b15tilo00an1n03x5 gen_filter_4__u_filter_filter_q_reg_gen_filter_7__u_filter_filter_q_reg_1212 (.o(net1212));
 b15tilo00an1n03x5 gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_7__u_filter_diff_ctr_q_reg_0__1213 (.o(net1213));
 b15tilo00an1n03x5 gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_7__u_filter_diff_ctr_q_reg_0__1214 (.o(net1214));
 b15tilo00an1n03x5 gen_filter_4__u_filter_stored_value_q_reg_1215 (.o(net1215));
 b15tilo00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_0__gen_filter_5__u_filter_diff_ctr_q_reg_1__1216 (.o(net1216));
 b15tilo00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_0__gen_filter_5__u_filter_diff_ctr_q_reg_1__1217 (.o(net1217));
 b15tilo00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_2__gen_filter_5__u_filter_diff_ctr_q_reg_3__1218 (.o(net1218));
 b15tilo00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_2__gen_filter_5__u_filter_diff_ctr_q_reg_3__1219 (.o(net1219));
 b15tilo00an1n03x5 gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_diff_ctr_q_reg_0__1220 (.o(net1220));
 b15tilo00an1n03x5 gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_diff_ctr_q_reg_0__1221 (.o(net1221));
 b15tilo00an1n03x5 gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_filter_q_reg_1222 (.o(net1222));
 b15tilo00an1n03x5 gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_filter_q_reg_1223 (.o(net1223));
 b15tilo00an1n03x5 gen_filter_5__u_filter_stored_value_q_reg_1224 (.o(net1224));
 b15tilo00an1n03x5 gen_filter_6__u_filter_diff_ctr_q_reg_1__gen_filter_6__u_filter_diff_ctr_q_reg_2__1225 (.o(net1225));
 b15tilo00an1n03x5 gen_filter_6__u_filter_diff_ctr_q_reg_1__gen_filter_6__u_filter_diff_ctr_q_reg_2__1226 (.o(net1226));
 b15tilo00an1n03x5 gen_filter_6__u_filter_diff_ctr_q_reg_3__gen_filter_15__u_filter_diff_ctr_q_reg_0__1227 (.o(net1227));
 b15tilo00an1n03x5 gen_filter_6__u_filter_diff_ctr_q_reg_3__gen_filter_15__u_filter_diff_ctr_q_reg_0__1228 (.o(net1228));
 b15tilo00an1n03x5 gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1229 (.o(net1229));
 b15tilo00an1n03x5 gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1230 (.o(net1230));
 b15tilo00an1n03x5 gen_filter_6__u_filter_stored_value_q_reg_1231 (.o(net1231));
 b15tilo00an1n03x5 gen_filter_7__u_filter_diff_ctr_q_reg_1__gen_filter_7__u_filter_diff_ctr_q_reg_2__1232 (.o(net1232));
 b15tilo00an1n03x5 gen_filter_7__u_filter_diff_ctr_q_reg_1__gen_filter_7__u_filter_diff_ctr_q_reg_2__1233 (.o(net1233));
 b15tilo00an1n03x5 gen_filter_7__u_filter_diff_ctr_q_reg_3__gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1234 (.o(net1234));
 b15tilo00an1n03x5 gen_filter_7__u_filter_diff_ctr_q_reg_3__gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1235 (.o(net1235));
 b15tilo00an1n03x5 gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_9__u_filter_diff_ctr_q_reg_0__1236 (.o(net1236));
 b15tilo00an1n03x5 gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_9__u_filter_diff_ctr_q_reg_0__1237 (.o(net1237));
 b15tilo00an1n03x5 gen_filter_7__u_filter_stored_value_q_reg_1238 (.o(net1238));
 b15tilo00an1n03x5 gen_filter_8__u_filter_diff_ctr_q_reg_1__gen_filter_8__u_filter_diff_ctr_q_reg_2__1239 (.o(net1239));
 b15tilo00an1n03x5 gen_filter_8__u_filter_diff_ctr_q_reg_1__gen_filter_8__u_filter_diff_ctr_q_reg_2__1240 (.o(net1240));
 b15tilo00an1n03x5 gen_filter_8__u_filter_diff_ctr_q_reg_3__gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1241 (.o(net1241));
 b15tilo00an1n03x5 gen_filter_8__u_filter_diff_ctr_q_reg_3__gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1242 (.o(net1242));
 b15tilo00an1n03x5 gen_filter_8__u_filter_filter_q_reg_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1243 (.o(net1243));
 b15tilo00an1n03x5 gen_filter_8__u_filter_filter_q_reg_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1244 (.o(net1244));
 b15tilo00an1n03x5 gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_diff_ctr_q_reg_2__1245 (.o(net1245));
 b15tilo00an1n03x5 gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_diff_ctr_q_reg_2__1246 (.o(net1246));
 b15tilo00an1n03x5 gen_filter_8__u_filter_stored_value_q_reg_1247 (.o(net1247));
 b15tilo00an1n03x5 gen_filter_9__u_filter_diff_ctr_q_reg_1__gen_filter_9__u_filter_diff_ctr_q_reg_2__1248 (.o(net1248));
 b15tilo00an1n03x5 gen_filter_9__u_filter_diff_ctr_q_reg_1__gen_filter_9__u_filter_diff_ctr_q_reg_2__1249 (.o(net1249));
 b15tilo00an1n03x5 gen_filter_9__u_filter_diff_ctr_q_reg_3__gen_filter_9__u_filter_filter_q_reg_1250 (.o(net1250));
 b15tilo00an1n03x5 gen_filter_9__u_filter_diff_ctr_q_reg_3__gen_filter_9__u_filter_filter_q_reg_1251 (.o(net1251));
 b15tilo00an1n03x5 gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1252 (.o(net1252));
 b15tilo00an1n03x5 gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1253 (.o(net1253));
 b15tilo00an1n03x5 gen_filter_9__u_filter_stored_value_q_reg_1254 (.o(net1254));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_10__intr_hw_intr_o_reg_11__1255 (.o(net1255));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_10__intr_hw_intr_o_reg_11__1256 (.o(net1256));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_12__intr_hw_intr_o_reg_14__1257 (.o(net1257));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_12__intr_hw_intr_o_reg_14__1258 (.o(net1258));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_15__intr_hw_intr_o_reg_25__1259 (.o(net1259));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_15__intr_hw_intr_o_reg_25__1260 (.o(net1260));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_16__intr_hw_intr_o_reg_17__1261 (.o(net1261));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_16__intr_hw_intr_o_reg_17__1262 (.o(net1262));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_18__intr_hw_intr_o_reg_19__1263 (.o(net1263));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_18__intr_hw_intr_o_reg_19__1264 (.o(net1264));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_1__intr_hw_intr_o_reg_2__1265 (.o(net1265));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_1__intr_hw_intr_o_reg_2__1266 (.o(net1266));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_20__intr_hw_intr_o_reg_21__1267 (.o(net1267));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_20__intr_hw_intr_o_reg_21__1268 (.o(net1268));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_22__intr_hw_intr_o_reg_23__1269 (.o(net1269));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_22__intr_hw_intr_o_reg_23__1270 (.o(net1270));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_24__intr_hw_intr_o_reg_26__1271 (.o(net1271));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_24__intr_hw_intr_o_reg_26__1272 (.o(net1272));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_27__intr_hw_intr_o_reg_28__1273 (.o(net1273));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_27__intr_hw_intr_o_reg_28__1274 (.o(net1274));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_29__intr_hw_intr_o_reg_30__1275 (.o(net1275));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_29__intr_hw_intr_o_reg_30__1276 (.o(net1276));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_31__u_reg_u_data_in_q_reg_1__1277 (.o(net1277));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_31__u_reg_u_data_in_q_reg_1__1278 (.o(net1278));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_3__intr_hw_intr_o_reg_4__1279 (.o(net1279));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_3__intr_hw_intr_o_reg_4__1280 (.o(net1280));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_5__intr_hw_intr_o_reg_6__1281 (.o(net1281));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_5__intr_hw_intr_o_reg_6__1282 (.o(net1282));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_7__intr_hw_intr_o_reg_8__1283 (.o(net1283));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_7__intr_hw_intr_o_reg_8__1284 (.o(net1284));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_9__intr_hw_intr_o_reg_13__1285 (.o(net1285));
 b15tilo00an1n03x5 intr_hw_intr_o_reg_9__intr_hw_intr_o_reg_13__1286 (.o(net1286));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_clk_gate_q_reg_0_latch_1287 (.o(net1287));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_clk_gate_q_reg_latch_1288 (.o(net1288));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_0__u_reg_u_ctrl_en_input_filter_q_reg_1__1289 (.o(net1289));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_0__u_reg_u_ctrl_en_input_filter_q_reg_1__1290 (.o(net1290));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_10__u_reg_u_ctrl_en_input_filter_q_reg_11__1291 (.o(net1291));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_10__u_reg_u_ctrl_en_input_filter_q_reg_11__1292 (.o(net1292));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_12__u_reg_u_ctrl_en_input_filter_q_reg_13__1293 (.o(net1293));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_12__u_reg_u_ctrl_en_input_filter_q_reg_13__1294 (.o(net1294));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_14__u_reg_u_ctrl_en_input_filter_q_reg_15__1295 (.o(net1295));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_14__u_reg_u_ctrl_en_input_filter_q_reg_15__1296 (.o(net1296));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_16__u_reg_u_ctrl_en_input_filter_q_reg_17__1297 (.o(net1297));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_16__u_reg_u_ctrl_en_input_filter_q_reg_17__1298 (.o(net1298));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_18__u_reg_u_ctrl_en_input_filter_q_reg_19__1299 (.o(net1299));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_18__u_reg_u_ctrl_en_input_filter_q_reg_19__1300 (.o(net1300));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_20__u_reg_u_ctrl_en_input_filter_q_reg_21__1301 (.o(net1301));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_20__u_reg_u_ctrl_en_input_filter_q_reg_21__1302 (.o(net1302));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_22__u_reg_u_ctrl_en_input_filter_q_reg_23__1303 (.o(net1303));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_22__u_reg_u_ctrl_en_input_filter_q_reg_23__1304 (.o(net1304));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_24__u_reg_u_ctrl_en_input_filter_q_reg_25__1305 (.o(net1305));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_24__u_reg_u_ctrl_en_input_filter_q_reg_25__1306 (.o(net1306));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_26__u_reg_u_ctrl_en_input_filter_q_reg_27__1307 (.o(net1307));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_26__u_reg_u_ctrl_en_input_filter_q_reg_27__1308 (.o(net1308));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_28__u_reg_u_ctrl_en_input_filter_q_reg_29__1309 (.o(net1309));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_28__u_reg_u_ctrl_en_input_filter_q_reg_29__1310 (.o(net1310));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_2__u_reg_u_ctrl_en_input_filter_q_reg_3__1311 (.o(net1311));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_2__u_reg_u_ctrl_en_input_filter_q_reg_3__1312 (.o(net1312));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_30__u_reg_u_ctrl_en_input_filter_q_reg_31__1313 (.o(net1313));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_30__u_reg_u_ctrl_en_input_filter_q_reg_31__1314 (.o(net1314));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_4__u_reg_u_ctrl_en_input_filter_q_reg_5__1315 (.o(net1315));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_4__u_reg_u_ctrl_en_input_filter_q_reg_5__1316 (.o(net1316));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_6__u_reg_u_ctrl_en_input_filter_q_reg_7__1317 (.o(net1317));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_6__u_reg_u_ctrl_en_input_filter_q_reg_7__1318 (.o(net1318));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_8__u_reg_u_ctrl_en_input_filter_q_reg_9__1319 (.o(net1319));
 b15tilo00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_8__u_reg_u_ctrl_en_input_filter_q_reg_9__1320 (.o(net1320));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_0__u_reg_u_data_in_q_reg_3__1321 (.o(net1321));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_0__u_reg_u_data_in_q_reg_3__1322 (.o(net1322));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_10__u_reg_u_data_in_q_reg_14__1323 (.o(net1323));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_10__u_reg_u_data_in_q_reg_14__1324 (.o(net1324));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_11__u_reg_u_data_in_q_reg_12__1325 (.o(net1325));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_11__u_reg_u_data_in_q_reg_12__1326 (.o(net1326));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_13__u_reg_u_reg_if_rspop_reg_1__1327 (.o(net1327));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_13__u_reg_u_reg_if_rspop_reg_1__1328 (.o(net1328));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_15__u_reg_u_data_in_q_reg_20__1329 (.o(net1329));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_15__u_reg_u_data_in_q_reg_20__1330 (.o(net1330));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_16__u_reg_u_data_in_q_reg_17__1331 (.o(net1331));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_16__u_reg_u_data_in_q_reg_17__1332 (.o(net1332));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_18__u_reg_u_data_in_q_reg_19__1333 (.o(net1333));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_18__u_reg_u_data_in_q_reg_19__1334 (.o(net1334));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_21__u_reg_u_data_in_q_reg_22__1335 (.o(net1335));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_21__u_reg_u_data_in_q_reg_22__1336 (.o(net1336));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_23__1337 (.o(net1337));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_24__u_reg_u_data_in_q_reg_25__1338 (.o(net1338));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_24__u_reg_u_data_in_q_reg_25__1339 (.o(net1339));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_26__1340 (.o(net1340));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_27__u_reg_u_data_in_q_reg_28__1341 (.o(net1341));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_27__u_reg_u_data_in_q_reg_28__1342 (.o(net1342));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_29__u_reg_u_data_in_q_reg_30__1343 (.o(net1343));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_29__u_reg_u_data_in_q_reg_30__1344 (.o(net1344));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_2__1345 (.o(net1345));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_31__1346 (.o(net1346));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_4__u_reg_u_data_in_q_reg_5__1347 (.o(net1347));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_4__u_reg_u_data_in_q_reg_5__1348 (.o(net1348));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_6__u_reg_u_data_in_q_reg_7__1349 (.o(net1349));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_6__u_reg_u_data_in_q_reg_7__1350 (.o(net1350));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_8__u_reg_u_data_in_q_reg_9__1351 (.o(net1351));
 b15tilo00an1n03x5 u_reg_u_data_in_q_reg_8__u_reg_u_data_in_q_reg_9__1352 (.o(net1352));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_clk_gate_q_reg_0_latch_1353 (.o(net1353));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_clk_gate_q_reg_latch_1354 (.o(net1354));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_0__u_reg_u_intr_ctrl_en_falling_q_reg_1__1355 (.o(net1355));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_0__u_reg_u_intr_ctrl_en_falling_q_reg_1__1356 (.o(net1356));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_10__u_reg_u_intr_ctrl_en_falling_q_reg_11__1357 (.o(net1357));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_10__u_reg_u_intr_ctrl_en_falling_q_reg_11__1358 (.o(net1358));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_12__u_reg_u_intr_ctrl_en_falling_q_reg_13__1359 (.o(net1359));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_12__u_reg_u_intr_ctrl_en_falling_q_reg_13__1360 (.o(net1360));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_14__u_reg_u_intr_ctrl_en_falling_q_reg_15__1361 (.o(net1361));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_14__u_reg_u_intr_ctrl_en_falling_q_reg_15__1362 (.o(net1362));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_16__u_reg_u_intr_ctrl_en_falling_q_reg_17__1363 (.o(net1363));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_16__u_reg_u_intr_ctrl_en_falling_q_reg_17__1364 (.o(net1364));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_18__u_reg_u_intr_ctrl_en_falling_q_reg_19__1365 (.o(net1365));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_18__u_reg_u_intr_ctrl_en_falling_q_reg_19__1366 (.o(net1366));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_20__u_reg_u_intr_ctrl_en_falling_q_reg_21__1367 (.o(net1367));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_20__u_reg_u_intr_ctrl_en_falling_q_reg_21__1368 (.o(net1368));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_22__u_reg_u_intr_ctrl_en_falling_q_reg_23__1369 (.o(net1369));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_22__u_reg_u_intr_ctrl_en_falling_q_reg_23__1370 (.o(net1370));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_24__u_reg_u_intr_ctrl_en_falling_q_reg_25__1371 (.o(net1371));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_24__u_reg_u_intr_ctrl_en_falling_q_reg_25__1372 (.o(net1372));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_26__u_reg_u_intr_ctrl_en_falling_q_reg_27__1373 (.o(net1373));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_26__u_reg_u_intr_ctrl_en_falling_q_reg_27__1374 (.o(net1374));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_28__u_reg_u_intr_ctrl_en_falling_q_reg_29__1375 (.o(net1375));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_28__u_reg_u_intr_ctrl_en_falling_q_reg_29__1376 (.o(net1376));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_2__u_reg_u_intr_ctrl_en_falling_q_reg_3__1377 (.o(net1377));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_2__u_reg_u_intr_ctrl_en_falling_q_reg_3__1378 (.o(net1378));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_30__u_reg_u_intr_ctrl_en_falling_q_reg_31__1379 (.o(net1379));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_30__u_reg_u_intr_ctrl_en_falling_q_reg_31__1380 (.o(net1380));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_4__u_reg_u_intr_ctrl_en_falling_q_reg_5__1381 (.o(net1381));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_4__u_reg_u_intr_ctrl_en_falling_q_reg_5__1382 (.o(net1382));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_6__u_reg_u_intr_ctrl_en_falling_q_reg_7__1383 (.o(net1383));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_6__u_reg_u_intr_ctrl_en_falling_q_reg_7__1384 (.o(net1384));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_8__u_reg_u_intr_ctrl_en_falling_q_reg_9__1385 (.o(net1385));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_8__u_reg_u_intr_ctrl_en_falling_q_reg_9__1386 (.o(net1386));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_clk_gate_q_reg_0_latch_1387 (.o(net1387));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_clk_gate_q_reg_latch_1388 (.o(net1388));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_0__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_1__1389 (.o(net1389));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_0__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_1__1390 (.o(net1390));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_10__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_11__1391 (.o(net1391));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_10__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_11__1392 (.o(net1392));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_12__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_13__1393 (.o(net1393));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_12__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_13__1394 (.o(net1394));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_14__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_15__1395 (.o(net1395));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_14__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_15__1396 (.o(net1396));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_16__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_17__1397 (.o(net1397));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_16__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_17__1398 (.o(net1398));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_18__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_19__1399 (.o(net1399));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_18__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_19__1400 (.o(net1400));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_20__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_21__1401 (.o(net1401));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_20__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_21__1402 (.o(net1402));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_22__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_23__1403 (.o(net1403));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_22__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_23__1404 (.o(net1404));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_24__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_25__1405 (.o(net1405));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_24__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_25__1406 (.o(net1406));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_26__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_27__1407 (.o(net1407));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_26__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_27__1408 (.o(net1408));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_28__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_29__1409 (.o(net1409));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_28__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_29__1410 (.o(net1410));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_2__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_3__1411 (.o(net1411));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_2__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_3__1412 (.o(net1412));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_30__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_31__1413 (.o(net1413));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_30__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_31__1414 (.o(net1414));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_4__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_5__1415 (.o(net1415));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_4__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_5__1416 (.o(net1416));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_6__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_7__1417 (.o(net1417));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_6__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_7__1418 (.o(net1418));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_8__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_9__1419 (.o(net1419));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_8__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_9__1420 (.o(net1420));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_clk_gate_q_reg_0_latch_1421 (.o(net1421));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_clk_gate_q_reg_latch_1422 (.o(net1422));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_0__u_reg_u_intr_ctrl_en_lvllow_q_reg_1__1423 (.o(net1423));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_0__u_reg_u_intr_ctrl_en_lvllow_q_reg_1__1424 (.o(net1424));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_10__u_reg_u_intr_ctrl_en_lvllow_q_reg_11__1425 (.o(net1425));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_10__u_reg_u_intr_ctrl_en_lvllow_q_reg_11__1426 (.o(net1426));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_12__u_reg_u_intr_ctrl_en_lvllow_q_reg_13__1427 (.o(net1427));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_12__u_reg_u_intr_ctrl_en_lvllow_q_reg_13__1428 (.o(net1428));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_14__u_reg_u_intr_ctrl_en_lvllow_q_reg_15__1429 (.o(net1429));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_14__u_reg_u_intr_ctrl_en_lvllow_q_reg_15__1430 (.o(net1430));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_16__u_reg_u_intr_ctrl_en_lvllow_q_reg_17__1431 (.o(net1431));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_16__u_reg_u_intr_ctrl_en_lvllow_q_reg_17__1432 (.o(net1432));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_18__u_reg_u_intr_ctrl_en_lvllow_q_reg_19__1433 (.o(net1433));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_18__u_reg_u_intr_ctrl_en_lvllow_q_reg_19__1434 (.o(net1434));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_20__u_reg_u_intr_ctrl_en_lvllow_q_reg_21__1435 (.o(net1435));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_20__u_reg_u_intr_ctrl_en_lvllow_q_reg_21__1436 (.o(net1436));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_22__u_reg_u_intr_ctrl_en_lvllow_q_reg_23__1437 (.o(net1437));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_22__u_reg_u_intr_ctrl_en_lvllow_q_reg_23__1438 (.o(net1438));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_24__u_reg_u_intr_ctrl_en_lvllow_q_reg_25__1439 (.o(net1439));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_24__u_reg_u_intr_ctrl_en_lvllow_q_reg_25__1440 (.o(net1440));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_26__u_reg_u_intr_ctrl_en_lvllow_q_reg_27__1441 (.o(net1441));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_26__u_reg_u_intr_ctrl_en_lvllow_q_reg_27__1442 (.o(net1442));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_28__u_reg_u_intr_ctrl_en_lvllow_q_reg_29__1443 (.o(net1443));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_28__u_reg_u_intr_ctrl_en_lvllow_q_reg_29__1444 (.o(net1444));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_2__u_reg_u_intr_ctrl_en_lvllow_q_reg_3__1445 (.o(net1445));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_2__u_reg_u_intr_ctrl_en_lvllow_q_reg_3__1446 (.o(net1446));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_30__u_reg_u_intr_ctrl_en_lvllow_q_reg_31__1447 (.o(net1447));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_30__u_reg_u_intr_ctrl_en_lvllow_q_reg_31__1448 (.o(net1448));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_4__u_reg_u_intr_ctrl_en_lvllow_q_reg_5__1449 (.o(net1449));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_4__u_reg_u_intr_ctrl_en_lvllow_q_reg_5__1450 (.o(net1450));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_6__u_reg_u_intr_ctrl_en_lvllow_q_reg_7__1451 (.o(net1451));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_6__u_reg_u_intr_ctrl_en_lvllow_q_reg_7__1452 (.o(net1452));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_8__u_reg_u_intr_ctrl_en_lvllow_q_reg_9__1453 (.o(net1453));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_8__u_reg_u_intr_ctrl_en_lvllow_q_reg_9__1454 (.o(net1454));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_clk_gate_q_reg_0_latch_1455 (.o(net1455));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_clk_gate_q_reg_latch_1456 (.o(net1456));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_0__u_reg_u_intr_ctrl_en_rising_q_reg_1__1457 (.o(net1457));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_0__u_reg_u_intr_ctrl_en_rising_q_reg_1__1458 (.o(net1458));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_10__u_reg_u_intr_ctrl_en_rising_q_reg_11__1459 (.o(net1459));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_10__u_reg_u_intr_ctrl_en_rising_q_reg_11__1460 (.o(net1460));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_12__u_reg_u_intr_ctrl_en_rising_q_reg_13__1461 (.o(net1461));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_12__u_reg_u_intr_ctrl_en_rising_q_reg_13__1462 (.o(net1462));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_14__u_reg_u_intr_ctrl_en_rising_q_reg_15__1463 (.o(net1463));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_14__u_reg_u_intr_ctrl_en_rising_q_reg_15__1464 (.o(net1464));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_16__u_reg_u_intr_ctrl_en_rising_q_reg_17__1465 (.o(net1465));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_16__u_reg_u_intr_ctrl_en_rising_q_reg_17__1466 (.o(net1466));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_18__u_reg_u_intr_ctrl_en_rising_q_reg_19__1467 (.o(net1467));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_18__u_reg_u_intr_ctrl_en_rising_q_reg_19__1468 (.o(net1468));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_20__u_reg_u_intr_ctrl_en_rising_q_reg_21__1469 (.o(net1469));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_20__u_reg_u_intr_ctrl_en_rising_q_reg_21__1470 (.o(net1470));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_22__u_reg_u_intr_ctrl_en_rising_q_reg_23__1471 (.o(net1471));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_22__u_reg_u_intr_ctrl_en_rising_q_reg_23__1472 (.o(net1472));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_24__u_reg_u_intr_ctrl_en_rising_q_reg_25__1473 (.o(net1473));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_24__u_reg_u_intr_ctrl_en_rising_q_reg_25__1474 (.o(net1474));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_26__u_reg_u_intr_ctrl_en_rising_q_reg_27__1475 (.o(net1475));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_26__u_reg_u_intr_ctrl_en_rising_q_reg_27__1476 (.o(net1476));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_28__u_reg_u_intr_ctrl_en_rising_q_reg_29__1477 (.o(net1477));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_28__u_reg_u_intr_ctrl_en_rising_q_reg_29__1478 (.o(net1478));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_2__u_reg_u_intr_ctrl_en_rising_q_reg_3__1479 (.o(net1479));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_2__u_reg_u_intr_ctrl_en_rising_q_reg_3__1480 (.o(net1480));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_30__u_reg_u_intr_ctrl_en_rising_q_reg_31__1481 (.o(net1481));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_30__u_reg_u_intr_ctrl_en_rising_q_reg_31__1482 (.o(net1482));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_4__u_reg_u_intr_ctrl_en_rising_q_reg_5__1483 (.o(net1483));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_4__u_reg_u_intr_ctrl_en_rising_q_reg_5__1484 (.o(net1484));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_6__u_reg_u_intr_ctrl_en_rising_q_reg_7__1485 (.o(net1485));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_6__u_reg_u_intr_ctrl_en_rising_q_reg_7__1486 (.o(net1486));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_8__u_reg_u_intr_ctrl_en_rising_q_reg_9__1487 (.o(net1487));
 b15tilo00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_8__u_reg_u_intr_ctrl_en_rising_q_reg_9__1488 (.o(net1488));
 b15tilo00an1n03x5 u_reg_u_intr_enable_clk_gate_q_reg_0_latch_1489 (.o(net1489));
 b15tilo00an1n03x5 u_reg_u_intr_enable_clk_gate_q_reg_latch_1490 (.o(net1490));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_0__u_reg_u_intr_enable_q_reg_1__1491 (.o(net1491));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_0__u_reg_u_intr_enable_q_reg_1__1492 (.o(net1492));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_10__u_reg_u_intr_enable_q_reg_11__1493 (.o(net1493));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_10__u_reg_u_intr_enable_q_reg_11__1494 (.o(net1494));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_12__u_reg_u_intr_enable_q_reg_13__1495 (.o(net1495));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_12__u_reg_u_intr_enable_q_reg_13__1496 (.o(net1496));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_14__u_reg_u_intr_enable_q_reg_15__1497 (.o(net1497));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_14__u_reg_u_intr_enable_q_reg_15__1498 (.o(net1498));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_16__u_reg_u_intr_enable_q_reg_17__1499 (.o(net1499));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_16__u_reg_u_intr_enable_q_reg_17__1500 (.o(net1500));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_18__u_reg_u_intr_enable_q_reg_19__1501 (.o(net1501));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_18__u_reg_u_intr_enable_q_reg_19__1502 (.o(net1502));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_20__u_reg_u_intr_enable_q_reg_21__1503 (.o(net1503));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_20__u_reg_u_intr_enable_q_reg_21__1504 (.o(net1504));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_22__u_reg_u_intr_enable_q_reg_23__1505 (.o(net1505));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_22__u_reg_u_intr_enable_q_reg_23__1506 (.o(net1506));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_24__u_reg_u_intr_enable_q_reg_25__1507 (.o(net1507));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_24__u_reg_u_intr_enable_q_reg_25__1508 (.o(net1508));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_26__u_reg_u_intr_enable_q_reg_27__1509 (.o(net1509));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_26__u_reg_u_intr_enable_q_reg_27__1510 (.o(net1510));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_28__u_reg_u_intr_enable_q_reg_29__1511 (.o(net1511));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_28__u_reg_u_intr_enable_q_reg_29__1512 (.o(net1512));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_2__u_reg_u_intr_enable_q_reg_3__1513 (.o(net1513));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_2__u_reg_u_intr_enable_q_reg_3__1514 (.o(net1514));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_30__u_reg_u_intr_enable_q_reg_31__1515 (.o(net1515));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_30__u_reg_u_intr_enable_q_reg_31__1516 (.o(net1516));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_4__u_reg_u_intr_enable_q_reg_5__1517 (.o(net1517));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_4__u_reg_u_intr_enable_q_reg_5__1518 (.o(net1518));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_6__u_reg_u_intr_enable_q_reg_7__1519 (.o(net1519));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_6__u_reg_u_intr_enable_q_reg_7__1520 (.o(net1520));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_8__u_reg_u_intr_enable_q_reg_9__1521 (.o(net1521));
 b15tilo00an1n03x5 u_reg_u_intr_enable_q_reg_8__u_reg_u_intr_enable_q_reg_9__1522 (.o(net1522));
 b15tilo00an1n03x5 u_reg_u_intr_state_clk_gate_q_reg_0_latch_1523 (.o(net1523));
 b15tilo00an1n03x5 u_reg_u_intr_state_clk_gate_q_reg_latch_1524 (.o(net1524));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_0__u_reg_u_intr_state_q_reg_1__1525 (.o(net1525));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_0__u_reg_u_intr_state_q_reg_1__1526 (.o(net1526));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_10__u_reg_u_intr_state_q_reg_11__1527 (.o(net1527));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_10__u_reg_u_intr_state_q_reg_11__1528 (.o(net1528));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_12__u_reg_u_intr_state_q_reg_13__1529 (.o(net1529));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_12__u_reg_u_intr_state_q_reg_13__1530 (.o(net1530));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_14__u_reg_u_intr_state_q_reg_15__1531 (.o(net1531));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_14__u_reg_u_intr_state_q_reg_15__1532 (.o(net1532));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_16__u_reg_u_intr_state_q_reg_17__1533 (.o(net1533));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_16__u_reg_u_intr_state_q_reg_17__1534 (.o(net1534));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_18__u_reg_u_intr_state_q_reg_19__1535 (.o(net1535));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_18__u_reg_u_intr_state_q_reg_19__1536 (.o(net1536));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_20__u_reg_u_intr_state_q_reg_21__1537 (.o(net1537));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_20__u_reg_u_intr_state_q_reg_21__1538 (.o(net1538));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_22__u_reg_u_intr_state_q_reg_23__1539 (.o(net1539));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_22__u_reg_u_intr_state_q_reg_23__1540 (.o(net1540));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_24__u_reg_u_intr_state_q_reg_25__1541 (.o(net1541));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_24__u_reg_u_intr_state_q_reg_25__1542 (.o(net1542));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_26__u_reg_u_intr_state_q_reg_27__1543 (.o(net1543));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_26__u_reg_u_intr_state_q_reg_27__1544 (.o(net1544));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_28__u_reg_u_intr_state_q_reg_29__1545 (.o(net1545));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_28__u_reg_u_intr_state_q_reg_29__1546 (.o(net1546));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_2__u_reg_u_intr_state_q_reg_3__1547 (.o(net1547));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_2__u_reg_u_intr_state_q_reg_3__1548 (.o(net1548));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_30__u_reg_u_intr_state_q_reg_31__1549 (.o(net1549));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_30__u_reg_u_intr_state_q_reg_31__1550 (.o(net1550));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_4__u_reg_u_intr_state_q_reg_5__1551 (.o(net1551));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_4__u_reg_u_intr_state_q_reg_5__1552 (.o(net1552));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_6__u_reg_u_intr_state_q_reg_7__1553 (.o(net1553));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_6__u_reg_u_intr_state_q_reg_7__1554 (.o(net1554));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_8__u_reg_u_intr_state_q_reg_9__1555 (.o(net1555));
 b15tilo00an1n03x5 u_reg_u_intr_state_q_reg_8__u_reg_u_intr_state_q_reg_9__1556 (.o(net1556));
 b15tilo00an1n03x5 u_reg_u_reg_if_clk_gate_rdata_reg_0_latch_1557 (.o(net1557));
 b15tilo00an1n03x5 u_reg_u_reg_if_clk_gate_rdata_reg_latch_1558 (.o(net1558));
 b15tilo00an1n03x5 u_reg_u_reg_if_clk_gate_reqid_reg_latch_1559 (.o(net1559));
 b15tilo00an1n03x5 u_reg_u_reg_if_error_reg_1560 (.o(net1560));
 b15tilo00an1n03x5 u_reg_u_reg_if_outstanding_reg_1561 (.o(net1561));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_0__u_reg_u_reg_if_rdata_reg_1__1562 (.o(net1562));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_0__u_reg_u_reg_if_rdata_reg_1__1563 (.o(net1563));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_10__u_reg_u_reg_if_rdata_reg_11__1564 (.o(net1564));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_10__u_reg_u_reg_if_rdata_reg_11__1565 (.o(net1565));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_12__u_reg_u_reg_if_rdata_reg_13__1566 (.o(net1566));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_12__u_reg_u_reg_if_rdata_reg_13__1567 (.o(net1567));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_14__u_reg_u_reg_if_rdata_reg_15__1568 (.o(net1568));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_14__u_reg_u_reg_if_rdata_reg_15__1569 (.o(net1569));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_16__u_reg_u_reg_if_rdata_reg_17__1570 (.o(net1570));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_16__u_reg_u_reg_if_rdata_reg_17__1571 (.o(net1571));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_18__u_reg_u_reg_if_rdata_reg_19__1572 (.o(net1572));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_18__u_reg_u_reg_if_rdata_reg_19__1573 (.o(net1573));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_20__u_reg_u_reg_if_rdata_reg_21__1574 (.o(net1574));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_20__u_reg_u_reg_if_rdata_reg_21__1575 (.o(net1575));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_22__u_reg_u_reg_if_rdata_reg_23__1576 (.o(net1576));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_22__u_reg_u_reg_if_rdata_reg_23__1577 (.o(net1577));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_24__u_reg_u_reg_if_rdata_reg_25__1578 (.o(net1578));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_24__u_reg_u_reg_if_rdata_reg_25__1579 (.o(net1579));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_26__u_reg_u_reg_if_rdata_reg_27__1580 (.o(net1580));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_26__u_reg_u_reg_if_rdata_reg_27__1581 (.o(net1581));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_28__u_reg_u_reg_if_rdata_reg_29__1582 (.o(net1582));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_28__u_reg_u_reg_if_rdata_reg_29__1583 (.o(net1583));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_2__u_reg_u_reg_if_rdata_reg_3__1584 (.o(net1584));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_2__u_reg_u_reg_if_rdata_reg_3__1585 (.o(net1585));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_30__u_reg_u_reg_if_rdata_reg_31__1586 (.o(net1586));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_30__u_reg_u_reg_if_rdata_reg_31__1587 (.o(net1587));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_4__u_reg_u_reg_if_rdata_reg_5__1588 (.o(net1588));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_4__u_reg_u_reg_if_rdata_reg_5__1589 (.o(net1589));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_6__u_reg_u_reg_if_rdata_reg_7__1590 (.o(net1590));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_6__u_reg_u_reg_if_rdata_reg_7__1591 (.o(net1591));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_8__u_reg_u_reg_if_rdata_reg_9__1592 (.o(net1592));
 b15tilo00an1n03x5 u_reg_u_reg_if_rdata_reg_8__u_reg_u_reg_if_rdata_reg_9__1593 (.o(net1593));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_reg_0__u_reg_u_reg_if_reqid_reg_1__1594 (.o(net1594));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_reg_0__u_reg_u_reg_if_reqid_reg_1__1595 (.o(net1595));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_reg_2__u_reg_u_reg_if_reqid_reg_3__1596 (.o(net1596));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_reg_2__u_reg_u_reg_if_reqid_reg_3__1597 (.o(net1597));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_reg_4__u_reg_u_reg_if_reqid_reg_5__1598 (.o(net1598));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_reg_4__u_reg_u_reg_if_reqid_reg_5__1599 (.o(net1599));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_reg_6__u_reg_u_reg_if_reqid_reg_7__1600 (.o(net1600));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqid_reg_6__u_reg_u_reg_if_reqid_reg_7__1601 (.o(net1601));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqsz_reg_0__1602 (.o(net1602));
 b15tilo00an1n03x5 u_reg_u_reg_if_reqsz_reg_1__1603 (.o(net1603));
 b15tilo00an1n03x5 u_reg_u_reg_if_rspop_reg_0__1604 (.o(net1604));
 b15tilo00an1n03x5 u_reg_u_reg_if_rspop_reg_2__1605 (.o(net1605));
 b15tihi00an1n03x5 U3327_1607 (.o(net1607));
 b15tihi00an1n03x5 U3329_1608 (.o(net1608));
 b15tihi00an1n03x5 U3331_1609 (.o(net1609));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_0__cio_gpio_en_q_reg_1__1610 (.o(net1610));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_10__cio_gpio_en_q_reg_11__1611 (.o(net1611));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_12__cio_gpio_en_q_reg_13__1612 (.o(net1612));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_14__cio_gpio_en_q_reg_15__1613 (.o(net1613));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_16__cio_gpio_en_q_reg_17__1614 (.o(net1614));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_18__cio_gpio_en_q_reg_19__1615 (.o(net1615));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_20__cio_gpio_en_q_reg_21__1616 (.o(net1616));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_22__cio_gpio_en_q_reg_23__1617 (.o(net1617));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_24__cio_gpio_en_q_reg_25__1618 (.o(net1618));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_26__cio_gpio_en_q_reg_27__1619 (.o(net1619));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_28__cio_gpio_en_q_reg_29__1620 (.o(net1620));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_2__cio_gpio_en_q_reg_3__1621 (.o(net1621));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_30__cio_gpio_en_q_reg_31__1622 (.o(net1622));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_4__cio_gpio_en_q_reg_5__1623 (.o(net1623));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_6__cio_gpio_en_q_reg_7__1624 (.o(net1624));
 b15tihi00an1n03x5 cio_gpio_en_q_reg_8__cio_gpio_en_q_reg_9__1625 (.o(net1625));
 b15tihi00an1n03x5 cio_gpio_q_reg_0__cio_gpio_q_reg_1__1626 (.o(net1626));
 b15tihi00an1n03x5 cio_gpio_q_reg_10__cio_gpio_q_reg_11__1627 (.o(net1627));
 b15tihi00an1n03x5 cio_gpio_q_reg_12__cio_gpio_q_reg_13__1628 (.o(net1628));
 b15tihi00an1n03x5 cio_gpio_q_reg_14__cio_gpio_q_reg_15__1629 (.o(net1629));
 b15tihi00an1n03x5 cio_gpio_q_reg_16__cio_gpio_q_reg_17__1630 (.o(net1630));
 b15tihi00an1n03x5 cio_gpio_q_reg_18__cio_gpio_q_reg_19__1631 (.o(net1631));
 b15tihi00an1n03x5 cio_gpio_q_reg_20__cio_gpio_q_reg_21__1632 (.o(net1632));
 b15tihi00an1n03x5 cio_gpio_q_reg_22__cio_gpio_q_reg_23__1633 (.o(net1633));
 b15tihi00an1n03x5 cio_gpio_q_reg_24__cio_gpio_q_reg_25__1634 (.o(net1634));
 b15tihi00an1n03x5 cio_gpio_q_reg_26__cio_gpio_q_reg_27__1635 (.o(net1635));
 b15tihi00an1n03x5 cio_gpio_q_reg_28__cio_gpio_q_reg_29__1636 (.o(net1636));
 b15tihi00an1n03x5 cio_gpio_q_reg_2__cio_gpio_q_reg_3__1637 (.o(net1637));
 b15tihi00an1n03x5 cio_gpio_q_reg_30__cio_gpio_q_reg_31__1638 (.o(net1638));
 b15tihi00an1n03x5 cio_gpio_q_reg_4__cio_gpio_q_reg_5__1639 (.o(net1639));
 b15tihi00an1n03x5 cio_gpio_q_reg_6__cio_gpio_q_reg_7__1640 (.o(net1640));
 b15tihi00an1n03x5 cio_gpio_q_reg_8__cio_gpio_q_reg_9__1641 (.o(net1641));
 b15tihi00an1n03x5 data_in_q_reg_0__data_in_q_reg_1__1642 (.o(net1642));
 b15tihi00an1n03x5 data_in_q_reg_10__data_in_q_reg_11__1643 (.o(net1643));
 b15tihi00an1n03x5 data_in_q_reg_12__data_in_q_reg_13__1644 (.o(net1644));
 b15tihi00an1n03x5 data_in_q_reg_14__data_in_q_reg_15__1645 (.o(net1645));
 b15tihi00an1n03x5 data_in_q_reg_16__data_in_q_reg_17__1646 (.o(net1646));
 b15tihi00an1n03x5 data_in_q_reg_18__data_in_q_reg_19__1647 (.o(net1647));
 b15tihi00an1n03x5 data_in_q_reg_20__data_in_q_reg_21__1648 (.o(net1648));
 b15tihi00an1n03x5 data_in_q_reg_22__data_in_q_reg_23__1649 (.o(net1649));
 b15tihi00an1n03x5 data_in_q_reg_24__data_in_q_reg_25__1650 (.o(net1650));
 b15tihi00an1n03x5 data_in_q_reg_26__data_in_q_reg_27__1651 (.o(net1651));
 b15tihi00an1n03x5 data_in_q_reg_28__data_in_q_reg_29__1652 (.o(net1652));
 b15tihi00an1n03x5 data_in_q_reg_2__data_in_q_reg_3__1653 (.o(net1653));
 b15tihi00an1n03x5 data_in_q_reg_30__data_in_q_reg_31__1654 (.o(net1654));
 b15tihi00an1n03x5 data_in_q_reg_4__data_in_q_reg_5__1655 (.o(net1655));
 b15tihi00an1n03x5 data_in_q_reg_6__data_in_q_reg_7__1656 (.o(net1656));
 b15tihi00an1n03x5 data_in_q_reg_8__data_in_q_reg_9__1657 (.o(net1657));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_alert_set_q_reg_gen_filter_5__u_filter_filter_q_reg_1658 (.o(net1658));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_alert_test_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_0__1659 (.o(net1659));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_ping_set_q_reg_gen_alert_tx_0__u_prim_alert_sender_state_q_reg_1__1660 (.o(net1660));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_state_q_reg_2__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_pq_reg_1661 (.o(net1661));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nq_reg_1662 (.o(net1662));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1663 (.o(net1663));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1664 (.o(net1664));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1665 (.o(net1665));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_0__1666 (.o(net1666));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q_reg_1__1667 (.o(net1667));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q_reg_gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pq_reg_1668 (.o(net1668));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nq_reg_1669 (.o(net1669));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1670 (.o(net1670));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1671 (.o(net1671));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1672 (.o(net1672));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_0__1673 (.o(net1673));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q_reg_1__1674 (.o(net1674));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q_reg_gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1675 (.o(net1675));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_0__u_filter_diff_ctr_q_reg_0__1676 (.o(net1676));
 b15tihi00an1n03x5 gen_alert_tx_0__u_prim_alert_sender_u_prim_flop_alert_u_secure_anchor_flop_gen_generic_u_impl_generic_q_o_reg_1__1677 (.o(net1677));
 b15tihi00an1n03x5 gen_filter_0__u_filter_diff_ctr_q_reg_1__gen_filter_0__u_filter_diff_ctr_q_reg_2__1678 (.o(net1678));
 b15tihi00an1n03x5 gen_filter_0__u_filter_diff_ctr_q_reg_3__gen_filter_0__u_filter_filter_q_reg_1679 (.o(net1679));
 b15tihi00an1n03x5 gen_filter_0__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_16__u_filter_diff_ctr_q_reg_0__1680 (.o(net1680));
 b15tihi00an1n03x5 gen_filter_0__u_filter_stored_value_q_reg_1681 (.o(net1681));
 b15tihi00an1n03x5 gen_filter_10__u_filter_diff_ctr_q_reg_0__gen_filter_10__u_filter_diff_ctr_q_reg_3__1682 (.o(net1682));
 b15tihi00an1n03x5 gen_filter_10__u_filter_diff_ctr_q_reg_1__gen_filter_10__u_filter_diff_ctr_q_reg_2__1683 (.o(net1683));
 b15tihi00an1n03x5 gen_filter_10__u_filter_filter_q_reg_gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1684 (.o(net1684));
 b15tihi00an1n03x5 gen_filter_10__u_filter_stored_value_q_reg_1685 (.o(net1685));
 b15tihi00an1n03x5 gen_filter_11__u_filter_diff_ctr_q_reg_0__gen_filter_11__u_filter_diff_ctr_q_reg_1__1686 (.o(net1686));
 b15tihi00an1n03x5 gen_filter_11__u_filter_diff_ctr_q_reg_3__gen_filter_11__u_filter_filter_q_reg_1687 (.o(net1687));
 b15tihi00an1n03x5 gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1688 (.o(net1688));
 b15tihi00an1n03x5 gen_filter_11__u_filter_stored_value_q_reg_1689 (.o(net1689));
 b15tihi00an1n03x5 gen_filter_12__u_filter_diff_ctr_q_reg_0__gen_filter_12__u_filter_diff_ctr_q_reg_1__1690 (.o(net1690));
 b15tihi00an1n03x5 gen_filter_12__u_filter_diff_ctr_q_reg_2__gen_filter_12__u_filter_diff_ctr_q_reg_3__1691 (.o(net1691));
 b15tihi00an1n03x5 gen_filter_12__u_filter_filter_q_reg_gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1692 (.o(net1692));
 b15tihi00an1n03x5 gen_filter_12__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_13__u_filter_diff_ctr_q_reg_0__1693 (.o(net1693));
 b15tihi00an1n03x5 gen_filter_12__u_filter_stored_value_q_reg_1694 (.o(net1694));
 b15tihi00an1n03x5 gen_filter_13__u_filter_diff_ctr_q_reg_1__gen_filter_13__u_filter_diff_ctr_q_reg_2__1695 (.o(net1695));
 b15tihi00an1n03x5 gen_filter_13__u_filter_diff_ctr_q_reg_3__gen_filter_13__u_filter_filter_q_reg_1696 (.o(net1696));
 b15tihi00an1n03x5 gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_13__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1697 (.o(net1697));
 b15tihi00an1n03x5 gen_filter_13__u_filter_stored_value_q_reg_1698 (.o(net1698));
 b15tihi00an1n03x5 gen_filter_14__u_filter_diff_ctr_q_reg_0__gen_filter_14__u_filter_diff_ctr_q_reg_1__1699 (.o(net1699));
 b15tihi00an1n03x5 gen_filter_14__u_filter_diff_ctr_q_reg_2__gen_filter_14__u_filter_diff_ctr_q_reg_3__1700 (.o(net1700));
 b15tihi00an1n03x5 gen_filter_14__u_filter_filter_q_reg_gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1701 (.o(net1701));
 b15tihi00an1n03x5 gen_filter_14__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1702 (.o(net1702));
 b15tihi00an1n03x5 gen_filter_14__u_filter_stored_value_q_reg_1703 (.o(net1703));
 b15tihi00an1n03x5 gen_filter_15__u_filter_diff_ctr_q_reg_1__gen_filter_15__u_filter_diff_ctr_q_reg_2__1704 (.o(net1704));
 b15tihi00an1n03x5 gen_filter_15__u_filter_diff_ctr_q_reg_3__gen_filter_15__u_filter_filter_q_reg_1705 (.o(net1705));
 b15tihi00an1n03x5 gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_15__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1706 (.o(net1706));
 b15tihi00an1n03x5 gen_filter_15__u_filter_stored_value_q_reg_1707 (.o(net1707));
 b15tihi00an1n03x5 gen_filter_16__u_filter_diff_ctr_q_reg_1__gen_filter_16__u_filter_diff_ctr_q_reg_2__1708 (.o(net1708));
 b15tihi00an1n03x5 gen_filter_16__u_filter_diff_ctr_q_reg_3__gen_filter_16__u_filter_filter_q_reg_1709 (.o(net1709));
 b15tihi00an1n03x5 gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_diff_ctr_q_reg_0__1710 (.o(net1710));
 b15tihi00an1n03x5 gen_filter_16__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_30__u_filter_diff_ctr_q_reg_0__1711 (.o(net1711));
 b15tihi00an1n03x5 gen_filter_16__u_filter_stored_value_q_reg_1712 (.o(net1712));
 b15tihi00an1n03x5 gen_filter_17__u_filter_diff_ctr_q_reg_1__gen_filter_17__u_filter_diff_ctr_q_reg_2__1713 (.o(net1713));
 b15tihi00an1n03x5 gen_filter_17__u_filter_diff_ctr_q_reg_3__gen_filter_17__u_filter_filter_q_reg_1714 (.o(net1714));
 b15tihi00an1n03x5 gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_17__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1715 (.o(net1715));
 b15tihi00an1n03x5 gen_filter_17__u_filter_stored_value_q_reg_1716 (.o(net1716));
 b15tihi00an1n03x5 gen_filter_18__u_filter_diff_ctr_q_reg_0__gen_filter_18__u_filter_diff_ctr_q_reg_1__1717 (.o(net1717));
 b15tihi00an1n03x5 gen_filter_18__u_filter_diff_ctr_q_reg_2__gen_filter_18__u_filter_diff_ctr_q_reg_3__1718 (.o(net1718));
 b15tihi00an1n03x5 gen_filter_18__u_filter_filter_q_reg_gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1719 (.o(net1719));
 b15tihi00an1n03x5 gen_filter_18__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_19__u_filter_diff_ctr_q_reg_0__1720 (.o(net1720));
 b15tihi00an1n03x5 gen_filter_18__u_filter_stored_value_q_reg_1721 (.o(net1721));
 b15tihi00an1n03x5 gen_filter_19__u_filter_diff_ctr_q_reg_1__gen_filter_19__u_filter_diff_ctr_q_reg_2__1722 (.o(net1722));
 b15tihi00an1n03x5 gen_filter_19__u_filter_diff_ctr_q_reg_3__gen_filter_19__u_filter_filter_q_reg_1723 (.o(net1723));
 b15tihi00an1n03x5 gen_filter_19__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_21__u_filter_diff_ctr_q_reg_0__1724 (.o(net1724));
 b15tihi00an1n03x5 gen_filter_19__u_filter_stored_value_q_reg_1725 (.o(net1725));
 b15tihi00an1n03x5 gen_filter_1__u_filter_diff_ctr_q_reg_0__gen_filter_1__u_filter_diff_ctr_q_reg_1__1726 (.o(net1726));
 b15tihi00an1n03x5 gen_filter_1__u_filter_diff_ctr_q_reg_2__gen_filter_1__u_filter_diff_ctr_q_reg_3__1727 (.o(net1727));
 b15tihi00an1n03x5 gen_filter_1__u_filter_filter_q_reg_gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1728 (.o(net1728));
 b15tihi00an1n03x5 gen_filter_1__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__intr_hw_intr_o_reg_0__1729 (.o(net1729));
 b15tihi00an1n03x5 gen_filter_1__u_filter_stored_value_q_reg_1730 (.o(net1730));
 b15tihi00an1n03x5 gen_filter_20__u_filter_diff_ctr_q_reg_0__gen_filter_20__u_filter_diff_ctr_q_reg_1__1731 (.o(net1731));
 b15tihi00an1n03x5 gen_filter_20__u_filter_diff_ctr_q_reg_2__gen_filter_20__u_filter_diff_ctr_q_reg_3__1732 (.o(net1732));
 b15tihi00an1n03x5 gen_filter_20__u_filter_filter_q_reg_gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1733 (.o(net1733));
 b15tihi00an1n03x5 gen_filter_20__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_diff_ctr_q_reg_0__1734 (.o(net1734));
 b15tihi00an1n03x5 gen_filter_20__u_filter_stored_value_q_reg_1735 (.o(net1735));
 b15tihi00an1n03x5 gen_filter_21__u_filter_diff_ctr_q_reg_1__gen_filter_21__u_filter_diff_ctr_q_reg_2__1736 (.o(net1736));
 b15tihi00an1n03x5 gen_filter_21__u_filter_diff_ctr_q_reg_3__gen_filter_21__u_filter_filter_q_reg_1737 (.o(net1737));
 b15tihi00an1n03x5 gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_21__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1738 (.o(net1738));
 b15tihi00an1n03x5 gen_filter_21__u_filter_stored_value_q_reg_1739 (.o(net1739));
 b15tihi00an1n03x5 gen_filter_22__u_filter_diff_ctr_q_reg_0__gen_filter_22__u_filter_diff_ctr_q_reg_1__1740 (.o(net1740));
 b15tihi00an1n03x5 gen_filter_22__u_filter_diff_ctr_q_reg_2__gen_filter_22__u_filter_diff_ctr_q_reg_3__1741 (.o(net1741));
 b15tihi00an1n03x5 gen_filter_22__u_filter_filter_q_reg_gen_filter_24__u_filter_diff_ctr_q_reg_0__1742 (.o(net1742));
 b15tihi00an1n03x5 gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_22__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1743 (.o(net1743));
 b15tihi00an1n03x5 gen_filter_22__u_filter_stored_value_q_reg_1744 (.o(net1744));
 b15tihi00an1n03x5 gen_filter_23__u_filter_diff_ctr_q_reg_1__gen_filter_23__u_filter_diff_ctr_q_reg_2__1745 (.o(net1745));
 b15tihi00an1n03x5 gen_filter_23__u_filter_diff_ctr_q_reg_3__gen_filter_23__u_filter_filter_q_reg_1746 (.o(net1746));
 b15tihi00an1n03x5 gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_23__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1747 (.o(net1747));
 b15tihi00an1n03x5 gen_filter_23__u_filter_stored_value_q_reg_1748 (.o(net1748));
 b15tihi00an1n03x5 gen_filter_24__u_filter_diff_ctr_q_reg_1__gen_filter_24__u_filter_diff_ctr_q_reg_3__1749 (.o(net1749));
 b15tihi00an1n03x5 gen_filter_24__u_filter_diff_ctr_q_reg_2__gen_filter_24__u_filter_filter_q_reg_1750 (.o(net1750));
 b15tihi00an1n03x5 gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_24__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1751 (.o(net1751));
 b15tihi00an1n03x5 gen_filter_24__u_filter_stored_value_q_reg_1752 (.o(net1752));
 b15tihi00an1n03x5 gen_filter_25__u_filter_diff_ctr_q_reg_0__gen_filter_25__u_filter_diff_ctr_q_reg_1__1753 (.o(net1753));
 b15tihi00an1n03x5 gen_filter_25__u_filter_diff_ctr_q_reg_2__gen_filter_25__u_filter_diff_ctr_q_reg_3__1754 (.o(net1754));
 b15tihi00an1n03x5 gen_filter_25__u_filter_filter_q_reg_1755 (.o(net1755));
 b15tihi00an1n03x5 gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_25__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1756 (.o(net1756));
 b15tihi00an1n03x5 gen_filter_25__u_filter_stored_value_q_reg_1757 (.o(net1757));
 b15tihi00an1n03x5 gen_filter_26__u_filter_diff_ctr_q_reg_0__gen_filter_26__u_filter_diff_ctr_q_reg_1__1758 (.o(net1758));
 b15tihi00an1n03x5 gen_filter_26__u_filter_diff_ctr_q_reg_2__gen_filter_26__u_filter_diff_ctr_q_reg_3__1759 (.o(net1759));
 b15tihi00an1n03x5 gen_filter_26__u_filter_filter_q_reg_gen_filter_31__u_filter_diff_ctr_q_reg_0__1760 (.o(net1760));
 b15tihi00an1n03x5 gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_diff_ctr_q_reg_0__1761 (.o(net1761));
 b15tihi00an1n03x5 gen_filter_26__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_31__u_filter_diff_ctr_q_reg_1__1762 (.o(net1762));
 b15tihi00an1n03x5 gen_filter_26__u_filter_stored_value_q_reg_1763 (.o(net1763));
 b15tihi00an1n03x5 gen_filter_27__u_filter_diff_ctr_q_reg_0__gen_filter_27__u_filter_diff_ctr_q_reg_1__1764 (.o(net1764));
 b15tihi00an1n03x5 gen_filter_27__u_filter_diff_ctr_q_reg_2__gen_filter_27__u_filter_diff_ctr_q_reg_3__1765 (.o(net1765));
 b15tihi00an1n03x5 gen_filter_27__u_filter_filter_q_reg_gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1766 (.o(net1766));
 b15tihi00an1n03x5 gen_filter_27__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_30__u_filter_diff_ctr_q_reg_1__1767 (.o(net1767));
 b15tihi00an1n03x5 gen_filter_27__u_filter_stored_value_q_reg_1768 (.o(net1768));
 b15tihi00an1n03x5 gen_filter_28__u_filter_diff_ctr_q_reg_1__gen_filter_28__u_filter_diff_ctr_q_reg_2__1769 (.o(net1769));
 b15tihi00an1n03x5 gen_filter_28__u_filter_diff_ctr_q_reg_3__gen_filter_28__u_filter_filter_q_reg_1770 (.o(net1770));
 b15tihi00an1n03x5 gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_28__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1771 (.o(net1771));
 b15tihi00an1n03x5 gen_filter_28__u_filter_stored_value_q_reg_1772 (.o(net1772));
 b15tihi00an1n03x5 gen_filter_29__u_filter_diff_ctr_q_reg_0__gen_filter_29__u_filter_diff_ctr_q_reg_1__1773 (.o(net1773));
 b15tihi00an1n03x5 gen_filter_29__u_filter_diff_ctr_q_reg_2__gen_filter_29__u_filter_diff_ctr_q_reg_3__1774 (.o(net1774));
 b15tihi00an1n03x5 gen_filter_29__u_filter_filter_q_reg_1775 (.o(net1775));
 b15tihi00an1n03x5 gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_29__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1776 (.o(net1776));
 b15tihi00an1n03x5 gen_filter_29__u_filter_stored_value_q_reg_1777 (.o(net1777));
 b15tihi00an1n03x5 gen_filter_2__u_filter_diff_ctr_q_reg_0__gen_filter_2__u_filter_diff_ctr_q_reg_1__1778 (.o(net1778));
 b15tihi00an1n03x5 gen_filter_2__u_filter_diff_ctr_q_reg_2__gen_filter_2__u_filter_diff_ctr_q_reg_3__1779 (.o(net1779));
 b15tihi00an1n03x5 gen_filter_2__u_filter_filter_q_reg_gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1780 (.o(net1780));
 b15tihi00an1n03x5 gen_filter_2__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_3__u_filter_diff_ctr_q_reg_0__1781 (.o(net1781));
 b15tihi00an1n03x5 gen_filter_2__u_filter_stored_value_q_reg_1782 (.o(net1782));
 b15tihi00an1n03x5 gen_filter_30__u_filter_diff_ctr_q_reg_2__gen_filter_30__u_filter_diff_ctr_q_reg_3__1783 (.o(net1783));
 b15tihi00an1n03x5 gen_filter_30__u_filter_filter_q_reg_gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1784 (.o(net1784));
 b15tihi00an1n03x5 gen_filter_30__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1785 (.o(net1785));
 b15tihi00an1n03x5 gen_filter_30__u_filter_stored_value_q_reg_1786 (.o(net1786));
 b15tihi00an1n03x5 gen_filter_31__u_filter_diff_ctr_q_reg_2__gen_filter_31__u_filter_diff_ctr_q_reg_3__1787 (.o(net1787));
 b15tihi00an1n03x5 gen_filter_31__u_filter_filter_q_reg_gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1788 (.o(net1788));
 b15tihi00an1n03x5 gen_filter_31__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__u_reg_err_q_reg_1789 (.o(net1789));
 b15tihi00an1n03x5 gen_filter_31__u_filter_stored_value_q_reg_1790 (.o(net1790));
 b15tihi00an1n03x5 gen_filter_3__u_filter_diff_ctr_q_reg_1__gen_filter_3__u_filter_diff_ctr_q_reg_2__1791 (.o(net1791));
 b15tihi00an1n03x5 gen_filter_3__u_filter_diff_ctr_q_reg_3__gen_filter_3__u_filter_filter_q_reg_1792 (.o(net1792));
 b15tihi00an1n03x5 gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_4__u_filter_diff_ctr_q_reg_1__1793 (.o(net1793));
 b15tihi00an1n03x5 gen_filter_3__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_8__u_filter_diff_ctr_q_reg_0__1794 (.o(net1794));
 b15tihi00an1n03x5 gen_filter_3__u_filter_stored_value_q_reg_1795 (.o(net1795));
 b15tihi00an1n03x5 gen_filter_4__u_filter_diff_ctr_q_reg_0__gen_filter_4__u_filter_diff_ctr_q_reg_2__1796 (.o(net1796));
 b15tihi00an1n03x5 gen_filter_4__u_filter_diff_ctr_q_reg_3__gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1797 (.o(net1797));
 b15tihi00an1n03x5 gen_filter_4__u_filter_filter_q_reg_gen_filter_7__u_filter_filter_q_reg_1798 (.o(net1798));
 b15tihi00an1n03x5 gen_filter_4__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_7__u_filter_diff_ctr_q_reg_0__1799 (.o(net1799));
 b15tihi00an1n03x5 gen_filter_4__u_filter_stored_value_q_reg_1800 (.o(net1800));
 b15tihi00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_0__gen_filter_5__u_filter_diff_ctr_q_reg_1__1801 (.o(net1801));
 b15tihi00an1n03x5 gen_filter_5__u_filter_diff_ctr_q_reg_2__gen_filter_5__u_filter_diff_ctr_q_reg_3__1802 (.o(net1802));
 b15tihi00an1n03x5 gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_diff_ctr_q_reg_0__1803 (.o(net1803));
 b15tihi00an1n03x5 gen_filter_5__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_filter_q_reg_1804 (.o(net1804));
 b15tihi00an1n03x5 gen_filter_5__u_filter_stored_value_q_reg_1805 (.o(net1805));
 b15tihi00an1n03x5 gen_filter_6__u_filter_diff_ctr_q_reg_1__gen_filter_6__u_filter_diff_ctr_q_reg_2__1806 (.o(net1806));
 b15tihi00an1n03x5 gen_filter_6__u_filter_diff_ctr_q_reg_3__gen_filter_15__u_filter_diff_ctr_q_reg_0__1807 (.o(net1807));
 b15tihi00an1n03x5 gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_6__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1808 (.o(net1808));
 b15tihi00an1n03x5 gen_filter_6__u_filter_stored_value_q_reg_1809 (.o(net1809));
 b15tihi00an1n03x5 gen_filter_7__u_filter_diff_ctr_q_reg_1__gen_filter_7__u_filter_diff_ctr_q_reg_2__1810 (.o(net1810));
 b15tihi00an1n03x5 gen_filter_7__u_filter_diff_ctr_q_reg_3__gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1811 (.o(net1811));
 b15tihi00an1n03x5 gen_filter_7__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_9__u_filter_diff_ctr_q_reg_0__1812 (.o(net1812));
 b15tihi00an1n03x5 gen_filter_7__u_filter_stored_value_q_reg_1813 (.o(net1813));
 b15tihi00an1n03x5 gen_filter_8__u_filter_diff_ctr_q_reg_1__gen_filter_8__u_filter_diff_ctr_q_reg_2__1814 (.o(net1814));
 b15tihi00an1n03x5 gen_filter_8__u_filter_diff_ctr_q_reg_3__gen_filter_10__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1815 (.o(net1815));
 b15tihi00an1n03x5 gen_filter_8__u_filter_filter_q_reg_gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__1816 (.o(net1816));
 b15tihi00an1n03x5 gen_filter_8__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_11__u_filter_diff_ctr_q_reg_2__1817 (.o(net1817));
 b15tihi00an1n03x5 gen_filter_8__u_filter_stored_value_q_reg_1818 (.o(net1818));
 b15tihi00an1n03x5 gen_filter_9__u_filter_diff_ctr_q_reg_1__gen_filter_9__u_filter_diff_ctr_q_reg_2__1819 (.o(net1819));
 b15tihi00an1n03x5 gen_filter_9__u_filter_diff_ctr_q_reg_3__gen_filter_9__u_filter_filter_q_reg_1820 (.o(net1820));
 b15tihi00an1n03x5 gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_1_gen_generic_u_impl_generic_q_o_reg_0__gen_filter_9__u_filter_gen_async_prim_flop_2sync_u_sync_2_gen_generic_u_impl_generic_q_o_reg_0__1821 (.o(net1821));
 b15tihi00an1n03x5 gen_filter_9__u_filter_stored_value_q_reg_1822 (.o(net1822));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_10__intr_hw_intr_o_reg_11__1823 (.o(net1823));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_12__intr_hw_intr_o_reg_14__1824 (.o(net1824));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_15__intr_hw_intr_o_reg_25__1825 (.o(net1825));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_16__intr_hw_intr_o_reg_17__1826 (.o(net1826));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_18__intr_hw_intr_o_reg_19__1827 (.o(net1827));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_1__intr_hw_intr_o_reg_2__1828 (.o(net1828));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_20__intr_hw_intr_o_reg_21__1829 (.o(net1829));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_22__intr_hw_intr_o_reg_23__1830 (.o(net1830));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_24__intr_hw_intr_o_reg_26__1831 (.o(net1831));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_27__intr_hw_intr_o_reg_28__1832 (.o(net1832));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_29__intr_hw_intr_o_reg_30__1833 (.o(net1833));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_31__u_reg_u_data_in_q_reg_1__1834 (.o(net1834));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_3__intr_hw_intr_o_reg_4__1835 (.o(net1835));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_5__intr_hw_intr_o_reg_6__1836 (.o(net1836));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_7__intr_hw_intr_o_reg_8__1837 (.o(net1837));
 b15tihi00an1n03x5 intr_hw_intr_o_reg_9__intr_hw_intr_o_reg_13__1838 (.o(net1838));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_0__u_reg_u_ctrl_en_input_filter_q_reg_1__1839 (.o(net1839));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_10__u_reg_u_ctrl_en_input_filter_q_reg_11__1840 (.o(net1840));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_12__u_reg_u_ctrl_en_input_filter_q_reg_13__1841 (.o(net1841));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_14__u_reg_u_ctrl_en_input_filter_q_reg_15__1842 (.o(net1842));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_16__u_reg_u_ctrl_en_input_filter_q_reg_17__1843 (.o(net1843));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_18__u_reg_u_ctrl_en_input_filter_q_reg_19__1844 (.o(net1844));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_20__u_reg_u_ctrl_en_input_filter_q_reg_21__1845 (.o(net1845));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_22__u_reg_u_ctrl_en_input_filter_q_reg_23__1846 (.o(net1846));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_24__u_reg_u_ctrl_en_input_filter_q_reg_25__1847 (.o(net1847));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_26__u_reg_u_ctrl_en_input_filter_q_reg_27__1848 (.o(net1848));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_28__u_reg_u_ctrl_en_input_filter_q_reg_29__1849 (.o(net1849));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_2__u_reg_u_ctrl_en_input_filter_q_reg_3__1850 (.o(net1850));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_30__u_reg_u_ctrl_en_input_filter_q_reg_31__1851 (.o(net1851));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_4__u_reg_u_ctrl_en_input_filter_q_reg_5__1852 (.o(net1852));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_6__u_reg_u_ctrl_en_input_filter_q_reg_7__1853 (.o(net1853));
 b15tihi00an1n03x5 u_reg_u_ctrl_en_input_filter_q_reg_8__u_reg_u_ctrl_en_input_filter_q_reg_9__1854 (.o(net1854));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_0__u_reg_u_data_in_q_reg_3__1855 (.o(net1855));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_10__u_reg_u_data_in_q_reg_14__1856 (.o(net1856));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_11__u_reg_u_data_in_q_reg_12__1857 (.o(net1857));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_13__u_reg_u_reg_if_rspop_reg_1__1858 (.o(net1858));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_15__u_reg_u_data_in_q_reg_20__1859 (.o(net1859));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_16__u_reg_u_data_in_q_reg_17__1860 (.o(net1860));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_18__u_reg_u_data_in_q_reg_19__1861 (.o(net1861));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_21__u_reg_u_data_in_q_reg_22__1862 (.o(net1862));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_23__1863 (.o(net1863));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_24__u_reg_u_data_in_q_reg_25__1864 (.o(net1864));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_26__1865 (.o(net1865));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_27__u_reg_u_data_in_q_reg_28__1866 (.o(net1866));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_29__u_reg_u_data_in_q_reg_30__1867 (.o(net1867));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_2__1868 (.o(net1868));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_31__1869 (.o(net1869));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_4__u_reg_u_data_in_q_reg_5__1870 (.o(net1870));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_6__u_reg_u_data_in_q_reg_7__1871 (.o(net1871));
 b15tihi00an1n03x5 u_reg_u_data_in_q_reg_8__u_reg_u_data_in_q_reg_9__1872 (.o(net1872));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_0__u_reg_u_intr_ctrl_en_falling_q_reg_1__1873 (.o(net1873));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_10__u_reg_u_intr_ctrl_en_falling_q_reg_11__1874 (.o(net1874));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_12__u_reg_u_intr_ctrl_en_falling_q_reg_13__1875 (.o(net1875));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_14__u_reg_u_intr_ctrl_en_falling_q_reg_15__1876 (.o(net1876));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_16__u_reg_u_intr_ctrl_en_falling_q_reg_17__1877 (.o(net1877));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_18__u_reg_u_intr_ctrl_en_falling_q_reg_19__1878 (.o(net1878));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_20__u_reg_u_intr_ctrl_en_falling_q_reg_21__1879 (.o(net1879));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_22__u_reg_u_intr_ctrl_en_falling_q_reg_23__1880 (.o(net1880));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_24__u_reg_u_intr_ctrl_en_falling_q_reg_25__1881 (.o(net1881));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_26__u_reg_u_intr_ctrl_en_falling_q_reg_27__1882 (.o(net1882));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_28__u_reg_u_intr_ctrl_en_falling_q_reg_29__1883 (.o(net1883));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_2__u_reg_u_intr_ctrl_en_falling_q_reg_3__1884 (.o(net1884));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_30__u_reg_u_intr_ctrl_en_falling_q_reg_31__1885 (.o(net1885));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_4__u_reg_u_intr_ctrl_en_falling_q_reg_5__1886 (.o(net1886));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_6__u_reg_u_intr_ctrl_en_falling_q_reg_7__1887 (.o(net1887));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_falling_q_reg_8__u_reg_u_intr_ctrl_en_falling_q_reg_9__1888 (.o(net1888));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_0__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_1__1889 (.o(net1889));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_10__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_11__1890 (.o(net1890));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_12__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_13__1891 (.o(net1891));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_14__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_15__1892 (.o(net1892));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_16__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_17__1893 (.o(net1893));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_18__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_19__1894 (.o(net1894));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_20__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_21__1895 (.o(net1895));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_22__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_23__1896 (.o(net1896));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_24__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_25__1897 (.o(net1897));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_26__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_27__1898 (.o(net1898));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_28__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_29__1899 (.o(net1899));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_2__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_3__1900 (.o(net1900));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_30__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_31__1901 (.o(net1901));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_4__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_5__1902 (.o(net1902));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_6__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_7__1903 (.o(net1903));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvlhigh_q_reg_8__u_reg_u_intr_ctrl_en_lvlhigh_q_reg_9__1904 (.o(net1904));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_0__u_reg_u_intr_ctrl_en_lvllow_q_reg_1__1905 (.o(net1905));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_10__u_reg_u_intr_ctrl_en_lvllow_q_reg_11__1906 (.o(net1906));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_12__u_reg_u_intr_ctrl_en_lvllow_q_reg_13__1907 (.o(net1907));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_14__u_reg_u_intr_ctrl_en_lvllow_q_reg_15__1908 (.o(net1908));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_16__u_reg_u_intr_ctrl_en_lvllow_q_reg_17__1909 (.o(net1909));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_18__u_reg_u_intr_ctrl_en_lvllow_q_reg_19__1910 (.o(net1910));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_20__u_reg_u_intr_ctrl_en_lvllow_q_reg_21__1911 (.o(net1911));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_22__u_reg_u_intr_ctrl_en_lvllow_q_reg_23__1912 (.o(net1912));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_24__u_reg_u_intr_ctrl_en_lvllow_q_reg_25__1913 (.o(net1913));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_26__u_reg_u_intr_ctrl_en_lvllow_q_reg_27__1914 (.o(net1914));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_28__u_reg_u_intr_ctrl_en_lvllow_q_reg_29__1915 (.o(net1915));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_2__u_reg_u_intr_ctrl_en_lvllow_q_reg_3__1916 (.o(net1916));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_30__u_reg_u_intr_ctrl_en_lvllow_q_reg_31__1917 (.o(net1917));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_4__u_reg_u_intr_ctrl_en_lvllow_q_reg_5__1918 (.o(net1918));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_6__u_reg_u_intr_ctrl_en_lvllow_q_reg_7__1919 (.o(net1919));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_lvllow_q_reg_8__u_reg_u_intr_ctrl_en_lvllow_q_reg_9__1920 (.o(net1920));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_0__u_reg_u_intr_ctrl_en_rising_q_reg_1__1921 (.o(net1921));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_10__u_reg_u_intr_ctrl_en_rising_q_reg_11__1922 (.o(net1922));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_12__u_reg_u_intr_ctrl_en_rising_q_reg_13__1923 (.o(net1923));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_14__u_reg_u_intr_ctrl_en_rising_q_reg_15__1924 (.o(net1924));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_16__u_reg_u_intr_ctrl_en_rising_q_reg_17__1925 (.o(net1925));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_18__u_reg_u_intr_ctrl_en_rising_q_reg_19__1926 (.o(net1926));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_20__u_reg_u_intr_ctrl_en_rising_q_reg_21__1927 (.o(net1927));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_22__u_reg_u_intr_ctrl_en_rising_q_reg_23__1928 (.o(net1928));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_24__u_reg_u_intr_ctrl_en_rising_q_reg_25__1929 (.o(net1929));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_26__u_reg_u_intr_ctrl_en_rising_q_reg_27__1930 (.o(net1930));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_28__u_reg_u_intr_ctrl_en_rising_q_reg_29__1931 (.o(net1931));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_2__u_reg_u_intr_ctrl_en_rising_q_reg_3__1932 (.o(net1932));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_30__u_reg_u_intr_ctrl_en_rising_q_reg_31__1933 (.o(net1933));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_4__u_reg_u_intr_ctrl_en_rising_q_reg_5__1934 (.o(net1934));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_6__u_reg_u_intr_ctrl_en_rising_q_reg_7__1935 (.o(net1935));
 b15tihi00an1n03x5 u_reg_u_intr_ctrl_en_rising_q_reg_8__u_reg_u_intr_ctrl_en_rising_q_reg_9__1936 (.o(net1936));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_0__u_reg_u_intr_enable_q_reg_1__1937 (.o(net1937));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_10__u_reg_u_intr_enable_q_reg_11__1938 (.o(net1938));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_12__u_reg_u_intr_enable_q_reg_13__1939 (.o(net1939));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_14__u_reg_u_intr_enable_q_reg_15__1940 (.o(net1940));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_16__u_reg_u_intr_enable_q_reg_17__1941 (.o(net1941));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_18__u_reg_u_intr_enable_q_reg_19__1942 (.o(net1942));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_20__u_reg_u_intr_enable_q_reg_21__1943 (.o(net1943));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_22__u_reg_u_intr_enable_q_reg_23__1944 (.o(net1944));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_24__u_reg_u_intr_enable_q_reg_25__1945 (.o(net1945));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_26__u_reg_u_intr_enable_q_reg_27__1946 (.o(net1946));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_28__u_reg_u_intr_enable_q_reg_29__1947 (.o(net1947));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_2__u_reg_u_intr_enable_q_reg_3__1948 (.o(net1948));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_30__u_reg_u_intr_enable_q_reg_31__1949 (.o(net1949));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_4__u_reg_u_intr_enable_q_reg_5__1950 (.o(net1950));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_6__u_reg_u_intr_enable_q_reg_7__1951 (.o(net1951));
 b15tihi00an1n03x5 u_reg_u_intr_enable_q_reg_8__u_reg_u_intr_enable_q_reg_9__1952 (.o(net1952));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_0__u_reg_u_intr_state_q_reg_1__1953 (.o(net1953));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_10__u_reg_u_intr_state_q_reg_11__1954 (.o(net1954));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_12__u_reg_u_intr_state_q_reg_13__1955 (.o(net1955));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_14__u_reg_u_intr_state_q_reg_15__1956 (.o(net1956));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_16__u_reg_u_intr_state_q_reg_17__1957 (.o(net1957));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_18__u_reg_u_intr_state_q_reg_19__1958 (.o(net1958));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_20__u_reg_u_intr_state_q_reg_21__1959 (.o(net1959));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_22__u_reg_u_intr_state_q_reg_23__1960 (.o(net1960));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_24__u_reg_u_intr_state_q_reg_25__1961 (.o(net1961));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_26__u_reg_u_intr_state_q_reg_27__1962 (.o(net1962));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_28__u_reg_u_intr_state_q_reg_29__1963 (.o(net1963));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_2__u_reg_u_intr_state_q_reg_3__1964 (.o(net1964));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_30__u_reg_u_intr_state_q_reg_31__1965 (.o(net1965));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_4__u_reg_u_intr_state_q_reg_5__1966 (.o(net1966));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_6__u_reg_u_intr_state_q_reg_7__1967 (.o(net1967));
 b15tihi00an1n03x5 u_reg_u_intr_state_q_reg_8__u_reg_u_intr_state_q_reg_9__1968 (.o(net1968));
 b15tihi00an1n03x5 u_reg_u_reg_if_error_reg_1969 (.o(net1969));
 b15tihi00an1n03x5 u_reg_u_reg_if_outstanding_reg_1970 (.o(net1970));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_0__u_reg_u_reg_if_rdata_reg_1__1971 (.o(net1971));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_10__u_reg_u_reg_if_rdata_reg_11__1972 (.o(net1972));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_12__u_reg_u_reg_if_rdata_reg_13__1973 (.o(net1973));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_14__u_reg_u_reg_if_rdata_reg_15__1974 (.o(net1974));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_16__u_reg_u_reg_if_rdata_reg_17__1975 (.o(net1975));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_18__u_reg_u_reg_if_rdata_reg_19__1976 (.o(net1976));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_20__u_reg_u_reg_if_rdata_reg_21__1977 (.o(net1977));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_22__u_reg_u_reg_if_rdata_reg_23__1978 (.o(net1978));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_24__u_reg_u_reg_if_rdata_reg_25__1979 (.o(net1979));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_26__u_reg_u_reg_if_rdata_reg_27__1980 (.o(net1980));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_28__u_reg_u_reg_if_rdata_reg_29__1981 (.o(net1981));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_2__u_reg_u_reg_if_rdata_reg_3__1982 (.o(net1982));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_30__u_reg_u_reg_if_rdata_reg_31__1983 (.o(net1983));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_4__u_reg_u_reg_if_rdata_reg_5__1984 (.o(net1984));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_6__u_reg_u_reg_if_rdata_reg_7__1985 (.o(net1985));
 b15tihi00an1n03x5 u_reg_u_reg_if_rdata_reg_8__u_reg_u_reg_if_rdata_reg_9__1986 (.o(net1986));
 b15tihi00an1n03x5 u_reg_u_reg_if_reqid_reg_0__u_reg_u_reg_if_reqid_reg_1__1987 (.o(net1987));
 b15tihi00an1n03x5 u_reg_u_reg_if_reqid_reg_2__u_reg_u_reg_if_reqid_reg_3__1988 (.o(net1988));
 b15tihi00an1n03x5 u_reg_u_reg_if_reqid_reg_4__u_reg_u_reg_if_reqid_reg_5__1989 (.o(net1989));
 b15tihi00an1n03x5 u_reg_u_reg_if_reqid_reg_6__u_reg_u_reg_if_reqid_reg_7__1990 (.o(net1990));
 b15tihi00an1n03x5 u_reg_u_reg_if_reqsz_reg_0__1991 (.o(net1991));
 b15tihi00an1n03x5 u_reg_u_reg_if_reqsz_reg_1__1992 (.o(net1992));
 b15tihi00an1n03x5 u_reg_u_reg_if_rspop_reg_0__1993 (.o(net1993));
 b15tihi00an1n03x5 u_reg_u_reg_if_rspop_reg_2__1994 (.o(net1994));
 b15cbf000an1n16x5 clkbuf_leaf_1_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_1_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_2_clk_i (.clk(net1996),
    .clkout(clknet_leaf_2_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_3_clk_i (.clk(net1998),
    .clkout(clknet_leaf_3_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_4_clk_i (.clk(net1998),
    .clkout(clknet_leaf_4_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_5_clk_i (.clk(net1997),
    .clkout(clknet_leaf_5_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_6_clk_i (.clk(net1997),
    .clkout(clknet_leaf_6_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_7_clk_i (.clk(clknet_1_1__leaf_clk_i),
    .clkout(clknet_leaf_7_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_8_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_8_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_9_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_9_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_10_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_10_clk_i));
 b15cbf000an1n16x5 clkbuf_leaf_11_clk_i (.clk(clknet_1_0__leaf_clk_i),
    .clkout(clknet_leaf_11_clk_i));
 b15cbf000an1n16x5 clkbuf_0_clk_i (.clk(net1995),
    .clkout(clknet_0_clk_i));
 b15cbf000an1n16x5 clkbuf_1_0__f_clk_i (.clk(clknet_0_clk_i),
    .clkout(clknet_1_0__leaf_clk_i));
 b15cbf000an1n16x5 clkbuf_1_1__f_clk_i (.clk(clknet_0_clk_i),
    .clkout(clknet_1_1__leaf_clk_i));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_reg_if_net2113 (.clk(u_reg_u_reg_if_net2113),
    .clkout(clknet_0_u_reg_u_reg_if_net2113));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_reg_if_net2113 (.clk(clknet_0_u_reg_u_reg_if_net2113),
    .clkout(clknet_1_0__leaf_u_reg_u_reg_if_net2113));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_reg_if_net2113 (.clk(clknet_0_u_reg_u_reg_if_net2113),
    .clkout(clknet_1_1__leaf_u_reg_u_reg_if_net2113));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_reg_if_net2119 (.clk(u_reg_u_reg_if_net2119),
    .clkout(clknet_0_u_reg_u_reg_if_net2119));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_reg_if_net2119 (.clk(clknet_0_u_reg_u_reg_if_net2119),
    .clkout(clknet_1_0__leaf_u_reg_u_reg_if_net2119));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_reg_if_net2119 (.clk(clknet_0_u_reg_u_reg_if_net2119),
    .clkout(clknet_1_1__leaf_u_reg_u_reg_if_net2119));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_reg_if_net2124 (.clk(u_reg_u_reg_if_net2124),
    .clkout(clknet_0_u_reg_u_reg_if_net2124));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_reg_if_net2124 (.clk(clknet_0_u_reg_u_reg_if_net2124),
    .clkout(clknet_1_0__leaf_u_reg_u_reg_if_net2124));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_reg_if_net2124 (.clk(clknet_0_u_reg_u_reg_if_net2124),
    .clkout(clknet_1_1__leaf_u_reg_u_reg_if_net2124));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_state_net2090 (.clk(u_reg_u_intr_state_net2090),
    .clkout(clknet_0_u_reg_u_intr_state_net2090));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_state_net2090 (.clk(clknet_0_u_reg_u_intr_state_net2090),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_state_net2090));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_state_net2090 (.clk(clknet_0_u_reg_u_intr_state_net2090),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_state_net2090));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_state_net2096 (.clk(u_reg_u_intr_state_net2096),
    .clkout(clknet_0_u_reg_u_intr_state_net2096));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_state_net2096 (.clk(clknet_0_u_reg_u_intr_state_net2096),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_state_net2096));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_state_net2096 (.clk(clknet_0_u_reg_u_intr_state_net2096),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_state_net2096));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_enable_net2067 (.clk(u_reg_u_intr_enable_net2067),
    .clkout(clknet_0_u_reg_u_intr_enable_net2067));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_enable_net2067 (.clk(clknet_0_u_reg_u_intr_enable_net2067),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_enable_net2067));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_enable_net2067 (.clk(clknet_0_u_reg_u_intr_enable_net2067),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_enable_net2067));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_enable_net2073 (.clk(u_reg_u_intr_enable_net2073),
    .clkout(clknet_0_u_reg_u_intr_enable_net2073));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_enable_net2073 (.clk(clknet_0_u_reg_u_intr_enable_net2073),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_enable_net2073));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_enable_net2073 (.clk(clknet_0_u_reg_u_intr_enable_net2073),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_enable_net2073));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_rising_net2067 (.clk(u_reg_u_intr_ctrl_en_rising_net2067),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_rising_net2067));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_rising_net2067 (.clk(clknet_0_u_reg_u_intr_ctrl_en_rising_net2067),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2067));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_rising_net2067 (.clk(clknet_0_u_reg_u_intr_ctrl_en_rising_net2067),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2067));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_rising_net2073 (.clk(u_reg_u_intr_ctrl_en_rising_net2073),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_rising_net2073));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_rising_net2073 (.clk(clknet_0_u_reg_u_intr_ctrl_en_rising_net2073),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_rising_net2073));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_rising_net2073 (.clk(clknet_0_u_reg_u_intr_ctrl_en_rising_net2073),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_rising_net2073));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_lvllow_net2067 (.clk(u_reg_u_intr_ctrl_en_lvllow_net2067),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2067));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_lvllow_net2067 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2067),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2067));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_lvllow_net2067 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2067),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2067));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_lvllow_net2073 (.clk(u_reg_u_intr_ctrl_en_lvllow_net2073),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2073));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_lvllow_net2073 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2073),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvllow_net2073));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_lvllow_net2073 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvllow_net2073),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvllow_net2073));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_lvlhigh_net2067 (.clk(u_reg_u_intr_ctrl_en_lvlhigh_net2067),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2067));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_lvlhigh_net2067 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2067),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2067));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_lvlhigh_net2067 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2067),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2067));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_lvlhigh_net2073 (.clk(u_reg_u_intr_ctrl_en_lvlhigh_net2073),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2073));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_lvlhigh_net2073 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2073),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2073));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_lvlhigh_net2073 (.clk(clknet_0_u_reg_u_intr_ctrl_en_lvlhigh_net2073),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_lvlhigh_net2073));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_falling_net2067 (.clk(u_reg_u_intr_ctrl_en_falling_net2067),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_falling_net2067));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_falling_net2067 (.clk(clknet_0_u_reg_u_intr_ctrl_en_falling_net2067),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2067));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_falling_net2067 (.clk(clknet_0_u_reg_u_intr_ctrl_en_falling_net2067),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2067));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_intr_ctrl_en_falling_net2073 (.clk(u_reg_u_intr_ctrl_en_falling_net2073),
    .clkout(clknet_0_u_reg_u_intr_ctrl_en_falling_net2073));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_intr_ctrl_en_falling_net2073 (.clk(clknet_0_u_reg_u_intr_ctrl_en_falling_net2073),
    .clkout(clknet_1_0__leaf_u_reg_u_intr_ctrl_en_falling_net2073));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_intr_ctrl_en_falling_net2073 (.clk(clknet_0_u_reg_u_intr_ctrl_en_falling_net2073),
    .clkout(clknet_1_1__leaf_u_reg_u_intr_ctrl_en_falling_net2073));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_ctrl_en_input_filter_net2067 (.clk(u_reg_u_ctrl_en_input_filter_net2067),
    .clkout(clknet_0_u_reg_u_ctrl_en_input_filter_net2067));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_ctrl_en_input_filter_net2067 (.clk(clknet_0_u_reg_u_ctrl_en_input_filter_net2067),
    .clkout(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2067));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_ctrl_en_input_filter_net2067 (.clk(clknet_0_u_reg_u_ctrl_en_input_filter_net2067),
    .clkout(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2067));
 b15cbf000an1n16x5 clkbuf_0_u_reg_u_ctrl_en_input_filter_net2073 (.clk(u_reg_u_ctrl_en_input_filter_net2073),
    .clkout(clknet_0_u_reg_u_ctrl_en_input_filter_net2073));
 b15cbf000an1n16x5 clkbuf_1_0__f_u_reg_u_ctrl_en_input_filter_net2073 (.clk(clknet_0_u_reg_u_ctrl_en_input_filter_net2073),
    .clkout(clknet_1_0__leaf_u_reg_u_ctrl_en_input_filter_net2073));
 b15cbf000an1n16x5 clkbuf_1_1__f_u_reg_u_ctrl_en_input_filter_net2073 (.clk(clknet_0_u_reg_u_ctrl_en_input_filter_net2073),
    .clkout(clknet_1_1__leaf_u_reg_u_ctrl_en_input_filter_net2073));
 b15cbf000an1n16x5 clkbuf_0_net2034 (.clk(net2034),
    .clkout(clknet_0_net2034));
 b15cbf000an1n16x5 clkbuf_1_0__f_net2034 (.clk(clknet_0_net2034),
    .clkout(clknet_1_0__leaf_net2034));
 b15cbf000an1n16x5 clkbuf_1_1__f_net2034 (.clk(clknet_0_net2034),
    .clkout(clknet_1_1__leaf_net2034));
 b15cbf000an1n16x5 clkbuf_0_net2040 (.clk(net2040),
    .clkout(clknet_0_net2040));
 b15cbf000an1n16x5 clkbuf_1_0__f_net2040 (.clk(clknet_0_net2040),
    .clkout(clknet_1_0__leaf_net2040));
 b15cbf000an1n16x5 clkbuf_1_1__f_net2040 (.clk(clknet_0_net2040),
    .clkout(clknet_1_1__leaf_net2040));
 b15cbf000an1n16x5 clkbuf_0_net2045 (.clk(net2045),
    .clkout(clknet_0_net2045));
 b15cbf000an1n16x5 clkbuf_1_0__f_net2045 (.clk(clknet_0_net2045),
    .clkout(clknet_1_0__leaf_net2045));
 b15cbf000an1n16x5 clkbuf_1_1__f_net2045 (.clk(clknet_0_net2045),
    .clkout(clknet_1_1__leaf_net2045));
 b15cbf000an1n16x5 clkbuf_0_net2050 (.clk(net2050),
    .clkout(clknet_0_net2050));
 b15cbf000an1n16x5 clkbuf_1_0__f_net2050 (.clk(clknet_0_net2050),
    .clkout(clknet_1_0__leaf_net2050));
 b15cbf000an1n16x5 clkbuf_1_1__f_net2050 (.clk(clknet_0_net2050),
    .clkout(clknet_1_1__leaf_net2050));
 b15bfn001ah1n32x5 wire1 (.a(clk_i),
    .o(net1995));
 b15bfn001ah1n24x5 max_length2 (.a(net1998),
    .o(net1996));
 b15bfn001ah1n24x5 wire3 (.a(net1998),
    .o(net1997));
 b15bfn001as1n24x5 max_length4 (.a(clknet_1_1__leaf_clk_i),
    .o(net1998));
 b15cbf034ar1n64x5 hold5 (.clk(net2011),
    .clkout(net1999));
 b15cbf034ar1n64x5 hold6 (.clk(net2000),
    .clkout(tl_o[1]));
 b15cbf034ar1n64x5 hold7 (.clk(net2025),
    .clkout(net2001));
 b15cbf034ar1n64x5 hold8 (.clk(net2002),
    .clkout(tl_o[58]));
 b15cbf034ar1n64x5 hold9 (.clk(net2570),
    .clkout(net2003));
 b15cbf034ar1n64x5 hold10 (.clk(net2004),
    .clkout(intr_gpio_o[0]));
 b15cbf034ar1n64x5 hold11 (.clk(net2572),
    .clkout(net2005));
 b15cbf034ar1n64x5 hold12 (.clk(net2006),
    .clkout(intr_gpio_o[25]));
 b15cbf034ar1n64x5 hold13 (.clk(net2039),
    .clkout(net2007));
 b15cbf034ar1n64x5 hold14 (.clk(net2008),
    .clkout(tl_o[64]));
 b15cbf034ar1n64x5 hold15 (.clk(net2574),
    .clkout(net2009));
 b15cbf034ar1n64x5 hold16 (.clk(net2010),
    .clkout(intr_gpio_o[15]));
 b15cbf034ar1n64x5 hold17 (.clk(net248),
    .clkout(net2011));
 b15cbf034ar1n64x5 hold18 (.clk(net1999),
    .clkout(net2012));
 b15cbf034ar1n64x5 hold19 (.clk(net239),
    .clkout(net2013));
 b15cbf034ar1n64x5 hold20 (.clk(net2014),
    .clkout(tl_o[11]));
 b15cbf034ar1n64x5 hold21 (.clk(net2576),
    .clkout(net2015));
 b15cbf034ar1n64x5 hold22 (.clk(net2016),
    .clkout(intr_gpio_o[11]));
 b15cbf034ar1n64x5 hold23 (.clk(net2580),
    .clkout(net2017));
 b15cbf034ar1n64x5 hold24 (.clk(net2018),
    .clkout(intr_gpio_o[1]));
 b15cbf034ar1n64x5 hold25 (.clk(net2081),
    .clkout(net2019));
 b15cbf034ar1n64x5 hold26 (.clk(net2020),
    .clkout(tl_o[65]));
 b15cbf034ar1n64x5 hold27 (.clk(net2578),
    .clkout(net2021));
 b15cbf034ar1n64x5 hold28 (.clk(net2022),
    .clkout(intr_gpio_o[10]));
 b15cbf034ar1n64x5 hold29 (.clk(net2586),
    .clkout(net2023));
 b15cbf034ar1n64x5 hold30 (.clk(net2024),
    .clkout(intr_gpio_o[2]));
 b15cbf034ar1n64x5 hold31 (.clk(net289),
    .clkout(net2025));
 b15cbf034ar1n64x5 hold32 (.clk(net2001),
    .clkout(net2026));
 b15cbf034ar1n64x5 hold33 (.clk(net241),
    .clkout(net2027));
 b15cbf034ar1n64x5 hold34 (.clk(net2584),
    .clkout(net2028));
 b15cbf034ar1n64x5 hold35 (.clk(net2029),
    .clkout(alert_tx_o[0]));
 b15cbf034ar1n64x5 hold36 (.clk(net2075),
    .clkout(net2030));
 b15cbf034ar1n64x5 hold37 (.clk(net2031),
    .clkout(tl_o[57]));
 b15cbf034ar1n64x5 hold38 (.clk(net2592),
    .clkout(net2032));
 b15cbf034ar1n64x5 hold39 (.clk(net2033),
    .clkout(intr_gpio_o[21]));
 b15cbf034ar1n64x5 hold40 (.clk(net2593),
    .clkout(net2035));
 b15cbf034ar1n64x5 hold41 (.clk(net2036),
    .clkout(intr_gpio_o[20]));
 b15cbf034ar1n64x5 hold42 (.clk(net2582),
    .clkout(net2037));
 b15cbf034ar1n64x5 hold43 (.clk(net2038),
    .clkout(alert_tx_o[1]));
 b15cbf034ar1n64x5 hold44 (.clk(net293),
    .clkout(net2039));
 b15cbf034ar1n64x5 hold45 (.clk(net2007),
    .clkout(net2041));
 b15cbf034ar1n64x5 hold46 (.clk(net240),
    .clkout(net2042));
 b15cbf034ar1n64x5 hold47 (.clk(net2043),
    .clkout(tl_o[12]));
 b15cbf034ar1n64x5 hold48 (.clk(net2588),
    .clkout(net2044));
 b15cbf034ar1n64x5 hold49 (.clk(net2046),
    .clkout(intr_gpio_o[28]));
 b15cbf034ar1n64x5 hold50 (.clk(net2590),
    .clkout(net2047));
 b15cbf034ar1n64x5 hold51 (.clk(net2048),
    .clkout(intr_gpio_o[27]));
 b15cbf034ar1n64x5 hold52 (.clk(net2598),
    .clkout(net2049));
 b15cbf034ar1n64x5 hold53 (.clk(net2051),
    .clkout(intr_gpio_o[23]));
 b15cbf034ar1n64x5 hold54 (.clk(net2599),
    .clkout(net2052));
 b15cbf034ar1n64x5 hold55 (.clk(net2053),
    .clkout(intr_gpio_o[22]));
 b15cbf034ar1n64x5 hold56 (.clk(net2080),
    .clkout(net2054));
 b15cbf034ar1n64x5 hold57 (.clk(net737),
    .clkout(net2055));
 b15cbf034ar1n64x5 hold58 (.clk(n2939),
    .clkout(net2056));
 b15cbf034ar1n64x5 hold59 (.clk(n2941),
    .clkout(net2057));
 b15cbf034ar1n64x5 hold60 (.clk(net298),
    .clkout(net2058));
 b15cbf034ar1n64x5 hold61 (.clk(net2606),
    .clkout(net2059));
 b15cbf034ar1n64x5 hold62 (.clk(net2060),
    .clkout(intr_gpio_o[8]));
 b15cbf034ar1n64x5 hold63 (.clk(net2594),
    .clkout(net2061));
 b15cbf034ar1n64x5 hold64 (.clk(net2062),
    .clkout(intr_gpio_o[4]));
 b15cbf034ar1n64x5 hold65 (.clk(net2600),
    .clkout(net2063));
 b15cbf034ar1n64x5 hold66 (.clk(net2064),
    .clkout(intr_gpio_o[18]));
 b15cbf034ar1n64x5 hold67 (.clk(net2596),
    .clkout(net2065));
 b15cbf034ar1n64x5 hold68 (.clk(net2066),
    .clkout(intr_gpio_o[3]));
 b15cbf034ar1n64x5 hold69 (.clk(net2608),
    .clkout(net2067));
 b15cbf034ar1n64x5 hold70 (.clk(net2068),
    .clkout(intr_gpio_o[13]));
 b15cbf034ar1n64x5 hold71 (.clk(net2601),
    .clkout(net2069));
 b15cbf034ar1n64x5 hold72 (.clk(net2070),
    .clkout(intr_gpio_o[6]));
 b15cbf034ar1n64x5 hold73 (.clk(net2602),
    .clkout(net2071));
 b15cbf034ar1n64x5 hold74 (.clk(net2072),
    .clkout(intr_gpio_o[5]));
 b15cbf034ar1n64x5 hold75 (.clk(net2604),
    .clkout(net2073));
 b15cbf034ar1n64x5 hold76 (.clk(net2074),
    .clkout(intr_gpio_o[7]));
 b15cbf034ar1n64x5 hold77 (.clk(net288),
    .clkout(net2075));
 b15cbf034ar1n64x5 hold78 (.clk(net2030),
    .clkout(net2076));
 b15cbf034ar1n64x5 hold79 (.clk(net238),
    .clkout(net2077));
 b15cbf034ar1n64x5 hold80 (.clk(net2609),
    .clkout(net2078));
 b15cbf034ar1n64x5 hold81 (.clk(net2079),
    .clkout(intr_gpio_o[9]));
 b15cbf034ar1n64x5 hold82 (.clk(net292),
    .clkout(net2080));
 b15cbf034ar1n64x5 hold83 (.clk(net294),
    .clkout(net2081));
 b15cbf034ar1n64x5 hold84 (.clk(net2019),
    .clkout(net2082));
 b15cbf034ar1n64x5 hold85 (.clk(net237),
    .clkout(net2083));
 b15cbf034ar1n64x5 hold86 (.clk(net2605),
    .clkout(net2084));
 b15cbf034ar1n64x5 hold87 (.clk(net2085),
    .clkout(intr_gpio_o[14]));
 b15cbf034ar1n64x5 hold88 (.clk(net2603),
    .clkout(net2086));
 b15cbf034ar1n64x5 hold89 (.clk(net2087),
    .clkout(intr_gpio_o[19]));
 b15cbf034ar1n64x5 hold90 (.clk(net2121),
    .clkout(net2088));
 b15cbf034ar1n64x5 hold91 (.clk(net2089),
    .clkout(tl_o[62]));
 b15cbf034ar1n64x5 hold92 (.clk(net2607),
    .clkout(net2090));
 b15cbf034ar1n64x5 hold93 (.clk(net2091),
    .clkout(intr_gpio_o[12]));
 b15cbf034ar1n64x5 hold94 (.clk(net2617),
    .clkout(net2092));
 b15cbf034ar1n64x5 hold95 (.clk(net2093),
    .clkout(tl_o[56]));
 b15cbf034ar1n64x5 hold96 (.clk(net2619),
    .clkout(net2094));
 b15cbf034ar1n64x5 hold97 (.clk(net2095),
    .clkout(tl_o[55]));
 b15cbf034ar1n64x5 hold98 (.clk(net2611),
    .clkout(net2096));
 b15cbf034ar1n64x5 hold99 (.clk(net2097),
    .clkout(intr_gpio_o[16]));
 b15cbf034ar1n64x5 hold100 (.clk(net2620),
    .clkout(net2098));
 b15cbf034ar1n64x5 hold101 (.clk(net2099),
    .clkout(tl_o[53]));
 b15cbf034ar1n64x5 hold102 (.clk(net2621),
    .clkout(net2100));
 b15cbf034ar1n64x5 hold103 (.clk(net2101),
    .clkout(tl_o[50]));
 b15cbf034ar1n64x5 hold104 (.clk(net2622),
    .clkout(net2102));
 b15cbf034ar1n64x5 hold105 (.clk(net2103),
    .clkout(tl_o[49]));
 b15cbf034ar1n64x5 hold106 (.clk(net2623),
    .clkout(net2104));
 b15cbf034ar1n64x5 hold107 (.clk(net2105),
    .clkout(tl_o[54]));
 b15cbf034ar1n64x5 hold108 (.clk(net2614),
    .clkout(net2106));
 b15cbf034ar1n64x5 hold109 (.clk(net2107),
    .clkout(intr_gpio_o[17]));
 b15cbf034ar1n64x5 hold110 (.clk(net2612),
    .clkout(net2108));
 b15cbf034ar1n64x5 hold111 (.clk(net2109),
    .clkout(intr_gpio_o[30]));
 b15cbf034ar1n64x5 hold112 (.clk(net2613),
    .clkout(net2110));
 b15cbf034ar1n64x5 hold113 (.clk(net2111),
    .clkout(intr_gpio_o[29]));
 b15cbf034ar1n64x5 hold114 (.clk(net2615),
    .clkout(net2112));
 b15cbf034ar1n64x5 hold115 (.clk(net2113),
    .clkout(intr_gpio_o[24]));
 b15cbf034ar1n64x5 hold116 (.clk(net247),
    .clkout(net2114));
 b15cbf034ar1n64x5 hold117 (.clk(net475),
    .clkout(net2115));
 b15cbf034ar1n64x5 hold118 (.clk(net2116),
    .clkout(tl_o[19]));
 b15cbf034ar1n64x5 hold119 (.clk(net2626),
    .clkout(net2117));
 b15cbf034ar1n64x5 hold120 (.clk(net2118),
    .clkout(tl_o[51]));
 b15cbf034ar1n64x5 hold121 (.clk(net2625),
    .clkout(net2119));
 b15cbf034ar1n64x5 hold122 (.clk(net2120),
    .clkout(tl_o[52]));
 b15cbf034ar1n64x5 hold123 (.clk(net291),
    .clkout(net2121));
 b15cbf034ar1n64x5 hold124 (.clk(net2088),
    .clkout(net2122));
 b15cbf034ar1n64x5 hold125 (.clk(net2610),
    .clkout(net2123));
 b15cbf034ar1n64x5 hold126 (.clk(net2124),
    .clkout(intr_gpio_o[31]));
 b15cbf034ar1n64x5 hold127 (.clk(net2618),
    .clkout(net2125));
 b15cbf034ar1n64x5 hold128 (.clk(net2126),
    .clkout(intr_gpio_o[26]));
 b15cbf034ar1n64x5 hold129 (.clk(net2628),
    .clkout(net2127));
 b15cbf034ar1n64x5 hold130 (.clk(net2128),
    .clkout(tl_o[22]));
 b15cbf034ar1n64x5 hold131 (.clk(net2616),
    .clkout(net2129));
 b15cbf034ar1n64x5 hold132 (.clk(net2130),
    .clkout(tl_o[30]));
 b15cbf034ar1n64x5 hold133 (.clk(net2635),
    .clkout(net2131));
 b15cbf034ar1n64x5 hold134 (.clk(net2132),
    .clkout(tl_o[37]));
 b15cbf034ar1n64x5 hold135 (.clk(net261),
    .clkout(net2133));
 b15cbf034ar1n64x5 hold136 (.clk(net497),
    .clkout(net2134));
 b15cbf034ar1n64x5 hold137 (.clk(net2135),
    .clkout(tl_o[31]));
 b15cbf034ar1n64x5 hold138 (.clk(net2298),
    .clkout(net2136));
 b15cbf034ar1n64x5 hold139 (.clk(n3013),
    .clkout(net2137));
 b15cbf034ar1n64x5 hold140 (.clk(net295),
    .clkout(net2138));
 b15cbf034ar1n64x5 hold141 (.clk(net2624),
    .clkout(net2139));
 b15cbf034ar1n64x5 hold142 (.clk(net2140),
    .clkout(tl_o[27]));
 b15cbf034ar1n64x5 hold143 (.clk(net2629),
    .clkout(net2141));
 b15cbf034ar1n64x5 hold144 (.clk(net2142),
    .clkout(tl_o[29]));
 b15cbf034ar1n64x5 hold145 (.clk(net2200),
    .clkout(net2143));
 b15cbf034ar1n64x5 hold146 (.clk(net506),
    .clkout(net2144));
 b15cbf034ar1n64x5 hold147 (.clk(net505),
    .clkout(net2145));
 b15cbf034ar1n64x5 hold148 (.clk(net2632),
    .clkout(net2146));
 b15cbf034ar1n64x5 hold149 (.clk(net2147),
    .clkout(tl_o[28]));
 b15cbf034ar1n64x5 hold150 (.clk(net271),
    .clkout(net2148));
 b15cbf034ar1n64x5 hold151 (.clk(net2149),
    .clkout(tl_o[40]));
 b15cbf034ar1n64x5 hold152 (.clk(net276),
    .clkout(net2150));
 b15cbf034ar1n64x5 hold153 (.clk(net2151),
    .clkout(tl_o[45]));
 b15cbf034ar1n64x5 hold154 (.clk(net145),
    .clkout(net2152));
 b15cbf034ar1n64x5 hold155 (.clk(net2153),
    .clkout(cio_gpio_en_o[13]));
 b15cbf034ar1n64x5 hold156 (.clk(net254),
    .clkout(net2154));
 b15cbf034ar1n64x5 hold157 (.clk(net461),
    .clkout(net2155));
 b15cbf034ar1n64x5 hold158 (.clk(net246),
    .clkout(net2156));
 b15cbf034ar1n64x5 hold159 (.clk(net477),
    .clkout(net2157));
 b15cbf034ar1n64x5 hold160 (.clk(net2158),
    .clkout(tl_o[18]));
 b15cbf034ar1n64x5 hold161 (.clk(u_reg_data_in_qs[29]),
    .clkout(net2159));
 b15cbf034ar1n64x5 hold162 (.clk(n3991),
    .clkout(net2160));
 b15cbf034ar1n64x5 hold163 (.clk(u_reg_u_reg_if_N43),
    .clkout(net2161));
 b15cbf034ar1n64x5 hold164 (.clk(net152),
    .clkout(net2162));
 b15cbf034ar1n64x5 hold165 (.clk(net2163),
    .clkout(cio_gpio_en_o[1]));
 b15cbf034ar1n64x5 hold166 (.clk(net250),
    .clkout(net2164));
 b15cbf034ar1n64x5 hold167 (.clk(net467),
    .clkout(net2165));
 b15cbf034ar1n64x5 hold168 (.clk(net252),
    .clkout(net2166));
 b15cbf034ar1n64x5 hold169 (.clk(net463),
    .clkout(net2167));
 b15cbf034ar1n64x5 hold170 (.clk(net2168),
    .clkout(tl_o[23]));
 b15cbf034ar1n64x5 hold171 (.clk(net167),
    .clkout(net2169));
 b15cbf034ar1n64x5 hold172 (.clk(net2170),
    .clkout(cio_gpio_en_o[4]));
 b15cbf034ar1n64x5 hold173 (.clk(net171),
    .clkout(net2171));
 b15cbf034ar1n64x5 hold174 (.clk(net2172),
    .clkout(cio_gpio_en_o[8]));
 b15cbf034ar1n64x5 hold175 (.clk(net142),
    .clkout(net2173));
 b15cbf034ar1n64x5 hold176 (.clk(net730),
    .clkout(net2174));
 b15cbf034ar1n64x5 hold177 (.clk(net275),
    .clkout(net2175));
 b15cbf034ar1n64x5 hold178 (.clk(net2176),
    .clkout(tl_o[44]));
 b15cbf034ar1n64x5 hold179 (.clk(net2285),
    .clkout(net2177));
 b15cbf034ar1n64x5 hold180 (.clk(n3009),
    .clkout(net2178));
 b15cbf034ar1n64x5 hold181 (.clk(net270),
    .clkout(net2179));
 b15cbf034ar1n64x5 hold182 (.clk(net253),
    .clkout(net2180));
 b15cbf034ar1n64x5 hold183 (.clk(net2181),
    .clkout(tl_o[24]));
 b15cbf034ar1n64x5 hold184 (.clk(net2184),
    .clkout(net2182));
 b15cbf034ar1n64x5 hold185 (.clk(net2183),
    .clkout(tl_o[34]));
 b15cbf034ar1n64x5 hold186 (.clk(net264),
    .clkout(net2184));
 b15cbf034ar1n64x5 hold187 (.clk(net296),
    .clkout(net2185));
 b15cbf034ar1n64x5 hold188 (.clk(net154),
    .clkout(net2186));
 b15cbf034ar1n64x5 hold189 (.clk(net2187),
    .clkout(cio_gpio_en_o[21]));
 b15cbf034ar1n64x5 hold190 (.clk(u_reg_data_in_qs[25]),
    .clkout(net2188));
 b15cbf034ar1n64x5 hold191 (.clk(n3952),
    .clkout(net2189));
 b15cbf034ar1n64x5 hold192 (.clk(u_reg_u_reg_if_N39),
    .clkout(net2190));
 b15cbf034ar1n64x5 hold193 (.clk(net274),
    .clkout(net2191));
 b15cbf034ar1n64x5 hold194 (.clk(net2192),
    .clkout(tl_o[43]));
 b15cbf034ar1n64x5 hold195 (.clk(u_reg_data_in_qs[31]),
    .clkout(net2193));
 b15cbf034ar1n64x5 hold196 (.clk(n3323),
    .clkout(net2194));
 b15cbf034ar1n64x5 hold197 (.clk(u_reg_u_reg_if_N45),
    .clkout(net2195));
 b15cbf034ar1n64x5 hold198 (.clk(net156),
    .clkout(net2196));
 b15cbf034ar1n64x5 hold199 (.clk(net2197),
    .clkout(cio_gpio_en_o[23]));
 b15cbf034ar1n64x5 hold200 (.clk(net170),
    .clkout(net2198));
 b15cbf034ar1n64x5 hold201 (.clk(net2199),
    .clkout(cio_gpio_en_o[7]));
 b15cbf034ar1n64x5 hold202 (.clk(net255),
    .clkout(net2200));
 b15cbf034ar1n64x5 hold203 (.clk(n3039),
    .clkout(net2201));
 b15cbf034ar1n64x5 hold204 (.clk(net290),
    .clkout(net2202));
 b15cbf034ar1n64x5 hold205 (.clk(u_reg_data_in_qs[10]),
    .clkout(net2203));
 b15cbf034ar1n64x5 hold206 (.clk(n3836),
    .clkout(net2204));
 b15cbf034ar1n64x5 hold207 (.clk(net262),
    .clkout(net2205));
 b15cbf034ar1n64x5 hold208 (.clk(net2206),
    .clkout(tl_o[32]));
 b15cbf034ar1n64x5 hold209 (.clk(net157),
    .clkout(net2207));
 b15cbf034ar1n64x5 hold210 (.clk(net710),
    .clkout(net2208));
 b15cbf034ar1n64x5 hold211 (.clk(net151),
    .clkout(net2209));
 b15cbf034ar1n64x5 hold212 (.clk(net716),
    .clkout(net2210));
 b15cbf034ar1n64x5 hold213 (.clk(u_reg_data_in_qs[26]),
    .clkout(net2211));
 b15cbf034ar1n64x5 hold214 (.clk(n3959),
    .clkout(net2212));
 b15cbf034ar1n64x5 hold215 (.clk(u_reg_u_reg_if_N40),
    .clkout(net2213));
 b15cbf034ar1n64x5 hold216 (.clk(net2229),
    .clkout(net2214));
 b15cbf034ar1n64x5 hold217 (.clk(n2957),
    .clkout(net2215));
 b15cbf034ar1n64x5 hold218 (.clk(n2960),
    .clkout(net2216));
 b15cbf034ar1n64x5 hold219 (.clk(net297),
    .clkout(net2217));
 b15cbf034ar1n64x5 hold220 (.clk(net272),
    .clkout(net2218));
 b15cbf034ar1n64x5 hold221 (.clk(net163),
    .clkout(net2219));
 b15cbf034ar1n64x5 hold222 (.clk(net278),
    .clkout(net2220));
 b15cbf034ar1n64x5 hold223 (.clk(net168),
    .clkout(net2221));
 b15cbf034ar1n64x5 hold224 (.clk(net169),
    .clkout(net2222));
 b15cbf034ar1n64x5 hold225 (.clk(net2223),
    .clkout(cio_gpio_en_o[6]));
 b15cbf034ar1n64x5 hold226 (.clk(net146),
    .clkout(net2224));
 b15cbf034ar1n64x5 hold227 (.clk(net727),
    .clkout(net2225));
 b15cbf034ar1n64x5 hold228 (.clk(net158),
    .clkout(net2226));
 b15cbf034ar1n64x5 hold229 (.clk(net707),
    .clkout(net2227));
 b15cbf034ar1n64x5 hold230 (.clk(net150),
    .clkout(net2228));
 b15cbf034ar1n64x5 hold231 (.clk(net245),
    .clkout(net2229));
 b15cbf034ar1n64x5 hold232 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_n_intq_0_),
    .clkout(net2230));
 b15cbf034ar1n64x5 hold233 (.clk(net155),
    .clkout(net2231));
 b15cbf034ar1n64x5 hold234 (.clk(net161),
    .clkout(net2232));
 b15cbf034ar1n64x5 hold235 (.clk(net703),
    .clkout(net2233));
 b15cbf034ar1n64x5 hold236 (.clk(net147),
    .clkout(net2234));
 b15cbf034ar1n64x5 hold237 (.clk(net725),
    .clkout(net2235));
 b15cbf034ar1n64x5 hold238 (.clk(u_reg_data_in_qs[18]),
    .clkout(net2236));
 b15cbf034ar1n64x5 hold239 (.clk(n3896),
    .clkout(net2237));
 b15cbf034ar1n64x5 hold240 (.clk(n3899),
    .clkout(net2238));
 b15cbf034ar1n64x5 hold241 (.clk(u_reg_u_reg_if_N32),
    .clkout(net2239));
 b15cbf034ar1n64x5 hold242 (.clk(u_reg_data_in_qs[16]),
    .clkout(net2240));
 b15cbf034ar1n64x5 hold243 (.clk(n3886),
    .clkout(net2241));
 b15cbf034ar1n64x5 hold244 (.clk(u_reg_u_reg_if_N30),
    .clkout(net2242));
 b15cbf034ar1n64x5 hold245 (.clk(net143),
    .clkout(net2243));
 b15cbf034ar1n64x5 hold246 (.clk(u_reg_data_in_qs[28]),
    .clkout(net2244));
 b15cbf034ar1n64x5 hold247 (.clk(n3971),
    .clkout(net2245));
 b15cbf034ar1n64x5 hold248 (.clk(u_reg_u_reg_if_N42),
    .clkout(net2246));
 b15cbf034ar1n64x5 hold249 (.clk(net141),
    .clkout(net2247));
 b15cbf034ar1n64x5 hold250 (.clk(net172),
    .clkout(net2248));
 b15cbf034ar1n64x5 hold251 (.clk(net694),
    .clkout(net2249));
 b15cbf034ar1n64x5 hold252 (.clk(net164),
    .clkout(net2250));
 b15cbf034ar1n64x5 hold253 (.clk(net166),
    .clkout(net2251));
 b15cbf034ar1n64x5 hold254 (.clk(net144),
    .clkout(net2252));
 b15cbf034ar1n64x5 hold255 (.clk(gen_filter_22__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2253));
 b15cbf034ar1n64x5 hold256 (.clk(gen_filter_29__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2254));
 b15cbf034ar1n64x5 hold257 (.clk(gen_filter_21__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2255));
 b15cbf034ar1n64x5 hold258 (.clk(gen_filter_27__u_filter_stored_value_q),
    .clkout(net2256));
 b15cbf034ar1n64x5 hold259 (.clk(net265),
    .clkout(net2257));
 b15cbf034ar1n64x5 hold260 (.clk(gen_filter_3__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2258));
 b15cbf034ar1n64x5 hold261 (.clk(gen_filter_6__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2259));
 b15cbf034ar1n64x5 hold262 (.clk(gen_filter_15__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2260));
 b15cbf034ar1n64x5 hold263 (.clk(gen_filter_25__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2261));
 b15cbf034ar1n64x5 hold264 (.clk(gen_filter_23__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2262));
 b15cbf034ar1n64x5 hold265 (.clk(gen_filter_24__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2263));
 b15cbf034ar1n64x5 hold266 (.clk(gen_filter_28__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2264));
 b15cbf034ar1n64x5 hold267 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_i_sync_p_intq_0_),
    .clkout(net2265));
 b15cbf034ar1n64x5 hold268 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_p_intq_0_),
    .clkout(net2266));
 b15cbf034ar1n64x5 hold269 (.clk(gen_filter_17__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2267));
 b15cbf034ar1n64x5 hold270 (.clk(gen_filter_13__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2268));
 b15cbf034ar1n64x5 hold271 (.clk(gen_filter_9__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2269));
 b15cbf034ar1n64x5 hold272 (.clk(gen_filter_11__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2270));
 b15cbf034ar1n64x5 hold273 (.clk(gen_filter_1__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2271));
 b15cbf034ar1n64x5 hold274 (.clk(gen_filter_18__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2272));
 b15cbf034ar1n64x5 hold275 (.clk(gen_filter_27__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2273));
 b15cbf034ar1n64x5 hold276 (.clk(net244),
    .clkout(net2274));
 b15cbf034ar1n64x5 hold277 (.clk(net511),
    .clkout(net2275));
 b15cbf034ar1n64x5 hold278 (.clk(net2303),
    .clkout(net2276));
 b15cbf034ar1n64x5 hold279 (.clk(net280),
    .clkout(net2277));
 b15cbf034ar1n64x5 hold280 (.clk(net268),
    .clkout(net2278));
 b15cbf034ar1n64x5 hold281 (.clk(u_reg_data_in_qs[17]),
    .clkout(net2279));
 b15cbf034ar1n64x5 hold282 (.clk(n3895),
    .clkout(net2280));
 b15cbf034ar1n64x5 hold283 (.clk(u_reg_u_reg_if_N31),
    .clkout(net2281));
 b15cbf034ar1n64x5 hold284 (.clk(u_reg_data_in_qs[23]),
    .clkout(net2282));
 b15cbf034ar1n64x5 hold285 (.clk(n3936),
    .clkout(net2283));
 b15cbf034ar1n64x5 hold286 (.clk(u_reg_u_reg_if_N37),
    .clkout(net2284));
 b15cbf034ar1n64x5 hold287 (.clk(net249),
    .clkout(net2285));
 b15cbf034ar1n64x5 hold288 (.clk(gen_filter_7__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2286));
 b15cbf034ar1n64x5 hold289 (.clk(reg2hw_intr_ctrl_en_rising__q__22_),
    .clkout(net2287));
 b15cbf034ar1n64x5 hold290 (.clk(n3924),
    .clkout(net2288));
 b15cbf034ar1n64x5 hold291 (.clk(u_reg_u_reg_if_N36),
    .clkout(net2289));
 b15cbf034ar1n64x5 hold292 (.clk(net153),
    .clkout(net2290));
 b15cbf034ar1n64x5 hold293 (.clk(gen_filter_4__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2291));
 b15cbf034ar1n64x5 hold294 (.clk(net263),
    .clkout(net2292));
 b15cbf034ar1n64x5 hold295 (.clk(net259),
    .clkout(net2293));
 b15cbf034ar1n64x5 hold296 (.clk(reg2hw_intr_ctrl_en_lvllow__q__19_),
    .clkout(net2294));
 b15cbf034ar1n64x5 hold297 (.clk(n3331),
    .clkout(net2295));
 b15cbf034ar1n64x5 hold298 (.clk(u_reg_u_reg_if_N33),
    .clkout(net2296));
 b15cbf034ar1n64x5 hold299 (.clk(net149),
    .clkout(net2297));
 b15cbf034ar1n64x5 hold300 (.clk(net269),
    .clkout(net2298));
 b15cbf034ar1n64x5 hold301 (.clk(gen_filter_16__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2299));
 b15cbf034ar1n64x5 hold302 (.clk(gen_filter_5__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2300));
 b15cbf034ar1n64x5 hold303 (.clk(gen_filter_14__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2301));
 b15cbf034ar1n64x5 hold304 (.clk(net180),
    .clkout(net2302));
 b15cbf034ar1n64x5 hold305 (.clk(net277),
    .clkout(net2303));
 b15cbf034ar1n64x5 hold306 (.clk(net162),
    .clkout(net2304));
 b15cbf034ar1n64x5 hold307 (.clk(rst_ni),
    .clkout(net2305));
 b15cbf034ar1n64x5 hold308 (.clk(u_reg_data_in_qs[2]),
    .clkout(net2306));
 b15cbf034ar1n64x5 hold309 (.clk(u_reg_u_reg_if_N16),
    .clkout(net2307));
 b15cbf034ar1n64x5 hold310 (.clk(net266),
    .clkout(net2308));
 b15cbf034ar1n64x5 hold311 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_i_sync_n_intq_0_),
    .clkout(net2309));
 b15cbf034ar1n64x5 hold312 (.clk(gen_filter_12__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2310));
 b15cbf034ar1n64x5 hold313 (.clk(net148),
    .clkout(net2311));
 b15cbf034ar1n64x5 hold314 (.clk(net273),
    .clkout(net2312));
 b15cbf034ar1n64x5 hold315 (.clk(net181),
    .clkout(net2313));
 b15cbf034ar1n64x5 hold316 (.clk(gen_filter_25__u_filter_stored_value_q),
    .clkout(net2314));
 b15cbf034ar1n64x5 hold317 (.clk(u_reg_data_in_qs[4]),
    .clkout(net2315));
 b15cbf034ar1n64x5 hold318 (.clk(net165),
    .clkout(net2316));
 b15cbf034ar1n64x5 hold319 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_state_q[0]),
    .clkout(net2317));
 b15cbf034ar1n64x5 hold320 (.clk(gen_alert_tx_0__u_prim_alert_sender_n1),
    .clkout(net2318));
 b15cbf034ar1n64x5 hold321 (.clk(gen_filter_24__u_filter_filter_q),
    .clkout(net2319));
 b15cbf034ar1n64x5 hold322 (.clk(gen_filter_24__u_filter_diff_ctr_d[1]),
    .clkout(net2320));
 b15cbf034ar1n64x5 hold323 (.clk(reg2hw_intr_ctrl_en_rising__q__21_),
    .clkout(net2321));
 b15cbf034ar1n64x5 hold324 (.clk(u_reg_u_reg_if_N35),
    .clkout(net2322));
 b15cbf034ar1n64x5 hold325 (.clk(gen_filter_24__u_filter_diff_ctr_q[3]),
    .clkout(net2323));
 b15cbf034ar1n64x5 hold326 (.clk(gen_filter_24__u_filter_diff_ctr_d[3]),
    .clkout(net2324));
 b15cbf034ar1n64x5 hold327 (.clk(gen_filter_2__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2325));
 b15cbf034ar1n64x5 hold328 (.clk(gen_filter_12__u_filter_filter_q),
    .clkout(net2326));
 b15cbf034ar1n64x5 hold329 (.clk(n2864),
    .clkout(net2327));
 b15cbf034ar1n64x5 hold330 (.clk(gen_filter_12__u_filter_diff_ctr_d[2]),
    .clkout(net2328));
 b15cbf034ar1n64x5 hold331 (.clk(gen_filter_13__u_filter_diff_ctr_q[0]),
    .clkout(net2329));
 b15cbf034ar1n64x5 hold332 (.clk(gen_filter_13__u_filter_diff_ctr_d[1]),
    .clkout(net2330));
 b15cbf034ar1n64x5 hold333 (.clk(gen_filter_16__u_filter_diff_ctr_q[2]),
    .clkout(net2331));
 b15cbf034ar1n64x5 hold334 (.clk(n2861),
    .clkout(net2332));
 b15cbf034ar1n64x5 hold335 (.clk(gen_filter_31__u_filter_stored_value_q),
    .clkout(net2333));
 b15cbf034ar1n64x5 hold336 (.clk(gen_filter_22__u_filter_diff_ctr_q[0]),
    .clkout(net2334));
 b15cbf034ar1n64x5 hold337 (.clk(n2684),
    .clkout(net2335));
 b15cbf034ar1n64x5 hold338 (.clk(gen_filter_22__u_filter_diff_ctr_d[3]),
    .clkout(net2336));
 b15cbf034ar1n64x5 hold339 (.clk(data_in_q[29]),
    .clkout(net2337));
 b15cbf034ar1n64x5 hold340 (.clk(u_reg_u_intr_state_wr_data[29]),
    .clkout(net2338));
 b15cbf034ar1n64x5 hold341 (.clk(reg2hw_intr_enable__q__11_),
    .clkout(net2339));
 b15cbf034ar1n64x5 hold342 (.clk(n3845),
    .clkout(net2340));
 b15cbf034ar1n64x5 hold343 (.clk(u_reg_u_reg_if_N25),
    .clkout(net2341));
 b15cbf034ar1n64x5 hold344 (.clk(u_reg_data_in_qs[27]),
    .clkout(net2342));
 b15cbf034ar1n64x5 hold345 (.clk(u_reg_u_reg_if_N41),
    .clkout(net2343));
 b15cbf034ar1n64x5 hold346 (.clk(gen_filter_12__u_filter_diff_ctr_q[3]),
    .clkout(net2344));
 b15cbf034ar1n64x5 hold347 (.clk(u_reg_data_in_qs[0]),
    .clkout(net2345));
 b15cbf034ar1n64x5 hold348 (.clk(net200),
    .clkout(net2346));
 b15cbf034ar1n64x5 hold349 (.clk(gen_filter_30__u_filter_stored_value_q),
    .clkout(net2347));
 b15cbf034ar1n64x5 hold350 (.clk(gen_filter_31__u_filter_filter_synced),
    .clkout(net2348));
 b15cbf034ar1n64x5 hold351 (.clk(gen_filter_19__u_filter_stored_value_q),
    .clkout(net2349));
 b15cbf034ar1n64x5 hold352 (.clk(gen_filter_12__u_filter_diff_ctr_q[0]),
    .clkout(net2350));
 b15cbf034ar1n64x5 hold353 (.clk(gen_filter_17__u_filter_filter_q),
    .clkout(net2351));
 b15cbf034ar1n64x5 hold354 (.clk(gen_filter_17__u_filter_diff_ctr_d[1]),
    .clkout(net2352));
 b15cbf034ar1n64x5 hold355 (.clk(gen_filter_18__u_filter_diff_ctr_q[3]),
    .clkout(net2353));
 b15cbf034ar1n64x5 hold356 (.clk(gen_filter_5__u_filter_stored_value_q),
    .clkout(net2354));
 b15cbf034ar1n64x5 hold357 (.clk(u_reg_u_data_in_wr_data[5]),
    .clkout(net2355));
 b15cbf034ar1n64x5 hold358 (.clk(gen_filter_30__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2356));
 b15cbf034ar1n64x5 hold359 (.clk(gen_filter_18__u_filter_diff_ctr_q[0]),
    .clkout(net2357));
 b15cbf034ar1n64x5 hold360 (.clk(gen_filter_19__u_filter_filter_q),
    .clkout(net2358));
 b15cbf034ar1n64x5 hold361 (.clk(gen_filter_19__u_filter_diff_ctr_d[0]),
    .clkout(net2359));
 b15cbf034ar1n64x5 hold362 (.clk(gen_filter_17__u_filter_diff_ctr_q[3]),
    .clkout(net2360));
 b15cbf034ar1n64x5 hold363 (.clk(gen_filter_17__u_filter_diff_ctr_d[2]),
    .clkout(net2361));
 b15cbf034ar1n64x5 hold364 (.clk(gen_filter_29__u_filter_filter_synced),
    .clkout(net2362));
 b15cbf034ar1n64x5 hold365 (.clk(gen_filter_13__u_filter_diff_ctr_q[2]),
    .clkout(net2363));
 b15cbf034ar1n64x5 hold366 (.clk(gen_filter_13__u_filter_diff_ctr_d[2]),
    .clkout(net2364));
 b15cbf034ar1n64x5 hold367 (.clk(gen_filter_30__u_filter_filter_q),
    .clkout(net2365));
 b15cbf034ar1n64x5 hold368 (.clk(gen_filter_30__u_filter_diff_ctr_d[0]),
    .clkout(net2366));
 b15cbf034ar1n64x5 hold369 (.clk(gen_filter_19__u_filter_diff_ctr_q[2]),
    .clkout(net2367));
 b15cbf034ar1n64x5 hold370 (.clk(gen_filter_16__u_filter_diff_ctr_q[3]),
    .clkout(net2368));
 b15cbf034ar1n64x5 hold371 (.clk(gen_filter_16__u_filter_diff_ctr_d[2]),
    .clkout(net2369));
 b15cbf034ar1n64x5 hold372 (.clk(u_reg_data_in_qs[30]),
    .clkout(net2370));
 b15cbf034ar1n64x5 hold373 (.clk(u_reg_u_reg_if_N44),
    .clkout(net2371));
 b15cbf034ar1n64x5 hold374 (.clk(gen_filter_11__u_filter_filter_q),
    .clkout(net2372));
 b15cbf034ar1n64x5 hold375 (.clk(gen_filter_11__u_filter_diff_ctr_d[3]),
    .clkout(net2373));
 b15cbf034ar1n64x5 hold376 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nd),
    .clkout(net2374));
 b15cbf034ar1n64x5 hold377 (.clk(gen_filter_23__u_filter_diff_ctr_q[2]),
    .clkout(net2375));
 b15cbf034ar1n64x5 hold378 (.clk(n2729),
    .clkout(net2376));
 b15cbf034ar1n64x5 hold379 (.clk(gen_filter_23__u_filter_diff_ctr_d[2]),
    .clkout(net2377));
 b15cbf034ar1n64x5 hold380 (.clk(gen_filter_13__u_filter_filter_q),
    .clkout(net2378));
 b15cbf034ar1n64x5 hold381 (.clk(gen_filter_22__u_filter_filter_q),
    .clkout(net2379));
 b15cbf034ar1n64x5 hold382 (.clk(n2706),
    .clkout(net2380));
 b15cbf034ar1n64x5 hold383 (.clk(gen_filter_11__u_filter_diff_ctr_q[3]),
    .clkout(net2381));
 b15cbf034ar1n64x5 hold384 (.clk(gen_filter_11__u_filter_diff_ctr_d[2]),
    .clkout(net2382));
 b15cbf034ar1n64x5 hold385 (.clk(gen_filter_22__u_filter_diff_ctr_q[1]),
    .clkout(net2383));
 b15cbf034ar1n64x5 hold386 (.clk(n2683),
    .clkout(net2384));
 b15cbf034ar1n64x5 hold387 (.clk(gen_filter_0__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2385));
 b15cbf034ar1n64x5 hold388 (.clk(gen_filter_0__u_filter_filter_q),
    .clkout(net2386));
 b15cbf034ar1n64x5 hold389 (.clk(gen_filter_0__u_filter_diff_ctr_d[0]),
    .clkout(net2387));
 b15cbf034ar1n64x5 hold390 (.clk(gen_filter_17__u_filter_diff_ctr_q[2]),
    .clkout(net2388));
 b15cbf034ar1n64x5 hold391 (.clk(n2903),
    .clkout(net2389));
 b15cbf034ar1n64x5 hold392 (.clk(gen_filter_20__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2390));
 b15cbf034ar1n64x5 hold393 (.clk(gen_filter_29__u_filter_diff_ctr_q[0]),
    .clkout(net2391));
 b15cbf034ar1n64x5 hold394 (.clk(gen_filter_29__u_filter_diff_ctr_d[0]),
    .clkout(net2392));
 b15cbf034ar1n64x5 hold395 (.clk(gen_filter_10__u_filter_diff_ctr_q[3]),
    .clkout(net2393));
 b15cbf034ar1n64x5 hold396 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_level_q),
    .clkout(net2394));
 b15cbf034ar1n64x5 hold397 (.clk(gen_filter_10__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2395));
 b15cbf034ar1n64x5 hold398 (.clk(gen_filter_2__u_filter_diff_ctr_q[1]),
    .clkout(net2396));
 b15cbf034ar1n64x5 hold399 (.clk(gen_filter_2__u_filter_diff_ctr_d[1]),
    .clkout(net2397));
 b15cbf034ar1n64x5 hold400 (.clk(gen_filter_6__u_filter_filter_q),
    .clkout(net2398));
 b15cbf034ar1n64x5 hold401 (.clk(gen_filter_6__u_filter_diff_ctr_d[1]),
    .clkout(net2399));
 b15cbf034ar1n64x5 hold402 (.clk(gen_filter_6__u_filter_diff_ctr_q[3]),
    .clkout(net2400));
 b15cbf034ar1n64x5 hold403 (.clk(gen_filter_6__u_filter_diff_ctr_d[0]),
    .clkout(net2401));
 b15cbf034ar1n64x5 hold404 (.clk(u_reg_data_in_qs[24]),
    .clkout(net2402));
 b15cbf034ar1n64x5 hold405 (.clk(u_reg_u_reg_if_N38),
    .clkout(net2403));
 b15cbf034ar1n64x5 hold406 (.clk(gen_filter_2__u_filter_diff_ctr_q[3]),
    .clkout(net2404));
 b15cbf034ar1n64x5 hold407 (.clk(gen_filter_2__u_filter_diff_ctr_d[3]),
    .clkout(net2405));
 b15cbf034ar1n64x5 hold408 (.clk(gen_filter_5__u_filter_diff_ctr_q[3]),
    .clkout(net2406));
 b15cbf034ar1n64x5 hold409 (.clk(n2818),
    .clkout(net2407));
 b15cbf034ar1n64x5 hold410 (.clk(gen_filter_5__u_filter_diff_ctr_d[1]),
    .clkout(net2408));
 b15cbf034ar1n64x5 hold411 (.clk(gen_filter_30__u_filter_diff_ctr_q[3]),
    .clkout(net2409));
 b15cbf034ar1n64x5 hold412 (.clk(gen_filter_29__u_filter_filter_q),
    .clkout(net2410));
 b15cbf034ar1n64x5 hold413 (.clk(gen_filter_29__u_filter_diff_ctr_d[2]),
    .clkout(net2411));
 b15cbf034ar1n64x5 hold414 (.clk(gen_filter_0__u_filter_diff_ctr_q[3]),
    .clkout(net2412));
 b15cbf034ar1n64x5 hold415 (.clk(n2807),
    .clkout(net2413));
 b15cbf034ar1n64x5 hold416 (.clk(gen_filter_14__u_filter_stored_value_q),
    .clkout(net2414));
 b15cbf034ar1n64x5 hold417 (.clk(gen_filter_5__u_filter_filter_q),
    .clkout(net2415));
 b15cbf034ar1n64x5 hold418 (.clk(gen_filter_5__u_filter_diff_ctr_d[0]),
    .clkout(net2416));
 b15cbf034ar1n64x5 hold419 (.clk(gen_filter_6__u_filter_diff_ctr_q[2]),
    .clkout(net2417));
 b15cbf034ar1n64x5 hold420 (.clk(n2692),
    .clkout(net2418));
 b15cbf034ar1n64x5 hold421 (.clk(gen_filter_6__u_filter_diff_ctr_d[2]),
    .clkout(net2419));
 b15cbf034ar1n64x5 hold422 (.clk(gen_filter_20__u_filter_diff_ctr_q[0]),
    .clkout(net2420));
 b15cbf034ar1n64x5 hold423 (.clk(gen_filter_20__u_filter_diff_ctr_d[0]),
    .clkout(net2421));
 b15cbf034ar1n64x5 hold424 (.clk(u_reg_data_in_qs[14]),
    .clkout(net2422));
 b15cbf034ar1n64x5 hold425 (.clk(u_reg_u_reg_if_N28),
    .clkout(net2423));
 b15cbf034ar1n64x5 hold426 (.clk(gen_filter_1__u_filter_diff_ctr_q[3]),
    .clkout(net2424));
 b15cbf034ar1n64x5 hold427 (.clk(gen_filter_1__u_filter_diff_ctr_d[3]),
    .clkout(net2425));
 b15cbf034ar1n64x5 hold428 (.clk(gen_filter_11__u_filter_diff_ctr_q[0]),
    .clkout(net2426));
 b15cbf034ar1n64x5 hold429 (.clk(gen_filter_16__u_filter_filter_q),
    .clkout(net2427));
 b15cbf034ar1n64x5 hold430 (.clk(data_in_q[28]),
    .clkout(net2428));
 b15cbf034ar1n64x5 hold431 (.clk(n3729),
    .clkout(net2429));
 b15cbf034ar1n64x5 hold432 (.clk(gen_filter_2__u_filter_diff_ctr_q[0]),
    .clkout(net2430));
 b15cbf034ar1n64x5 hold433 (.clk(gen_filter_2__u_filter_diff_ctr_d[0]),
    .clkout(net2431));
 b15cbf034ar1n64x5 hold434 (.clk(gen_filter_25__u_filter_diff_ctr_q[2]),
    .clkout(net2432));
 b15cbf034ar1n64x5 hold435 (.clk(n3995),
    .clkout(net2433));
 b15cbf034ar1n64x5 hold436 (.clk(gen_filter_25__u_filter_diff_ctr_d[2]),
    .clkout(net2434));
 b15cbf034ar1n64x5 hold437 (.clk(gen_filter_20__u_filter_diff_ctr_q[3]),
    .clkout(net2435));
 b15cbf034ar1n64x5 hold438 (.clk(n2923),
    .clkout(net2436));
 b15cbf034ar1n64x5 hold439 (.clk(gen_filter_20__u_filter_diff_ctr_d[1]),
    .clkout(net2437));
 b15cbf034ar1n64x5 hold440 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_level_q),
    .clkout(net2438));
 b15cbf034ar1n64x5 hold441 (.clk(gen_alert_tx_0__u_prim_alert_sender_ack_level),
    .clkout(net2439));
 b15cbf034ar1n64x5 hold442 (.clk(gen_filter_27__u_filter_diff_ctr_q[3]),
    .clkout(net2440));
 b15cbf034ar1n64x5 hold443 (.clk(gen_filter_27__u_filter_diff_ctr_d[2]),
    .clkout(net2441));
 b15cbf034ar1n64x5 hold444 (.clk(gen_filter_29__u_filter_diff_ctr_q[3]),
    .clkout(net2442));
 b15cbf034ar1n64x5 hold445 (.clk(gen_alert_tx_0__u_prim_alert_sender_ping_set_q),
    .clkout(net2443));
 b15cbf034ar1n64x5 hold446 (.clk(gen_alert_tx_0__u_prim_alert_sender_ping_set_d),
    .clkout(net2444));
 b15cbf034ar1n64x5 hold447 (.clk(u_reg_data_in_qs[13]),
    .clkout(net2445));
 b15cbf034ar1n64x5 hold448 (.clk(u_reg_err_q),
    .clkout(net2446));
 b15cbf034ar1n64x5 hold449 (.clk(gen_filter_5__u_filter_diff_ctr_q[2]),
    .clkout(net2447));
 b15cbf034ar1n64x5 hold450 (.clk(n2731),
    .clkout(net2448));
 b15cbf034ar1n64x5 hold451 (.clk(gen_filter_27__u_filter_filter_q),
    .clkout(net2449));
 b15cbf034ar1n64x5 hold452 (.clk(gen_filter_1__u_filter_diff_ctr_q[1]),
    .clkout(net2450));
 b15cbf034ar1n64x5 hold453 (.clk(gen_filter_1__u_filter_diff_ctr_d[1]),
    .clkout(net2451));
 b15cbf034ar1n64x5 hold454 (.clk(gen_filter_20__u_filter_diff_ctr_q[2]),
    .clkout(net2452));
 b15cbf034ar1n64x5 hold455 (.clk(n2725),
    .clkout(net2453));
 b15cbf034ar1n64x5 hold456 (.clk(gen_filter_28__u_filter_filter_q),
    .clkout(net2454));
 b15cbf034ar1n64x5 hold457 (.clk(gen_filter_28__u_filter_diff_ctr_d[3]),
    .clkout(net2455));
 b15cbf034ar1n64x5 hold458 (.clk(gen_filter_8__u_filter_filter_synced),
    .clkout(net2456));
 b15cbf034ar1n64x5 hold459 (.clk(gen_filter_24__u_filter_stored_value_q),
    .clkout(net2457));
 b15cbf034ar1n64x5 hold460 (.clk(gen_filter_27__u_filter_diff_ctr_q[1]),
    .clkout(net2458));
 b15cbf034ar1n64x5 hold461 (.clk(gen_filter_27__u_filter_diff_ctr_d[1]),
    .clkout(net2459));
 b15cbf034ar1n64x5 hold462 (.clk(gen_filter_16__u_filter_diff_ctr_q[1]),
    .clkout(net2460));
 b15cbf034ar1n64x5 hold463 (.clk(gen_filter_16__u_filter_diff_ctr_d[1]),
    .clkout(net2461));
 b15cbf034ar1n64x5 hold464 (.clk(gen_filter_14__u_filter_diff_ctr_q[2]),
    .clkout(net2462));
 b15cbf034ar1n64x5 hold465 (.clk(n2776),
    .clkout(net2463));
 b15cbf034ar1n64x5 hold466 (.clk(gen_filter_14__u_filter_diff_ctr_d[0]),
    .clkout(net2464));
 b15cbf034ar1n64x5 hold467 (.clk(gen_filter_2__u_filter_stored_value_q),
    .clkout(net2465));
 b15cbf034ar1n64x5 hold468 (.clk(reg2hw_intr_state__q__6_),
    .clkout(net2466));
 b15cbf034ar1n64x5 hold469 (.clk(gen_filter_21__u_filter_diff_ctr_q[2]),
    .clkout(net2467));
 b15cbf034ar1n64x5 hold470 (.clk(n2709),
    .clkout(net2468));
 b15cbf034ar1n64x5 hold471 (.clk(gen_filter_21__u_filter_diff_ctr_d[2]),
    .clkout(net2469));
 b15cbf034ar1n64x5 hold472 (.clk(data_in_q[27]),
    .clkout(net2470));
 b15cbf034ar1n64x5 hold473 (.clk(gen_filter_29__u_filter_diff_ctr_q[1]),
    .clkout(net2471));
 b15cbf034ar1n64x5 hold474 (.clk(n2757),
    .clkout(net2472));
 b15cbf034ar1n64x5 hold475 (.clk(gen_filter_17__u_filter_diff_ctr_q[0]),
    .clkout(net2473));
 b15cbf034ar1n64x5 hold476 (.clk(gen_filter_19__u_filter_diff_ctr_q[3]),
    .clkout(net2474));
 b15cbf034ar1n64x5 hold477 (.clk(gen_filter_19__u_filter_diff_ctr_d[1]),
    .clkout(net2475));
 b15cbf034ar1n64x5 hold478 (.clk(gen_filter_30__u_filter_diff_ctr_q[2]),
    .clkout(net2476));
 b15cbf034ar1n64x5 hold479 (.clk(gen_filter_14__u_filter_diff_ctr_q[3]),
    .clkout(net2477));
 b15cbf034ar1n64x5 hold480 (.clk(net159),
    .clkout(net2478));
 b15cbf034ar1n64x5 hold481 (.clk(gen_filter_26__u_filter_filter_q),
    .clkout(net2479));
 b15cbf034ar1n64x5 hold482 (.clk(gen_filter_26__u_filter_diff_ctr_d[3]),
    .clkout(net2480));
 b15cbf034ar1n64x5 hold483 (.clk(gen_filter_8__u_filter_gen_async_prim_flop_2sync_intq_0_),
    .clkout(net2481));
 b15cbf034ar1n64x5 hold484 (.clk(reg2hw_intr_state__q__9_),
    .clkout(net2482));
 b15cbf034ar1n64x5 hold485 (.clk(intr_hw_N23),
    .clkout(net2483));
 b15cbf034ar1n64x5 hold486 (.clk(reg2hw_intr_enable__q__8_),
    .clkout(net2484));
 b15cbf034ar1n64x5 hold487 (.clk(gen_filter_3__u_filter_filter_q),
    .clkout(net2485));
 b15cbf034ar1n64x5 hold488 (.clk(gen_filter_3__u_filter_diff_ctr_d[1]),
    .clkout(net2486));
 b15cbf034ar1n64x5 hold489 (.clk(gen_filter_1__u_filter_diff_ctr_q[2]),
    .clkout(net2487));
 b15cbf034ar1n64x5 hold490 (.clk(gen_filter_1__u_filter_diff_ctr_d[2]),
    .clkout(net2488));
 b15cbf034ar1n64x5 hold491 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ack_gen_async_diff_nd),
    .clkout(net2489));
 b15cbf034ar1n64x5 hold492 (.clk(gen_filter_9__u_filter_filter_q),
    .clkout(net2490));
 b15cbf034ar1n64x5 hold493 (.clk(gen_filter_9__u_filter_diff_ctr_d[3]),
    .clkout(net2491));
 b15cbf034ar1n64x5 hold494 (.clk(gen_filter_8__u_filter_diff_ctr_q[2]),
    .clkout(net2492));
 b15cbf034ar1n64x5 hold495 (.clk(n2762),
    .clkout(net2493));
 b15cbf034ar1n64x5 hold496 (.clk(gen_filter_8__u_filter_diff_ctr_d[1]),
    .clkout(net2494));
 b15cbf034ar1n64x5 hold497 (.clk(reg2hw_intr_state__q__25_),
    .clkout(net2495));
 b15cbf034ar1n64x5 hold498 (.clk(u_reg_u_intr_state_wr_data[25]),
    .clkout(net2496));
 b15cbf034ar1n64x5 hold499 (.clk(gen_filter_12__u_filter_diff_ctr_q[1]),
    .clkout(net2497));
 b15cbf034ar1n64x5 hold500 (.clk(reg2hw_ctrl_en_input_filter__q__8_),
    .clkout(net2498));
 b15cbf034ar1n64x5 hold501 (.clk(gen_filter_1__u_filter_diff_ctr_q[0]),
    .clkout(net2499));
 b15cbf034ar1n64x5 hold502 (.clk(gen_filter_1__u_filter_diff_ctr_d[0]),
    .clkout(net2500));
 b15cbf034ar1n64x5 hold503 (.clk(gen_filter_22__u_filter_filter_synced),
    .clkout(net2501));
 b15cbf034ar1n64x5 hold504 (.clk(data_in_q[17]),
    .clkout(net2502));
 b15cbf034ar1n64x5 hold505 (.clk(gen_filter_4__u_filter_diff_ctr_q[2]),
    .clkout(net2503));
 b15cbf034ar1n64x5 hold506 (.clk(gen_filter_4__u_filter_diff_ctr_d[2]),
    .clkout(net2504));
 b15cbf034ar1n64x5 hold507 (.clk(data_in_q[16]),
    .clkout(net2505));
 b15cbf034ar1n64x5 hold508 (.clk(gen_filter_0__u_filter_diff_ctr_q[2]),
    .clkout(net2506));
 b15cbf034ar1n64x5 hold509 (.clk(n2736),
    .clkout(net2507));
 b15cbf034ar1n64x5 hold510 (.clk(gen_filter_0__u_filter_diff_ctr_d[2]),
    .clkout(net2508));
 b15cbf034ar1n64x5 hold511 (.clk(gen_filter_25__u_filter_diff_ctr_q[0]),
    .clkout(net2509));
 b15cbf034ar1n64x5 hold512 (.clk(gen_filter_22__u_filter_diff_ctr_q[0]),
    .clkout(net2510));
 b15cbf034ar1n64x5 hold513 (.clk(gen_filter_3__u_filter_diff_ctr_q[3]),
    .clkout(net2511));
 b15cbf034ar1n64x5 hold514 (.clk(gen_filter_2__u_filter_diff_ctr_q[2]),
    .clkout(net2512));
 b15cbf034ar1n64x5 hold515 (.clk(n2845),
    .clkout(net2513));
 b15cbf034ar1n64x5 hold516 (.clk(gen_filter_2__u_filter_diff_ctr_d[2]),
    .clkout(net2514));
 b15cbf034ar1n64x5 hold517 (.clk(gen_filter_15__u_filter_diff_ctr_q[2]),
    .clkout(net2515));
 b15cbf034ar1n64x5 hold518 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_pd),
    .clkout(net2516));
 b15cbf034ar1n64x5 hold519 (.clk(gen_filter_16__u_filter_diff_ctr_q[0]),
    .clkout(net2517));
 b15cbf034ar1n64x5 hold520 (.clk(reg2hw_intr_ctrl_en_lvllow__q__20_),
    .clkout(net2518));
 b15cbf034ar1n64x5 hold521 (.clk(reg2hw_intr_enable__q__7_),
    .clkout(net2519));
 b15cbf034ar1n64x5 hold522 (.clk(reg2hw_intr_enable__q__14_),
    .clkout(net2520));
 b15cbf034ar1n64x5 hold523 (.clk(reg2hw_intr_state__q__1_),
    .clkout(net2521));
 b15cbf034ar1n64x5 hold524 (.clk(gen_filter_26__u_filter_diff_ctr_q[3]),
    .clkout(net2522));
 b15cbf034ar1n64x5 hold525 (.clk(n2790),
    .clkout(net2523));
 b15cbf034ar1n64x5 hold526 (.clk(gen_filter_26__u_filter_diff_ctr_d[1]),
    .clkout(net2524));
 b15cbf034ar1n64x5 hold527 (.clk(gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .clkout(net2525));
 b15cbf034ar1n64x5 hold528 (.clk(gen_filter_27__u_filter_diff_ctr_q[0]),
    .clkout(net2526));
 b15cbf034ar1n64x5 hold529 (.clk(gen_filter_21__u_filter_filter_q),
    .clkout(net2527));
 b15cbf034ar1n64x5 hold530 (.clk(gen_filter_23__u_filter_filter_q),
    .clkout(net2528));
 b15cbf034ar1n64x5 hold531 (.clk(gen_filter_23__u_filter_diff_ctr_d[1]),
    .clkout(net2529));
 b15cbf034ar1n64x5 hold532 (.clk(net174),
    .clkout(net2530));
 b15cbf034ar1n64x5 hold533 (.clk(gen_filter_4__u_filter_filter_q),
    .clkout(net2531));
 b15cbf034ar1n64x5 hold534 (.clk(gen_filter_4__u_filter_diff_ctr_d[0]),
    .clkout(net2532));
 b15cbf034ar1n64x5 hold535 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_diff_nd),
    .clkout(net2533));
 b15cbf034ar1n64x5 hold536 (.clk(gen_filter_8__u_filter_diff_ctr_q[3]),
    .clkout(net2534));
 b15cbf034ar1n64x5 hold537 (.clk(gen_filter_31__u_filter_diff_ctr_q[2]),
    .clkout(net2535));
 b15cbf034ar1n64x5 hold538 (.clk(gen_filter_31__u_filter_diff_ctr_d[2]),
    .clkout(net2536));
 b15cbf034ar1n64x5 hold539 (.clk(gen_filter_7__u_filter_filter_q),
    .clkout(net2537));
 b15cbf034ar1n64x5 hold540 (.clk(gen_filter_7__u_filter_diff_ctr_d[1]),
    .clkout(net2538));
 b15cbf034ar1n64x5 hold541 (.clk(data_in_q[9]),
    .clkout(net2539));
 b15cbf034ar1n64x5 hold542 (.clk(gen_filter_28__u_filter_stored_value_q),
    .clkout(net2540));
 b15cbf034ar1n64x5 hold543 (.clk(gen_filter_21__u_filter_filter_synced),
    .clkout(net2541));
 b15cbf034ar1n64x5 hold544 (.clk(reg2hw_intr_ctrl_en_rising__q__3_),
    .clkout(net2542));
 b15cbf034ar1n64x5 hold545 (.clk(gen_filter_28__u_filter_diff_ctr_q[2]),
    .clkout(net2543));
 b15cbf034ar1n64x5 hold546 (.clk(n2783),
    .clkout(net2544));
 b15cbf034ar1n64x5 hold547 (.clk(gen_filter_17__u_filter_filter_synced),
    .clkout(net2545));
 b15cbf034ar1n64x5 hold548 (.clk(gen_filter_7__u_filter_diff_ctr_q[3]),
    .clkout(net2546));
 b15cbf034ar1n64x5 hold549 (.clk(gen_filter_0__u_filter_filter_synced),
    .clkout(net2547));
 b15cbf034ar1n64x5 hold550 (.clk(net160),
    .clkout(net2548));
 b15cbf034ar1n64x5 hold551 (.clk(tl_i[42]),
    .clkout(net2549));
 b15cbf034ar1n64x5 hold552 (.clk(gen_filter_28__u_filter_diff_ctr_q[3]),
    .clkout(net2550));
 b15cbf034ar1n64x5 hold553 (.clk(gen_filter_12__u_filter_diff_ctr_q[2]),
    .clkout(net2551));
 b15cbf034ar1n64x5 hold554 (.clk(gen_filter_21__u_filter_diff_ctr_q[3]),
    .clkout(net2552));
 b15cbf034ar1n64x5 hold555 (.clk(gen_filter_26__u_filter_diff_ctr_q[0]),
    .clkout(net2553));
 b15cbf034ar1n64x5 hold556 (.clk(gen_filter_11__u_filter_diff_ctr_q[1]),
    .clkout(net2554));
 b15cbf034ar1n64x5 hold557 (.clk(gen_filter_11__u_filter_filter_synced),
    .clkout(net2555));
 b15cbf034ar1n64x5 hold558 (.clk(gen_filter_7__u_filter_diff_ctr_q[2]),
    .clkout(net2556));
 b15cbf034ar1n64x5 hold559 (.clk(reg2hw_intr_state__q__24_),
    .clkout(net2557));
 b15cbf034ar1n64x5 hold560 (.clk(gen_filter_7__u_filter_diff_ctr_q[1]),
    .clkout(net2558));
 b15cbf034ar1n64x5 hold561 (.clk(reg2hw_intr_state__q__5_),
    .clkout(net2559));
 b15cbf034ar1n64x5 hold562 (.clk(data_in_q[8]),
    .clkout(net2560));
 b15cbf034ar1n64x5 hold563 (.clk(gen_filter_31__u_filter_diff_ctr_q[3]),
    .clkout(net2561));
 b15cbf034ar1n64x5 hold564 (.clk(reg2hw_intr_enable__q__1_),
    .clkout(net2562));
 b15cbf034ar1n64x5 hold565 (.clk(reg2hw_intr_state__q__4_),
    .clkout(net2563));
 b15cbf034ar1n64x5 hold566 (.clk(gen_alert_tx_0__u_prim_alert_sender_u_decode_ping_gen_async_state_q[1]),
    .clkout(net2564));
 b15cbf034ar1n64x5 hold567 (.clk(reg2hw_ctrl_en_input_filter__q__6_),
    .clkout(net2565));
 b15cbf034ar1n64x5 hold568 (.clk(gen_filter_11__u_filter_diff_ctr_q[2]),
    .clkout(net2566));
 b15cbf034ar1n64x5 hold569 (.clk(gen_filter_9__u_filter_stored_value_q),
    .clkout(net2567));
 b15cbf034ar1n64x5 hold570 (.clk(gen_filter_10__u_filter_stored_value_q),
    .clkout(net2568));
 b15cbf034ar1n64x5 hold571 (.clk(reg2hw_intr_state__q__22_),
    .clkout(net2569));
 b15cbf034ar1n64x5 hold572 (.clk(net205),
    .clkout(net2570));
 b15cbf034ar1n64x5 hold573 (.clk(net2003),
    .clkout(net2571));
 b15cbf034ar1n64x5 hold574 (.clk(net222),
    .clkout(net2572));
 b15cbf034ar1n64x5 hold575 (.clk(net2005),
    .clkout(net2573));
 b15cbf034ar1n64x5 hold576 (.clk(net211),
    .clkout(net2574));
 b15cbf034ar1n64x5 hold577 (.clk(net2009),
    .clkout(net2575));
 b15cbf034ar1n64x5 hold578 (.clk(net207),
    .clkout(net2576));
 b15cbf034ar1n64x5 hold579 (.clk(net2015),
    .clkout(net2577));
 b15cbf034ar1n64x5 hold580 (.clk(net206),
    .clkout(net2578));
 b15cbf034ar1n64x5 hold581 (.clk(net2021),
    .clkout(net2579));
 b15cbf034ar1n64x5 hold582 (.clk(net216),
    .clkout(net2580));
 b15cbf034ar1n64x5 hold583 (.clk(net2017),
    .clkout(net2581));
 b15cbf034ar1n64x5 hold584 (.clk(net140),
    .clkout(net2582));
 b15cbf034ar1n64x5 hold585 (.clk(net2037),
    .clkout(net2583));
 b15cbf034ar1n64x5 hold586 (.clk(net139),
    .clkout(net2584));
 b15cbf034ar1n64x5 hold587 (.clk(net2028),
    .clkout(net2585));
 b15cbf034ar1n64x5 hold588 (.clk(net227),
    .clkout(net2586));
 b15cbf034ar1n64x5 hold589 (.clk(net2023),
    .clkout(net2587));
 b15cbf034ar1n64x5 hold590 (.clk(net225),
    .clkout(net2588));
 b15cbf034ar1n64x5 hold591 (.clk(net2044),
    .clkout(net2589));
 b15cbf034ar1n64x5 hold592 (.clk(net224),
    .clkout(net2590));
 b15cbf034ar1n64x5 hold593 (.clk(net2047),
    .clkout(net2591));
 b15cbf034ar1n64x5 hold594 (.clk(net218),
    .clkout(net2592));
 b15cbf034ar1n64x5 hold595 (.clk(net217),
    .clkout(net2593));
 b15cbf034ar1n64x5 hold596 (.clk(net231),
    .clkout(net2594));
 b15cbf034ar1n64x5 hold597 (.clk(net2061),
    .clkout(net2595));
 b15cbf034ar1n64x5 hold598 (.clk(net230),
    .clkout(net2596));
 b15cbf034ar1n64x5 hold599 (.clk(net2065),
    .clkout(net2597));
 b15cbf034ar1n64x5 hold600 (.clk(net220),
    .clkout(net2598));
 b15cbf034ar1n64x5 hold601 (.clk(net219),
    .clkout(net2599));
 b15cbf034ar1n64x5 hold602 (.clk(net214),
    .clkout(net2600));
 b15cbf034ar1n64x5 hold603 (.clk(net233),
    .clkout(net2601));
 b15cbf034ar1n64x5 hold604 (.clk(net232),
    .clkout(net2602));
 b15cbf034ar1n64x5 hold605 (.clk(net215),
    .clkout(net2603));
 b15cbf034ar1n64x5 hold606 (.clk(net234),
    .clkout(net2604));
 b15cbf034ar1n64x5 hold607 (.clk(net210),
    .clkout(net2605));
 b15cbf034ar1n64x5 hold608 (.clk(net235),
    .clkout(net2606));
 b15cbf034ar1n64x5 hold609 (.clk(net208),
    .clkout(net2607));
 b15cbf034ar1n64x5 hold610 (.clk(net209),
    .clkout(net2608));
 b15cbf034ar1n64x5 hold611 (.clk(net236),
    .clkout(net2609));
 b15cbf034ar1n64x5 hold612 (.clk(net229),
    .clkout(net2610));
 b15cbf034ar1n64x5 hold613 (.clk(net212),
    .clkout(net2611));
 b15cbf034ar1n64x5 hold614 (.clk(net228),
    .clkout(net2612));
 b15cbf034ar1n64x5 hold615 (.clk(net226),
    .clkout(net2613));
 b15cbf034ar1n64x5 hold616 (.clk(net213),
    .clkout(net2614));
 b15cbf034ar1n64x5 hold617 (.clk(net221),
    .clkout(net2615));
 b15cbf034ar1n64x5 hold618 (.clk(net260),
    .clkout(net2616));
 b15cbf034ar1n64x5 hold619 (.clk(net287),
    .clkout(net2617));
 b15cbf034ar1n64x5 hold620 (.clk(net223),
    .clkout(net2618));
 b15cbf034ar1n64x5 hold621 (.clk(net286),
    .clkout(net2619));
 b15cbf034ar1n64x5 hold622 (.clk(net284),
    .clkout(net2620));
 b15cbf034ar1n64x5 hold623 (.clk(net281),
    .clkout(net2621));
 b15cbf034ar1n64x5 hold624 (.clk(net279),
    .clkout(net2622));
 b15cbf034ar1n64x5 hold625 (.clk(net285),
    .clkout(net2623));
 b15cbf034ar1n64x5 hold626 (.clk(net256),
    .clkout(net2624));
 b15cbf034ar1n64x5 hold627 (.clk(net283),
    .clkout(net2625));
 b15cbf034ar1n64x5 hold628 (.clk(net282),
    .clkout(net2626));
 b15cbf034ar1n64x5 hold629 (.clk(gen_filter_13__u_filter_diff_ctr_q[0]),
    .clkout(net2627));
 b15cbf034ar1n64x5 hold630 (.clk(net251),
    .clkout(net2628));
 b15cbf034ar1n64x5 hold631 (.clk(net258),
    .clkout(net2629));
 b15cbf034ar1n64x5 hold632 (.clk(gen_filter_31__u_filter_diff_ctr_q[2]),
    .clkout(net2630));
 b15cbf034ar1n64x5 hold633 (.clk(gen_filter_31__u_filter_diff_ctr_d[3]),
    .clkout(net2631));
 b15cbf034ar1n64x5 hold634 (.clk(net257),
    .clkout(net2632));
 b15cbf034ar1n64x5 hold635 (.clk(gen_filter_19__u_filter_diff_ctr_q[3]),
    .clkout(net2633));
 b15cbf034ar1n64x5 hold636 (.clk(net156),
    .clkout(net2634));
 b15cbf034ar1n64x5 hold637 (.clk(net267),
    .clkout(net2635));
 b15cbf034ar1n64x5 hold638 (.clk(gen_alert_tx_0__u_prim_alert_sender_state_q[0]),
    .clkout(net2636));
 b15cbf034ar1n64x5 hold639 (.clk(gen_filter_12__u_filter_diff_ctr_q[2]),
    .clkout(net2637));
 b15cbf034ar1n64x5 hold640 (.clk(reg2hw_intr_state__q__5_),
    .clkout(net2638));
 b15cbf034ar1n64x5 hold641 (.clk(gen_filter_29__u_filter_diff_ctr_q[0]),
    .clkout(net2639));
 b15zdnd11an1n64x5 FILLER_0_8 ();
 b15zdnd11an1n64x5 FILLER_0_72 ();
 b15zdnd11an1n08x5 FILLER_0_136 ();
 b15zdnd11an1n64x5 FILLER_0_186 ();
 b15zdnd11an1n64x5 FILLER_0_250 ();
 b15zdnd11an1n64x5 FILLER_0_314 ();
 b15zdnd11an1n64x5 FILLER_0_378 ();
 b15zdnd11an1n08x5 FILLER_0_442 ();
 b15zdnd11an1n04x5 FILLER_0_450 ();
 b15zdnd11an1n16x5 FILLER_0_459 ();
 b15zdnd00an1n02x5 FILLER_0_475 ();
 b15zdnd00an1n01x5 FILLER_0_477 ();
 b15zdnd11an1n04x5 FILLER_0_482 ();
 b15zdnd11an1n32x5 FILLER_0_528 ();
 b15zdnd11an1n16x5 FILLER_0_560 ();
 b15zdnd11an1n04x5 FILLER_0_576 ();
 b15zdnd11an1n04x5 FILLER_0_584 ();
 b15zdnd11an1n04x5 FILLER_0_630 ();
 b15zdnd11an1n08x5 FILLER_0_638 ();
 b15zdnd11an1n04x5 FILLER_0_646 ();
 b15zdnd00an1n01x5 FILLER_0_650 ();
 b15zdnd11an1n04x5 FILLER_0_655 ();
 b15zdnd11an1n04x5 FILLER_0_663 ();
 b15zdnd00an1n02x5 FILLER_0_667 ();
 b15zdnd00an1n01x5 FILLER_0_669 ();
 b15zdnd11an1n04x5 FILLER_0_712 ();
 b15zdnd00an1n02x5 FILLER_0_716 ();
 b15zdnd11an1n04x5 FILLER_0_726 ();
 b15zdnd11an1n08x5 FILLER_0_734 ();
 b15zdnd11an1n04x5 FILLER_0_742 ();
 b15zdnd00an1n01x5 FILLER_0_746 ();
 b15zdnd11an1n04x5 FILLER_0_789 ();
 b15zdnd11an1n04x5 FILLER_0_835 ();
 b15zdnd11an1n04x5 FILLER_0_881 ();
 b15zdnd11an1n08x5 FILLER_0_889 ();
 b15zdnd11an1n04x5 FILLER_0_897 ();
 b15zdnd11an1n04x5 FILLER_0_905 ();
 b15zdnd11an1n04x5 FILLER_0_913 ();
 b15zdnd11an1n04x5 FILLER_0_959 ();
 b15zdnd11an1n04x5 FILLER_0_1005 ();
 b15zdnd11an1n32x5 FILLER_0_1051 ();
 b15zdnd11an1n08x5 FILLER_0_1083 ();
 b15zdnd00an1n02x5 FILLER_0_1091 ();
 b15zdnd11an1n08x5 FILLER_0_1135 ();
 b15zdnd11an1n04x5 FILLER_0_1143 ();
 b15zdnd00an1n01x5 FILLER_0_1147 ();
 b15zdnd11an1n04x5 FILLER_0_1190 ();
 b15zdnd11an1n08x5 FILLER_0_1214 ();
 b15zdnd11an1n04x5 FILLER_0_1222 ();
 b15zdnd11an1n32x5 FILLER_0_1230 ();
 b15zdnd00an1n02x5 FILLER_0_1262 ();
 b15zdnd11an1n64x5 FILLER_0_1268 ();
 b15zdnd00an1n02x5 FILLER_0_1332 ();
 b15zdnd00an1n01x5 FILLER_0_1334 ();
 b15zdnd11an1n32x5 FILLER_0_1339 ();
 b15zdnd11an1n04x5 FILLER_0_1371 ();
 b15zdnd00an1n01x5 FILLER_0_1375 ();
 b15zdnd11an1n04x5 FILLER_0_1380 ();
 b15zdnd11an1n08x5 FILLER_0_1388 ();
 b15zdnd00an1n02x5 FILLER_0_1396 ();
 b15zdnd00an1n01x5 FILLER_0_1398 ();
 b15zdnd11an1n04x5 FILLER_0_1403 ();
 b15zdnd11an1n16x5 FILLER_0_1411 ();
 b15zdnd11an1n08x5 FILLER_0_1427 ();
 b15zdnd00an1n01x5 FILLER_0_1435 ();
 b15zdnd11an1n04x5 FILLER_0_1444 ();
 b15zdnd00an1n02x5 FILLER_0_1448 ();
 b15zdnd11an1n04x5 FILLER_0_1454 ();
 b15zdnd11an1n16x5 FILLER_0_1500 ();
 b15zdnd11an1n08x5 FILLER_0_1516 ();
 b15zdnd11an1n16x5 FILLER_0_1531 ();
 b15zdnd11an1n04x5 FILLER_0_1547 ();
 b15zdnd00an1n02x5 FILLER_0_1551 ();
 b15zdnd00an1n01x5 FILLER_0_1553 ();
 b15zdnd11an1n04x5 FILLER_0_1558 ();
 b15zdnd11an1n32x5 FILLER_0_1566 ();
 b15zdnd11an1n08x5 FILLER_0_1598 ();
 b15zdnd11an1n04x5 FILLER_0_1606 ();
 b15zdnd00an1n02x5 FILLER_0_1610 ();
 b15zdnd00an1n01x5 FILLER_0_1612 ();
 b15zdnd11an1n64x5 FILLER_0_1617 ();
 b15zdnd11an1n64x5 FILLER_0_1681 ();
 b15zdnd11an1n64x5 FILLER_0_1745 ();
 b15zdnd11an1n64x5 FILLER_0_1809 ();
 b15zdnd11an1n64x5 FILLER_0_1873 ();
 b15zdnd11an1n64x5 FILLER_0_1937 ();
 b15zdnd11an1n64x5 FILLER_0_2001 ();
 b15zdnd11an1n64x5 FILLER_0_2065 ();
 b15zdnd11an1n16x5 FILLER_0_2129 ();
 b15zdnd11an1n08x5 FILLER_0_2145 ();
 b15zdnd00an1n01x5 FILLER_0_2153 ();
 b15zdnd11an1n64x5 FILLER_0_2162 ();
 b15zdnd11an1n32x5 FILLER_0_2226 ();
 b15zdnd11an1n16x5 FILLER_0_2258 ();
 b15zdnd00an1n02x5 FILLER_0_2274 ();
 b15zdnd11an1n64x5 FILLER_1_0 ();
 b15zdnd11an1n64x5 FILLER_1_64 ();
 b15zdnd11an1n16x5 FILLER_1_128 ();
 b15zdnd00an1n02x5 FILLER_1_144 ();
 b15zdnd00an1n01x5 FILLER_1_146 ();
 b15zdnd11an1n64x5 FILLER_1_161 ();
 b15zdnd11an1n64x5 FILLER_1_225 ();
 b15zdnd11an1n64x5 FILLER_1_289 ();
 b15zdnd11an1n64x5 FILLER_1_353 ();
 b15zdnd11an1n64x5 FILLER_1_417 ();
 b15zdnd11an1n64x5 FILLER_1_481 ();
 b15zdnd11an1n64x5 FILLER_1_545 ();
 b15zdnd11an1n16x5 FILLER_1_609 ();
 b15zdnd11an1n08x5 FILLER_1_625 ();
 b15zdnd00an1n02x5 FILLER_1_633 ();
 b15zdnd11an1n04x5 FILLER_1_677 ();
 b15zdnd11an1n16x5 FILLER_1_685 ();
 b15zdnd00an1n01x5 FILLER_1_701 ();
 b15zdnd11an1n04x5 FILLER_1_744 ();
 b15zdnd00an1n02x5 FILLER_1_748 ();
 b15zdnd11an1n16x5 FILLER_1_754 ();
 b15zdnd11an1n08x5 FILLER_1_770 ();
 b15zdnd11an1n04x5 FILLER_1_778 ();
 b15zdnd11an1n04x5 FILLER_1_824 ();
 b15zdnd11an1n08x5 FILLER_1_870 ();
 b15zdnd00an1n02x5 FILLER_1_878 ();
 b15zdnd00an1n01x5 FILLER_1_880 ();
 b15zdnd11an1n04x5 FILLER_1_923 ();
 b15zdnd00an1n02x5 FILLER_1_927 ();
 b15zdnd11an1n08x5 FILLER_1_971 ();
 b15zdnd00an1n02x5 FILLER_1_979 ();
 b15zdnd11an1n08x5 FILLER_1_987 ();
 b15zdnd00an1n02x5 FILLER_1_995 ();
 b15zdnd00an1n01x5 FILLER_1_997 ();
 b15zdnd11an1n04x5 FILLER_1_1002 ();
 b15zdnd11an1n32x5 FILLER_1_1048 ();
 b15zdnd11an1n08x5 FILLER_1_1080 ();
 b15zdnd11an1n04x5 FILLER_1_1088 ();
 b15zdnd00an1n02x5 FILLER_1_1092 ();
 b15zdnd00an1n01x5 FILLER_1_1094 ();
 b15zdnd11an1n16x5 FILLER_1_1099 ();
 b15zdnd11an1n08x5 FILLER_1_1115 ();
 b15zdnd11an1n16x5 FILLER_1_1127 ();
 b15zdnd11an1n08x5 FILLER_1_1143 ();
 b15zdnd11an1n04x5 FILLER_1_1151 ();
 b15zdnd00an1n01x5 FILLER_1_1155 ();
 b15zdnd11an1n04x5 FILLER_1_1160 ();
 b15zdnd11an1n08x5 FILLER_1_1168 ();
 b15zdnd00an1n02x5 FILLER_1_1176 ();
 b15zdnd00an1n01x5 FILLER_1_1178 ();
 b15zdnd11an1n64x5 FILLER_1_1221 ();
 b15zdnd11an1n64x5 FILLER_1_1285 ();
 b15zdnd11an1n32x5 FILLER_1_1349 ();
 b15zdnd11an1n16x5 FILLER_1_1381 ();
 b15zdnd11an1n04x5 FILLER_1_1397 ();
 b15zdnd00an1n01x5 FILLER_1_1401 ();
 b15zdnd11an1n64x5 FILLER_1_1444 ();
 b15zdnd11an1n64x5 FILLER_1_1508 ();
 b15zdnd11an1n08x5 FILLER_1_1572 ();
 b15zdnd11an1n64x5 FILLER_1_1584 ();
 b15zdnd11an1n64x5 FILLER_1_1648 ();
 b15zdnd11an1n64x5 FILLER_1_1712 ();
 b15zdnd11an1n64x5 FILLER_1_1776 ();
 b15zdnd11an1n64x5 FILLER_1_1840 ();
 b15zdnd11an1n64x5 FILLER_1_1904 ();
 b15zdnd11an1n64x5 FILLER_1_1968 ();
 b15zdnd11an1n64x5 FILLER_1_2032 ();
 b15zdnd11an1n64x5 FILLER_1_2096 ();
 b15zdnd11an1n64x5 FILLER_1_2160 ();
 b15zdnd11an1n32x5 FILLER_1_2224 ();
 b15zdnd11an1n16x5 FILLER_1_2256 ();
 b15zdnd11an1n08x5 FILLER_1_2272 ();
 b15zdnd11an1n04x5 FILLER_1_2280 ();
 b15zdnd11an1n64x5 FILLER_2_8 ();
 b15zdnd11an1n64x5 FILLER_2_72 ();
 b15zdnd11an1n64x5 FILLER_2_136 ();
 b15zdnd11an1n64x5 FILLER_2_200 ();
 b15zdnd11an1n64x5 FILLER_2_264 ();
 b15zdnd11an1n64x5 FILLER_2_328 ();
 b15zdnd11an1n64x5 FILLER_2_392 ();
 b15zdnd11an1n64x5 FILLER_2_456 ();
 b15zdnd11an1n64x5 FILLER_2_520 ();
 b15zdnd11an1n64x5 FILLER_2_584 ();
 b15zdnd11an1n16x5 FILLER_2_648 ();
 b15zdnd11an1n04x5 FILLER_2_668 ();
 b15zdnd00an1n02x5 FILLER_2_672 ();
 b15zdnd11an1n16x5 FILLER_2_678 ();
 b15zdnd11an1n04x5 FILLER_2_694 ();
 b15zdnd00an1n02x5 FILLER_2_698 ();
 b15zdnd00an1n01x5 FILLER_2_700 ();
 b15zdnd11an1n04x5 FILLER_2_705 ();
 b15zdnd00an1n02x5 FILLER_2_709 ();
 b15zdnd00an1n02x5 FILLER_2_715 ();
 b15zdnd00an1n01x5 FILLER_2_717 ();
 b15zdnd11an1n32x5 FILLER_2_726 ();
 b15zdnd11an1n16x5 FILLER_2_758 ();
 b15zdnd11an1n08x5 FILLER_2_774 ();
 b15zdnd00an1n02x5 FILLER_2_782 ();
 b15zdnd00an1n01x5 FILLER_2_784 ();
 b15zdnd11an1n04x5 FILLER_2_789 ();
 b15zdnd00an1n01x5 FILLER_2_793 ();
 b15zdnd11an1n16x5 FILLER_2_798 ();
 b15zdnd11an1n04x5 FILLER_2_814 ();
 b15zdnd11an1n04x5 FILLER_2_822 ();
 b15zdnd00an1n01x5 FILLER_2_826 ();
 b15zdnd11an1n32x5 FILLER_2_869 ();
 b15zdnd11an1n08x5 FILLER_2_901 ();
 b15zdnd11an1n04x5 FILLER_2_909 ();
 b15zdnd00an1n01x5 FILLER_2_913 ();
 b15zdnd11an1n04x5 FILLER_2_918 ();
 b15zdnd11an1n16x5 FILLER_2_926 ();
 b15zdnd11an1n04x5 FILLER_2_946 ();
 b15zdnd00an1n02x5 FILLER_2_950 ();
 b15zdnd00an1n01x5 FILLER_2_952 ();
 b15zdnd11an1n04x5 FILLER_2_957 ();
 b15zdnd11an1n04x5 FILLER_2_965 ();
 b15zdnd11an1n04x5 FILLER_2_973 ();
 b15zdnd11an1n04x5 FILLER_2_981 ();
 b15zdnd11an1n04x5 FILLER_2_989 ();
 b15zdnd11an1n04x5 FILLER_2_997 ();
 b15zdnd11an1n64x5 FILLER_2_1043 ();
 b15zdnd11an1n64x5 FILLER_2_1107 ();
 b15zdnd11an1n04x5 FILLER_2_1171 ();
 b15zdnd11an1n08x5 FILLER_2_1195 ();
 b15zdnd00an1n02x5 FILLER_2_1203 ();
 b15zdnd11an1n04x5 FILLER_2_1209 ();
 b15zdnd00an1n02x5 FILLER_2_1213 ();
 b15zdnd11an1n64x5 FILLER_2_1229 ();
 b15zdnd11an1n64x5 FILLER_2_1293 ();
 b15zdnd11an1n32x5 FILLER_2_1357 ();
 b15zdnd11an1n16x5 FILLER_2_1389 ();
 b15zdnd11an1n04x5 FILLER_2_1405 ();
 b15zdnd00an1n01x5 FILLER_2_1409 ();
 b15zdnd11an1n64x5 FILLER_2_1452 ();
 b15zdnd11an1n64x5 FILLER_2_1516 ();
 b15zdnd11an1n64x5 FILLER_2_1580 ();
 b15zdnd11an1n64x5 FILLER_2_1644 ();
 b15zdnd11an1n64x5 FILLER_2_1708 ();
 b15zdnd11an1n64x5 FILLER_2_1772 ();
 b15zdnd11an1n64x5 FILLER_2_1836 ();
 b15zdnd11an1n64x5 FILLER_2_1900 ();
 b15zdnd11an1n64x5 FILLER_2_1964 ();
 b15zdnd11an1n64x5 FILLER_2_2028 ();
 b15zdnd11an1n32x5 FILLER_2_2092 ();
 b15zdnd11an1n16x5 FILLER_2_2124 ();
 b15zdnd11an1n08x5 FILLER_2_2140 ();
 b15zdnd11an1n04x5 FILLER_2_2148 ();
 b15zdnd00an1n02x5 FILLER_2_2152 ();
 b15zdnd11an1n64x5 FILLER_2_2162 ();
 b15zdnd11an1n32x5 FILLER_2_2226 ();
 b15zdnd11an1n16x5 FILLER_2_2258 ();
 b15zdnd00an1n02x5 FILLER_2_2274 ();
 b15zdnd11an1n64x5 FILLER_3_0 ();
 b15zdnd11an1n64x5 FILLER_3_64 ();
 b15zdnd11an1n64x5 FILLER_3_128 ();
 b15zdnd11an1n64x5 FILLER_3_192 ();
 b15zdnd11an1n64x5 FILLER_3_256 ();
 b15zdnd11an1n64x5 FILLER_3_320 ();
 b15zdnd11an1n64x5 FILLER_3_384 ();
 b15zdnd11an1n64x5 FILLER_3_448 ();
 b15zdnd11an1n64x5 FILLER_3_512 ();
 b15zdnd11an1n64x5 FILLER_3_576 ();
 b15zdnd11an1n64x5 FILLER_3_640 ();
 b15zdnd11an1n64x5 FILLER_3_704 ();
 b15zdnd11an1n32x5 FILLER_3_768 ();
 b15zdnd11an1n16x5 FILLER_3_800 ();
 b15zdnd11an1n08x5 FILLER_3_816 ();
 b15zdnd00an1n02x5 FILLER_3_824 ();
 b15zdnd11an1n04x5 FILLER_3_830 ();
 b15zdnd11an1n04x5 FILLER_3_838 ();
 b15zdnd11an1n04x5 FILLER_3_846 ();
 b15zdnd11an1n04x5 FILLER_3_854 ();
 b15zdnd00an1n01x5 FILLER_3_858 ();
 b15zdnd11an1n64x5 FILLER_3_863 ();
 b15zdnd11an1n16x5 FILLER_3_927 ();
 b15zdnd11an1n08x5 FILLER_3_943 ();
 b15zdnd00an1n02x5 FILLER_3_951 ();
 b15zdnd11an1n08x5 FILLER_3_984 ();
 b15zdnd11an1n04x5 FILLER_3_996 ();
 b15zdnd11an1n64x5 FILLER_3_1042 ();
 b15zdnd11an1n64x5 FILLER_3_1106 ();
 b15zdnd11an1n08x5 FILLER_3_1170 ();
 b15zdnd00an1n02x5 FILLER_3_1178 ();
 b15zdnd00an1n01x5 FILLER_3_1180 ();
 b15zdnd11an1n64x5 FILLER_3_1201 ();
 b15zdnd11an1n64x5 FILLER_3_1265 ();
 b15zdnd11an1n64x5 FILLER_3_1329 ();
 b15zdnd11an1n64x5 FILLER_3_1393 ();
 b15zdnd11an1n64x5 FILLER_3_1457 ();
 b15zdnd11an1n64x5 FILLER_3_1521 ();
 b15zdnd11an1n64x5 FILLER_3_1585 ();
 b15zdnd11an1n64x5 FILLER_3_1649 ();
 b15zdnd11an1n64x5 FILLER_3_1713 ();
 b15zdnd11an1n64x5 FILLER_3_1777 ();
 b15zdnd11an1n64x5 FILLER_3_1841 ();
 b15zdnd11an1n64x5 FILLER_3_1905 ();
 b15zdnd11an1n64x5 FILLER_3_1969 ();
 b15zdnd11an1n64x5 FILLER_3_2033 ();
 b15zdnd11an1n64x5 FILLER_3_2097 ();
 b15zdnd11an1n64x5 FILLER_3_2161 ();
 b15zdnd11an1n32x5 FILLER_3_2225 ();
 b15zdnd11an1n16x5 FILLER_3_2257 ();
 b15zdnd11an1n08x5 FILLER_3_2273 ();
 b15zdnd00an1n02x5 FILLER_3_2281 ();
 b15zdnd00an1n01x5 FILLER_3_2283 ();
 b15zdnd11an1n64x5 FILLER_4_8 ();
 b15zdnd11an1n64x5 FILLER_4_72 ();
 b15zdnd11an1n64x5 FILLER_4_136 ();
 b15zdnd11an1n64x5 FILLER_4_200 ();
 b15zdnd11an1n64x5 FILLER_4_264 ();
 b15zdnd11an1n64x5 FILLER_4_328 ();
 b15zdnd11an1n64x5 FILLER_4_392 ();
 b15zdnd11an1n64x5 FILLER_4_456 ();
 b15zdnd11an1n64x5 FILLER_4_520 ();
 b15zdnd11an1n64x5 FILLER_4_584 ();
 b15zdnd11an1n64x5 FILLER_4_648 ();
 b15zdnd11an1n04x5 FILLER_4_712 ();
 b15zdnd00an1n02x5 FILLER_4_716 ();
 b15zdnd11an1n32x5 FILLER_4_726 ();
 b15zdnd11an1n04x5 FILLER_4_758 ();
 b15zdnd11an1n64x5 FILLER_4_804 ();
 b15zdnd11an1n32x5 FILLER_4_868 ();
 b15zdnd11an1n08x5 FILLER_4_900 ();
 b15zdnd00an1n01x5 FILLER_4_908 ();
 b15zdnd11an1n04x5 FILLER_4_951 ();
 b15zdnd00an1n02x5 FILLER_4_955 ();
 b15zdnd00an1n01x5 FILLER_4_957 ();
 b15zdnd11an1n04x5 FILLER_4_962 ();
 b15zdnd00an1n01x5 FILLER_4_966 ();
 b15zdnd11an1n04x5 FILLER_4_971 ();
 b15zdnd11an1n04x5 FILLER_4_979 ();
 b15zdnd11an1n64x5 FILLER_4_1025 ();
 b15zdnd11an1n64x5 FILLER_4_1089 ();
 b15zdnd11an1n64x5 FILLER_4_1153 ();
 b15zdnd11an1n64x5 FILLER_4_1217 ();
 b15zdnd11an1n64x5 FILLER_4_1281 ();
 b15zdnd11an1n64x5 FILLER_4_1345 ();
 b15zdnd11an1n64x5 FILLER_4_1409 ();
 b15zdnd11an1n64x5 FILLER_4_1481 ();
 b15zdnd11an1n64x5 FILLER_4_1545 ();
 b15zdnd11an1n64x5 FILLER_4_1609 ();
 b15zdnd11an1n64x5 FILLER_4_1673 ();
 b15zdnd11an1n64x5 FILLER_4_1737 ();
 b15zdnd11an1n64x5 FILLER_4_1801 ();
 b15zdnd11an1n64x5 FILLER_4_1865 ();
 b15zdnd11an1n64x5 FILLER_4_1929 ();
 b15zdnd11an1n64x5 FILLER_4_1993 ();
 b15zdnd11an1n64x5 FILLER_4_2057 ();
 b15zdnd11an1n32x5 FILLER_4_2121 ();
 b15zdnd00an1n01x5 FILLER_4_2153 ();
 b15zdnd11an1n64x5 FILLER_4_2162 ();
 b15zdnd11an1n32x5 FILLER_4_2226 ();
 b15zdnd11an1n16x5 FILLER_4_2258 ();
 b15zdnd00an1n02x5 FILLER_4_2274 ();
 b15zdnd11an1n64x5 FILLER_5_0 ();
 b15zdnd11an1n64x5 FILLER_5_64 ();
 b15zdnd11an1n64x5 FILLER_5_128 ();
 b15zdnd11an1n64x5 FILLER_5_192 ();
 b15zdnd11an1n64x5 FILLER_5_256 ();
 b15zdnd11an1n64x5 FILLER_5_320 ();
 b15zdnd11an1n64x5 FILLER_5_384 ();
 b15zdnd11an1n64x5 FILLER_5_448 ();
 b15zdnd11an1n64x5 FILLER_5_512 ();
 b15zdnd11an1n64x5 FILLER_5_576 ();
 b15zdnd11an1n64x5 FILLER_5_640 ();
 b15zdnd11an1n16x5 FILLER_5_704 ();
 b15zdnd11an1n08x5 FILLER_5_720 ();
 b15zdnd11an1n04x5 FILLER_5_728 ();
 b15zdnd00an1n02x5 FILLER_5_732 ();
 b15zdnd00an1n01x5 FILLER_5_734 ();
 b15zdnd11an1n16x5 FILLER_5_777 ();
 b15zdnd00an1n02x5 FILLER_5_793 ();
 b15zdnd00an1n01x5 FILLER_5_795 ();
 b15zdnd11an1n16x5 FILLER_5_838 ();
 b15zdnd11an1n04x5 FILLER_5_854 ();
 b15zdnd00an1n01x5 FILLER_5_858 ();
 b15zdnd11an1n32x5 FILLER_5_864 ();
 b15zdnd11an1n16x5 FILLER_5_896 ();
 b15zdnd11an1n08x5 FILLER_5_912 ();
 b15zdnd11an1n04x5 FILLER_5_920 ();
 b15zdnd11an1n08x5 FILLER_5_966 ();
 b15zdnd11an1n04x5 FILLER_5_974 ();
 b15zdnd11an1n04x5 FILLER_5_1020 ();
 b15zdnd00an1n02x5 FILLER_5_1024 ();
 b15zdnd11an1n64x5 FILLER_5_1068 ();
 b15zdnd11an1n64x5 FILLER_5_1132 ();
 b15zdnd11an1n64x5 FILLER_5_1196 ();
 b15zdnd11an1n64x5 FILLER_5_1260 ();
 b15zdnd11an1n64x5 FILLER_5_1324 ();
 b15zdnd11an1n64x5 FILLER_5_1388 ();
 b15zdnd11an1n64x5 FILLER_5_1452 ();
 b15zdnd11an1n64x5 FILLER_5_1516 ();
 b15zdnd11an1n64x5 FILLER_5_1580 ();
 b15zdnd11an1n64x5 FILLER_5_1644 ();
 b15zdnd11an1n64x5 FILLER_5_1708 ();
 b15zdnd11an1n64x5 FILLER_5_1772 ();
 b15zdnd11an1n64x5 FILLER_5_1836 ();
 b15zdnd11an1n64x5 FILLER_5_1900 ();
 b15zdnd11an1n64x5 FILLER_5_1964 ();
 b15zdnd11an1n64x5 FILLER_5_2028 ();
 b15zdnd11an1n64x5 FILLER_5_2092 ();
 b15zdnd11an1n64x5 FILLER_5_2156 ();
 b15zdnd11an1n64x5 FILLER_5_2220 ();
 b15zdnd11an1n64x5 FILLER_6_8 ();
 b15zdnd11an1n64x5 FILLER_6_72 ();
 b15zdnd11an1n64x5 FILLER_6_136 ();
 b15zdnd11an1n64x5 FILLER_6_200 ();
 b15zdnd11an1n64x5 FILLER_6_264 ();
 b15zdnd11an1n64x5 FILLER_6_328 ();
 b15zdnd11an1n64x5 FILLER_6_392 ();
 b15zdnd11an1n64x5 FILLER_6_456 ();
 b15zdnd11an1n64x5 FILLER_6_520 ();
 b15zdnd11an1n64x5 FILLER_6_584 ();
 b15zdnd11an1n64x5 FILLER_6_648 ();
 b15zdnd11an1n04x5 FILLER_6_712 ();
 b15zdnd00an1n02x5 FILLER_6_716 ();
 b15zdnd11an1n64x5 FILLER_6_726 ();
 b15zdnd11an1n32x5 FILLER_6_790 ();
 b15zdnd11an1n04x5 FILLER_6_822 ();
 b15zdnd11an1n08x5 FILLER_6_868 ();
 b15zdnd11an1n04x5 FILLER_6_876 ();
 b15zdnd00an1n02x5 FILLER_6_880 ();
 b15zdnd11an1n04x5 FILLER_6_924 ();
 b15zdnd11an1n08x5 FILLER_6_932 ();
 b15zdnd11an1n04x5 FILLER_6_940 ();
 b15zdnd00an1n02x5 FILLER_6_944 ();
 b15zdnd11an1n04x5 FILLER_6_954 ();
 b15zdnd11an1n32x5 FILLER_6_1003 ();
 b15zdnd11an1n16x5 FILLER_6_1035 ();
 b15zdnd00an1n01x5 FILLER_6_1051 ();
 b15zdnd11an1n64x5 FILLER_6_1094 ();
 b15zdnd11an1n64x5 FILLER_6_1158 ();
 b15zdnd11an1n64x5 FILLER_6_1222 ();
 b15zdnd11an1n64x5 FILLER_6_1286 ();
 b15zdnd11an1n64x5 FILLER_6_1350 ();
 b15zdnd11an1n64x5 FILLER_6_1414 ();
 b15zdnd11an1n64x5 FILLER_6_1478 ();
 b15zdnd11an1n64x5 FILLER_6_1542 ();
 b15zdnd11an1n64x5 FILLER_6_1606 ();
 b15zdnd11an1n64x5 FILLER_6_1670 ();
 b15zdnd11an1n64x5 FILLER_6_1734 ();
 b15zdnd11an1n64x5 FILLER_6_1798 ();
 b15zdnd11an1n64x5 FILLER_6_1862 ();
 b15zdnd11an1n64x5 FILLER_6_1926 ();
 b15zdnd11an1n64x5 FILLER_6_1990 ();
 b15zdnd11an1n64x5 FILLER_6_2054 ();
 b15zdnd11an1n32x5 FILLER_6_2118 ();
 b15zdnd11an1n04x5 FILLER_6_2150 ();
 b15zdnd11an1n64x5 FILLER_6_2162 ();
 b15zdnd11an1n32x5 FILLER_6_2226 ();
 b15zdnd11an1n16x5 FILLER_6_2258 ();
 b15zdnd00an1n02x5 FILLER_6_2274 ();
 b15zdnd11an1n64x5 FILLER_7_0 ();
 b15zdnd11an1n32x5 FILLER_7_64 ();
 b15zdnd11an1n08x5 FILLER_7_96 ();
 b15zdnd11an1n04x5 FILLER_7_104 ();
 b15zdnd00an1n01x5 FILLER_7_108 ();
 b15zdnd11an1n16x5 FILLER_7_112 ();
 b15zdnd11an1n64x5 FILLER_7_131 ();
 b15zdnd11an1n64x5 FILLER_7_195 ();
 b15zdnd11an1n64x5 FILLER_7_259 ();
 b15zdnd11an1n04x5 FILLER_7_323 ();
 b15zdnd11an1n64x5 FILLER_7_330 ();
 b15zdnd11an1n16x5 FILLER_7_394 ();
 b15zdnd11an1n08x5 FILLER_7_410 ();
 b15zdnd11an1n04x5 FILLER_7_418 ();
 b15zdnd00an1n02x5 FILLER_7_422 ();
 b15zdnd11an1n16x5 FILLER_7_428 ();
 b15zdnd11an1n04x5 FILLER_7_444 ();
 b15zdnd00an1n01x5 FILLER_7_448 ();
 b15zdnd11an1n64x5 FILLER_7_455 ();
 b15zdnd11an1n64x5 FILLER_7_519 ();
 b15zdnd11an1n64x5 FILLER_7_583 ();
 b15zdnd11an1n32x5 FILLER_7_647 ();
 b15zdnd11an1n16x5 FILLER_7_679 ();
 b15zdnd00an1n02x5 FILLER_7_695 ();
 b15zdnd11an1n64x5 FILLER_7_704 ();
 b15zdnd11an1n32x5 FILLER_7_768 ();
 b15zdnd11an1n08x5 FILLER_7_800 ();
 b15zdnd11an1n04x5 FILLER_7_808 ();
 b15zdnd00an1n02x5 FILLER_7_812 ();
 b15zdnd00an1n01x5 FILLER_7_814 ();
 b15zdnd11an1n04x5 FILLER_7_835 ();
 b15zdnd11an1n04x5 FILLER_7_881 ();
 b15zdnd11an1n04x5 FILLER_7_916 ();
 b15zdnd11an1n04x5 FILLER_7_927 ();
 b15zdnd00an1n02x5 FILLER_7_931 ();
 b15zdnd00an1n01x5 FILLER_7_933 ();
 b15zdnd11an1n04x5 FILLER_7_943 ();
 b15zdnd00an1n02x5 FILLER_7_947 ();
 b15zdnd11an1n08x5 FILLER_7_991 ();
 b15zdnd11an1n04x5 FILLER_7_999 ();
 b15zdnd11an1n04x5 FILLER_7_1045 ();
 b15zdnd00an1n01x5 FILLER_7_1049 ();
 b15zdnd11an1n64x5 FILLER_7_1092 ();
 b15zdnd11an1n32x5 FILLER_7_1156 ();
 b15zdnd11an1n08x5 FILLER_7_1188 ();
 b15zdnd00an1n01x5 FILLER_7_1196 ();
 b15zdnd11an1n64x5 FILLER_7_1239 ();
 b15zdnd11an1n64x5 FILLER_7_1303 ();
 b15zdnd11an1n64x5 FILLER_7_1367 ();
 b15zdnd11an1n64x5 FILLER_7_1431 ();
 b15zdnd11an1n64x5 FILLER_7_1495 ();
 b15zdnd11an1n64x5 FILLER_7_1559 ();
 b15zdnd11an1n64x5 FILLER_7_1623 ();
 b15zdnd11an1n64x5 FILLER_7_1687 ();
 b15zdnd11an1n64x5 FILLER_7_1751 ();
 b15zdnd11an1n64x5 FILLER_7_1815 ();
 b15zdnd11an1n32x5 FILLER_7_1879 ();
 b15zdnd11an1n08x5 FILLER_7_1911 ();
 b15zdnd11an1n64x5 FILLER_7_1922 ();
 b15zdnd11an1n64x5 FILLER_7_1986 ();
 b15zdnd11an1n64x5 FILLER_7_2050 ();
 b15zdnd11an1n64x5 FILLER_7_2114 ();
 b15zdnd11an1n64x5 FILLER_7_2178 ();
 b15zdnd11an1n32x5 FILLER_7_2242 ();
 b15zdnd11an1n08x5 FILLER_7_2274 ();
 b15zdnd00an1n02x5 FILLER_7_2282 ();
 b15zdnd11an1n64x5 FILLER_8_8 ();
 b15zdnd11an1n32x5 FILLER_8_72 ();
 b15zdnd11an1n04x5 FILLER_8_104 ();
 b15zdnd00an1n02x5 FILLER_8_108 ();
 b15zdnd11an1n08x5 FILLER_8_113 ();
 b15zdnd11an1n04x5 FILLER_8_121 ();
 b15zdnd00an1n01x5 FILLER_8_125 ();
 b15zdnd11an1n64x5 FILLER_8_129 ();
 b15zdnd11an1n64x5 FILLER_8_193 ();
 b15zdnd11an1n64x5 FILLER_8_257 ();
 b15zdnd11an1n08x5 FILLER_8_321 ();
 b15zdnd00an1n02x5 FILLER_8_329 ();
 b15zdnd11an1n64x5 FILLER_8_334 ();
 b15zdnd00an1n02x5 FILLER_8_398 ();
 b15zdnd11an1n04x5 FILLER_8_404 ();
 b15zdnd00an1n02x5 FILLER_8_408 ();
 b15zdnd11an1n04x5 FILLER_8_413 ();
 b15zdnd11an1n08x5 FILLER_8_432 ();
 b15zdnd00an1n02x5 FILLER_8_440 ();
 b15zdnd00an1n01x5 FILLER_8_442 ();
 b15zdnd11an1n64x5 FILLER_8_474 ();
 b15zdnd11an1n16x5 FILLER_8_538 ();
 b15zdnd00an1n01x5 FILLER_8_554 ();
 b15zdnd11an1n16x5 FILLER_8_586 ();
 b15zdnd11an1n08x5 FILLER_8_602 ();
 b15zdnd11an1n04x5 FILLER_8_610 ();
 b15zdnd00an1n02x5 FILLER_8_614 ();
 b15zdnd11an1n16x5 FILLER_8_641 ();
 b15zdnd11an1n04x5 FILLER_8_657 ();
 b15zdnd00an1n02x5 FILLER_8_661 ();
 b15zdnd11an1n16x5 FILLER_8_683 ();
 b15zdnd00an1n01x5 FILLER_8_699 ();
 b15zdnd11an1n04x5 FILLER_8_714 ();
 b15zdnd11an1n16x5 FILLER_8_726 ();
 b15zdnd11an1n08x5 FILLER_8_742 ();
 b15zdnd11an1n04x5 FILLER_8_750 ();
 b15zdnd00an1n02x5 FILLER_8_754 ();
 b15zdnd00an1n01x5 FILLER_8_756 ();
 b15zdnd11an1n08x5 FILLER_8_799 ();
 b15zdnd11an1n04x5 FILLER_8_807 ();
 b15zdnd00an1n01x5 FILLER_8_811 ();
 b15zdnd11an1n04x5 FILLER_8_836 ();
 b15zdnd11an1n08x5 FILLER_8_845 ();
 b15zdnd00an1n02x5 FILLER_8_853 ();
 b15zdnd00an1n01x5 FILLER_8_855 ();
 b15zdnd11an1n04x5 FILLER_8_901 ();
 b15zdnd11an1n04x5 FILLER_8_947 ();
 b15zdnd00an1n02x5 FILLER_8_951 ();
 b15zdnd11an1n04x5 FILLER_8_957 ();
 b15zdnd11an1n04x5 FILLER_8_1006 ();
 b15zdnd11an1n04x5 FILLER_8_1017 ();
 b15zdnd11an1n04x5 FILLER_8_1028 ();
 b15zdnd11an1n08x5 FILLER_8_1040 ();
 b15zdnd11an1n04x5 FILLER_8_1048 ();
 b15zdnd11an1n16x5 FILLER_8_1060 ();
 b15zdnd11an1n08x5 FILLER_8_1076 ();
 b15zdnd11an1n04x5 FILLER_8_1084 ();
 b15zdnd11an1n64x5 FILLER_8_1133 ();
 b15zdnd11an1n16x5 FILLER_8_1197 ();
 b15zdnd11an1n08x5 FILLER_8_1213 ();
 b15zdnd11an1n04x5 FILLER_8_1221 ();
 b15zdnd11an1n16x5 FILLER_8_1270 ();
 b15zdnd11an1n08x5 FILLER_8_1286 ();
 b15zdnd11an1n04x5 FILLER_8_1294 ();
 b15zdnd00an1n02x5 FILLER_8_1298 ();
 b15zdnd11an1n16x5 FILLER_8_1314 ();
 b15zdnd11an1n04x5 FILLER_8_1330 ();
 b15zdnd00an1n01x5 FILLER_8_1334 ();
 b15zdnd11an1n64x5 FILLER_8_1355 ();
 b15zdnd11an1n64x5 FILLER_8_1419 ();
 b15zdnd11an1n64x5 FILLER_8_1483 ();
 b15zdnd11an1n64x5 FILLER_8_1547 ();
 b15zdnd11an1n64x5 FILLER_8_1611 ();
 b15zdnd11an1n64x5 FILLER_8_1675 ();
 b15zdnd11an1n64x5 FILLER_8_1739 ();
 b15zdnd11an1n64x5 FILLER_8_1803 ();
 b15zdnd11an1n32x5 FILLER_8_1867 ();
 b15zdnd11an1n08x5 FILLER_8_1899 ();
 b15zdnd11an1n04x5 FILLER_8_1907 ();
 b15zdnd00an1n02x5 FILLER_8_1911 ();
 b15zdnd11an1n04x5 FILLER_8_1916 ();
 b15zdnd11an1n64x5 FILLER_8_1927 ();
 b15zdnd11an1n64x5 FILLER_8_1991 ();
 b15zdnd11an1n64x5 FILLER_8_2055 ();
 b15zdnd11an1n32x5 FILLER_8_2119 ();
 b15zdnd00an1n02x5 FILLER_8_2151 ();
 b15zdnd00an1n01x5 FILLER_8_2153 ();
 b15zdnd11an1n64x5 FILLER_8_2162 ();
 b15zdnd11an1n32x5 FILLER_8_2226 ();
 b15zdnd11an1n16x5 FILLER_8_2258 ();
 b15zdnd00an1n02x5 FILLER_8_2274 ();
 b15zdnd11an1n64x5 FILLER_9_0 ();
 b15zdnd11an1n64x5 FILLER_9_64 ();
 b15zdnd11an1n64x5 FILLER_9_128 ();
 b15zdnd11an1n64x5 FILLER_9_192 ();
 b15zdnd11an1n64x5 FILLER_9_256 ();
 b15zdnd11an1n64x5 FILLER_9_320 ();
 b15zdnd11an1n16x5 FILLER_9_384 ();
 b15zdnd00an1n02x5 FILLER_9_400 ();
 b15zdnd11an1n04x5 FILLER_9_407 ();
 b15zdnd11an1n04x5 FILLER_9_424 ();
 b15zdnd11an1n04x5 FILLER_9_437 ();
 b15zdnd11an1n08x5 FILLER_9_448 ();
 b15zdnd00an1n02x5 FILLER_9_456 ();
 b15zdnd00an1n01x5 FILLER_9_458 ();
 b15zdnd11an1n04x5 FILLER_9_462 ();
 b15zdnd11an1n64x5 FILLER_9_475 ();
 b15zdnd11an1n64x5 FILLER_9_539 ();
 b15zdnd11an1n16x5 FILLER_9_603 ();
 b15zdnd00an1n02x5 FILLER_9_619 ();
 b15zdnd00an1n01x5 FILLER_9_621 ();
 b15zdnd11an1n04x5 FILLER_9_628 ();
 b15zdnd00an1n02x5 FILLER_9_632 ();
 b15zdnd11an1n04x5 FILLER_9_679 ();
 b15zdnd11an1n64x5 FILLER_9_690 ();
 b15zdnd11an1n16x5 FILLER_9_754 ();
 b15zdnd11an1n08x5 FILLER_9_770 ();
 b15zdnd11an1n08x5 FILLER_9_784 ();
 b15zdnd11an1n04x5 FILLER_9_792 ();
 b15zdnd00an1n01x5 FILLER_9_796 ();
 b15zdnd11an1n04x5 FILLER_9_839 ();
 b15zdnd00an1n02x5 FILLER_9_843 ();
 b15zdnd11an1n08x5 FILLER_9_887 ();
 b15zdnd00an1n02x5 FILLER_9_895 ();
 b15zdnd11an1n08x5 FILLER_9_904 ();
 b15zdnd00an1n01x5 FILLER_9_912 ();
 b15zdnd11an1n04x5 FILLER_9_955 ();
 b15zdnd11an1n04x5 FILLER_9_1001 ();
 b15zdnd11an1n08x5 FILLER_9_1047 ();
 b15zdnd00an1n02x5 FILLER_9_1055 ();
 b15zdnd00an1n01x5 FILLER_9_1057 ();
 b15zdnd11an1n64x5 FILLER_9_1100 ();
 b15zdnd11an1n16x5 FILLER_9_1164 ();
 b15zdnd11an1n08x5 FILLER_9_1180 ();
 b15zdnd00an1n01x5 FILLER_9_1188 ();
 b15zdnd11an1n16x5 FILLER_9_1206 ();
 b15zdnd11an1n04x5 FILLER_9_1222 ();
 b15zdnd00an1n02x5 FILLER_9_1226 ();
 b15zdnd00an1n01x5 FILLER_9_1228 ();
 b15zdnd11an1n04x5 FILLER_9_1236 ();
 b15zdnd11an1n04x5 FILLER_9_1285 ();
 b15zdnd00an1n02x5 FILLER_9_1289 ();
 b15zdnd00an1n01x5 FILLER_9_1291 ();
 b15zdnd11an1n04x5 FILLER_9_1295 ();
 b15zdnd11an1n32x5 FILLER_9_1326 ();
 b15zdnd11an1n16x5 FILLER_9_1358 ();
 b15zdnd11an1n08x5 FILLER_9_1374 ();
 b15zdnd11an1n04x5 FILLER_9_1382 ();
 b15zdnd00an1n01x5 FILLER_9_1386 ();
 b15zdnd11an1n64x5 FILLER_9_1413 ();
 b15zdnd11an1n64x5 FILLER_9_1477 ();
 b15zdnd11an1n64x5 FILLER_9_1541 ();
 b15zdnd11an1n64x5 FILLER_9_1605 ();
 b15zdnd11an1n64x5 FILLER_9_1669 ();
 b15zdnd11an1n64x5 FILLER_9_1733 ();
 b15zdnd11an1n32x5 FILLER_9_1797 ();
 b15zdnd11an1n16x5 FILLER_9_1829 ();
 b15zdnd11an1n08x5 FILLER_9_1845 ();
 b15zdnd11an1n16x5 FILLER_9_1884 ();
 b15zdnd11an1n08x5 FILLER_9_1900 ();
 b15zdnd00an1n02x5 FILLER_9_1908 ();
 b15zdnd00an1n01x5 FILLER_9_1910 ();
 b15zdnd11an1n16x5 FILLER_9_1925 ();
 b15zdnd00an1n01x5 FILLER_9_1941 ();
 b15zdnd11an1n64x5 FILLER_9_1945 ();
 b15zdnd11an1n64x5 FILLER_9_2009 ();
 b15zdnd11an1n64x5 FILLER_9_2073 ();
 b15zdnd11an1n64x5 FILLER_9_2137 ();
 b15zdnd11an1n64x5 FILLER_9_2201 ();
 b15zdnd11an1n16x5 FILLER_9_2265 ();
 b15zdnd00an1n02x5 FILLER_9_2281 ();
 b15zdnd00an1n01x5 FILLER_9_2283 ();
 b15zdnd11an1n64x5 FILLER_10_8 ();
 b15zdnd11an1n64x5 FILLER_10_72 ();
 b15zdnd11an1n64x5 FILLER_10_136 ();
 b15zdnd11an1n64x5 FILLER_10_200 ();
 b15zdnd11an1n64x5 FILLER_10_264 ();
 b15zdnd11an1n64x5 FILLER_10_328 ();
 b15zdnd11an1n08x5 FILLER_10_392 ();
 b15zdnd11an1n04x5 FILLER_10_400 ();
 b15zdnd00an1n02x5 FILLER_10_404 ();
 b15zdnd00an1n01x5 FILLER_10_406 ();
 b15zdnd11an1n04x5 FILLER_10_412 ();
 b15zdnd11an1n04x5 FILLER_10_458 ();
 b15zdnd11an1n64x5 FILLER_10_468 ();
 b15zdnd11an1n32x5 FILLER_10_532 ();
 b15zdnd11an1n08x5 FILLER_10_564 ();
 b15zdnd11an1n04x5 FILLER_10_587 ();
 b15zdnd11an1n32x5 FILLER_10_643 ();
 b15zdnd11an1n08x5 FILLER_10_675 ();
 b15zdnd00an1n02x5 FILLER_10_683 ();
 b15zdnd00an1n01x5 FILLER_10_685 ();
 b15zdnd11an1n16x5 FILLER_10_698 ();
 b15zdnd11an1n04x5 FILLER_10_714 ();
 b15zdnd11an1n32x5 FILLER_10_726 ();
 b15zdnd11an1n08x5 FILLER_10_758 ();
 b15zdnd11an1n04x5 FILLER_10_769 ();
 b15zdnd11an1n16x5 FILLER_10_776 ();
 b15zdnd11an1n08x5 FILLER_10_792 ();
 b15zdnd11an1n04x5 FILLER_10_800 ();
 b15zdnd00an1n02x5 FILLER_10_804 ();
 b15zdnd00an1n01x5 FILLER_10_806 ();
 b15zdnd11an1n32x5 FILLER_10_812 ();
 b15zdnd11an1n04x5 FILLER_10_844 ();
 b15zdnd00an1n02x5 FILLER_10_848 ();
 b15zdnd11an1n04x5 FILLER_10_902 ();
 b15zdnd00an1n02x5 FILLER_10_906 ();
 b15zdnd11an1n04x5 FILLER_10_939 ();
 b15zdnd11an1n08x5 FILLER_10_988 ();
 b15zdnd11an1n04x5 FILLER_10_996 ();
 b15zdnd11an1n16x5 FILLER_10_1042 ();
 b15zdnd00an1n02x5 FILLER_10_1058 ();
 b15zdnd00an1n01x5 FILLER_10_1060 ();
 b15zdnd11an1n08x5 FILLER_10_1068 ();
 b15zdnd00an1n02x5 FILLER_10_1076 ();
 b15zdnd11an1n64x5 FILLER_10_1120 ();
 b15zdnd11an1n16x5 FILLER_10_1184 ();
 b15zdnd00an1n02x5 FILLER_10_1200 ();
 b15zdnd00an1n01x5 FILLER_10_1202 ();
 b15zdnd11an1n04x5 FILLER_10_1206 ();
 b15zdnd11an1n16x5 FILLER_10_1213 ();
 b15zdnd11an1n04x5 FILLER_10_1229 ();
 b15zdnd11an1n04x5 FILLER_10_1275 ();
 b15zdnd11an1n32x5 FILLER_10_1299 ();
 b15zdnd11an1n16x5 FILLER_10_1331 ();
 b15zdnd11an1n08x5 FILLER_10_1347 ();
 b15zdnd11an1n04x5 FILLER_10_1355 ();
 b15zdnd00an1n02x5 FILLER_10_1359 ();
 b15zdnd11an1n04x5 FILLER_10_1364 ();
 b15zdnd11an1n04x5 FILLER_10_1371 ();
 b15zdnd11an1n64x5 FILLER_10_1392 ();
 b15zdnd11an1n64x5 FILLER_10_1456 ();
 b15zdnd11an1n32x5 FILLER_10_1520 ();
 b15zdnd11an1n16x5 FILLER_10_1552 ();
 b15zdnd11an1n08x5 FILLER_10_1568 ();
 b15zdnd00an1n02x5 FILLER_10_1576 ();
 b15zdnd00an1n01x5 FILLER_10_1578 ();
 b15zdnd11an1n64x5 FILLER_10_1582 ();
 b15zdnd00an1n01x5 FILLER_10_1646 ();
 b15zdnd11an1n64x5 FILLER_10_1651 ();
 b15zdnd11an1n64x5 FILLER_10_1715 ();
 b15zdnd11an1n64x5 FILLER_10_1779 ();
 b15zdnd11an1n32x5 FILLER_10_1843 ();
 b15zdnd11an1n16x5 FILLER_10_1875 ();
 b15zdnd11an1n08x5 FILLER_10_1891 ();
 b15zdnd00an1n01x5 FILLER_10_1899 ();
 b15zdnd11an1n04x5 FILLER_10_1910 ();
 b15zdnd00an1n02x5 FILLER_10_1914 ();
 b15zdnd11an1n08x5 FILLER_10_1928 ();
 b15zdnd00an1n02x5 FILLER_10_1936 ();
 b15zdnd11an1n64x5 FILLER_10_1943 ();
 b15zdnd11an1n64x5 FILLER_10_2007 ();
 b15zdnd11an1n64x5 FILLER_10_2071 ();
 b15zdnd11an1n16x5 FILLER_10_2135 ();
 b15zdnd00an1n02x5 FILLER_10_2151 ();
 b15zdnd00an1n01x5 FILLER_10_2153 ();
 b15zdnd11an1n64x5 FILLER_10_2162 ();
 b15zdnd11an1n32x5 FILLER_10_2226 ();
 b15zdnd11an1n16x5 FILLER_10_2258 ();
 b15zdnd00an1n02x5 FILLER_10_2274 ();
 b15zdnd11an1n64x5 FILLER_11_0 ();
 b15zdnd11an1n64x5 FILLER_11_64 ();
 b15zdnd11an1n64x5 FILLER_11_128 ();
 b15zdnd11an1n64x5 FILLER_11_192 ();
 b15zdnd11an1n64x5 FILLER_11_256 ();
 b15zdnd11an1n64x5 FILLER_11_320 ();
 b15zdnd11an1n32x5 FILLER_11_384 ();
 b15zdnd00an1n01x5 FILLER_11_416 ();
 b15zdnd11an1n64x5 FILLER_11_423 ();
 b15zdnd11an1n64x5 FILLER_11_487 ();
 b15zdnd11an1n32x5 FILLER_11_551 ();
 b15zdnd11an1n16x5 FILLER_11_583 ();
 b15zdnd11an1n08x5 FILLER_11_599 ();
 b15zdnd11an1n04x5 FILLER_11_607 ();
 b15zdnd11an1n04x5 FILLER_11_614 ();
 b15zdnd11an1n04x5 FILLER_11_621 ();
 b15zdnd11an1n64x5 FILLER_11_628 ();
 b15zdnd11an1n08x5 FILLER_11_692 ();
 b15zdnd11an1n04x5 FILLER_11_700 ();
 b15zdnd00an1n02x5 FILLER_11_704 ();
 b15zdnd00an1n01x5 FILLER_11_706 ();
 b15zdnd11an1n32x5 FILLER_11_714 ();
 b15zdnd11an1n32x5 FILLER_11_798 ();
 b15zdnd11an1n16x5 FILLER_11_830 ();
 b15zdnd11an1n04x5 FILLER_11_877 ();
 b15zdnd11an1n08x5 FILLER_11_888 ();
 b15zdnd00an1n02x5 FILLER_11_896 ();
 b15zdnd11an1n04x5 FILLER_11_940 ();
 b15zdnd11an1n04x5 FILLER_11_951 ();
 b15zdnd00an1n01x5 FILLER_11_955 ();
 b15zdnd11an1n32x5 FILLER_11_1008 ();
 b15zdnd11an1n16x5 FILLER_11_1040 ();
 b15zdnd00an1n01x5 FILLER_11_1056 ();
 b15zdnd11an1n04x5 FILLER_11_1099 ();
 b15zdnd11an1n64x5 FILLER_11_1106 ();
 b15zdnd11an1n08x5 FILLER_11_1170 ();
 b15zdnd11an1n04x5 FILLER_11_1178 ();
 b15zdnd00an1n02x5 FILLER_11_1182 ();
 b15zdnd00an1n01x5 FILLER_11_1184 ();
 b15zdnd11an1n04x5 FILLER_11_1237 ();
 b15zdnd00an1n01x5 FILLER_11_1241 ();
 b15zdnd11an1n08x5 FILLER_11_1273 ();
 b15zdnd00an1n02x5 FILLER_11_1281 ();
 b15zdnd00an1n01x5 FILLER_11_1283 ();
 b15zdnd11an1n04x5 FILLER_11_1304 ();
 b15zdnd11an1n16x5 FILLER_11_1314 ();
 b15zdnd11an1n08x5 FILLER_11_1330 ();
 b15zdnd11an1n04x5 FILLER_11_1338 ();
 b15zdnd00an1n01x5 FILLER_11_1342 ();
 b15zdnd11an1n64x5 FILLER_11_1395 ();
 b15zdnd11an1n64x5 FILLER_11_1459 ();
 b15zdnd11an1n16x5 FILLER_11_1523 ();
 b15zdnd11an1n08x5 FILLER_11_1539 ();
 b15zdnd11an1n04x5 FILLER_11_1547 ();
 b15zdnd00an1n02x5 FILLER_11_1551 ();
 b15zdnd11an1n64x5 FILLER_11_1605 ();
 b15zdnd11an1n64x5 FILLER_11_1669 ();
 b15zdnd11an1n64x5 FILLER_11_1733 ();
 b15zdnd11an1n64x5 FILLER_11_1797 ();
 b15zdnd11an1n32x5 FILLER_11_1861 ();
 b15zdnd11an1n16x5 FILLER_11_1893 ();
 b15zdnd11an1n04x5 FILLER_11_1909 ();
 b15zdnd00an1n02x5 FILLER_11_1913 ();
 b15zdnd11an1n16x5 FILLER_11_1957 ();
 b15zdnd11an1n04x5 FILLER_11_1973 ();
 b15zdnd00an1n01x5 FILLER_11_1977 ();
 b15zdnd11an1n64x5 FILLER_11_1981 ();
 b15zdnd11an1n64x5 FILLER_11_2045 ();
 b15zdnd11an1n64x5 FILLER_11_2109 ();
 b15zdnd11an1n64x5 FILLER_11_2173 ();
 b15zdnd11an1n32x5 FILLER_11_2237 ();
 b15zdnd11an1n08x5 FILLER_11_2269 ();
 b15zdnd11an1n04x5 FILLER_11_2277 ();
 b15zdnd00an1n02x5 FILLER_11_2281 ();
 b15zdnd00an1n01x5 FILLER_11_2283 ();
 b15zdnd11an1n64x5 FILLER_12_8 ();
 b15zdnd11an1n64x5 FILLER_12_72 ();
 b15zdnd11an1n64x5 FILLER_12_136 ();
 b15zdnd11an1n64x5 FILLER_12_200 ();
 b15zdnd11an1n64x5 FILLER_12_264 ();
 b15zdnd11an1n64x5 FILLER_12_328 ();
 b15zdnd11an1n64x5 FILLER_12_392 ();
 b15zdnd11an1n64x5 FILLER_12_456 ();
 b15zdnd11an1n64x5 FILLER_12_520 ();
 b15zdnd11an1n16x5 FILLER_12_584 ();
 b15zdnd11an1n08x5 FILLER_12_600 ();
 b15zdnd00an1n02x5 FILLER_12_608 ();
 b15zdnd11an1n04x5 FILLER_12_613 ();
 b15zdnd11an1n64x5 FILLER_12_623 ();
 b15zdnd11an1n16x5 FILLER_12_687 ();
 b15zdnd11an1n08x5 FILLER_12_703 ();
 b15zdnd11an1n04x5 FILLER_12_711 ();
 b15zdnd00an1n02x5 FILLER_12_715 ();
 b15zdnd00an1n01x5 FILLER_12_717 ();
 b15zdnd00an1n02x5 FILLER_12_726 ();
 b15zdnd11an1n04x5 FILLER_12_770 ();
 b15zdnd11an1n08x5 FILLER_12_777 ();
 b15zdnd11an1n32x5 FILLER_12_792 ();
 b15zdnd11an1n16x5 FILLER_12_824 ();
 b15zdnd11an1n04x5 FILLER_12_840 ();
 b15zdnd00an1n02x5 FILLER_12_844 ();
 b15zdnd00an1n01x5 FILLER_12_846 ();
 b15zdnd11an1n32x5 FILLER_12_899 ();
 b15zdnd11an1n04x5 FILLER_12_931 ();
 b15zdnd00an1n02x5 FILLER_12_935 ();
 b15zdnd11an1n04x5 FILLER_12_979 ();
 b15zdnd11an1n04x5 FILLER_12_990 ();
 b15zdnd11an1n04x5 FILLER_12_1001 ();
 b15zdnd11an1n32x5 FILLER_12_1008 ();
 b15zdnd11an1n08x5 FILLER_12_1040 ();
 b15zdnd11an1n04x5 FILLER_12_1048 ();
 b15zdnd11an1n64x5 FILLER_12_1104 ();
 b15zdnd11an1n32x5 FILLER_12_1168 ();
 b15zdnd11an1n08x5 FILLER_12_1200 ();
 b15zdnd00an1n02x5 FILLER_12_1208 ();
 b15zdnd11an1n32x5 FILLER_12_1213 ();
 b15zdnd11an1n16x5 FILLER_12_1245 ();
 b15zdnd11an1n08x5 FILLER_12_1261 ();
 b15zdnd11an1n04x5 FILLER_12_1269 ();
 b15zdnd11an1n64x5 FILLER_12_1284 ();
 b15zdnd11an1n04x5 FILLER_12_1348 ();
 b15zdnd00an1n02x5 FILLER_12_1352 ();
 b15zdnd00an1n01x5 FILLER_12_1354 ();
 b15zdnd11an1n04x5 FILLER_12_1364 ();
 b15zdnd11an1n32x5 FILLER_12_1371 ();
 b15zdnd11an1n16x5 FILLER_12_1403 ();
 b15zdnd11an1n08x5 FILLER_12_1419 ();
 b15zdnd11an1n64x5 FILLER_12_1430 ();
 b15zdnd11an1n64x5 FILLER_12_1494 ();
 b15zdnd11an1n08x5 FILLER_12_1558 ();
 b15zdnd11an1n04x5 FILLER_12_1566 ();
 b15zdnd00an1n01x5 FILLER_12_1570 ();
 b15zdnd11an1n04x5 FILLER_12_1574 ();
 b15zdnd11an1n64x5 FILLER_12_1581 ();
 b15zdnd11an1n64x5 FILLER_12_1645 ();
 b15zdnd11an1n64x5 FILLER_12_1709 ();
 b15zdnd11an1n64x5 FILLER_12_1773 ();
 b15zdnd11an1n64x5 FILLER_12_1837 ();
 b15zdnd00an1n02x5 FILLER_12_1901 ();
 b15zdnd00an1n01x5 FILLER_12_1903 ();
 b15zdnd11an1n08x5 FILLER_12_1908 ();
 b15zdnd00an1n02x5 FILLER_12_1916 ();
 b15zdnd11an1n04x5 FILLER_12_1921 ();
 b15zdnd11an1n04x5 FILLER_12_1934 ();
 b15zdnd11an1n04x5 FILLER_12_1944 ();
 b15zdnd11an1n16x5 FILLER_12_1953 ();
 b15zdnd11an1n64x5 FILLER_12_2011 ();
 b15zdnd11an1n64x5 FILLER_12_2075 ();
 b15zdnd11an1n08x5 FILLER_12_2139 ();
 b15zdnd11an1n04x5 FILLER_12_2147 ();
 b15zdnd00an1n02x5 FILLER_12_2151 ();
 b15zdnd00an1n01x5 FILLER_12_2153 ();
 b15zdnd11an1n64x5 FILLER_12_2162 ();
 b15zdnd11an1n32x5 FILLER_12_2226 ();
 b15zdnd11an1n16x5 FILLER_12_2258 ();
 b15zdnd00an1n02x5 FILLER_12_2274 ();
 b15zdnd11an1n64x5 FILLER_13_0 ();
 b15zdnd11an1n64x5 FILLER_13_64 ();
 b15zdnd11an1n64x5 FILLER_13_128 ();
 b15zdnd11an1n64x5 FILLER_13_192 ();
 b15zdnd11an1n64x5 FILLER_13_256 ();
 b15zdnd11an1n64x5 FILLER_13_320 ();
 b15zdnd11an1n16x5 FILLER_13_384 ();
 b15zdnd11an1n08x5 FILLER_13_400 ();
 b15zdnd00an1n01x5 FILLER_13_408 ();
 b15zdnd11an1n32x5 FILLER_13_451 ();
 b15zdnd11an1n08x5 FILLER_13_483 ();
 b15zdnd00an1n02x5 FILLER_13_491 ();
 b15zdnd00an1n01x5 FILLER_13_493 ();
 b15zdnd11an1n64x5 FILLER_13_498 ();
 b15zdnd11an1n16x5 FILLER_13_562 ();
 b15zdnd11an1n04x5 FILLER_13_578 ();
 b15zdnd00an1n01x5 FILLER_13_582 ();
 b15zdnd11an1n64x5 FILLER_13_635 ();
 b15zdnd11an1n08x5 FILLER_13_699 ();
 b15zdnd00an1n01x5 FILLER_13_707 ();
 b15zdnd11an1n32x5 FILLER_13_715 ();
 b15zdnd11an1n16x5 FILLER_13_747 ();
 b15zdnd11an1n04x5 FILLER_13_763 ();
 b15zdnd00an1n01x5 FILLER_13_767 ();
 b15zdnd11an1n32x5 FILLER_13_810 ();
 b15zdnd11an1n16x5 FILLER_13_842 ();
 b15zdnd11an1n08x5 FILLER_13_858 ();
 b15zdnd11an1n04x5 FILLER_13_869 ();
 b15zdnd11an1n04x5 FILLER_13_876 ();
 b15zdnd11an1n04x5 FILLER_13_883 ();
 b15zdnd00an1n01x5 FILLER_13_887 ();
 b15zdnd11an1n32x5 FILLER_13_891 ();
 b15zdnd11an1n16x5 FILLER_13_923 ();
 b15zdnd11an1n04x5 FILLER_13_939 ();
 b15zdnd11an1n08x5 FILLER_13_949 ();
 b15zdnd00an1n02x5 FILLER_13_957 ();
 b15zdnd11an1n32x5 FILLER_13_1001 ();
 b15zdnd11an1n16x5 FILLER_13_1033 ();
 b15zdnd11an1n32x5 FILLER_13_1091 ();
 b15zdnd11an1n04x5 FILLER_13_1126 ();
 b15zdnd00an1n02x5 FILLER_13_1130 ();
 b15zdnd00an1n01x5 FILLER_13_1132 ();
 b15zdnd11an1n64x5 FILLER_13_1136 ();
 b15zdnd11an1n64x5 FILLER_13_1200 ();
 b15zdnd11an1n64x5 FILLER_13_1264 ();
 b15zdnd11an1n64x5 FILLER_13_1328 ();
 b15zdnd11an1n08x5 FILLER_13_1392 ();
 b15zdnd00an1n01x5 FILLER_13_1400 ();
 b15zdnd11an1n64x5 FILLER_13_1453 ();
 b15zdnd11an1n32x5 FILLER_13_1517 ();
 b15zdnd11an1n16x5 FILLER_13_1549 ();
 b15zdnd11an1n04x5 FILLER_13_1565 ();
 b15zdnd00an1n02x5 FILLER_13_1569 ();
 b15zdnd00an1n01x5 FILLER_13_1571 ();
 b15zdnd11an1n08x5 FILLER_13_1614 ();
 b15zdnd11an1n04x5 FILLER_13_1622 ();
 b15zdnd00an1n02x5 FILLER_13_1626 ();
 b15zdnd00an1n01x5 FILLER_13_1628 ();
 b15zdnd11an1n64x5 FILLER_13_1656 ();
 b15zdnd11an1n04x5 FILLER_13_1720 ();
 b15zdnd00an1n02x5 FILLER_13_1724 ();
 b15zdnd11an1n64x5 FILLER_13_1778 ();
 b15zdnd11an1n32x5 FILLER_13_1842 ();
 b15zdnd11an1n16x5 FILLER_13_1874 ();
 b15zdnd11an1n08x5 FILLER_13_1890 ();
 b15zdnd11an1n04x5 FILLER_13_1898 ();
 b15zdnd11an1n16x5 FILLER_13_1909 ();
 b15zdnd11an1n08x5 FILLER_13_1925 ();
 b15zdnd11an1n04x5 FILLER_13_1933 ();
 b15zdnd00an1n02x5 FILLER_13_1937 ();
 b15zdnd00an1n01x5 FILLER_13_1939 ();
 b15zdnd11an1n04x5 FILLER_13_1982 ();
 b15zdnd11an1n04x5 FILLER_13_1989 ();
 b15zdnd11an1n64x5 FILLER_13_1996 ();
 b15zdnd11an1n64x5 FILLER_13_2060 ();
 b15zdnd11an1n64x5 FILLER_13_2124 ();
 b15zdnd11an1n64x5 FILLER_13_2188 ();
 b15zdnd11an1n32x5 FILLER_13_2252 ();
 b15zdnd11an1n64x5 FILLER_14_8 ();
 b15zdnd11an1n64x5 FILLER_14_72 ();
 b15zdnd11an1n64x5 FILLER_14_136 ();
 b15zdnd11an1n64x5 FILLER_14_200 ();
 b15zdnd11an1n64x5 FILLER_14_264 ();
 b15zdnd11an1n64x5 FILLER_14_328 ();
 b15zdnd11an1n32x5 FILLER_14_392 ();
 b15zdnd11an1n08x5 FILLER_14_466 ();
 b15zdnd11an1n04x5 FILLER_14_474 ();
 b15zdnd00an1n02x5 FILLER_14_478 ();
 b15zdnd00an1n01x5 FILLER_14_480 ();
 b15zdnd11an1n64x5 FILLER_14_495 ();
 b15zdnd11an1n32x5 FILLER_14_559 ();
 b15zdnd11an1n08x5 FILLER_14_591 ();
 b15zdnd00an1n02x5 FILLER_14_599 ();
 b15zdnd11an1n04x5 FILLER_14_604 ();
 b15zdnd11an1n32x5 FILLER_14_611 ();
 b15zdnd11an1n16x5 FILLER_14_643 ();
 b15zdnd11an1n08x5 FILLER_14_659 ();
 b15zdnd11an1n04x5 FILLER_14_667 ();
 b15zdnd00an1n02x5 FILLER_14_671 ();
 b15zdnd00an1n01x5 FILLER_14_673 ();
 b15zdnd11an1n32x5 FILLER_14_682 ();
 b15zdnd11an1n04x5 FILLER_14_714 ();
 b15zdnd11an1n32x5 FILLER_14_726 ();
 b15zdnd11an1n64x5 FILLER_14_778 ();
 b15zdnd11an1n32x5 FILLER_14_842 ();
 b15zdnd11an1n04x5 FILLER_14_877 ();
 b15zdnd11an1n64x5 FILLER_14_884 ();
 b15zdnd11an1n08x5 FILLER_14_948 ();
 b15zdnd00an1n01x5 FILLER_14_956 ();
 b15zdnd11an1n08x5 FILLER_14_964 ();
 b15zdnd00an1n02x5 FILLER_14_972 ();
 b15zdnd11an1n04x5 FILLER_14_981 ();
 b15zdnd11an1n64x5 FILLER_14_988 ();
 b15zdnd11an1n16x5 FILLER_14_1052 ();
 b15zdnd00an1n02x5 FILLER_14_1068 ();
 b15zdnd00an1n01x5 FILLER_14_1070 ();
 b15zdnd11an1n04x5 FILLER_14_1074 ();
 b15zdnd11an1n08x5 FILLER_14_1081 ();
 b15zdnd11an1n04x5 FILLER_14_1089 ();
 b15zdnd00an1n02x5 FILLER_14_1093 ();
 b15zdnd00an1n01x5 FILLER_14_1095 ();
 b15zdnd11an1n64x5 FILLER_14_1148 ();
 b15zdnd11an1n64x5 FILLER_14_1212 ();
 b15zdnd11an1n64x5 FILLER_14_1276 ();
 b15zdnd11an1n64x5 FILLER_14_1340 ();
 b15zdnd11an1n08x5 FILLER_14_1404 ();
 b15zdnd11an1n04x5 FILLER_14_1412 ();
 b15zdnd00an1n01x5 FILLER_14_1416 ();
 b15zdnd11an1n64x5 FILLER_14_1459 ();
 b15zdnd11an1n64x5 FILLER_14_1523 ();
 b15zdnd11an1n64x5 FILLER_14_1587 ();
 b15zdnd11an1n32x5 FILLER_14_1651 ();
 b15zdnd11an1n16x5 FILLER_14_1683 ();
 b15zdnd11an1n04x5 FILLER_14_1699 ();
 b15zdnd00an1n02x5 FILLER_14_1703 ();
 b15zdnd00an1n01x5 FILLER_14_1705 ();
 b15zdnd11an1n32x5 FILLER_14_1709 ();
 b15zdnd11an1n04x5 FILLER_14_1741 ();
 b15zdnd11an1n04x5 FILLER_14_1748 ();
 b15zdnd11an1n04x5 FILLER_14_1755 ();
 b15zdnd11an1n64x5 FILLER_14_1762 ();
 b15zdnd11an1n64x5 FILLER_14_1826 ();
 b15zdnd11an1n64x5 FILLER_14_1890 ();
 b15zdnd00an1n01x5 FILLER_14_1954 ();
 b15zdnd11an1n64x5 FILLER_14_2007 ();
 b15zdnd11an1n64x5 FILLER_14_2071 ();
 b15zdnd11an1n16x5 FILLER_14_2135 ();
 b15zdnd00an1n02x5 FILLER_14_2151 ();
 b15zdnd00an1n01x5 FILLER_14_2153 ();
 b15zdnd11an1n64x5 FILLER_14_2162 ();
 b15zdnd11an1n32x5 FILLER_14_2226 ();
 b15zdnd11an1n16x5 FILLER_14_2258 ();
 b15zdnd00an1n02x5 FILLER_14_2274 ();
 b15zdnd11an1n64x5 FILLER_15_0 ();
 b15zdnd11an1n64x5 FILLER_15_64 ();
 b15zdnd11an1n64x5 FILLER_15_128 ();
 b15zdnd11an1n64x5 FILLER_15_192 ();
 b15zdnd11an1n64x5 FILLER_15_256 ();
 b15zdnd11an1n64x5 FILLER_15_320 ();
 b15zdnd11an1n64x5 FILLER_15_384 ();
 b15zdnd11an1n32x5 FILLER_15_448 ();
 b15zdnd00an1n01x5 FILLER_15_480 ();
 b15zdnd11an1n32x5 FILLER_15_523 ();
 b15zdnd11an1n08x5 FILLER_15_555 ();
 b15zdnd00an1n01x5 FILLER_15_563 ();
 b15zdnd11an1n64x5 FILLER_15_606 ();
 b15zdnd11an1n16x5 FILLER_15_670 ();
 b15zdnd11an1n08x5 FILLER_15_686 ();
 b15zdnd00an1n02x5 FILLER_15_694 ();
 b15zdnd11an1n64x5 FILLER_15_702 ();
 b15zdnd11an1n64x5 FILLER_15_766 ();
 b15zdnd11an1n64x5 FILLER_15_830 ();
 b15zdnd11an1n64x5 FILLER_15_894 ();
 b15zdnd11an1n04x5 FILLER_15_958 ();
 b15zdnd00an1n01x5 FILLER_15_962 ();
 b15zdnd11an1n08x5 FILLER_15_969 ();
 b15zdnd00an1n02x5 FILLER_15_977 ();
 b15zdnd11an1n64x5 FILLER_15_982 ();
 b15zdnd11an1n64x5 FILLER_15_1046 ();
 b15zdnd11an1n08x5 FILLER_15_1110 ();
 b15zdnd00an1n01x5 FILLER_15_1118 ();
 b15zdnd11an1n64x5 FILLER_15_1122 ();
 b15zdnd11an1n64x5 FILLER_15_1186 ();
 b15zdnd11an1n64x5 FILLER_15_1250 ();
 b15zdnd11an1n32x5 FILLER_15_1314 ();
 b15zdnd11an1n16x5 FILLER_15_1346 ();
 b15zdnd11an1n08x5 FILLER_15_1362 ();
 b15zdnd11an1n16x5 FILLER_15_1390 ();
 b15zdnd11an1n08x5 FILLER_15_1406 ();
 b15zdnd11an1n04x5 FILLER_15_1414 ();
 b15zdnd00an1n01x5 FILLER_15_1418 ();
 b15zdnd11an1n04x5 FILLER_15_1422 ();
 b15zdnd11an1n04x5 FILLER_15_1429 ();
 b15zdnd11an1n64x5 FILLER_15_1441 ();
 b15zdnd11an1n08x5 FILLER_15_1505 ();
 b15zdnd11an1n04x5 FILLER_15_1513 ();
 b15zdnd00an1n02x5 FILLER_15_1517 ();
 b15zdnd00an1n01x5 FILLER_15_1519 ();
 b15zdnd11an1n64x5 FILLER_15_1572 ();
 b15zdnd11an1n32x5 FILLER_15_1636 ();
 b15zdnd11an1n04x5 FILLER_15_1668 ();
 b15zdnd00an1n01x5 FILLER_15_1672 ();
 b15zdnd11an1n64x5 FILLER_15_1713 ();
 b15zdnd11an1n64x5 FILLER_15_1777 ();
 b15zdnd11an1n64x5 FILLER_15_1841 ();
 b15zdnd11an1n64x5 FILLER_15_1905 ();
 b15zdnd11an1n64x5 FILLER_15_1969 ();
 b15zdnd11an1n64x5 FILLER_15_2033 ();
 b15zdnd11an1n64x5 FILLER_15_2097 ();
 b15zdnd11an1n64x5 FILLER_15_2161 ();
 b15zdnd11an1n32x5 FILLER_15_2225 ();
 b15zdnd11an1n16x5 FILLER_15_2257 ();
 b15zdnd11an1n08x5 FILLER_15_2273 ();
 b15zdnd00an1n02x5 FILLER_15_2281 ();
 b15zdnd00an1n01x5 FILLER_15_2283 ();
 b15zdnd11an1n64x5 FILLER_16_8 ();
 b15zdnd11an1n64x5 FILLER_16_72 ();
 b15zdnd11an1n64x5 FILLER_16_136 ();
 b15zdnd11an1n32x5 FILLER_16_200 ();
 b15zdnd11an1n16x5 FILLER_16_232 ();
 b15zdnd00an1n01x5 FILLER_16_248 ();
 b15zdnd11an1n64x5 FILLER_16_294 ();
 b15zdnd11an1n32x5 FILLER_16_358 ();
 b15zdnd11an1n08x5 FILLER_16_390 ();
 b15zdnd11an1n04x5 FILLER_16_398 ();
 b15zdnd00an1n02x5 FILLER_16_402 ();
 b15zdnd11an1n64x5 FILLER_16_407 ();
 b15zdnd11an1n64x5 FILLER_16_471 ();
 b15zdnd11an1n64x5 FILLER_16_535 ();
 b15zdnd11an1n32x5 FILLER_16_599 ();
 b15zdnd11an1n16x5 FILLER_16_631 ();
 b15zdnd00an1n02x5 FILLER_16_647 ();
 b15zdnd11an1n32x5 FILLER_16_656 ();
 b15zdnd11an1n16x5 FILLER_16_688 ();
 b15zdnd11an1n08x5 FILLER_16_704 ();
 b15zdnd11an1n04x5 FILLER_16_712 ();
 b15zdnd00an1n02x5 FILLER_16_716 ();
 b15zdnd11an1n64x5 FILLER_16_726 ();
 b15zdnd11an1n64x5 FILLER_16_790 ();
 b15zdnd11an1n64x5 FILLER_16_854 ();
 b15zdnd11an1n64x5 FILLER_16_918 ();
 b15zdnd11an1n64x5 FILLER_16_982 ();
 b15zdnd11an1n64x5 FILLER_16_1046 ();
 b15zdnd11an1n64x5 FILLER_16_1110 ();
 b15zdnd11an1n64x5 FILLER_16_1174 ();
 b15zdnd11an1n64x5 FILLER_16_1238 ();
 b15zdnd11an1n64x5 FILLER_16_1302 ();
 b15zdnd11an1n32x5 FILLER_16_1366 ();
 b15zdnd00an1n02x5 FILLER_16_1398 ();
 b15zdnd11an1n64x5 FILLER_16_1442 ();
 b15zdnd11an1n32x5 FILLER_16_1506 ();
 b15zdnd11an1n04x5 FILLER_16_1538 ();
 b15zdnd00an1n01x5 FILLER_16_1542 ();
 b15zdnd11an1n04x5 FILLER_16_1546 ();
 b15zdnd11an1n64x5 FILLER_16_1553 ();
 b15zdnd11an1n16x5 FILLER_16_1617 ();
 b15zdnd11an1n04x5 FILLER_16_1633 ();
 b15zdnd11an1n32x5 FILLER_16_1663 ();
 b15zdnd11an1n16x5 FILLER_16_1695 ();
 b15zdnd11an1n64x5 FILLER_16_1714 ();
 b15zdnd11an1n64x5 FILLER_16_1778 ();
 b15zdnd11an1n64x5 FILLER_16_1842 ();
 b15zdnd11an1n64x5 FILLER_16_1906 ();
 b15zdnd11an1n64x5 FILLER_16_1970 ();
 b15zdnd11an1n64x5 FILLER_16_2034 ();
 b15zdnd11an1n32x5 FILLER_16_2098 ();
 b15zdnd11an1n16x5 FILLER_16_2130 ();
 b15zdnd11an1n08x5 FILLER_16_2146 ();
 b15zdnd11an1n64x5 FILLER_16_2162 ();
 b15zdnd11an1n32x5 FILLER_16_2226 ();
 b15zdnd11an1n16x5 FILLER_16_2258 ();
 b15zdnd00an1n02x5 FILLER_16_2274 ();
 b15zdnd11an1n64x5 FILLER_17_0 ();
 b15zdnd11an1n64x5 FILLER_17_64 ();
 b15zdnd11an1n64x5 FILLER_17_128 ();
 b15zdnd11an1n64x5 FILLER_17_192 ();
 b15zdnd11an1n64x5 FILLER_17_256 ();
 b15zdnd11an1n32x5 FILLER_17_320 ();
 b15zdnd11an1n16x5 FILLER_17_352 ();
 b15zdnd11an1n08x5 FILLER_17_368 ();
 b15zdnd00an1n01x5 FILLER_17_376 ();
 b15zdnd11an1n64x5 FILLER_17_429 ();
 b15zdnd11an1n32x5 FILLER_17_493 ();
 b15zdnd11an1n04x5 FILLER_17_525 ();
 b15zdnd00an1n02x5 FILLER_17_529 ();
 b15zdnd11an1n64x5 FILLER_17_534 ();
 b15zdnd11an1n32x5 FILLER_17_598 ();
 b15zdnd11an1n04x5 FILLER_17_630 ();
 b15zdnd11an1n32x5 FILLER_17_651 ();
 b15zdnd11an1n16x5 FILLER_17_683 ();
 b15zdnd11an1n64x5 FILLER_17_741 ();
 b15zdnd11an1n64x5 FILLER_17_805 ();
 b15zdnd11an1n08x5 FILLER_17_869 ();
 b15zdnd11an1n04x5 FILLER_17_877 ();
 b15zdnd11an1n32x5 FILLER_17_923 ();
 b15zdnd11an1n04x5 FILLER_17_955 ();
 b15zdnd00an1n02x5 FILLER_17_959 ();
 b15zdnd11an1n04x5 FILLER_17_1003 ();
 b15zdnd00an1n02x5 FILLER_17_1007 ();
 b15zdnd11an1n64x5 FILLER_17_1051 ();
 b15zdnd11an1n32x5 FILLER_17_1115 ();
 b15zdnd11an1n16x5 FILLER_17_1147 ();
 b15zdnd00an1n01x5 FILLER_17_1163 ();
 b15zdnd11an1n64x5 FILLER_17_1184 ();
 b15zdnd11an1n64x5 FILLER_17_1248 ();
 b15zdnd11an1n32x5 FILLER_17_1312 ();
 b15zdnd11an1n16x5 FILLER_17_1344 ();
 b15zdnd11an1n08x5 FILLER_17_1360 ();
 b15zdnd11an1n64x5 FILLER_17_1410 ();
 b15zdnd11an1n64x5 FILLER_17_1474 ();
 b15zdnd00an1n01x5 FILLER_17_1538 ();
 b15zdnd11an1n64x5 FILLER_17_1542 ();
 b15zdnd11an1n64x5 FILLER_17_1606 ();
 b15zdnd11an1n64x5 FILLER_17_1670 ();
 b15zdnd11an1n64x5 FILLER_17_1734 ();
 b15zdnd11an1n64x5 FILLER_17_1798 ();
 b15zdnd11an1n32x5 FILLER_17_1862 ();
 b15zdnd11an1n16x5 FILLER_17_1894 ();
 b15zdnd00an1n01x5 FILLER_17_1910 ();
 b15zdnd11an1n64x5 FILLER_17_1953 ();
 b15zdnd11an1n64x5 FILLER_17_2017 ();
 b15zdnd11an1n64x5 FILLER_17_2081 ();
 b15zdnd11an1n64x5 FILLER_17_2145 ();
 b15zdnd11an1n64x5 FILLER_17_2209 ();
 b15zdnd11an1n08x5 FILLER_17_2273 ();
 b15zdnd00an1n02x5 FILLER_17_2281 ();
 b15zdnd00an1n01x5 FILLER_17_2283 ();
 b15zdnd11an1n64x5 FILLER_18_8 ();
 b15zdnd11an1n64x5 FILLER_18_72 ();
 b15zdnd11an1n64x5 FILLER_18_136 ();
 b15zdnd11an1n64x5 FILLER_18_200 ();
 b15zdnd11an1n64x5 FILLER_18_264 ();
 b15zdnd11an1n64x5 FILLER_18_328 ();
 b15zdnd11an1n04x5 FILLER_18_392 ();
 b15zdnd11an1n04x5 FILLER_18_399 ();
 b15zdnd11an1n64x5 FILLER_18_406 ();
 b15zdnd11an1n32x5 FILLER_18_470 ();
 b15zdnd00an1n02x5 FILLER_18_502 ();
 b15zdnd11an1n64x5 FILLER_18_556 ();
 b15zdnd11an1n16x5 FILLER_18_620 ();
 b15zdnd11an1n08x5 FILLER_18_636 ();
 b15zdnd11an1n04x5 FILLER_18_644 ();
 b15zdnd00an1n01x5 FILLER_18_648 ();
 b15zdnd11an1n16x5 FILLER_18_691 ();
 b15zdnd11an1n08x5 FILLER_18_707 ();
 b15zdnd00an1n02x5 FILLER_18_715 ();
 b15zdnd00an1n01x5 FILLER_18_717 ();
 b15zdnd11an1n32x5 FILLER_18_726 ();
 b15zdnd00an1n02x5 FILLER_18_758 ();
 b15zdnd00an1n01x5 FILLER_18_760 ();
 b15zdnd11an1n64x5 FILLER_18_773 ();
 b15zdnd11an1n64x5 FILLER_18_837 ();
 b15zdnd11an1n64x5 FILLER_18_901 ();
 b15zdnd11an1n64x5 FILLER_18_965 ();
 b15zdnd11an1n64x5 FILLER_18_1029 ();
 b15zdnd11an1n32x5 FILLER_18_1093 ();
 b15zdnd11an1n08x5 FILLER_18_1125 ();
 b15zdnd11an1n64x5 FILLER_18_1153 ();
 b15zdnd11an1n64x5 FILLER_18_1217 ();
 b15zdnd11an1n64x5 FILLER_18_1281 ();
 b15zdnd11an1n64x5 FILLER_18_1345 ();
 b15zdnd11an1n64x5 FILLER_18_1451 ();
 b15zdnd11an1n64x5 FILLER_18_1515 ();
 b15zdnd11an1n64x5 FILLER_18_1579 ();
 b15zdnd11an1n16x5 FILLER_18_1643 ();
 b15zdnd11an1n08x5 FILLER_18_1659 ();
 b15zdnd11an1n04x5 FILLER_18_1667 ();
 b15zdnd00an1n02x5 FILLER_18_1671 ();
 b15zdnd11an1n64x5 FILLER_18_1715 ();
 b15zdnd11an1n64x5 FILLER_18_1779 ();
 b15zdnd11an1n64x5 FILLER_18_1843 ();
 b15zdnd11an1n64x5 FILLER_18_1907 ();
 b15zdnd11an1n64x5 FILLER_18_1971 ();
 b15zdnd11an1n64x5 FILLER_18_2035 ();
 b15zdnd11an1n32x5 FILLER_18_2099 ();
 b15zdnd11an1n16x5 FILLER_18_2131 ();
 b15zdnd11an1n04x5 FILLER_18_2147 ();
 b15zdnd00an1n02x5 FILLER_18_2151 ();
 b15zdnd00an1n01x5 FILLER_18_2153 ();
 b15zdnd11an1n64x5 FILLER_18_2162 ();
 b15zdnd11an1n32x5 FILLER_18_2226 ();
 b15zdnd11an1n16x5 FILLER_18_2258 ();
 b15zdnd00an1n02x5 FILLER_18_2274 ();
 b15zdnd11an1n64x5 FILLER_19_0 ();
 b15zdnd11an1n64x5 FILLER_19_64 ();
 b15zdnd11an1n64x5 FILLER_19_128 ();
 b15zdnd11an1n64x5 FILLER_19_192 ();
 b15zdnd11an1n64x5 FILLER_19_256 ();
 b15zdnd11an1n64x5 FILLER_19_320 ();
 b15zdnd11an1n64x5 FILLER_19_384 ();
 b15zdnd11an1n64x5 FILLER_19_448 ();
 b15zdnd11an1n16x5 FILLER_19_512 ();
 b15zdnd00an1n02x5 FILLER_19_528 ();
 b15zdnd11an1n04x5 FILLER_19_533 ();
 b15zdnd11an1n32x5 FILLER_19_540 ();
 b15zdnd11an1n16x5 FILLER_19_572 ();
 b15zdnd11an1n08x5 FILLER_19_588 ();
 b15zdnd11an1n04x5 FILLER_19_596 ();
 b15zdnd11an1n04x5 FILLER_19_642 ();
 b15zdnd11an1n64x5 FILLER_19_688 ();
 b15zdnd11an1n64x5 FILLER_19_752 ();
 b15zdnd11an1n16x5 FILLER_19_816 ();
 b15zdnd11an1n08x5 FILLER_19_832 ();
 b15zdnd00an1n02x5 FILLER_19_840 ();
 b15zdnd11an1n64x5 FILLER_19_884 ();
 b15zdnd11an1n32x5 FILLER_19_948 ();
 b15zdnd11an1n16x5 FILLER_19_980 ();
 b15zdnd11an1n08x5 FILLER_19_996 ();
 b15zdnd11an1n32x5 FILLER_19_1046 ();
 b15zdnd11an1n16x5 FILLER_19_1078 ();
 b15zdnd11an1n08x5 FILLER_19_1094 ();
 b15zdnd11an1n04x5 FILLER_19_1102 ();
 b15zdnd11an1n08x5 FILLER_19_1148 ();
 b15zdnd11an1n04x5 FILLER_19_1156 ();
 b15zdnd11an1n64x5 FILLER_19_1202 ();
 b15zdnd11an1n64x5 FILLER_19_1266 ();
 b15zdnd11an1n32x5 FILLER_19_1330 ();
 b15zdnd11an1n16x5 FILLER_19_1362 ();
 b15zdnd11an1n08x5 FILLER_19_1378 ();
 b15zdnd11an1n04x5 FILLER_19_1386 ();
 b15zdnd00an1n02x5 FILLER_19_1390 ();
 b15zdnd11an1n08x5 FILLER_19_1412 ();
 b15zdnd00an1n01x5 FILLER_19_1420 ();
 b15zdnd11an1n64x5 FILLER_19_1435 ();
 b15zdnd11an1n64x5 FILLER_19_1499 ();
 b15zdnd11an1n64x5 FILLER_19_1563 ();
 b15zdnd11an1n64x5 FILLER_19_1627 ();
 b15zdnd11an1n32x5 FILLER_19_1691 ();
 b15zdnd11an1n08x5 FILLER_19_1723 ();
 b15zdnd11an1n04x5 FILLER_19_1731 ();
 b15zdnd00an1n02x5 FILLER_19_1735 ();
 b15zdnd00an1n01x5 FILLER_19_1737 ();
 b15zdnd11an1n64x5 FILLER_19_1755 ();
 b15zdnd11an1n64x5 FILLER_19_1819 ();
 b15zdnd11an1n64x5 FILLER_19_1883 ();
 b15zdnd11an1n64x5 FILLER_19_1947 ();
 b15zdnd11an1n64x5 FILLER_19_2011 ();
 b15zdnd11an1n64x5 FILLER_19_2075 ();
 b15zdnd11an1n64x5 FILLER_19_2139 ();
 b15zdnd11an1n64x5 FILLER_19_2203 ();
 b15zdnd11an1n16x5 FILLER_19_2267 ();
 b15zdnd00an1n01x5 FILLER_19_2283 ();
 b15zdnd11an1n64x5 FILLER_20_8 ();
 b15zdnd11an1n64x5 FILLER_20_72 ();
 b15zdnd11an1n64x5 FILLER_20_136 ();
 b15zdnd11an1n64x5 FILLER_20_200 ();
 b15zdnd11an1n64x5 FILLER_20_264 ();
 b15zdnd11an1n64x5 FILLER_20_328 ();
 b15zdnd11an1n64x5 FILLER_20_392 ();
 b15zdnd11an1n64x5 FILLER_20_456 ();
 b15zdnd11an1n64x5 FILLER_20_520 ();
 b15zdnd11an1n64x5 FILLER_20_584 ();
 b15zdnd11an1n64x5 FILLER_20_648 ();
 b15zdnd11an1n04x5 FILLER_20_712 ();
 b15zdnd00an1n02x5 FILLER_20_716 ();
 b15zdnd11an1n32x5 FILLER_20_726 ();
 b15zdnd11an1n16x5 FILLER_20_758 ();
 b15zdnd11an1n08x5 FILLER_20_774 ();
 b15zdnd11an1n04x5 FILLER_20_782 ();
 b15zdnd00an1n02x5 FILLER_20_786 ();
 b15zdnd11an1n64x5 FILLER_20_830 ();
 b15zdnd11an1n64x5 FILLER_20_894 ();
 b15zdnd11an1n32x5 FILLER_20_958 ();
 b15zdnd11an1n16x5 FILLER_20_990 ();
 b15zdnd11an1n04x5 FILLER_20_1006 ();
 b15zdnd00an1n01x5 FILLER_20_1010 ();
 b15zdnd11an1n64x5 FILLER_20_1053 ();
 b15zdnd11an1n64x5 FILLER_20_1117 ();
 b15zdnd11an1n64x5 FILLER_20_1181 ();
 b15zdnd11an1n64x5 FILLER_20_1245 ();
 b15zdnd11an1n64x5 FILLER_20_1309 ();
 b15zdnd11an1n32x5 FILLER_20_1373 ();
 b15zdnd11an1n04x5 FILLER_20_1405 ();
 b15zdnd11an1n04x5 FILLER_20_1451 ();
 b15zdnd00an1n02x5 FILLER_20_1455 ();
 b15zdnd11an1n64x5 FILLER_20_1499 ();
 b15zdnd11an1n64x5 FILLER_20_1563 ();
 b15zdnd11an1n64x5 FILLER_20_1627 ();
 b15zdnd11an1n32x5 FILLER_20_1691 ();
 b15zdnd11an1n16x5 FILLER_20_1723 ();
 b15zdnd00an1n01x5 FILLER_20_1739 ();
 b15zdnd11an1n64x5 FILLER_20_1746 ();
 b15zdnd11an1n64x5 FILLER_20_1810 ();
 b15zdnd11an1n64x5 FILLER_20_1874 ();
 b15zdnd11an1n64x5 FILLER_20_1938 ();
 b15zdnd11an1n64x5 FILLER_20_2002 ();
 b15zdnd11an1n64x5 FILLER_20_2066 ();
 b15zdnd11an1n16x5 FILLER_20_2130 ();
 b15zdnd11an1n08x5 FILLER_20_2146 ();
 b15zdnd11an1n64x5 FILLER_20_2162 ();
 b15zdnd11an1n32x5 FILLER_20_2226 ();
 b15zdnd11an1n16x5 FILLER_20_2258 ();
 b15zdnd00an1n02x5 FILLER_20_2274 ();
 b15zdnd11an1n64x5 FILLER_21_0 ();
 b15zdnd11an1n64x5 FILLER_21_64 ();
 b15zdnd11an1n64x5 FILLER_21_128 ();
 b15zdnd11an1n64x5 FILLER_21_192 ();
 b15zdnd11an1n64x5 FILLER_21_256 ();
 b15zdnd11an1n64x5 FILLER_21_320 ();
 b15zdnd11an1n64x5 FILLER_21_384 ();
 b15zdnd11an1n64x5 FILLER_21_448 ();
 b15zdnd11an1n64x5 FILLER_21_512 ();
 b15zdnd11an1n64x5 FILLER_21_576 ();
 b15zdnd11an1n64x5 FILLER_21_640 ();
 b15zdnd11an1n64x5 FILLER_21_704 ();
 b15zdnd11an1n64x5 FILLER_21_768 ();
 b15zdnd11an1n64x5 FILLER_21_832 ();
 b15zdnd11an1n64x5 FILLER_21_896 ();
 b15zdnd11an1n16x5 FILLER_21_960 ();
 b15zdnd11an1n08x5 FILLER_21_976 ();
 b15zdnd11an1n04x5 FILLER_21_984 ();
 b15zdnd11an1n64x5 FILLER_21_997 ();
 b15zdnd11an1n64x5 FILLER_21_1061 ();
 b15zdnd11an1n64x5 FILLER_21_1125 ();
 b15zdnd11an1n64x5 FILLER_21_1189 ();
 b15zdnd11an1n64x5 FILLER_21_1253 ();
 b15zdnd11an1n64x5 FILLER_21_1317 ();
 b15zdnd11an1n64x5 FILLER_21_1381 ();
 b15zdnd11an1n64x5 FILLER_21_1445 ();
 b15zdnd11an1n64x5 FILLER_21_1509 ();
 b15zdnd11an1n64x5 FILLER_21_1573 ();
 b15zdnd11an1n08x5 FILLER_21_1637 ();
 b15zdnd00an1n02x5 FILLER_21_1645 ();
 b15zdnd00an1n01x5 FILLER_21_1647 ();
 b15zdnd11an1n08x5 FILLER_21_1651 ();
 b15zdnd11an1n04x5 FILLER_21_1659 ();
 b15zdnd00an1n02x5 FILLER_21_1663 ();
 b15zdnd00an1n01x5 FILLER_21_1665 ();
 b15zdnd11an1n64x5 FILLER_21_1672 ();
 b15zdnd11an1n64x5 FILLER_21_1736 ();
 b15zdnd11an1n64x5 FILLER_21_1800 ();
 b15zdnd11an1n32x5 FILLER_21_1864 ();
 b15zdnd11an1n16x5 FILLER_21_1896 ();
 b15zdnd11an1n08x5 FILLER_21_1912 ();
 b15zdnd11an1n64x5 FILLER_21_1923 ();
 b15zdnd11an1n64x5 FILLER_21_1987 ();
 b15zdnd11an1n64x5 FILLER_21_2051 ();
 b15zdnd11an1n64x5 FILLER_21_2115 ();
 b15zdnd11an1n64x5 FILLER_21_2179 ();
 b15zdnd11an1n32x5 FILLER_21_2243 ();
 b15zdnd11an1n08x5 FILLER_21_2275 ();
 b15zdnd00an1n01x5 FILLER_21_2283 ();
 b15zdnd11an1n64x5 FILLER_22_8 ();
 b15zdnd11an1n64x5 FILLER_22_72 ();
 b15zdnd11an1n64x5 FILLER_22_136 ();
 b15zdnd11an1n64x5 FILLER_22_200 ();
 b15zdnd11an1n64x5 FILLER_22_264 ();
 b15zdnd11an1n64x5 FILLER_22_328 ();
 b15zdnd11an1n64x5 FILLER_22_392 ();
 b15zdnd11an1n64x5 FILLER_22_456 ();
 b15zdnd11an1n64x5 FILLER_22_520 ();
 b15zdnd11an1n64x5 FILLER_22_584 ();
 b15zdnd11an1n64x5 FILLER_22_648 ();
 b15zdnd11an1n04x5 FILLER_22_712 ();
 b15zdnd00an1n02x5 FILLER_22_716 ();
 b15zdnd11an1n32x5 FILLER_22_726 ();
 b15zdnd11an1n16x5 FILLER_22_758 ();
 b15zdnd11an1n04x5 FILLER_22_774 ();
 b15zdnd11an1n64x5 FILLER_22_820 ();
 b15zdnd11an1n32x5 FILLER_22_884 ();
 b15zdnd11an1n16x5 FILLER_22_916 ();
 b15zdnd11an1n08x5 FILLER_22_932 ();
 b15zdnd11an1n04x5 FILLER_22_940 ();
 b15zdnd00an1n01x5 FILLER_22_944 ();
 b15zdnd11an1n32x5 FILLER_22_987 ();
 b15zdnd11an1n16x5 FILLER_22_1019 ();
 b15zdnd00an1n02x5 FILLER_22_1035 ();
 b15zdnd11an1n64x5 FILLER_22_1079 ();
 b15zdnd11an1n64x5 FILLER_22_1143 ();
 b15zdnd11an1n64x5 FILLER_22_1207 ();
 b15zdnd11an1n64x5 FILLER_22_1271 ();
 b15zdnd11an1n08x5 FILLER_22_1335 ();
 b15zdnd00an1n02x5 FILLER_22_1343 ();
 b15zdnd00an1n01x5 FILLER_22_1345 ();
 b15zdnd11an1n64x5 FILLER_22_1366 ();
 b15zdnd11an1n64x5 FILLER_22_1430 ();
 b15zdnd11an1n64x5 FILLER_22_1494 ();
 b15zdnd11an1n64x5 FILLER_22_1558 ();
 b15zdnd11an1n16x5 FILLER_22_1622 ();
 b15zdnd11an1n04x5 FILLER_22_1638 ();
 b15zdnd00an1n02x5 FILLER_22_1642 ();
 b15zdnd00an1n01x5 FILLER_22_1644 ();
 b15zdnd11an1n32x5 FILLER_22_1666 ();
 b15zdnd11an1n16x5 FILLER_22_1698 ();
 b15zdnd11an1n08x5 FILLER_22_1714 ();
 b15zdnd11an1n64x5 FILLER_22_1746 ();
 b15zdnd11an1n64x5 FILLER_22_1810 ();
 b15zdnd11an1n32x5 FILLER_22_1874 ();
 b15zdnd11an1n08x5 FILLER_22_1906 ();
 b15zdnd11an1n04x5 FILLER_22_1914 ();
 b15zdnd00an1n02x5 FILLER_22_1918 ();
 b15zdnd11an1n64x5 FILLER_22_1923 ();
 b15zdnd11an1n64x5 FILLER_22_1987 ();
 b15zdnd11an1n64x5 FILLER_22_2051 ();
 b15zdnd11an1n32x5 FILLER_22_2115 ();
 b15zdnd11an1n04x5 FILLER_22_2147 ();
 b15zdnd00an1n02x5 FILLER_22_2151 ();
 b15zdnd00an1n01x5 FILLER_22_2153 ();
 b15zdnd11an1n64x5 FILLER_22_2162 ();
 b15zdnd11an1n32x5 FILLER_22_2226 ();
 b15zdnd11an1n16x5 FILLER_22_2258 ();
 b15zdnd00an1n02x5 FILLER_22_2274 ();
 b15zdnd11an1n64x5 FILLER_23_0 ();
 b15zdnd11an1n64x5 FILLER_23_64 ();
 b15zdnd11an1n64x5 FILLER_23_128 ();
 b15zdnd11an1n64x5 FILLER_23_192 ();
 b15zdnd11an1n64x5 FILLER_23_256 ();
 b15zdnd11an1n64x5 FILLER_23_320 ();
 b15zdnd11an1n64x5 FILLER_23_384 ();
 b15zdnd11an1n64x5 FILLER_23_448 ();
 b15zdnd11an1n64x5 FILLER_23_512 ();
 b15zdnd11an1n64x5 FILLER_23_576 ();
 b15zdnd11an1n64x5 FILLER_23_640 ();
 b15zdnd11an1n64x5 FILLER_23_704 ();
 b15zdnd11an1n64x5 FILLER_23_768 ();
 b15zdnd11an1n64x5 FILLER_23_832 ();
 b15zdnd11an1n32x5 FILLER_23_896 ();
 b15zdnd11an1n16x5 FILLER_23_928 ();
 b15zdnd11an1n08x5 FILLER_23_944 ();
 b15zdnd11an1n04x5 FILLER_23_952 ();
 b15zdnd00an1n02x5 FILLER_23_956 ();
 b15zdnd11an1n64x5 FILLER_23_1000 ();
 b15zdnd11an1n64x5 FILLER_23_1064 ();
 b15zdnd11an1n64x5 FILLER_23_1128 ();
 b15zdnd11an1n64x5 FILLER_23_1192 ();
 b15zdnd11an1n64x5 FILLER_23_1256 ();
 b15zdnd11an1n64x5 FILLER_23_1320 ();
 b15zdnd11an1n64x5 FILLER_23_1384 ();
 b15zdnd11an1n16x5 FILLER_23_1448 ();
 b15zdnd11an1n08x5 FILLER_23_1464 ();
 b15zdnd00an1n02x5 FILLER_23_1472 ();
 b15zdnd11an1n64x5 FILLER_23_1483 ();
 b15zdnd11an1n64x5 FILLER_23_1547 ();
 b15zdnd11an1n08x5 FILLER_23_1611 ();
 b15zdnd00an1n02x5 FILLER_23_1619 ();
 b15zdnd11an1n64x5 FILLER_23_1673 ();
 b15zdnd11an1n64x5 FILLER_23_1737 ();
 b15zdnd11an1n64x5 FILLER_23_1801 ();
 b15zdnd11an1n16x5 FILLER_23_1865 ();
 b15zdnd11an1n08x5 FILLER_23_1881 ();
 b15zdnd11an1n04x5 FILLER_23_1889 ();
 b15zdnd00an1n02x5 FILLER_23_1893 ();
 b15zdnd11an1n64x5 FILLER_23_1947 ();
 b15zdnd11an1n64x5 FILLER_23_2011 ();
 b15zdnd11an1n64x5 FILLER_23_2075 ();
 b15zdnd11an1n64x5 FILLER_23_2139 ();
 b15zdnd11an1n64x5 FILLER_23_2203 ();
 b15zdnd11an1n16x5 FILLER_23_2267 ();
 b15zdnd00an1n01x5 FILLER_23_2283 ();
 b15zdnd11an1n64x5 FILLER_24_8 ();
 b15zdnd11an1n64x5 FILLER_24_72 ();
 b15zdnd11an1n64x5 FILLER_24_136 ();
 b15zdnd11an1n64x5 FILLER_24_200 ();
 b15zdnd11an1n64x5 FILLER_24_264 ();
 b15zdnd11an1n64x5 FILLER_24_328 ();
 b15zdnd11an1n64x5 FILLER_24_392 ();
 b15zdnd11an1n64x5 FILLER_24_456 ();
 b15zdnd11an1n16x5 FILLER_24_520 ();
 b15zdnd11an1n04x5 FILLER_24_536 ();
 b15zdnd11an1n64x5 FILLER_24_582 ();
 b15zdnd11an1n32x5 FILLER_24_646 ();
 b15zdnd11an1n08x5 FILLER_24_678 ();
 b15zdnd11an1n04x5 FILLER_24_686 ();
 b15zdnd00an1n02x5 FILLER_24_690 ();
 b15zdnd00an1n01x5 FILLER_24_692 ();
 b15zdnd11an1n16x5 FILLER_24_696 ();
 b15zdnd11an1n04x5 FILLER_24_712 ();
 b15zdnd00an1n02x5 FILLER_24_716 ();
 b15zdnd11an1n64x5 FILLER_24_726 ();
 b15zdnd11an1n32x5 FILLER_24_790 ();
 b15zdnd11an1n16x5 FILLER_24_822 ();
 b15zdnd00an1n02x5 FILLER_24_838 ();
 b15zdnd11an1n64x5 FILLER_24_882 ();
 b15zdnd11an1n64x5 FILLER_24_946 ();
 b15zdnd11an1n64x5 FILLER_24_1010 ();
 b15zdnd11an1n08x5 FILLER_24_1074 ();
 b15zdnd11an1n04x5 FILLER_24_1082 ();
 b15zdnd00an1n01x5 FILLER_24_1086 ();
 b15zdnd11an1n64x5 FILLER_24_1090 ();
 b15zdnd11an1n64x5 FILLER_24_1154 ();
 b15zdnd11an1n64x5 FILLER_24_1218 ();
 b15zdnd11an1n64x5 FILLER_24_1282 ();
 b15zdnd11an1n64x5 FILLER_24_1346 ();
 b15zdnd11an1n64x5 FILLER_24_1410 ();
 b15zdnd11an1n64x5 FILLER_24_1474 ();
 b15zdnd11an1n64x5 FILLER_24_1538 ();
 b15zdnd11an1n32x5 FILLER_24_1602 ();
 b15zdnd11an1n08x5 FILLER_24_1634 ();
 b15zdnd11an1n04x5 FILLER_24_1642 ();
 b15zdnd11an1n64x5 FILLER_24_1649 ();
 b15zdnd11an1n64x5 FILLER_24_1713 ();
 b15zdnd11an1n64x5 FILLER_24_1777 ();
 b15zdnd11an1n64x5 FILLER_24_1841 ();
 b15zdnd11an1n08x5 FILLER_24_1905 ();
 b15zdnd11an1n04x5 FILLER_24_1913 ();
 b15zdnd00an1n02x5 FILLER_24_1917 ();
 b15zdnd00an1n01x5 FILLER_24_1919 ();
 b15zdnd11an1n64x5 FILLER_24_1923 ();
 b15zdnd11an1n64x5 FILLER_24_1987 ();
 b15zdnd11an1n64x5 FILLER_24_2051 ();
 b15zdnd11an1n32x5 FILLER_24_2115 ();
 b15zdnd11an1n04x5 FILLER_24_2147 ();
 b15zdnd00an1n02x5 FILLER_24_2151 ();
 b15zdnd00an1n01x5 FILLER_24_2153 ();
 b15zdnd11an1n64x5 FILLER_24_2162 ();
 b15zdnd11an1n32x5 FILLER_24_2226 ();
 b15zdnd11an1n16x5 FILLER_24_2258 ();
 b15zdnd00an1n02x5 FILLER_24_2274 ();
 b15zdnd11an1n64x5 FILLER_25_0 ();
 b15zdnd11an1n64x5 FILLER_25_64 ();
 b15zdnd11an1n64x5 FILLER_25_128 ();
 b15zdnd11an1n64x5 FILLER_25_192 ();
 b15zdnd11an1n64x5 FILLER_25_256 ();
 b15zdnd11an1n64x5 FILLER_25_320 ();
 b15zdnd11an1n64x5 FILLER_25_384 ();
 b15zdnd11an1n64x5 FILLER_25_448 ();
 b15zdnd11an1n64x5 FILLER_25_512 ();
 b15zdnd11an1n64x5 FILLER_25_576 ();
 b15zdnd11an1n16x5 FILLER_25_640 ();
 b15zdnd11an1n08x5 FILLER_25_656 ();
 b15zdnd00an1n02x5 FILLER_25_664 ();
 b15zdnd11an1n64x5 FILLER_25_718 ();
 b15zdnd11an1n04x5 FILLER_25_782 ();
 b15zdnd00an1n01x5 FILLER_25_786 ();
 b15zdnd11an1n32x5 FILLER_25_818 ();
 b15zdnd11an1n16x5 FILLER_25_850 ();
 b15zdnd11an1n04x5 FILLER_25_866 ();
 b15zdnd00an1n02x5 FILLER_25_870 ();
 b15zdnd11an1n16x5 FILLER_25_880 ();
 b15zdnd11an1n08x5 FILLER_25_896 ();
 b15zdnd00an1n01x5 FILLER_25_904 ();
 b15zdnd11an1n32x5 FILLER_25_914 ();
 b15zdnd00an1n01x5 FILLER_25_946 ();
 b15zdnd11an1n64x5 FILLER_25_962 ();
 b15zdnd11an1n16x5 FILLER_25_1026 ();
 b15zdnd00an1n01x5 FILLER_25_1042 ();
 b15zdnd11an1n08x5 FILLER_25_1050 ();
 b15zdnd00an1n02x5 FILLER_25_1058 ();
 b15zdnd11an1n64x5 FILLER_25_1112 ();
 b15zdnd11an1n64x5 FILLER_25_1176 ();
 b15zdnd11an1n64x5 FILLER_25_1240 ();
 b15zdnd11an1n64x5 FILLER_25_1304 ();
 b15zdnd11an1n64x5 FILLER_25_1368 ();
 b15zdnd11an1n64x5 FILLER_25_1432 ();
 b15zdnd11an1n64x5 FILLER_25_1496 ();
 b15zdnd11an1n64x5 FILLER_25_1560 ();
 b15zdnd11an1n16x5 FILLER_25_1624 ();
 b15zdnd11an1n04x5 FILLER_25_1640 ();
 b15zdnd00an1n02x5 FILLER_25_1644 ();
 b15zdnd00an1n01x5 FILLER_25_1646 ();
 b15zdnd11an1n64x5 FILLER_25_1650 ();
 b15zdnd11an1n64x5 FILLER_25_1714 ();
 b15zdnd11an1n64x5 FILLER_25_1778 ();
 b15zdnd11an1n64x5 FILLER_25_1842 ();
 b15zdnd11an1n64x5 FILLER_25_1906 ();
 b15zdnd11an1n64x5 FILLER_25_1970 ();
 b15zdnd11an1n64x5 FILLER_25_2034 ();
 b15zdnd11an1n64x5 FILLER_25_2098 ();
 b15zdnd11an1n64x5 FILLER_25_2162 ();
 b15zdnd11an1n32x5 FILLER_25_2226 ();
 b15zdnd11an1n16x5 FILLER_25_2258 ();
 b15zdnd11an1n08x5 FILLER_25_2274 ();
 b15zdnd00an1n02x5 FILLER_25_2282 ();
 b15zdnd11an1n64x5 FILLER_26_8 ();
 b15zdnd11an1n64x5 FILLER_26_72 ();
 b15zdnd11an1n64x5 FILLER_26_136 ();
 b15zdnd11an1n64x5 FILLER_26_200 ();
 b15zdnd11an1n64x5 FILLER_26_264 ();
 b15zdnd11an1n64x5 FILLER_26_328 ();
 b15zdnd11an1n64x5 FILLER_26_392 ();
 b15zdnd11an1n64x5 FILLER_26_456 ();
 b15zdnd11an1n64x5 FILLER_26_520 ();
 b15zdnd11an1n64x5 FILLER_26_584 ();
 b15zdnd11an1n32x5 FILLER_26_648 ();
 b15zdnd00an1n02x5 FILLER_26_680 ();
 b15zdnd00an1n01x5 FILLER_26_682 ();
 b15zdnd11an1n04x5 FILLER_26_686 ();
 b15zdnd00an1n02x5 FILLER_26_690 ();
 b15zdnd11an1n08x5 FILLER_26_695 ();
 b15zdnd11an1n04x5 FILLER_26_703 ();
 b15zdnd00an1n02x5 FILLER_26_707 ();
 b15zdnd00an1n02x5 FILLER_26_716 ();
 b15zdnd11an1n64x5 FILLER_26_726 ();
 b15zdnd11an1n64x5 FILLER_26_790 ();
 b15zdnd11an1n32x5 FILLER_26_854 ();
 b15zdnd11an1n08x5 FILLER_26_886 ();
 b15zdnd00an1n02x5 FILLER_26_894 ();
 b15zdnd11an1n64x5 FILLER_26_938 ();
 b15zdnd11an1n64x5 FILLER_26_1002 ();
 b15zdnd11an1n08x5 FILLER_26_1066 ();
 b15zdnd11an1n04x5 FILLER_26_1074 ();
 b15zdnd00an1n01x5 FILLER_26_1078 ();
 b15zdnd11an1n04x5 FILLER_26_1082 ();
 b15zdnd11an1n04x5 FILLER_26_1089 ();
 b15zdnd00an1n02x5 FILLER_26_1093 ();
 b15zdnd11an1n04x5 FILLER_26_1102 ();
 b15zdnd11an1n64x5 FILLER_26_1148 ();
 b15zdnd11an1n64x5 FILLER_26_1212 ();
 b15zdnd11an1n64x5 FILLER_26_1276 ();
 b15zdnd11an1n64x5 FILLER_26_1340 ();
 b15zdnd11an1n64x5 FILLER_26_1404 ();
 b15zdnd11an1n64x5 FILLER_26_1468 ();
 b15zdnd11an1n64x5 FILLER_26_1532 ();
 b15zdnd11an1n64x5 FILLER_26_1596 ();
 b15zdnd11an1n64x5 FILLER_26_1660 ();
 b15zdnd11an1n64x5 FILLER_26_1724 ();
 b15zdnd11an1n64x5 FILLER_26_1788 ();
 b15zdnd11an1n64x5 FILLER_26_1852 ();
 b15zdnd11an1n64x5 FILLER_26_1916 ();
 b15zdnd11an1n64x5 FILLER_26_1980 ();
 b15zdnd11an1n64x5 FILLER_26_2044 ();
 b15zdnd11an1n32x5 FILLER_26_2108 ();
 b15zdnd11an1n08x5 FILLER_26_2140 ();
 b15zdnd11an1n04x5 FILLER_26_2148 ();
 b15zdnd00an1n02x5 FILLER_26_2152 ();
 b15zdnd11an1n64x5 FILLER_26_2162 ();
 b15zdnd11an1n32x5 FILLER_26_2226 ();
 b15zdnd11an1n16x5 FILLER_26_2258 ();
 b15zdnd00an1n02x5 FILLER_26_2274 ();
 b15zdnd11an1n64x5 FILLER_27_0 ();
 b15zdnd11an1n64x5 FILLER_27_64 ();
 b15zdnd11an1n64x5 FILLER_27_128 ();
 b15zdnd11an1n64x5 FILLER_27_192 ();
 b15zdnd11an1n64x5 FILLER_27_256 ();
 b15zdnd11an1n64x5 FILLER_27_320 ();
 b15zdnd11an1n08x5 FILLER_27_384 ();
 b15zdnd11an1n04x5 FILLER_27_392 ();
 b15zdnd00an1n02x5 FILLER_27_396 ();
 b15zdnd00an1n01x5 FILLER_27_398 ();
 b15zdnd11an1n04x5 FILLER_27_439 ();
 b15zdnd11an1n64x5 FILLER_27_446 ();
 b15zdnd11an1n64x5 FILLER_27_510 ();
 b15zdnd11an1n64x5 FILLER_27_574 ();
 b15zdnd11an1n04x5 FILLER_27_638 ();
 b15zdnd00an1n01x5 FILLER_27_642 ();
 b15zdnd11an1n64x5 FILLER_27_685 ();
 b15zdnd11an1n64x5 FILLER_27_749 ();
 b15zdnd11an1n64x5 FILLER_27_813 ();
 b15zdnd11an1n64x5 FILLER_27_877 ();
 b15zdnd11an1n16x5 FILLER_27_941 ();
 b15zdnd11an1n04x5 FILLER_27_957 ();
 b15zdnd00an1n02x5 FILLER_27_961 ();
 b15zdnd00an1n01x5 FILLER_27_963 ();
 b15zdnd11an1n64x5 FILLER_27_973 ();
 b15zdnd11an1n32x5 FILLER_27_1037 ();
 b15zdnd11an1n08x5 FILLER_27_1069 ();
 b15zdnd00an1n02x5 FILLER_27_1077 ();
 b15zdnd00an1n01x5 FILLER_27_1079 ();
 b15zdnd11an1n64x5 FILLER_27_1100 ();
 b15zdnd11an1n64x5 FILLER_27_1164 ();
 b15zdnd11an1n64x5 FILLER_27_1228 ();
 b15zdnd11an1n64x5 FILLER_27_1292 ();
 b15zdnd11an1n32x5 FILLER_27_1356 ();
 b15zdnd11an1n16x5 FILLER_27_1388 ();
 b15zdnd00an1n02x5 FILLER_27_1404 ();
 b15zdnd11an1n64x5 FILLER_27_1423 ();
 b15zdnd11an1n64x5 FILLER_27_1487 ();
 b15zdnd11an1n64x5 FILLER_27_1551 ();
 b15zdnd11an1n64x5 FILLER_27_1615 ();
 b15zdnd11an1n64x5 FILLER_27_1679 ();
 b15zdnd11an1n64x5 FILLER_27_1743 ();
 b15zdnd11an1n64x5 FILLER_27_1807 ();
 b15zdnd11an1n64x5 FILLER_27_1871 ();
 b15zdnd11an1n64x5 FILLER_27_1935 ();
 b15zdnd11an1n64x5 FILLER_27_1999 ();
 b15zdnd11an1n64x5 FILLER_27_2063 ();
 b15zdnd11an1n64x5 FILLER_27_2127 ();
 b15zdnd11an1n64x5 FILLER_27_2191 ();
 b15zdnd11an1n16x5 FILLER_27_2255 ();
 b15zdnd11an1n08x5 FILLER_27_2271 ();
 b15zdnd11an1n04x5 FILLER_27_2279 ();
 b15zdnd00an1n01x5 FILLER_27_2283 ();
 b15zdnd11an1n64x5 FILLER_28_8 ();
 b15zdnd11an1n64x5 FILLER_28_72 ();
 b15zdnd11an1n64x5 FILLER_28_136 ();
 b15zdnd11an1n32x5 FILLER_28_200 ();
 b15zdnd00an1n01x5 FILLER_28_232 ();
 b15zdnd11an1n04x5 FILLER_28_264 ();
 b15zdnd00an1n02x5 FILLER_28_268 ();
 b15zdnd00an1n01x5 FILLER_28_270 ();
 b15zdnd11an1n64x5 FILLER_28_302 ();
 b15zdnd11an1n64x5 FILLER_28_366 ();
 b15zdnd00an1n01x5 FILLER_28_430 ();
 b15zdnd11an1n64x5 FILLER_28_434 ();
 b15zdnd11an1n16x5 FILLER_28_498 ();
 b15zdnd11an1n08x5 FILLER_28_514 ();
 b15zdnd11an1n64x5 FILLER_28_525 ();
 b15zdnd11an1n64x5 FILLER_28_589 ();
 b15zdnd11an1n64x5 FILLER_28_653 ();
 b15zdnd00an1n01x5 FILLER_28_717 ();
 b15zdnd11an1n64x5 FILLER_28_726 ();
 b15zdnd11an1n32x5 FILLER_28_790 ();
 b15zdnd11an1n08x5 FILLER_28_822 ();
 b15zdnd11an1n64x5 FILLER_28_863 ();
 b15zdnd11an1n64x5 FILLER_28_927 ();
 b15zdnd11an1n64x5 FILLER_28_991 ();
 b15zdnd11an1n32x5 FILLER_28_1055 ();
 b15zdnd11an1n16x5 FILLER_28_1087 ();
 b15zdnd11an1n08x5 FILLER_28_1103 ();
 b15zdnd11an1n08x5 FILLER_28_1153 ();
 b15zdnd00an1n01x5 FILLER_28_1161 ();
 b15zdnd11an1n16x5 FILLER_28_1204 ();
 b15zdnd11an1n64x5 FILLER_28_1227 ();
 b15zdnd11an1n64x5 FILLER_28_1291 ();
 b15zdnd11an1n64x5 FILLER_28_1355 ();
 b15zdnd11an1n64x5 FILLER_28_1419 ();
 b15zdnd11an1n64x5 FILLER_28_1483 ();
 b15zdnd11an1n64x5 FILLER_28_1547 ();
 b15zdnd11an1n64x5 FILLER_28_1611 ();
 b15zdnd11an1n64x5 FILLER_28_1675 ();
 b15zdnd11an1n64x5 FILLER_28_1739 ();
 b15zdnd11an1n64x5 FILLER_28_1803 ();
 b15zdnd11an1n64x5 FILLER_28_1867 ();
 b15zdnd11an1n64x5 FILLER_28_1931 ();
 b15zdnd11an1n64x5 FILLER_28_1995 ();
 b15zdnd11an1n64x5 FILLER_28_2059 ();
 b15zdnd11an1n16x5 FILLER_28_2123 ();
 b15zdnd11an1n08x5 FILLER_28_2139 ();
 b15zdnd11an1n04x5 FILLER_28_2147 ();
 b15zdnd00an1n02x5 FILLER_28_2151 ();
 b15zdnd00an1n01x5 FILLER_28_2153 ();
 b15zdnd11an1n64x5 FILLER_28_2162 ();
 b15zdnd11an1n32x5 FILLER_28_2226 ();
 b15zdnd11an1n16x5 FILLER_28_2258 ();
 b15zdnd00an1n02x5 FILLER_28_2274 ();
 b15zdnd11an1n64x5 FILLER_29_0 ();
 b15zdnd11an1n64x5 FILLER_29_64 ();
 b15zdnd11an1n64x5 FILLER_29_128 ();
 b15zdnd11an1n64x5 FILLER_29_192 ();
 b15zdnd11an1n64x5 FILLER_29_256 ();
 b15zdnd11an1n64x5 FILLER_29_320 ();
 b15zdnd11an1n32x5 FILLER_29_384 ();
 b15zdnd00an1n01x5 FILLER_29_416 ();
 b15zdnd11an1n32x5 FILLER_29_448 ();
 b15zdnd11an1n16x5 FILLER_29_480 ();
 b15zdnd11an1n08x5 FILLER_29_496 ();
 b15zdnd11an1n04x5 FILLER_29_504 ();
 b15zdnd00an1n02x5 FILLER_29_508 ();
 b15zdnd00an1n01x5 FILLER_29_510 ();
 b15zdnd11an1n64x5 FILLER_29_553 ();
 b15zdnd11an1n64x5 FILLER_29_617 ();
 b15zdnd11an1n64x5 FILLER_29_681 ();
 b15zdnd11an1n64x5 FILLER_29_745 ();
 b15zdnd11an1n16x5 FILLER_29_809 ();
 b15zdnd11an1n08x5 FILLER_29_825 ();
 b15zdnd11an1n04x5 FILLER_29_836 ();
 b15zdnd11an1n64x5 FILLER_29_867 ();
 b15zdnd11an1n64x5 FILLER_29_931 ();
 b15zdnd11an1n64x5 FILLER_29_995 ();
 b15zdnd11an1n64x5 FILLER_29_1059 ();
 b15zdnd11an1n64x5 FILLER_29_1123 ();
 b15zdnd11an1n32x5 FILLER_29_1187 ();
 b15zdnd11an1n04x5 FILLER_29_1219 ();
 b15zdnd00an1n01x5 FILLER_29_1223 ();
 b15zdnd11an1n64x5 FILLER_29_1244 ();
 b15zdnd11an1n64x5 FILLER_29_1308 ();
 b15zdnd11an1n32x5 FILLER_29_1372 ();
 b15zdnd11an1n04x5 FILLER_29_1404 ();
 b15zdnd00an1n02x5 FILLER_29_1408 ();
 b15zdnd11an1n04x5 FILLER_29_1452 ();
 b15zdnd00an1n02x5 FILLER_29_1456 ();
 b15zdnd11an1n64x5 FILLER_29_1500 ();
 b15zdnd11an1n64x5 FILLER_29_1564 ();
 b15zdnd11an1n64x5 FILLER_29_1628 ();
 b15zdnd11an1n64x5 FILLER_29_1692 ();
 b15zdnd11an1n64x5 FILLER_29_1756 ();
 b15zdnd11an1n64x5 FILLER_29_1820 ();
 b15zdnd11an1n64x5 FILLER_29_1884 ();
 b15zdnd11an1n64x5 FILLER_29_1948 ();
 b15zdnd11an1n64x5 FILLER_29_2012 ();
 b15zdnd11an1n64x5 FILLER_29_2076 ();
 b15zdnd11an1n64x5 FILLER_29_2140 ();
 b15zdnd11an1n64x5 FILLER_29_2204 ();
 b15zdnd11an1n16x5 FILLER_29_2268 ();
 b15zdnd11an1n64x5 FILLER_30_8 ();
 b15zdnd11an1n64x5 FILLER_30_72 ();
 b15zdnd11an1n64x5 FILLER_30_136 ();
 b15zdnd11an1n64x5 FILLER_30_200 ();
 b15zdnd11an1n64x5 FILLER_30_264 ();
 b15zdnd11an1n64x5 FILLER_30_328 ();
 b15zdnd11an1n64x5 FILLER_30_392 ();
 b15zdnd11an1n32x5 FILLER_30_456 ();
 b15zdnd11an1n04x5 FILLER_30_488 ();
 b15zdnd00an1n02x5 FILLER_30_492 ();
 b15zdnd00an1n01x5 FILLER_30_494 ();
 b15zdnd11an1n64x5 FILLER_30_547 ();
 b15zdnd11an1n64x5 FILLER_30_611 ();
 b15zdnd11an1n32x5 FILLER_30_675 ();
 b15zdnd11an1n08x5 FILLER_30_707 ();
 b15zdnd00an1n02x5 FILLER_30_715 ();
 b15zdnd00an1n01x5 FILLER_30_717 ();
 b15zdnd11an1n64x5 FILLER_30_726 ();
 b15zdnd11an1n64x5 FILLER_30_790 ();
 b15zdnd11an1n64x5 FILLER_30_854 ();
 b15zdnd11an1n64x5 FILLER_30_918 ();
 b15zdnd11an1n64x5 FILLER_30_982 ();
 b15zdnd11an1n64x5 FILLER_30_1046 ();
 b15zdnd11an1n64x5 FILLER_30_1110 ();
 b15zdnd11an1n64x5 FILLER_30_1174 ();
 b15zdnd00an1n02x5 FILLER_30_1238 ();
 b15zdnd00an1n01x5 FILLER_30_1240 ();
 b15zdnd11an1n64x5 FILLER_30_1244 ();
 b15zdnd11an1n64x5 FILLER_30_1308 ();
 b15zdnd11an1n64x5 FILLER_30_1372 ();
 b15zdnd11an1n64x5 FILLER_30_1436 ();
 b15zdnd11an1n64x5 FILLER_30_1500 ();
 b15zdnd11an1n64x5 FILLER_30_1564 ();
 b15zdnd11an1n64x5 FILLER_30_1628 ();
 b15zdnd11an1n64x5 FILLER_30_1692 ();
 b15zdnd11an1n64x5 FILLER_30_1756 ();
 b15zdnd11an1n16x5 FILLER_30_1820 ();
 b15zdnd11an1n08x5 FILLER_30_1836 ();
 b15zdnd11an1n64x5 FILLER_30_1848 ();
 b15zdnd11an1n64x5 FILLER_30_1912 ();
 b15zdnd11an1n64x5 FILLER_30_1976 ();
 b15zdnd11an1n64x5 FILLER_30_2040 ();
 b15zdnd11an1n32x5 FILLER_30_2104 ();
 b15zdnd11an1n16x5 FILLER_30_2136 ();
 b15zdnd00an1n02x5 FILLER_30_2152 ();
 b15zdnd11an1n64x5 FILLER_30_2162 ();
 b15zdnd11an1n32x5 FILLER_30_2226 ();
 b15zdnd11an1n16x5 FILLER_30_2258 ();
 b15zdnd00an1n02x5 FILLER_30_2274 ();
 b15zdnd11an1n64x5 FILLER_31_0 ();
 b15zdnd11an1n64x5 FILLER_31_64 ();
 b15zdnd11an1n64x5 FILLER_31_128 ();
 b15zdnd11an1n16x5 FILLER_31_192 ();
 b15zdnd11an1n08x5 FILLER_31_208 ();
 b15zdnd11an1n04x5 FILLER_31_216 ();
 b15zdnd00an1n02x5 FILLER_31_220 ();
 b15zdnd00an1n01x5 FILLER_31_222 ();
 b15zdnd11an1n64x5 FILLER_31_248 ();
 b15zdnd11an1n64x5 FILLER_31_312 ();
 b15zdnd11an1n64x5 FILLER_31_376 ();
 b15zdnd11an1n16x5 FILLER_31_440 ();
 b15zdnd11an1n04x5 FILLER_31_456 ();
 b15zdnd00an1n02x5 FILLER_31_460 ();
 b15zdnd11an1n04x5 FILLER_31_482 ();
 b15zdnd11an1n16x5 FILLER_31_489 ();
 b15zdnd11an1n08x5 FILLER_31_505 ();
 b15zdnd11an1n04x5 FILLER_31_516 ();
 b15zdnd11an1n64x5 FILLER_31_523 ();
 b15zdnd11an1n64x5 FILLER_31_587 ();
 b15zdnd11an1n64x5 FILLER_31_651 ();
 b15zdnd11an1n64x5 FILLER_31_715 ();
 b15zdnd11an1n64x5 FILLER_31_779 ();
 b15zdnd11an1n32x5 FILLER_31_843 ();
 b15zdnd11an1n08x5 FILLER_31_875 ();
 b15zdnd11an1n04x5 FILLER_31_883 ();
 b15zdnd00an1n02x5 FILLER_31_887 ();
 b15zdnd00an1n01x5 FILLER_31_889 ();
 b15zdnd11an1n64x5 FILLER_31_932 ();
 b15zdnd11an1n64x5 FILLER_31_996 ();
 b15zdnd11an1n64x5 FILLER_31_1060 ();
 b15zdnd11an1n08x5 FILLER_31_1124 ();
 b15zdnd00an1n02x5 FILLER_31_1132 ();
 b15zdnd00an1n01x5 FILLER_31_1134 ();
 b15zdnd11an1n64x5 FILLER_31_1149 ();
 b15zdnd11an1n04x5 FILLER_31_1213 ();
 b15zdnd00an1n02x5 FILLER_31_1217 ();
 b15zdnd11an1n04x5 FILLER_31_1230 ();
 b15zdnd00an1n01x5 FILLER_31_1234 ();
 b15zdnd11an1n04x5 FILLER_31_1244 ();
 b15zdnd00an1n02x5 FILLER_31_1248 ();
 b15zdnd11an1n64x5 FILLER_31_1253 ();
 b15zdnd11an1n32x5 FILLER_31_1317 ();
 b15zdnd11an1n16x5 FILLER_31_1349 ();
 b15zdnd00an1n01x5 FILLER_31_1365 ();
 b15zdnd11an1n04x5 FILLER_31_1369 ();
 b15zdnd11an1n64x5 FILLER_31_1376 ();
 b15zdnd11an1n16x5 FILLER_31_1440 ();
 b15zdnd11an1n08x5 FILLER_31_1456 ();
 b15zdnd00an1n02x5 FILLER_31_1464 ();
 b15zdnd11an1n64x5 FILLER_31_1478 ();
 b15zdnd11an1n64x5 FILLER_31_1542 ();
 b15zdnd11an1n64x5 FILLER_31_1606 ();
 b15zdnd11an1n64x5 FILLER_31_1670 ();
 b15zdnd00an1n02x5 FILLER_31_1734 ();
 b15zdnd00an1n01x5 FILLER_31_1736 ();
 b15zdnd11an1n64x5 FILLER_31_1741 ();
 b15zdnd11an1n32x5 FILLER_31_1805 ();
 b15zdnd11an1n16x5 FILLER_31_1837 ();
 b15zdnd11an1n08x5 FILLER_31_1853 ();
 b15zdnd11an1n04x5 FILLER_31_1861 ();
 b15zdnd00an1n02x5 FILLER_31_1865 ();
 b15zdnd00an1n01x5 FILLER_31_1867 ();
 b15zdnd11an1n16x5 FILLER_31_1875 ();
 b15zdnd11an1n08x5 FILLER_31_1891 ();
 b15zdnd11an1n04x5 FILLER_31_1899 ();
 b15zdnd00an1n01x5 FILLER_31_1903 ();
 b15zdnd11an1n64x5 FILLER_31_1928 ();
 b15zdnd11an1n64x5 FILLER_31_1992 ();
 b15zdnd11an1n64x5 FILLER_31_2056 ();
 b15zdnd11an1n64x5 FILLER_31_2120 ();
 b15zdnd11an1n64x5 FILLER_31_2184 ();
 b15zdnd11an1n32x5 FILLER_31_2248 ();
 b15zdnd11an1n04x5 FILLER_31_2280 ();
 b15zdnd11an1n64x5 FILLER_32_8 ();
 b15zdnd11an1n64x5 FILLER_32_72 ();
 b15zdnd11an1n64x5 FILLER_32_136 ();
 b15zdnd11an1n64x5 FILLER_32_200 ();
 b15zdnd11an1n64x5 FILLER_32_264 ();
 b15zdnd11an1n64x5 FILLER_32_328 ();
 b15zdnd11an1n32x5 FILLER_32_392 ();
 b15zdnd11an1n16x5 FILLER_32_424 ();
 b15zdnd11an1n04x5 FILLER_32_440 ();
 b15zdnd00an1n02x5 FILLER_32_444 ();
 b15zdnd11an1n64x5 FILLER_32_453 ();
 b15zdnd11an1n64x5 FILLER_32_517 ();
 b15zdnd11an1n32x5 FILLER_32_581 ();
 b15zdnd11an1n16x5 FILLER_32_613 ();
 b15zdnd11an1n04x5 FILLER_32_629 ();
 b15zdnd00an1n01x5 FILLER_32_633 ();
 b15zdnd11an1n32x5 FILLER_32_659 ();
 b15zdnd11an1n16x5 FILLER_32_691 ();
 b15zdnd11an1n08x5 FILLER_32_707 ();
 b15zdnd00an1n02x5 FILLER_32_715 ();
 b15zdnd00an1n01x5 FILLER_32_717 ();
 b15zdnd11an1n64x5 FILLER_32_726 ();
 b15zdnd11an1n64x5 FILLER_32_790 ();
 b15zdnd11an1n16x5 FILLER_32_854 ();
 b15zdnd11an1n04x5 FILLER_32_870 ();
 b15zdnd11an1n64x5 FILLER_32_926 ();
 b15zdnd11an1n64x5 FILLER_32_990 ();
 b15zdnd11an1n64x5 FILLER_32_1054 ();
 b15zdnd11an1n64x5 FILLER_32_1118 ();
 b15zdnd11an1n32x5 FILLER_32_1182 ();
 b15zdnd11an1n04x5 FILLER_32_1214 ();
 b15zdnd00an1n01x5 FILLER_32_1218 ();
 b15zdnd11an1n64x5 FILLER_32_1263 ();
 b15zdnd11an1n16x5 FILLER_32_1327 ();
 b15zdnd11an1n04x5 FILLER_32_1343 ();
 b15zdnd00an1n01x5 FILLER_32_1347 ();
 b15zdnd11an1n64x5 FILLER_32_1400 ();
 b15zdnd11an1n64x5 FILLER_32_1464 ();
 b15zdnd11an1n64x5 FILLER_32_1528 ();
 b15zdnd11an1n32x5 FILLER_32_1592 ();
 b15zdnd11an1n16x5 FILLER_32_1624 ();
 b15zdnd11an1n04x5 FILLER_32_1640 ();
 b15zdnd11an1n64x5 FILLER_32_1652 ();
 b15zdnd11an1n64x5 FILLER_32_1716 ();
 b15zdnd11an1n64x5 FILLER_32_1780 ();
 b15zdnd11an1n64x5 FILLER_32_1844 ();
 b15zdnd11an1n08x5 FILLER_32_1908 ();
 b15zdnd11an1n04x5 FILLER_32_1916 ();
 b15zdnd11an1n64x5 FILLER_32_1927 ();
 b15zdnd11an1n64x5 FILLER_32_1991 ();
 b15zdnd11an1n64x5 FILLER_32_2055 ();
 b15zdnd11an1n32x5 FILLER_32_2119 ();
 b15zdnd00an1n02x5 FILLER_32_2151 ();
 b15zdnd00an1n01x5 FILLER_32_2153 ();
 b15zdnd11an1n64x5 FILLER_32_2162 ();
 b15zdnd11an1n32x5 FILLER_32_2226 ();
 b15zdnd11an1n16x5 FILLER_32_2258 ();
 b15zdnd00an1n02x5 FILLER_32_2274 ();
 b15zdnd11an1n64x5 FILLER_33_0 ();
 b15zdnd11an1n64x5 FILLER_33_64 ();
 b15zdnd11an1n64x5 FILLER_33_128 ();
 b15zdnd11an1n64x5 FILLER_33_192 ();
 b15zdnd11an1n64x5 FILLER_33_256 ();
 b15zdnd11an1n64x5 FILLER_33_320 ();
 b15zdnd11an1n64x5 FILLER_33_384 ();
 b15zdnd11an1n64x5 FILLER_33_448 ();
 b15zdnd11an1n64x5 FILLER_33_512 ();
 b15zdnd11an1n64x5 FILLER_33_576 ();
 b15zdnd11an1n16x5 FILLER_33_640 ();
 b15zdnd00an1n02x5 FILLER_33_656 ();
 b15zdnd11an1n64x5 FILLER_33_666 ();
 b15zdnd11an1n64x5 FILLER_33_730 ();
 b15zdnd11an1n64x5 FILLER_33_794 ();
 b15zdnd11an1n32x5 FILLER_33_858 ();
 b15zdnd00an1n02x5 FILLER_33_890 ();
 b15zdnd00an1n01x5 FILLER_33_892 ();
 b15zdnd11an1n04x5 FILLER_33_896 ();
 b15zdnd11an1n04x5 FILLER_33_903 ();
 b15zdnd11an1n64x5 FILLER_33_959 ();
 b15zdnd11an1n32x5 FILLER_33_1023 ();
 b15zdnd11an1n04x5 FILLER_33_1055 ();
 b15zdnd00an1n01x5 FILLER_33_1059 ();
 b15zdnd11an1n64x5 FILLER_33_1078 ();
 b15zdnd11an1n64x5 FILLER_33_1142 ();
 b15zdnd11an1n32x5 FILLER_33_1206 ();
 b15zdnd11an1n16x5 FILLER_33_1238 ();
 b15zdnd11an1n64x5 FILLER_33_1257 ();
 b15zdnd11an1n32x5 FILLER_33_1321 ();
 b15zdnd11an1n16x5 FILLER_33_1353 ();
 b15zdnd11an1n04x5 FILLER_33_1369 ();
 b15zdnd11an1n64x5 FILLER_33_1376 ();
 b15zdnd11an1n64x5 FILLER_33_1440 ();
 b15zdnd11an1n64x5 FILLER_33_1504 ();
 b15zdnd11an1n64x5 FILLER_33_1568 ();
 b15zdnd11an1n64x5 FILLER_33_1632 ();
 b15zdnd11an1n64x5 FILLER_33_1696 ();
 b15zdnd11an1n16x5 FILLER_33_1760 ();
 b15zdnd11an1n08x5 FILLER_33_1776 ();
 b15zdnd00an1n01x5 FILLER_33_1784 ();
 b15zdnd11an1n08x5 FILLER_33_1827 ();
 b15zdnd00an1n01x5 FILLER_33_1835 ();
 b15zdnd11an1n08x5 FILLER_33_1840 ();
 b15zdnd00an1n02x5 FILLER_33_1848 ();
 b15zdnd11an1n64x5 FILLER_33_1854 ();
 b15zdnd11an1n32x5 FILLER_33_1918 ();
 b15zdnd11an1n16x5 FILLER_33_1950 ();
 b15zdnd11an1n64x5 FILLER_33_1983 ();
 b15zdnd11an1n64x5 FILLER_33_2047 ();
 b15zdnd11an1n64x5 FILLER_33_2111 ();
 b15zdnd11an1n64x5 FILLER_33_2175 ();
 b15zdnd11an1n32x5 FILLER_33_2239 ();
 b15zdnd11an1n08x5 FILLER_33_2271 ();
 b15zdnd11an1n04x5 FILLER_33_2279 ();
 b15zdnd00an1n01x5 FILLER_33_2283 ();
 b15zdnd11an1n64x5 FILLER_34_8 ();
 b15zdnd11an1n64x5 FILLER_34_72 ();
 b15zdnd11an1n64x5 FILLER_34_136 ();
 b15zdnd11an1n64x5 FILLER_34_200 ();
 b15zdnd11an1n64x5 FILLER_34_264 ();
 b15zdnd11an1n64x5 FILLER_34_328 ();
 b15zdnd11an1n64x5 FILLER_34_392 ();
 b15zdnd11an1n64x5 FILLER_34_456 ();
 b15zdnd11an1n16x5 FILLER_34_520 ();
 b15zdnd00an1n01x5 FILLER_34_536 ();
 b15zdnd11an1n64x5 FILLER_34_541 ();
 b15zdnd11an1n32x5 FILLER_34_605 ();
 b15zdnd11an1n16x5 FILLER_34_637 ();
 b15zdnd11an1n08x5 FILLER_34_653 ();
 b15zdnd11an1n32x5 FILLER_34_664 ();
 b15zdnd11an1n16x5 FILLER_34_696 ();
 b15zdnd11an1n04x5 FILLER_34_712 ();
 b15zdnd00an1n02x5 FILLER_34_716 ();
 b15zdnd11an1n08x5 FILLER_34_726 ();
 b15zdnd11an1n04x5 FILLER_34_734 ();
 b15zdnd00an1n02x5 FILLER_34_738 ();
 b15zdnd00an1n01x5 FILLER_34_740 ();
 b15zdnd11an1n64x5 FILLER_34_753 ();
 b15zdnd11an1n64x5 FILLER_34_817 ();
 b15zdnd11an1n16x5 FILLER_34_881 ();
 b15zdnd00an1n02x5 FILLER_34_897 ();
 b15zdnd00an1n01x5 FILLER_34_899 ();
 b15zdnd11an1n16x5 FILLER_34_903 ();
 b15zdnd11an1n08x5 FILLER_34_919 ();
 b15zdnd00an1n02x5 FILLER_34_927 ();
 b15zdnd00an1n01x5 FILLER_34_929 ();
 b15zdnd11an1n04x5 FILLER_34_933 ();
 b15zdnd11an1n04x5 FILLER_34_940 ();
 b15zdnd11an1n64x5 FILLER_34_947 ();
 b15zdnd11an1n08x5 FILLER_34_1011 ();
 b15zdnd00an1n01x5 FILLER_34_1019 ();
 b15zdnd11an1n64x5 FILLER_34_1040 ();
 b15zdnd11an1n64x5 FILLER_34_1104 ();
 b15zdnd11an1n64x5 FILLER_34_1168 ();
 b15zdnd11an1n64x5 FILLER_34_1232 ();
 b15zdnd11an1n64x5 FILLER_34_1296 ();
 b15zdnd11an1n64x5 FILLER_34_1360 ();
 b15zdnd11an1n16x5 FILLER_34_1424 ();
 b15zdnd11an1n04x5 FILLER_34_1440 ();
 b15zdnd11an1n64x5 FILLER_34_1461 ();
 b15zdnd11an1n64x5 FILLER_34_1525 ();
 b15zdnd11an1n64x5 FILLER_34_1589 ();
 b15zdnd11an1n64x5 FILLER_34_1653 ();
 b15zdnd11an1n64x5 FILLER_34_1717 ();
 b15zdnd11an1n64x5 FILLER_34_1781 ();
 b15zdnd11an1n64x5 FILLER_34_1845 ();
 b15zdnd11an1n64x5 FILLER_34_1909 ();
 b15zdnd11an1n64x5 FILLER_34_1973 ();
 b15zdnd11an1n08x5 FILLER_34_2037 ();
 b15zdnd00an1n02x5 FILLER_34_2045 ();
 b15zdnd00an1n01x5 FILLER_34_2047 ();
 b15zdnd11an1n64x5 FILLER_34_2055 ();
 b15zdnd11an1n32x5 FILLER_34_2119 ();
 b15zdnd00an1n02x5 FILLER_34_2151 ();
 b15zdnd00an1n01x5 FILLER_34_2153 ();
 b15zdnd11an1n64x5 FILLER_34_2162 ();
 b15zdnd11an1n32x5 FILLER_34_2226 ();
 b15zdnd11an1n16x5 FILLER_34_2258 ();
 b15zdnd00an1n02x5 FILLER_34_2274 ();
 b15zdnd11an1n64x5 FILLER_35_0 ();
 b15zdnd11an1n64x5 FILLER_35_64 ();
 b15zdnd11an1n64x5 FILLER_35_128 ();
 b15zdnd11an1n64x5 FILLER_35_192 ();
 b15zdnd11an1n64x5 FILLER_35_256 ();
 b15zdnd11an1n32x5 FILLER_35_320 ();
 b15zdnd11an1n04x5 FILLER_35_352 ();
 b15zdnd00an1n01x5 FILLER_35_356 ();
 b15zdnd11an1n64x5 FILLER_35_388 ();
 b15zdnd11an1n64x5 FILLER_35_452 ();
 b15zdnd11an1n64x5 FILLER_35_516 ();
 b15zdnd11an1n32x5 FILLER_35_580 ();
 b15zdnd11an1n16x5 FILLER_35_612 ();
 b15zdnd11an1n04x5 FILLER_35_628 ();
 b15zdnd00an1n02x5 FILLER_35_632 ();
 b15zdnd11an1n64x5 FILLER_35_686 ();
 b15zdnd11an1n64x5 FILLER_35_750 ();
 b15zdnd11an1n64x5 FILLER_35_814 ();
 b15zdnd11an1n32x5 FILLER_35_878 ();
 b15zdnd00an1n02x5 FILLER_35_910 ();
 b15zdnd00an1n01x5 FILLER_35_912 ();
 b15zdnd11an1n32x5 FILLER_35_937 ();
 b15zdnd11an1n16x5 FILLER_35_969 ();
 b15zdnd00an1n02x5 FILLER_35_985 ();
 b15zdnd00an1n01x5 FILLER_35_987 ();
 b15zdnd11an1n64x5 FILLER_35_1030 ();
 b15zdnd11an1n64x5 FILLER_35_1094 ();
 b15zdnd11an1n64x5 FILLER_35_1158 ();
 b15zdnd11an1n64x5 FILLER_35_1222 ();
 b15zdnd11an1n64x5 FILLER_35_1286 ();
 b15zdnd11an1n64x5 FILLER_35_1350 ();
 b15zdnd11an1n32x5 FILLER_35_1414 ();
 b15zdnd11an1n04x5 FILLER_35_1446 ();
 b15zdnd11an1n64x5 FILLER_35_1462 ();
 b15zdnd11an1n64x5 FILLER_35_1526 ();
 b15zdnd11an1n64x5 FILLER_35_1590 ();
 b15zdnd11an1n64x5 FILLER_35_1654 ();
 b15zdnd11an1n64x5 FILLER_35_1718 ();
 b15zdnd11an1n64x5 FILLER_35_1782 ();
 b15zdnd11an1n64x5 FILLER_35_1846 ();
 b15zdnd11an1n64x5 FILLER_35_1910 ();
 b15zdnd11an1n64x5 FILLER_35_1974 ();
 b15zdnd11an1n16x5 FILLER_35_2038 ();
 b15zdnd11an1n04x5 FILLER_35_2054 ();
 b15zdnd00an1n02x5 FILLER_35_2058 ();
 b15zdnd11an1n64x5 FILLER_35_2074 ();
 b15zdnd11an1n64x5 FILLER_35_2138 ();
 b15zdnd11an1n64x5 FILLER_35_2202 ();
 b15zdnd11an1n16x5 FILLER_35_2266 ();
 b15zdnd00an1n02x5 FILLER_35_2282 ();
 b15zdnd11an1n64x5 FILLER_36_8 ();
 b15zdnd11an1n64x5 FILLER_36_72 ();
 b15zdnd11an1n64x5 FILLER_36_136 ();
 b15zdnd11an1n64x5 FILLER_36_200 ();
 b15zdnd11an1n64x5 FILLER_36_264 ();
 b15zdnd11an1n32x5 FILLER_36_328 ();
 b15zdnd11an1n64x5 FILLER_36_378 ();
 b15zdnd11an1n64x5 FILLER_36_442 ();
 b15zdnd11an1n64x5 FILLER_36_506 ();
 b15zdnd11an1n08x5 FILLER_36_570 ();
 b15zdnd11an1n04x5 FILLER_36_578 ();
 b15zdnd11an1n04x5 FILLER_36_624 ();
 b15zdnd00an1n01x5 FILLER_36_628 ();
 b15zdnd11an1n32x5 FILLER_36_671 ();
 b15zdnd11an1n08x5 FILLER_36_703 ();
 b15zdnd11an1n04x5 FILLER_36_711 ();
 b15zdnd00an1n02x5 FILLER_36_715 ();
 b15zdnd00an1n01x5 FILLER_36_717 ();
 b15zdnd11an1n64x5 FILLER_36_726 ();
 b15zdnd11an1n64x5 FILLER_36_790 ();
 b15zdnd11an1n08x5 FILLER_36_854 ();
 b15zdnd11an1n04x5 FILLER_36_862 ();
 b15zdnd11an1n64x5 FILLER_36_874 ();
 b15zdnd11an1n32x5 FILLER_36_938 ();
 b15zdnd11an1n16x5 FILLER_36_970 ();
 b15zdnd11an1n08x5 FILLER_36_986 ();
 b15zdnd00an1n01x5 FILLER_36_994 ();
 b15zdnd11an1n64x5 FILLER_36_998 ();
 b15zdnd11an1n32x5 FILLER_36_1062 ();
 b15zdnd11an1n16x5 FILLER_36_1094 ();
 b15zdnd00an1n02x5 FILLER_36_1110 ();
 b15zdnd11an1n32x5 FILLER_36_1164 ();
 b15zdnd11an1n16x5 FILLER_36_1196 ();
 b15zdnd11an1n08x5 FILLER_36_1212 ();
 b15zdnd11an1n64x5 FILLER_36_1223 ();
 b15zdnd11an1n64x5 FILLER_36_1287 ();
 b15zdnd11an1n64x5 FILLER_36_1351 ();
 b15zdnd11an1n64x5 FILLER_36_1415 ();
 b15zdnd11an1n64x5 FILLER_36_1479 ();
 b15zdnd11an1n64x5 FILLER_36_1543 ();
 b15zdnd11an1n64x5 FILLER_36_1607 ();
 b15zdnd11an1n64x5 FILLER_36_1671 ();
 b15zdnd11an1n64x5 FILLER_36_1735 ();
 b15zdnd11an1n64x5 FILLER_36_1799 ();
 b15zdnd11an1n64x5 FILLER_36_1863 ();
 b15zdnd11an1n16x5 FILLER_36_1927 ();
 b15zdnd11an1n08x5 FILLER_36_1943 ();
 b15zdnd11an1n64x5 FILLER_36_1993 ();
 b15zdnd00an1n02x5 FILLER_36_2057 ();
 b15zdnd00an1n01x5 FILLER_36_2059 ();
 b15zdnd11an1n04x5 FILLER_36_2080 ();
 b15zdnd11an1n32x5 FILLER_36_2095 ();
 b15zdnd11an1n16x5 FILLER_36_2127 ();
 b15zdnd11an1n08x5 FILLER_36_2143 ();
 b15zdnd00an1n02x5 FILLER_36_2151 ();
 b15zdnd00an1n01x5 FILLER_36_2153 ();
 b15zdnd11an1n64x5 FILLER_36_2162 ();
 b15zdnd11an1n32x5 FILLER_36_2226 ();
 b15zdnd11an1n16x5 FILLER_36_2258 ();
 b15zdnd00an1n02x5 FILLER_36_2274 ();
 b15zdnd11an1n64x5 FILLER_37_0 ();
 b15zdnd11an1n64x5 FILLER_37_64 ();
 b15zdnd11an1n64x5 FILLER_37_128 ();
 b15zdnd11an1n64x5 FILLER_37_192 ();
 b15zdnd11an1n64x5 FILLER_37_256 ();
 b15zdnd11an1n16x5 FILLER_37_320 ();
 b15zdnd11an1n08x5 FILLER_37_336 ();
 b15zdnd00an1n02x5 FILLER_37_344 ();
 b15zdnd11an1n64x5 FILLER_37_349 ();
 b15zdnd11an1n32x5 FILLER_37_413 ();
 b15zdnd11an1n16x5 FILLER_37_445 ();
 b15zdnd11an1n08x5 FILLER_37_461 ();
 b15zdnd11an1n04x5 FILLER_37_469 ();
 b15zdnd00an1n02x5 FILLER_37_473 ();
 b15zdnd11an1n64x5 FILLER_37_492 ();
 b15zdnd11an1n32x5 FILLER_37_556 ();
 b15zdnd11an1n04x5 FILLER_37_588 ();
 b15zdnd00an1n02x5 FILLER_37_592 ();
 b15zdnd00an1n01x5 FILLER_37_594 ();
 b15zdnd11an1n32x5 FILLER_37_600 ();
 b15zdnd11an1n16x5 FILLER_37_632 ();
 b15zdnd11an1n04x5 FILLER_37_648 ();
 b15zdnd11an1n04x5 FILLER_37_655 ();
 b15zdnd11an1n64x5 FILLER_37_662 ();
 b15zdnd11an1n64x5 FILLER_37_726 ();
 b15zdnd11an1n08x5 FILLER_37_790 ();
 b15zdnd11an1n04x5 FILLER_37_798 ();
 b15zdnd00an1n02x5 FILLER_37_802 ();
 b15zdnd00an1n01x5 FILLER_37_804 ();
 b15zdnd11an1n64x5 FILLER_37_857 ();
 b15zdnd11an1n32x5 FILLER_37_921 ();
 b15zdnd11an1n08x5 FILLER_37_953 ();
 b15zdnd11an1n04x5 FILLER_37_961 ();
 b15zdnd00an1n02x5 FILLER_37_965 ();
 b15zdnd00an1n01x5 FILLER_37_967 ();
 b15zdnd11an1n64x5 FILLER_37_1020 ();
 b15zdnd11an1n32x5 FILLER_37_1084 ();
 b15zdnd11an1n16x5 FILLER_37_1116 ();
 b15zdnd11an1n04x5 FILLER_37_1135 ();
 b15zdnd11an1n64x5 FILLER_37_1142 ();
 b15zdnd11an1n32x5 FILLER_37_1206 ();
 b15zdnd11an1n08x5 FILLER_37_1238 ();
 b15zdnd11an1n04x5 FILLER_37_1249 ();
 b15zdnd11an1n64x5 FILLER_37_1256 ();
 b15zdnd11an1n64x5 FILLER_37_1320 ();
 b15zdnd11an1n32x5 FILLER_37_1384 ();
 b15zdnd11an1n08x5 FILLER_37_1416 ();
 b15zdnd11an1n04x5 FILLER_37_1424 ();
 b15zdnd00an1n02x5 FILLER_37_1428 ();
 b15zdnd11an1n64x5 FILLER_37_1433 ();
 b15zdnd11an1n64x5 FILLER_37_1497 ();
 b15zdnd11an1n64x5 FILLER_37_1561 ();
 b15zdnd11an1n64x5 FILLER_37_1625 ();
 b15zdnd11an1n64x5 FILLER_37_1689 ();
 b15zdnd11an1n64x5 FILLER_37_1753 ();
 b15zdnd11an1n64x5 FILLER_37_1817 ();
 b15zdnd11an1n64x5 FILLER_37_1881 ();
 b15zdnd11an1n64x5 FILLER_37_1945 ();
 b15zdnd11an1n64x5 FILLER_37_2009 ();
 b15zdnd11an1n64x5 FILLER_37_2073 ();
 b15zdnd11an1n64x5 FILLER_37_2137 ();
 b15zdnd11an1n64x5 FILLER_37_2201 ();
 b15zdnd11an1n16x5 FILLER_37_2265 ();
 b15zdnd00an1n02x5 FILLER_37_2281 ();
 b15zdnd00an1n01x5 FILLER_37_2283 ();
 b15zdnd11an1n64x5 FILLER_38_8 ();
 b15zdnd11an1n64x5 FILLER_38_72 ();
 b15zdnd11an1n64x5 FILLER_38_136 ();
 b15zdnd11an1n16x5 FILLER_38_200 ();
 b15zdnd00an1n02x5 FILLER_38_216 ();
 b15zdnd11an1n04x5 FILLER_38_221 ();
 b15zdnd11an1n16x5 FILLER_38_228 ();
 b15zdnd00an1n02x5 FILLER_38_244 ();
 b15zdnd11an1n32x5 FILLER_38_266 ();
 b15zdnd11an1n16x5 FILLER_38_298 ();
 b15zdnd11an1n04x5 FILLER_38_314 ();
 b15zdnd00an1n01x5 FILLER_38_318 ();
 b15zdnd11an1n64x5 FILLER_38_371 ();
 b15zdnd11an1n64x5 FILLER_38_435 ();
 b15zdnd11an1n64x5 FILLER_38_499 ();
 b15zdnd11an1n04x5 FILLER_38_563 ();
 b15zdnd11an1n64x5 FILLER_38_598 ();
 b15zdnd11an1n32x5 FILLER_38_662 ();
 b15zdnd11an1n16x5 FILLER_38_694 ();
 b15zdnd11an1n08x5 FILLER_38_710 ();
 b15zdnd11an1n64x5 FILLER_38_726 ();
 b15zdnd11an1n32x5 FILLER_38_790 ();
 b15zdnd00an1n02x5 FILLER_38_822 ();
 b15zdnd00an1n01x5 FILLER_38_824 ();
 b15zdnd11an1n04x5 FILLER_38_828 ();
 b15zdnd11an1n16x5 FILLER_38_835 ();
 b15zdnd00an1n01x5 FILLER_38_851 ();
 b15zdnd11an1n64x5 FILLER_38_894 ();
 b15zdnd11an1n16x5 FILLER_38_958 ();
 b15zdnd11an1n08x5 FILLER_38_974 ();
 b15zdnd00an1n02x5 FILLER_38_982 ();
 b15zdnd11an1n04x5 FILLER_38_987 ();
 b15zdnd00an1n02x5 FILLER_38_991 ();
 b15zdnd00an1n01x5 FILLER_38_993 ();
 b15zdnd11an1n04x5 FILLER_38_997 ();
 b15zdnd00an1n01x5 FILLER_38_1001 ();
 b15zdnd11an1n04x5 FILLER_38_1009 ();
 b15zdnd11an1n64x5 FILLER_38_1055 ();
 b15zdnd11an1n16x5 FILLER_38_1119 ();
 b15zdnd00an1n02x5 FILLER_38_1135 ();
 b15zdnd00an1n01x5 FILLER_38_1137 ();
 b15zdnd11an1n64x5 FILLER_38_1141 ();
 b15zdnd11an1n16x5 FILLER_38_1205 ();
 b15zdnd11an1n04x5 FILLER_38_1221 ();
 b15zdnd00an1n02x5 FILLER_38_1225 ();
 b15zdnd11an1n64x5 FILLER_38_1279 ();
 b15zdnd11an1n64x5 FILLER_38_1343 ();
 b15zdnd11an1n64x5 FILLER_38_1459 ();
 b15zdnd11an1n16x5 FILLER_38_1523 ();
 b15zdnd11an1n08x5 FILLER_38_1539 ();
 b15zdnd11an1n04x5 FILLER_38_1547 ();
 b15zdnd00an1n02x5 FILLER_38_1551 ();
 b15zdnd00an1n01x5 FILLER_38_1553 ();
 b15zdnd11an1n32x5 FILLER_38_1606 ();
 b15zdnd11an1n16x5 FILLER_38_1638 ();
 b15zdnd11an1n04x5 FILLER_38_1654 ();
 b15zdnd00an1n02x5 FILLER_38_1658 ();
 b15zdnd00an1n01x5 FILLER_38_1660 ();
 b15zdnd11an1n64x5 FILLER_38_1669 ();
 b15zdnd11an1n64x5 FILLER_38_1733 ();
 b15zdnd11an1n64x5 FILLER_38_1797 ();
 b15zdnd11an1n64x5 FILLER_38_1861 ();
 b15zdnd11an1n32x5 FILLER_38_1925 ();
 b15zdnd11an1n16x5 FILLER_38_1957 ();
 b15zdnd11an1n04x5 FILLER_38_1973 ();
 b15zdnd00an1n02x5 FILLER_38_1977 ();
 b15zdnd11an1n64x5 FILLER_38_2031 ();
 b15zdnd11an1n32x5 FILLER_38_2095 ();
 b15zdnd11an1n16x5 FILLER_38_2127 ();
 b15zdnd11an1n08x5 FILLER_38_2143 ();
 b15zdnd00an1n02x5 FILLER_38_2151 ();
 b15zdnd00an1n01x5 FILLER_38_2153 ();
 b15zdnd11an1n64x5 FILLER_38_2162 ();
 b15zdnd11an1n32x5 FILLER_38_2226 ();
 b15zdnd11an1n16x5 FILLER_38_2258 ();
 b15zdnd00an1n02x5 FILLER_38_2274 ();
 b15zdnd11an1n64x5 FILLER_39_0 ();
 b15zdnd11an1n64x5 FILLER_39_64 ();
 b15zdnd11an1n64x5 FILLER_39_128 ();
 b15zdnd11an1n04x5 FILLER_39_192 ();
 b15zdnd00an1n02x5 FILLER_39_196 ();
 b15zdnd00an1n01x5 FILLER_39_198 ();
 b15zdnd11an1n64x5 FILLER_39_251 ();
 b15zdnd11an1n16x5 FILLER_39_315 ();
 b15zdnd11an1n04x5 FILLER_39_331 ();
 b15zdnd00an1n02x5 FILLER_39_335 ();
 b15zdnd11an1n04x5 FILLER_39_340 ();
 b15zdnd11an1n64x5 FILLER_39_347 ();
 b15zdnd11an1n64x5 FILLER_39_411 ();
 b15zdnd11an1n64x5 FILLER_39_475 ();
 b15zdnd11an1n32x5 FILLER_39_539 ();
 b15zdnd11an1n16x5 FILLER_39_571 ();
 b15zdnd11an1n08x5 FILLER_39_587 ();
 b15zdnd11an1n04x5 FILLER_39_595 ();
 b15zdnd00an1n01x5 FILLER_39_599 ();
 b15zdnd11an1n64x5 FILLER_39_625 ();
 b15zdnd11an1n64x5 FILLER_39_689 ();
 b15zdnd11an1n64x5 FILLER_39_753 ();
 b15zdnd11an1n08x5 FILLER_39_817 ();
 b15zdnd11an1n16x5 FILLER_39_828 ();
 b15zdnd11an1n04x5 FILLER_39_844 ();
 b15zdnd11an1n32x5 FILLER_39_855 ();
 b15zdnd11an1n08x5 FILLER_39_887 ();
 b15zdnd11an1n04x5 FILLER_39_895 ();
 b15zdnd00an1n02x5 FILLER_39_899 ();
 b15zdnd11an1n64x5 FILLER_39_943 ();
 b15zdnd11an1n32x5 FILLER_39_1007 ();
 b15zdnd00an1n02x5 FILLER_39_1039 ();
 b15zdnd11an1n04x5 FILLER_39_1044 ();
 b15zdnd11an1n64x5 FILLER_39_1051 ();
 b15zdnd11an1n64x5 FILLER_39_1115 ();
 b15zdnd11an1n64x5 FILLER_39_1179 ();
 b15zdnd11an1n04x5 FILLER_39_1243 ();
 b15zdnd00an1n02x5 FILLER_39_1247 ();
 b15zdnd11an1n64x5 FILLER_39_1252 ();
 b15zdnd11an1n64x5 FILLER_39_1316 ();
 b15zdnd11an1n32x5 FILLER_39_1380 ();
 b15zdnd11an1n16x5 FILLER_39_1412 ();
 b15zdnd11an1n04x5 FILLER_39_1431 ();
 b15zdnd11an1n64x5 FILLER_39_1438 ();
 b15zdnd11an1n64x5 FILLER_39_1502 ();
 b15zdnd11an1n04x5 FILLER_39_1566 ();
 b15zdnd00an1n02x5 FILLER_39_1570 ();
 b15zdnd00an1n01x5 FILLER_39_1572 ();
 b15zdnd11an1n04x5 FILLER_39_1576 ();
 b15zdnd11an1n04x5 FILLER_39_1583 ();
 b15zdnd11an1n64x5 FILLER_39_1590 ();
 b15zdnd11an1n32x5 FILLER_39_1654 ();
 b15zdnd11an1n16x5 FILLER_39_1686 ();
 b15zdnd11an1n04x5 FILLER_39_1702 ();
 b15zdnd00an1n02x5 FILLER_39_1706 ();
 b15zdnd11an1n04x5 FILLER_39_1711 ();
 b15zdnd11an1n64x5 FILLER_39_1718 ();
 b15zdnd11an1n64x5 FILLER_39_1782 ();
 b15zdnd11an1n64x5 FILLER_39_1846 ();
 b15zdnd11an1n64x5 FILLER_39_1910 ();
 b15zdnd11an1n16x5 FILLER_39_1974 ();
 b15zdnd11an1n08x5 FILLER_39_1990 ();
 b15zdnd11an1n04x5 FILLER_39_1998 ();
 b15zdnd00an1n02x5 FILLER_39_2002 ();
 b15zdnd11an1n04x5 FILLER_39_2007 ();
 b15zdnd11an1n64x5 FILLER_39_2014 ();
 b15zdnd11an1n64x5 FILLER_39_2078 ();
 b15zdnd11an1n64x5 FILLER_39_2142 ();
 b15zdnd11an1n64x5 FILLER_39_2206 ();
 b15zdnd11an1n08x5 FILLER_39_2270 ();
 b15zdnd11an1n04x5 FILLER_39_2278 ();
 b15zdnd00an1n02x5 FILLER_39_2282 ();
 b15zdnd11an1n64x5 FILLER_40_8 ();
 b15zdnd11an1n64x5 FILLER_40_72 ();
 b15zdnd11an1n64x5 FILLER_40_136 ();
 b15zdnd11an1n16x5 FILLER_40_200 ();
 b15zdnd11an1n04x5 FILLER_40_216 ();
 b15zdnd00an1n01x5 FILLER_40_220 ();
 b15zdnd11an1n16x5 FILLER_40_224 ();
 b15zdnd00an1n02x5 FILLER_40_240 ();
 b15zdnd00an1n01x5 FILLER_40_242 ();
 b15zdnd11an1n04x5 FILLER_40_269 ();
 b15zdnd11an1n64x5 FILLER_40_287 ();
 b15zdnd11an1n64x5 FILLER_40_351 ();
 b15zdnd11an1n16x5 FILLER_40_415 ();
 b15zdnd00an1n02x5 FILLER_40_431 ();
 b15zdnd00an1n01x5 FILLER_40_433 ();
 b15zdnd11an1n04x5 FILLER_40_438 ();
 b15zdnd11an1n64x5 FILLER_40_449 ();
 b15zdnd11an1n64x5 FILLER_40_513 ();
 b15zdnd11an1n64x5 FILLER_40_577 ();
 b15zdnd11an1n64x5 FILLER_40_641 ();
 b15zdnd11an1n08x5 FILLER_40_705 ();
 b15zdnd11an1n04x5 FILLER_40_713 ();
 b15zdnd00an1n01x5 FILLER_40_717 ();
 b15zdnd11an1n64x5 FILLER_40_726 ();
 b15zdnd11an1n32x5 FILLER_40_790 ();
 b15zdnd11an1n16x5 FILLER_40_822 ();
 b15zdnd11an1n08x5 FILLER_40_838 ();
 b15zdnd00an1n02x5 FILLER_40_846 ();
 b15zdnd11an1n32x5 FILLER_40_851 ();
 b15zdnd11an1n04x5 FILLER_40_883 ();
 b15zdnd11an1n64x5 FILLER_40_929 ();
 b15zdnd11an1n32x5 FILLER_40_993 ();
 b15zdnd00an1n02x5 FILLER_40_1025 ();
 b15zdnd11an1n64x5 FILLER_40_1071 ();
 b15zdnd11an1n32x5 FILLER_40_1135 ();
 b15zdnd11an1n16x5 FILLER_40_1167 ();
 b15zdnd11an1n08x5 FILLER_40_1183 ();
 b15zdnd11an1n04x5 FILLER_40_1191 ();
 b15zdnd00an1n02x5 FILLER_40_1195 ();
 b15zdnd11an1n04x5 FILLER_40_1218 ();
 b15zdnd11an1n64x5 FILLER_40_1232 ();
 b15zdnd11an1n32x5 FILLER_40_1296 ();
 b15zdnd11an1n16x5 FILLER_40_1328 ();
 b15zdnd11an1n04x5 FILLER_40_1344 ();
 b15zdnd11an1n64x5 FILLER_40_1354 ();
 b15zdnd11an1n64x5 FILLER_40_1418 ();
 b15zdnd11an1n08x5 FILLER_40_1482 ();
 b15zdnd11an1n04x5 FILLER_40_1490 ();
 b15zdnd00an1n01x5 FILLER_40_1494 ();
 b15zdnd11an1n64x5 FILLER_40_1502 ();
 b15zdnd11an1n64x5 FILLER_40_1566 ();
 b15zdnd11an1n32x5 FILLER_40_1630 ();
 b15zdnd11an1n16x5 FILLER_40_1662 ();
 b15zdnd11an1n08x5 FILLER_40_1678 ();
 b15zdnd11an1n04x5 FILLER_40_1686 ();
 b15zdnd11an1n64x5 FILLER_40_1742 ();
 b15zdnd11an1n64x5 FILLER_40_1806 ();
 b15zdnd11an1n64x5 FILLER_40_1870 ();
 b15zdnd11an1n64x5 FILLER_40_1934 ();
 b15zdnd11an1n04x5 FILLER_40_1998 ();
 b15zdnd00an1n02x5 FILLER_40_2002 ();
 b15zdnd00an1n01x5 FILLER_40_2004 ();
 b15zdnd11an1n64x5 FILLER_40_2008 ();
 b15zdnd11an1n64x5 FILLER_40_2072 ();
 b15zdnd11an1n16x5 FILLER_40_2136 ();
 b15zdnd00an1n02x5 FILLER_40_2152 ();
 b15zdnd11an1n64x5 FILLER_40_2162 ();
 b15zdnd11an1n32x5 FILLER_40_2226 ();
 b15zdnd11an1n16x5 FILLER_40_2258 ();
 b15zdnd00an1n02x5 FILLER_40_2274 ();
 b15zdnd11an1n64x5 FILLER_41_0 ();
 b15zdnd11an1n64x5 FILLER_41_64 ();
 b15zdnd11an1n64x5 FILLER_41_128 ();
 b15zdnd11an1n08x5 FILLER_41_192 ();
 b15zdnd11an1n04x5 FILLER_41_200 ();
 b15zdnd00an1n02x5 FILLER_41_204 ();
 b15zdnd11an1n16x5 FILLER_41_226 ();
 b15zdnd11an1n04x5 FILLER_41_242 ();
 b15zdnd00an1n01x5 FILLER_41_246 ();
 b15zdnd11an1n64x5 FILLER_41_289 ();
 b15zdnd11an1n16x5 FILLER_41_353 ();
 b15zdnd11an1n32x5 FILLER_41_411 ();
 b15zdnd11an1n64x5 FILLER_41_474 ();
 b15zdnd00an1n02x5 FILLER_41_538 ();
 b15zdnd11an1n04x5 FILLER_41_561 ();
 b15zdnd00an1n01x5 FILLER_41_565 ();
 b15zdnd11an1n32x5 FILLER_41_591 ();
 b15zdnd11an1n16x5 FILLER_41_623 ();
 b15zdnd11an1n08x5 FILLER_41_639 ();
 b15zdnd11an1n64x5 FILLER_41_655 ();
 b15zdnd11an1n64x5 FILLER_41_719 ();
 b15zdnd11an1n32x5 FILLER_41_783 ();
 b15zdnd11an1n04x5 FILLER_41_815 ();
 b15zdnd00an1n02x5 FILLER_41_819 ();
 b15zdnd11an1n64x5 FILLER_41_873 ();
 b15zdnd11an1n64x5 FILLER_41_937 ();
 b15zdnd11an1n32x5 FILLER_41_1001 ();
 b15zdnd11an1n16x5 FILLER_41_1033 ();
 b15zdnd11an1n64x5 FILLER_41_1052 ();
 b15zdnd11an1n64x5 FILLER_41_1116 ();
 b15zdnd11an1n64x5 FILLER_41_1180 ();
 b15zdnd11an1n16x5 FILLER_41_1244 ();
 b15zdnd00an1n02x5 FILLER_41_1260 ();
 b15zdnd00an1n01x5 FILLER_41_1262 ();
 b15zdnd11an1n64x5 FILLER_41_1266 ();
 b15zdnd11an1n64x5 FILLER_41_1330 ();
 b15zdnd11an1n32x5 FILLER_41_1394 ();
 b15zdnd11an1n04x5 FILLER_41_1426 ();
 b15zdnd00an1n02x5 FILLER_41_1430 ();
 b15zdnd11an1n64x5 FILLER_41_1441 ();
 b15zdnd11an1n16x5 FILLER_41_1505 ();
 b15zdnd11an1n04x5 FILLER_41_1521 ();
 b15zdnd00an1n01x5 FILLER_41_1525 ();
 b15zdnd11an1n64x5 FILLER_41_1540 ();
 b15zdnd11an1n64x5 FILLER_41_1604 ();
 b15zdnd11an1n32x5 FILLER_41_1668 ();
 b15zdnd11an1n08x5 FILLER_41_1700 ();
 b15zdnd11an1n04x5 FILLER_41_1708 ();
 b15zdnd00an1n02x5 FILLER_41_1712 ();
 b15zdnd00an1n01x5 FILLER_41_1714 ();
 b15zdnd11an1n64x5 FILLER_41_1718 ();
 b15zdnd11an1n64x5 FILLER_41_1782 ();
 b15zdnd11an1n64x5 FILLER_41_1846 ();
 b15zdnd11an1n64x5 FILLER_41_1910 ();
 b15zdnd11an1n64x5 FILLER_41_1974 ();
 b15zdnd11an1n64x5 FILLER_41_2038 ();
 b15zdnd11an1n64x5 FILLER_41_2102 ();
 b15zdnd11an1n64x5 FILLER_41_2166 ();
 b15zdnd11an1n32x5 FILLER_41_2230 ();
 b15zdnd11an1n16x5 FILLER_41_2262 ();
 b15zdnd11an1n04x5 FILLER_41_2278 ();
 b15zdnd00an1n02x5 FILLER_41_2282 ();
 b15zdnd11an1n64x5 FILLER_42_8 ();
 b15zdnd11an1n64x5 FILLER_42_72 ();
 b15zdnd11an1n64x5 FILLER_42_136 ();
 b15zdnd11an1n16x5 FILLER_42_200 ();
 b15zdnd11an1n08x5 FILLER_42_216 ();
 b15zdnd00an1n01x5 FILLER_42_224 ();
 b15zdnd11an1n64x5 FILLER_42_250 ();
 b15zdnd11an1n32x5 FILLER_42_314 ();
 b15zdnd11an1n08x5 FILLER_42_346 ();
 b15zdnd11an1n04x5 FILLER_42_354 ();
 b15zdnd00an1n02x5 FILLER_42_358 ();
 b15zdnd11an1n64x5 FILLER_42_375 ();
 b15zdnd11an1n64x5 FILLER_42_439 ();
 b15zdnd11an1n32x5 FILLER_42_503 ();
 b15zdnd11an1n16x5 FILLER_42_535 ();
 b15zdnd11an1n08x5 FILLER_42_551 ();
 b15zdnd11an1n04x5 FILLER_42_559 ();
 b15zdnd00an1n01x5 FILLER_42_563 ();
 b15zdnd11an1n32x5 FILLER_42_595 ();
 b15zdnd11an1n04x5 FILLER_42_627 ();
 b15zdnd00an1n01x5 FILLER_42_631 ();
 b15zdnd11an1n32x5 FILLER_42_659 ();
 b15zdnd11an1n16x5 FILLER_42_691 ();
 b15zdnd11an1n08x5 FILLER_42_707 ();
 b15zdnd00an1n02x5 FILLER_42_715 ();
 b15zdnd00an1n01x5 FILLER_42_717 ();
 b15zdnd11an1n32x5 FILLER_42_726 ();
 b15zdnd11an1n16x5 FILLER_42_758 ();
 b15zdnd11an1n08x5 FILLER_42_774 ();
 b15zdnd00an1n02x5 FILLER_42_782 ();
 b15zdnd00an1n01x5 FILLER_42_784 ();
 b15zdnd11an1n32x5 FILLER_42_800 ();
 b15zdnd11an1n08x5 FILLER_42_832 ();
 b15zdnd11an1n04x5 FILLER_42_843 ();
 b15zdnd11an1n32x5 FILLER_42_850 ();
 b15zdnd11an1n64x5 FILLER_42_924 ();
 b15zdnd11an1n64x5 FILLER_42_988 ();
 b15zdnd11an1n64x5 FILLER_42_1052 ();
 b15zdnd11an1n64x5 FILLER_42_1116 ();
 b15zdnd11an1n64x5 FILLER_42_1180 ();
 b15zdnd11an1n64x5 FILLER_42_1244 ();
 b15zdnd11an1n64x5 FILLER_42_1308 ();
 b15zdnd00an1n02x5 FILLER_42_1372 ();
 b15zdnd00an1n01x5 FILLER_42_1374 ();
 b15zdnd11an1n64x5 FILLER_42_1391 ();
 b15zdnd11an1n64x5 FILLER_42_1455 ();
 b15zdnd11an1n64x5 FILLER_42_1519 ();
 b15zdnd11an1n64x5 FILLER_42_1583 ();
 b15zdnd11an1n64x5 FILLER_42_1647 ();
 b15zdnd11an1n08x5 FILLER_42_1711 ();
 b15zdnd00an1n01x5 FILLER_42_1719 ();
 b15zdnd11an1n64x5 FILLER_42_1726 ();
 b15zdnd11an1n64x5 FILLER_42_1790 ();
 b15zdnd11an1n64x5 FILLER_42_1854 ();
 b15zdnd11an1n64x5 FILLER_42_1918 ();
 b15zdnd11an1n64x5 FILLER_42_1982 ();
 b15zdnd11an1n64x5 FILLER_42_2046 ();
 b15zdnd11an1n32x5 FILLER_42_2110 ();
 b15zdnd11an1n08x5 FILLER_42_2142 ();
 b15zdnd11an1n04x5 FILLER_42_2150 ();
 b15zdnd11an1n64x5 FILLER_42_2162 ();
 b15zdnd11an1n32x5 FILLER_42_2226 ();
 b15zdnd11an1n16x5 FILLER_42_2258 ();
 b15zdnd00an1n02x5 FILLER_42_2274 ();
 b15zdnd11an1n64x5 FILLER_43_0 ();
 b15zdnd11an1n64x5 FILLER_43_64 ();
 b15zdnd11an1n64x5 FILLER_43_128 ();
 b15zdnd11an1n16x5 FILLER_43_192 ();
 b15zdnd11an1n64x5 FILLER_43_250 ();
 b15zdnd11an1n08x5 FILLER_43_314 ();
 b15zdnd11an1n04x5 FILLER_43_322 ();
 b15zdnd00an1n02x5 FILLER_43_326 ();
 b15zdnd11an1n64x5 FILLER_43_370 ();
 b15zdnd11an1n32x5 FILLER_43_434 ();
 b15zdnd11an1n64x5 FILLER_43_497 ();
 b15zdnd11an1n16x5 FILLER_43_561 ();
 b15zdnd11an1n08x5 FILLER_43_577 ();
 b15zdnd11an1n64x5 FILLER_43_594 ();
 b15zdnd11an1n04x5 FILLER_43_658 ();
 b15zdnd11an1n16x5 FILLER_43_669 ();
 b15zdnd11an1n64x5 FILLER_43_725 ();
 b15zdnd11an1n16x5 FILLER_43_789 ();
 b15zdnd11an1n08x5 FILLER_43_805 ();
 b15zdnd11an1n04x5 FILLER_43_813 ();
 b15zdnd00an1n02x5 FILLER_43_817 ();
 b15zdnd11an1n64x5 FILLER_43_861 ();
 b15zdnd11an1n64x5 FILLER_43_925 ();
 b15zdnd11an1n64x5 FILLER_43_989 ();
 b15zdnd11an1n64x5 FILLER_43_1053 ();
 b15zdnd11an1n64x5 FILLER_43_1117 ();
 b15zdnd11an1n64x5 FILLER_43_1181 ();
 b15zdnd11an1n64x5 FILLER_43_1245 ();
 b15zdnd11an1n64x5 FILLER_43_1309 ();
 b15zdnd11an1n08x5 FILLER_43_1373 ();
 b15zdnd11an1n04x5 FILLER_43_1381 ();
 b15zdnd00an1n01x5 FILLER_43_1385 ();
 b15zdnd11an1n64x5 FILLER_43_1403 ();
 b15zdnd11an1n64x5 FILLER_43_1467 ();
 b15zdnd11an1n64x5 FILLER_43_1531 ();
 b15zdnd11an1n64x5 FILLER_43_1595 ();
 b15zdnd11an1n64x5 FILLER_43_1659 ();
 b15zdnd11an1n64x5 FILLER_43_1723 ();
 b15zdnd11an1n32x5 FILLER_43_1787 ();
 b15zdnd00an1n02x5 FILLER_43_1819 ();
 b15zdnd00an1n01x5 FILLER_43_1821 ();
 b15zdnd11an1n64x5 FILLER_43_1836 ();
 b15zdnd11an1n64x5 FILLER_43_1900 ();
 b15zdnd11an1n64x5 FILLER_43_1964 ();
 b15zdnd11an1n64x5 FILLER_43_2028 ();
 b15zdnd11an1n64x5 FILLER_43_2092 ();
 b15zdnd11an1n64x5 FILLER_43_2156 ();
 b15zdnd11an1n64x5 FILLER_43_2220 ();
 b15zdnd11an1n64x5 FILLER_44_8 ();
 b15zdnd11an1n64x5 FILLER_44_72 ();
 b15zdnd11an1n64x5 FILLER_44_136 ();
 b15zdnd11an1n32x5 FILLER_44_200 ();
 b15zdnd11an1n16x5 FILLER_44_232 ();
 b15zdnd11an1n04x5 FILLER_44_248 ();
 b15zdnd00an1n01x5 FILLER_44_252 ();
 b15zdnd11an1n64x5 FILLER_44_267 ();
 b15zdnd11an1n64x5 FILLER_44_331 ();
 b15zdnd11an1n64x5 FILLER_44_395 ();
 b15zdnd11an1n64x5 FILLER_44_459 ();
 b15zdnd11an1n64x5 FILLER_44_523 ();
 b15zdnd11an1n64x5 FILLER_44_587 ();
 b15zdnd11an1n16x5 FILLER_44_651 ();
 b15zdnd11an1n08x5 FILLER_44_667 ();
 b15zdnd11an1n04x5 FILLER_44_675 ();
 b15zdnd00an1n01x5 FILLER_44_679 ();
 b15zdnd11an1n04x5 FILLER_44_711 ();
 b15zdnd00an1n02x5 FILLER_44_715 ();
 b15zdnd00an1n01x5 FILLER_44_717 ();
 b15zdnd11an1n64x5 FILLER_44_726 ();
 b15zdnd11an1n64x5 FILLER_44_790 ();
 b15zdnd11an1n64x5 FILLER_44_854 ();
 b15zdnd11an1n64x5 FILLER_44_918 ();
 b15zdnd11an1n64x5 FILLER_44_982 ();
 b15zdnd11an1n64x5 FILLER_44_1046 ();
 b15zdnd11an1n32x5 FILLER_44_1110 ();
 b15zdnd11an1n16x5 FILLER_44_1142 ();
 b15zdnd11an1n04x5 FILLER_44_1158 ();
 b15zdnd00an1n02x5 FILLER_44_1162 ();
 b15zdnd00an1n01x5 FILLER_44_1164 ();
 b15zdnd11an1n64x5 FILLER_44_1207 ();
 b15zdnd11an1n64x5 FILLER_44_1271 ();
 b15zdnd11an1n32x5 FILLER_44_1335 ();
 b15zdnd11an1n16x5 FILLER_44_1367 ();
 b15zdnd11an1n64x5 FILLER_44_1435 ();
 b15zdnd11an1n64x5 FILLER_44_1499 ();
 b15zdnd00an1n02x5 FILLER_44_1563 ();
 b15zdnd00an1n01x5 FILLER_44_1565 ();
 b15zdnd11an1n32x5 FILLER_44_1593 ();
 b15zdnd11an1n16x5 FILLER_44_1625 ();
 b15zdnd11an1n08x5 FILLER_44_1641 ();
 b15zdnd11an1n04x5 FILLER_44_1649 ();
 b15zdnd00an1n01x5 FILLER_44_1653 ();
 b15zdnd11an1n32x5 FILLER_44_1663 ();
 b15zdnd11an1n04x5 FILLER_44_1695 ();
 b15zdnd00an1n02x5 FILLER_44_1699 ();
 b15zdnd11an1n04x5 FILLER_44_1704 ();
 b15zdnd11an1n64x5 FILLER_44_1711 ();
 b15zdnd11an1n64x5 FILLER_44_1775 ();
 b15zdnd11an1n64x5 FILLER_44_1839 ();
 b15zdnd11an1n64x5 FILLER_44_1903 ();
 b15zdnd11an1n64x5 FILLER_44_1967 ();
 b15zdnd11an1n04x5 FILLER_44_2031 ();
 b15zdnd11an1n64x5 FILLER_44_2049 ();
 b15zdnd11an1n32x5 FILLER_44_2113 ();
 b15zdnd11an1n08x5 FILLER_44_2145 ();
 b15zdnd00an1n01x5 FILLER_44_2153 ();
 b15zdnd11an1n64x5 FILLER_44_2162 ();
 b15zdnd11an1n32x5 FILLER_44_2226 ();
 b15zdnd11an1n16x5 FILLER_44_2258 ();
 b15zdnd00an1n02x5 FILLER_44_2274 ();
 b15zdnd11an1n64x5 FILLER_45_0 ();
 b15zdnd11an1n64x5 FILLER_45_64 ();
 b15zdnd11an1n64x5 FILLER_45_128 ();
 b15zdnd11an1n64x5 FILLER_45_192 ();
 b15zdnd11an1n64x5 FILLER_45_256 ();
 b15zdnd11an1n64x5 FILLER_45_320 ();
 b15zdnd11an1n64x5 FILLER_45_384 ();
 b15zdnd11an1n64x5 FILLER_45_448 ();
 b15zdnd11an1n32x5 FILLER_45_512 ();
 b15zdnd11an1n04x5 FILLER_45_544 ();
 b15zdnd00an1n02x5 FILLER_45_548 ();
 b15zdnd11an1n64x5 FILLER_45_556 ();
 b15zdnd11an1n64x5 FILLER_45_620 ();
 b15zdnd11an1n64x5 FILLER_45_684 ();
 b15zdnd11an1n64x5 FILLER_45_748 ();
 b15zdnd11an1n64x5 FILLER_45_812 ();
 b15zdnd11an1n64x5 FILLER_45_876 ();
 b15zdnd11an1n64x5 FILLER_45_940 ();
 b15zdnd11an1n64x5 FILLER_45_1004 ();
 b15zdnd11an1n64x5 FILLER_45_1068 ();
 b15zdnd11an1n64x5 FILLER_45_1132 ();
 b15zdnd11an1n64x5 FILLER_45_1196 ();
 b15zdnd11an1n64x5 FILLER_45_1260 ();
 b15zdnd11an1n64x5 FILLER_45_1324 ();
 b15zdnd11an1n08x5 FILLER_45_1388 ();
 b15zdnd00an1n02x5 FILLER_45_1396 ();
 b15zdnd00an1n01x5 FILLER_45_1398 ();
 b15zdnd11an1n04x5 FILLER_45_1402 ();
 b15zdnd11an1n04x5 FILLER_45_1409 ();
 b15zdnd11an1n08x5 FILLER_45_1416 ();
 b15zdnd00an1n02x5 FILLER_45_1424 ();
 b15zdnd00an1n01x5 FILLER_45_1426 ();
 b15zdnd11an1n04x5 FILLER_45_1434 ();
 b15zdnd00an1n02x5 FILLER_45_1438 ();
 b15zdnd11an1n64x5 FILLER_45_1447 ();
 b15zdnd11an1n32x5 FILLER_45_1511 ();
 b15zdnd11an1n16x5 FILLER_45_1543 ();
 b15zdnd11an1n08x5 FILLER_45_1559 ();
 b15zdnd11an1n16x5 FILLER_45_1570 ();
 b15zdnd00an1n02x5 FILLER_45_1586 ();
 b15zdnd11an1n04x5 FILLER_45_1591 ();
 b15zdnd11an1n16x5 FILLER_45_1598 ();
 b15zdnd11an1n08x5 FILLER_45_1614 ();
 b15zdnd11an1n04x5 FILLER_45_1622 ();
 b15zdnd00an1n01x5 FILLER_45_1626 ();
 b15zdnd11an1n16x5 FILLER_45_1636 ();
 b15zdnd00an1n02x5 FILLER_45_1652 ();
 b15zdnd00an1n01x5 FILLER_45_1654 ();
 b15zdnd11an1n32x5 FILLER_45_1664 ();
 b15zdnd11an1n04x5 FILLER_45_1696 ();
 b15zdnd11an1n04x5 FILLER_45_1703 ();
 b15zdnd11an1n04x5 FILLER_45_1710 ();
 b15zdnd11an1n64x5 FILLER_45_1717 ();
 b15zdnd11an1n64x5 FILLER_45_1781 ();
 b15zdnd11an1n64x5 FILLER_45_1845 ();
 b15zdnd11an1n64x5 FILLER_45_1909 ();
 b15zdnd11an1n64x5 FILLER_45_1973 ();
 b15zdnd11an1n64x5 FILLER_45_2037 ();
 b15zdnd11an1n64x5 FILLER_45_2101 ();
 b15zdnd11an1n64x5 FILLER_45_2165 ();
 b15zdnd11an1n32x5 FILLER_45_2229 ();
 b15zdnd11an1n16x5 FILLER_45_2261 ();
 b15zdnd11an1n04x5 FILLER_45_2277 ();
 b15zdnd00an1n02x5 FILLER_45_2281 ();
 b15zdnd00an1n01x5 FILLER_45_2283 ();
 b15zdnd11an1n64x5 FILLER_46_8 ();
 b15zdnd11an1n64x5 FILLER_46_72 ();
 b15zdnd11an1n32x5 FILLER_46_136 ();
 b15zdnd11an1n16x5 FILLER_46_168 ();
 b15zdnd11an1n04x5 FILLER_46_184 ();
 b15zdnd00an1n02x5 FILLER_46_188 ();
 b15zdnd11an1n64x5 FILLER_46_193 ();
 b15zdnd11an1n64x5 FILLER_46_257 ();
 b15zdnd11an1n08x5 FILLER_46_321 ();
 b15zdnd00an1n02x5 FILLER_46_329 ();
 b15zdnd00an1n01x5 FILLER_46_331 ();
 b15zdnd11an1n64x5 FILLER_46_337 ();
 b15zdnd11an1n64x5 FILLER_46_401 ();
 b15zdnd11an1n64x5 FILLER_46_465 ();
 b15zdnd11an1n32x5 FILLER_46_529 ();
 b15zdnd11an1n08x5 FILLER_46_561 ();
 b15zdnd11an1n04x5 FILLER_46_569 ();
 b15zdnd00an1n02x5 FILLER_46_573 ();
 b15zdnd00an1n01x5 FILLER_46_575 ();
 b15zdnd11an1n64x5 FILLER_46_607 ();
 b15zdnd11an1n32x5 FILLER_46_671 ();
 b15zdnd11an1n08x5 FILLER_46_703 ();
 b15zdnd11an1n04x5 FILLER_46_711 ();
 b15zdnd00an1n02x5 FILLER_46_715 ();
 b15zdnd00an1n01x5 FILLER_46_717 ();
 b15zdnd11an1n64x5 FILLER_46_726 ();
 b15zdnd11an1n64x5 FILLER_46_790 ();
 b15zdnd11an1n64x5 FILLER_46_854 ();
 b15zdnd11an1n64x5 FILLER_46_918 ();
 b15zdnd11an1n64x5 FILLER_46_982 ();
 b15zdnd11an1n64x5 FILLER_46_1046 ();
 b15zdnd11an1n64x5 FILLER_46_1110 ();
 b15zdnd11an1n64x5 FILLER_46_1174 ();
 b15zdnd11an1n64x5 FILLER_46_1238 ();
 b15zdnd11an1n32x5 FILLER_46_1302 ();
 b15zdnd11an1n16x5 FILLER_46_1334 ();
 b15zdnd11an1n08x5 FILLER_46_1350 ();
 b15zdnd11an1n04x5 FILLER_46_1358 ();
 b15zdnd11an1n04x5 FILLER_46_1368 ();
 b15zdnd00an1n02x5 FILLER_46_1372 ();
 b15zdnd00an1n01x5 FILLER_46_1374 ();
 b15zdnd11an1n08x5 FILLER_46_1417 ();
 b15zdnd11an1n04x5 FILLER_46_1425 ();
 b15zdnd00an1n02x5 FILLER_46_1429 ();
 b15zdnd11an1n64x5 FILLER_46_1473 ();
 b15zdnd11an1n16x5 FILLER_46_1537 ();
 b15zdnd11an1n08x5 FILLER_46_1553 ();
 b15zdnd00an1n02x5 FILLER_46_1561 ();
 b15zdnd11an1n32x5 FILLER_46_1615 ();
 b15zdnd11an1n16x5 FILLER_46_1647 ();
 b15zdnd11an1n04x5 FILLER_46_1663 ();
 b15zdnd00an1n02x5 FILLER_46_1667 ();
 b15zdnd00an1n01x5 FILLER_46_1669 ();
 b15zdnd11an1n04x5 FILLER_46_1677 ();
 b15zdnd11an1n04x5 FILLER_46_1733 ();
 b15zdnd11an1n64x5 FILLER_46_1740 ();
 b15zdnd11an1n64x5 FILLER_46_1804 ();
 b15zdnd11an1n64x5 FILLER_46_1868 ();
 b15zdnd11an1n64x5 FILLER_46_1932 ();
 b15zdnd11an1n64x5 FILLER_46_1996 ();
 b15zdnd11an1n32x5 FILLER_46_2060 ();
 b15zdnd11an1n04x5 FILLER_46_2092 ();
 b15zdnd00an1n02x5 FILLER_46_2096 ();
 b15zdnd00an1n01x5 FILLER_46_2098 ();
 b15zdnd11an1n16x5 FILLER_46_2111 ();
 b15zdnd11an1n08x5 FILLER_46_2127 ();
 b15zdnd11an1n04x5 FILLER_46_2147 ();
 b15zdnd00an1n02x5 FILLER_46_2151 ();
 b15zdnd00an1n01x5 FILLER_46_2153 ();
 b15zdnd11an1n32x5 FILLER_46_2162 ();
 b15zdnd11an1n08x5 FILLER_46_2194 ();
 b15zdnd00an1n01x5 FILLER_46_2202 ();
 b15zdnd11an1n64x5 FILLER_46_2212 ();
 b15zdnd11an1n64x5 FILLER_47_0 ();
 b15zdnd11an1n64x5 FILLER_47_64 ();
 b15zdnd11an1n64x5 FILLER_47_128 ();
 b15zdnd00an1n01x5 FILLER_47_192 ();
 b15zdnd11an1n64x5 FILLER_47_198 ();
 b15zdnd11an1n64x5 FILLER_47_262 ();
 b15zdnd11an1n04x5 FILLER_47_326 ();
 b15zdnd00an1n02x5 FILLER_47_330 ();
 b15zdnd00an1n01x5 FILLER_47_332 ();
 b15zdnd11an1n64x5 FILLER_47_336 ();
 b15zdnd11an1n64x5 FILLER_47_400 ();
 b15zdnd11an1n16x5 FILLER_47_464 ();
 b15zdnd11an1n08x5 FILLER_47_480 ();
 b15zdnd11an1n04x5 FILLER_47_488 ();
 b15zdnd00an1n02x5 FILLER_47_492 ();
 b15zdnd11an1n08x5 FILLER_47_536 ();
 b15zdnd11an1n04x5 FILLER_47_544 ();
 b15zdnd00an1n01x5 FILLER_47_548 ();
 b15zdnd11an1n64x5 FILLER_47_556 ();
 b15zdnd11an1n64x5 FILLER_47_620 ();
 b15zdnd11an1n64x5 FILLER_47_684 ();
 b15zdnd11an1n64x5 FILLER_47_748 ();
 b15zdnd11an1n64x5 FILLER_47_812 ();
 b15zdnd11an1n64x5 FILLER_47_876 ();
 b15zdnd11an1n64x5 FILLER_47_940 ();
 b15zdnd11an1n64x5 FILLER_47_1004 ();
 b15zdnd11an1n16x5 FILLER_47_1068 ();
 b15zdnd11an1n08x5 FILLER_47_1084 ();
 b15zdnd00an1n02x5 FILLER_47_1092 ();
 b15zdnd00an1n01x5 FILLER_47_1094 ();
 b15zdnd11an1n64x5 FILLER_47_1137 ();
 b15zdnd11an1n64x5 FILLER_47_1201 ();
 b15zdnd11an1n64x5 FILLER_47_1265 ();
 b15zdnd11an1n64x5 FILLER_47_1329 ();
 b15zdnd11an1n64x5 FILLER_47_1393 ();
 b15zdnd11an1n64x5 FILLER_47_1457 ();
 b15zdnd11an1n32x5 FILLER_47_1521 ();
 b15zdnd11an1n16x5 FILLER_47_1553 ();
 b15zdnd11an1n04x5 FILLER_47_1569 ();
 b15zdnd11an1n04x5 FILLER_47_1576 ();
 b15zdnd11an1n04x5 FILLER_47_1583 ();
 b15zdnd11an1n04x5 FILLER_47_1590 ();
 b15zdnd11an1n64x5 FILLER_47_1597 ();
 b15zdnd11an1n16x5 FILLER_47_1661 ();
 b15zdnd00an1n02x5 FILLER_47_1677 ();
 b15zdnd00an1n01x5 FILLER_47_1679 ();
 b15zdnd11an1n64x5 FILLER_47_1732 ();
 b15zdnd11an1n64x5 FILLER_47_1796 ();
 b15zdnd11an1n64x5 FILLER_47_1860 ();
 b15zdnd11an1n64x5 FILLER_47_1924 ();
 b15zdnd11an1n64x5 FILLER_47_1988 ();
 b15zdnd11an1n64x5 FILLER_47_2052 ();
 b15zdnd11an1n64x5 FILLER_47_2116 ();
 b15zdnd11an1n64x5 FILLER_47_2180 ();
 b15zdnd11an1n32x5 FILLER_47_2244 ();
 b15zdnd11an1n08x5 FILLER_47_2276 ();
 b15zdnd11an1n64x5 FILLER_48_8 ();
 b15zdnd11an1n64x5 FILLER_48_72 ();
 b15zdnd11an1n32x5 FILLER_48_136 ();
 b15zdnd11an1n16x5 FILLER_48_168 ();
 b15zdnd11an1n08x5 FILLER_48_184 ();
 b15zdnd00an1n02x5 FILLER_48_192 ();
 b15zdnd00an1n01x5 FILLER_48_194 ();
 b15zdnd11an1n64x5 FILLER_48_237 ();
 b15zdnd11an1n64x5 FILLER_48_301 ();
 b15zdnd11an1n64x5 FILLER_48_365 ();
 b15zdnd11an1n64x5 FILLER_48_429 ();
 b15zdnd11an1n32x5 FILLER_48_493 ();
 b15zdnd00an1n02x5 FILLER_48_525 ();
 b15zdnd11an1n64x5 FILLER_48_558 ();
 b15zdnd11an1n32x5 FILLER_48_622 ();
 b15zdnd11an1n16x5 FILLER_48_654 ();
 b15zdnd11an1n08x5 FILLER_48_670 ();
 b15zdnd11an1n04x5 FILLER_48_678 ();
 b15zdnd00an1n02x5 FILLER_48_682 ();
 b15zdnd00an1n01x5 FILLER_48_684 ();
 b15zdnd00an1n02x5 FILLER_48_716 ();
 b15zdnd11an1n64x5 FILLER_48_726 ();
 b15zdnd11an1n64x5 FILLER_48_790 ();
 b15zdnd11an1n64x5 FILLER_48_854 ();
 b15zdnd11an1n64x5 FILLER_48_918 ();
 b15zdnd11an1n64x5 FILLER_48_982 ();
 b15zdnd11an1n64x5 FILLER_48_1046 ();
 b15zdnd11an1n64x5 FILLER_48_1110 ();
 b15zdnd11an1n64x5 FILLER_48_1174 ();
 b15zdnd11an1n04x5 FILLER_48_1238 ();
 b15zdnd11an1n64x5 FILLER_48_1265 ();
 b15zdnd11an1n64x5 FILLER_48_1329 ();
 b15zdnd11an1n64x5 FILLER_48_1393 ();
 b15zdnd11an1n64x5 FILLER_48_1457 ();
 b15zdnd00an1n02x5 FILLER_48_1521 ();
 b15zdnd11an1n16x5 FILLER_48_1535 ();
 b15zdnd00an1n02x5 FILLER_48_1551 ();
 b15zdnd11an1n64x5 FILLER_48_1605 ();
 b15zdnd11an1n08x5 FILLER_48_1669 ();
 b15zdnd11an1n04x5 FILLER_48_1677 ();
 b15zdnd00an1n02x5 FILLER_48_1681 ();
 b15zdnd00an1n01x5 FILLER_48_1683 ();
 b15zdnd11an1n64x5 FILLER_48_1736 ();
 b15zdnd11an1n32x5 FILLER_48_1800 ();
 b15zdnd11an1n16x5 FILLER_48_1832 ();
 b15zdnd00an1n02x5 FILLER_48_1848 ();
 b15zdnd11an1n64x5 FILLER_48_1853 ();
 b15zdnd11an1n64x5 FILLER_48_1917 ();
 b15zdnd11an1n64x5 FILLER_48_1981 ();
 b15zdnd11an1n64x5 FILLER_48_2045 ();
 b15zdnd11an1n32x5 FILLER_48_2109 ();
 b15zdnd11an1n08x5 FILLER_48_2141 ();
 b15zdnd11an1n04x5 FILLER_48_2149 ();
 b15zdnd00an1n01x5 FILLER_48_2153 ();
 b15zdnd11an1n64x5 FILLER_48_2162 ();
 b15zdnd11an1n32x5 FILLER_48_2226 ();
 b15zdnd11an1n16x5 FILLER_48_2258 ();
 b15zdnd00an1n02x5 FILLER_48_2274 ();
 b15zdnd11an1n64x5 FILLER_49_0 ();
 b15zdnd11an1n64x5 FILLER_49_64 ();
 b15zdnd11an1n64x5 FILLER_49_128 ();
 b15zdnd11an1n64x5 FILLER_49_192 ();
 b15zdnd11an1n64x5 FILLER_49_256 ();
 b15zdnd11an1n64x5 FILLER_49_320 ();
 b15zdnd11an1n64x5 FILLER_49_384 ();
 b15zdnd11an1n64x5 FILLER_49_448 ();
 b15zdnd11an1n64x5 FILLER_49_512 ();
 b15zdnd11an1n32x5 FILLER_49_576 ();
 b15zdnd11an1n04x5 FILLER_49_608 ();
 b15zdnd00an1n02x5 FILLER_49_612 ();
 b15zdnd11an1n32x5 FILLER_49_656 ();
 b15zdnd11an1n16x5 FILLER_49_688 ();
 b15zdnd00an1n02x5 FILLER_49_704 ();
 b15zdnd11an1n64x5 FILLER_49_748 ();
 b15zdnd11an1n64x5 FILLER_49_812 ();
 b15zdnd11an1n64x5 FILLER_49_876 ();
 b15zdnd11an1n64x5 FILLER_49_940 ();
 b15zdnd11an1n64x5 FILLER_49_1004 ();
 b15zdnd11an1n64x5 FILLER_49_1068 ();
 b15zdnd11an1n64x5 FILLER_49_1132 ();
 b15zdnd11an1n64x5 FILLER_49_1196 ();
 b15zdnd11an1n64x5 FILLER_49_1260 ();
 b15zdnd11an1n64x5 FILLER_49_1324 ();
 b15zdnd11an1n64x5 FILLER_49_1388 ();
 b15zdnd11an1n32x5 FILLER_49_1452 ();
 b15zdnd11an1n08x5 FILLER_49_1484 ();
 b15zdnd11an1n32x5 FILLER_49_1500 ();
 b15zdnd11an1n16x5 FILLER_49_1532 ();
 b15zdnd11an1n04x5 FILLER_49_1548 ();
 b15zdnd00an1n01x5 FILLER_49_1552 ();
 b15zdnd11an1n64x5 FILLER_49_1605 ();
 b15zdnd11an1n16x5 FILLER_49_1669 ();
 b15zdnd11an1n08x5 FILLER_49_1685 ();
 b15zdnd11an1n04x5 FILLER_49_1693 ();
 b15zdnd00an1n02x5 FILLER_49_1697 ();
 b15zdnd00an1n01x5 FILLER_49_1699 ();
 b15zdnd11an1n04x5 FILLER_49_1703 ();
 b15zdnd11an1n64x5 FILLER_49_1710 ();
 b15zdnd11an1n64x5 FILLER_49_1774 ();
 b15zdnd11an1n08x5 FILLER_49_1838 ();
 b15zdnd00an1n02x5 FILLER_49_1846 ();
 b15zdnd00an1n01x5 FILLER_49_1848 ();
 b15zdnd11an1n64x5 FILLER_49_1852 ();
 b15zdnd11an1n32x5 FILLER_49_1916 ();
 b15zdnd11an1n08x5 FILLER_49_1948 ();
 b15zdnd11an1n04x5 FILLER_49_1956 ();
 b15zdnd00an1n01x5 FILLER_49_1960 ();
 b15zdnd11an1n64x5 FILLER_49_1964 ();
 b15zdnd11an1n64x5 FILLER_49_2028 ();
 b15zdnd11an1n64x5 FILLER_49_2092 ();
 b15zdnd11an1n64x5 FILLER_49_2156 ();
 b15zdnd11an1n64x5 FILLER_49_2220 ();
 b15zdnd11an1n64x5 FILLER_50_8 ();
 b15zdnd11an1n64x5 FILLER_50_72 ();
 b15zdnd11an1n64x5 FILLER_50_136 ();
 b15zdnd11an1n64x5 FILLER_50_200 ();
 b15zdnd11an1n64x5 FILLER_50_264 ();
 b15zdnd11an1n64x5 FILLER_50_370 ();
 b15zdnd11an1n64x5 FILLER_50_434 ();
 b15zdnd11an1n16x5 FILLER_50_498 ();
 b15zdnd11an1n08x5 FILLER_50_514 ();
 b15zdnd11an1n04x5 FILLER_50_522 ();
 b15zdnd11an1n32x5 FILLER_50_568 ();
 b15zdnd11an1n08x5 FILLER_50_600 ();
 b15zdnd11an1n64x5 FILLER_50_611 ();
 b15zdnd11an1n16x5 FILLER_50_675 ();
 b15zdnd00an1n02x5 FILLER_50_716 ();
 b15zdnd11an1n64x5 FILLER_50_726 ();
 b15zdnd11an1n64x5 FILLER_50_790 ();
 b15zdnd11an1n64x5 FILLER_50_854 ();
 b15zdnd11an1n64x5 FILLER_50_918 ();
 b15zdnd11an1n64x5 FILLER_50_982 ();
 b15zdnd11an1n64x5 FILLER_50_1046 ();
 b15zdnd11an1n16x5 FILLER_50_1110 ();
 b15zdnd11an1n08x5 FILLER_50_1126 ();
 b15zdnd11an1n64x5 FILLER_50_1162 ();
 b15zdnd11an1n64x5 FILLER_50_1226 ();
 b15zdnd11an1n64x5 FILLER_50_1290 ();
 b15zdnd11an1n64x5 FILLER_50_1354 ();
 b15zdnd11an1n64x5 FILLER_50_1418 ();
 b15zdnd11an1n64x5 FILLER_50_1482 ();
 b15zdnd11an1n16x5 FILLER_50_1546 ();
 b15zdnd11an1n08x5 FILLER_50_1562 ();
 b15zdnd00an1n01x5 FILLER_50_1570 ();
 b15zdnd11an1n04x5 FILLER_50_1574 ();
 b15zdnd11an1n64x5 FILLER_50_1581 ();
 b15zdnd11an1n32x5 FILLER_50_1645 ();
 b15zdnd11an1n16x5 FILLER_50_1677 ();
 b15zdnd11an1n08x5 FILLER_50_1693 ();
 b15zdnd11an1n64x5 FILLER_50_1704 ();
 b15zdnd11an1n32x5 FILLER_50_1768 ();
 b15zdnd11an1n16x5 FILLER_50_1800 ();
 b15zdnd11an1n08x5 FILLER_50_1816 ();
 b15zdnd11an1n64x5 FILLER_50_1876 ();
 b15zdnd11an1n16x5 FILLER_50_1940 ();
 b15zdnd11an1n04x5 FILLER_50_1956 ();
 b15zdnd00an1n02x5 FILLER_50_1960 ();
 b15zdnd11an1n64x5 FILLER_50_1965 ();
 b15zdnd11an1n08x5 FILLER_50_2029 ();
 b15zdnd11an1n64x5 FILLER_50_2041 ();
 b15zdnd11an1n32x5 FILLER_50_2105 ();
 b15zdnd11an1n16x5 FILLER_50_2137 ();
 b15zdnd00an1n01x5 FILLER_50_2153 ();
 b15zdnd11an1n64x5 FILLER_50_2162 ();
 b15zdnd11an1n32x5 FILLER_50_2226 ();
 b15zdnd11an1n16x5 FILLER_50_2258 ();
 b15zdnd00an1n02x5 FILLER_50_2274 ();
 b15zdnd11an1n64x5 FILLER_51_0 ();
 b15zdnd11an1n64x5 FILLER_51_64 ();
 b15zdnd11an1n64x5 FILLER_51_128 ();
 b15zdnd11an1n64x5 FILLER_51_192 ();
 b15zdnd11an1n64x5 FILLER_51_256 ();
 b15zdnd11an1n64x5 FILLER_51_320 ();
 b15zdnd11an1n64x5 FILLER_51_384 ();
 b15zdnd11an1n64x5 FILLER_51_448 ();
 b15zdnd11an1n64x5 FILLER_51_512 ();
 b15zdnd11an1n04x5 FILLER_51_576 ();
 b15zdnd00an1n01x5 FILLER_51_580 ();
 b15zdnd11an1n64x5 FILLER_51_633 ();
 b15zdnd11an1n64x5 FILLER_51_697 ();
 b15zdnd11an1n64x5 FILLER_51_761 ();
 b15zdnd11an1n08x5 FILLER_51_825 ();
 b15zdnd11an1n04x5 FILLER_51_833 ();
 b15zdnd00an1n02x5 FILLER_51_837 ();
 b15zdnd11an1n64x5 FILLER_51_847 ();
 b15zdnd11an1n64x5 FILLER_51_911 ();
 b15zdnd11an1n32x5 FILLER_51_975 ();
 b15zdnd11an1n04x5 FILLER_51_1007 ();
 b15zdnd00an1n02x5 FILLER_51_1011 ();
 b15zdnd00an1n01x5 FILLER_51_1013 ();
 b15zdnd11an1n64x5 FILLER_51_1056 ();
 b15zdnd11an1n16x5 FILLER_51_1120 ();
 b15zdnd11an1n08x5 FILLER_51_1136 ();
 b15zdnd11an1n04x5 FILLER_51_1144 ();
 b15zdnd00an1n02x5 FILLER_51_1148 ();
 b15zdnd11an1n04x5 FILLER_51_1153 ();
 b15zdnd11an1n64x5 FILLER_51_1160 ();
 b15zdnd11an1n64x5 FILLER_51_1224 ();
 b15zdnd11an1n64x5 FILLER_51_1288 ();
 b15zdnd11an1n64x5 FILLER_51_1352 ();
 b15zdnd11an1n64x5 FILLER_51_1416 ();
 b15zdnd11an1n64x5 FILLER_51_1480 ();
 b15zdnd11an1n32x5 FILLER_51_1544 ();
 b15zdnd00an1n01x5 FILLER_51_1576 ();
 b15zdnd11an1n64x5 FILLER_51_1580 ();
 b15zdnd11an1n64x5 FILLER_51_1644 ();
 b15zdnd11an1n16x5 FILLER_51_1708 ();
 b15zdnd11an1n08x5 FILLER_51_1724 ();
 b15zdnd00an1n02x5 FILLER_51_1732 ();
 b15zdnd11an1n32x5 FILLER_51_1776 ();
 b15zdnd11an1n16x5 FILLER_51_1808 ();
 b15zdnd00an1n02x5 FILLER_51_1824 ();
 b15zdnd11an1n32x5 FILLER_51_1878 ();
 b15zdnd11an1n16x5 FILLER_51_1910 ();
 b15zdnd11an1n08x5 FILLER_51_1926 ();
 b15zdnd00an1n02x5 FILLER_51_1934 ();
 b15zdnd00an1n01x5 FILLER_51_1936 ();
 b15zdnd11an1n64x5 FILLER_51_1989 ();
 b15zdnd11an1n64x5 FILLER_51_2053 ();
 b15zdnd11an1n64x5 FILLER_51_2117 ();
 b15zdnd11an1n64x5 FILLER_51_2181 ();
 b15zdnd11an1n32x5 FILLER_51_2245 ();
 b15zdnd11an1n04x5 FILLER_51_2277 ();
 b15zdnd00an1n02x5 FILLER_51_2281 ();
 b15zdnd00an1n01x5 FILLER_51_2283 ();
 b15zdnd11an1n64x5 FILLER_52_8 ();
 b15zdnd11an1n64x5 FILLER_52_72 ();
 b15zdnd11an1n64x5 FILLER_52_136 ();
 b15zdnd11an1n64x5 FILLER_52_200 ();
 b15zdnd11an1n64x5 FILLER_52_264 ();
 b15zdnd11an1n64x5 FILLER_52_328 ();
 b15zdnd11an1n64x5 FILLER_52_392 ();
 b15zdnd11an1n64x5 FILLER_52_456 ();
 b15zdnd11an1n64x5 FILLER_52_520 ();
 b15zdnd11an1n16x5 FILLER_52_584 ();
 b15zdnd11an1n04x5 FILLER_52_603 ();
 b15zdnd11an1n64x5 FILLER_52_610 ();
 b15zdnd11an1n32x5 FILLER_52_674 ();
 b15zdnd11an1n08x5 FILLER_52_706 ();
 b15zdnd11an1n04x5 FILLER_52_714 ();
 b15zdnd11an1n64x5 FILLER_52_726 ();
 b15zdnd11an1n64x5 FILLER_52_790 ();
 b15zdnd11an1n08x5 FILLER_52_854 ();
 b15zdnd00an1n02x5 FILLER_52_862 ();
 b15zdnd00an1n01x5 FILLER_52_864 ();
 b15zdnd11an1n32x5 FILLER_52_907 ();
 b15zdnd11an1n08x5 FILLER_52_939 ();
 b15zdnd11an1n04x5 FILLER_52_947 ();
 b15zdnd11an1n64x5 FILLER_52_955 ();
 b15zdnd11an1n64x5 FILLER_52_1019 ();
 b15zdnd11an1n64x5 FILLER_52_1083 ();
 b15zdnd11an1n64x5 FILLER_52_1147 ();
 b15zdnd11an1n64x5 FILLER_52_1211 ();
 b15zdnd11an1n64x5 FILLER_52_1275 ();
 b15zdnd11an1n16x5 FILLER_52_1339 ();
 b15zdnd00an1n02x5 FILLER_52_1355 ();
 b15zdnd00an1n01x5 FILLER_52_1357 ();
 b15zdnd11an1n64x5 FILLER_52_1361 ();
 b15zdnd11an1n64x5 FILLER_52_1425 ();
 b15zdnd11an1n64x5 FILLER_52_1489 ();
 b15zdnd11an1n64x5 FILLER_52_1553 ();
 b15zdnd11an1n64x5 FILLER_52_1617 ();
 b15zdnd11an1n64x5 FILLER_52_1681 ();
 b15zdnd11an1n64x5 FILLER_52_1745 ();
 b15zdnd11an1n32x5 FILLER_52_1809 ();
 b15zdnd00an1n02x5 FILLER_52_1841 ();
 b15zdnd00an1n01x5 FILLER_52_1843 ();
 b15zdnd11an1n04x5 FILLER_52_1847 ();
 b15zdnd11an1n04x5 FILLER_52_1854 ();
 b15zdnd11an1n64x5 FILLER_52_1861 ();
 b15zdnd11an1n32x5 FILLER_52_1925 ();
 b15zdnd11an1n04x5 FILLER_52_1957 ();
 b15zdnd00an1n01x5 FILLER_52_1961 ();
 b15zdnd11an1n64x5 FILLER_52_1965 ();
 b15zdnd11an1n64x5 FILLER_52_2029 ();
 b15zdnd11an1n32x5 FILLER_52_2093 ();
 b15zdnd11an1n16x5 FILLER_52_2125 ();
 b15zdnd11an1n08x5 FILLER_52_2141 ();
 b15zdnd11an1n04x5 FILLER_52_2149 ();
 b15zdnd00an1n01x5 FILLER_52_2153 ();
 b15zdnd11an1n64x5 FILLER_52_2162 ();
 b15zdnd11an1n32x5 FILLER_52_2226 ();
 b15zdnd11an1n16x5 FILLER_52_2258 ();
 b15zdnd00an1n02x5 FILLER_52_2274 ();
 b15zdnd11an1n64x5 FILLER_53_0 ();
 b15zdnd11an1n64x5 FILLER_53_64 ();
 b15zdnd11an1n64x5 FILLER_53_128 ();
 b15zdnd11an1n64x5 FILLER_53_192 ();
 b15zdnd11an1n64x5 FILLER_53_256 ();
 b15zdnd11an1n64x5 FILLER_53_320 ();
 b15zdnd11an1n64x5 FILLER_53_384 ();
 b15zdnd11an1n16x5 FILLER_53_448 ();
 b15zdnd11an1n08x5 FILLER_53_464 ();
 b15zdnd00an1n02x5 FILLER_53_472 ();
 b15zdnd00an1n01x5 FILLER_53_474 ();
 b15zdnd11an1n64x5 FILLER_53_500 ();
 b15zdnd11an1n32x5 FILLER_53_564 ();
 b15zdnd11an1n04x5 FILLER_53_596 ();
 b15zdnd11an1n08x5 FILLER_53_618 ();
 b15zdnd00an1n02x5 FILLER_53_626 ();
 b15zdnd11an1n64x5 FILLER_53_670 ();
 b15zdnd11an1n64x5 FILLER_53_734 ();
 b15zdnd11an1n64x5 FILLER_53_798 ();
 b15zdnd11an1n64x5 FILLER_53_862 ();
 b15zdnd11an1n64x5 FILLER_53_926 ();
 b15zdnd11an1n32x5 FILLER_53_990 ();
 b15zdnd11an1n08x5 FILLER_53_1022 ();
 b15zdnd11an1n04x5 FILLER_53_1030 ();
 b15zdnd00an1n01x5 FILLER_53_1034 ();
 b15zdnd11an1n64x5 FILLER_53_1039 ();
 b15zdnd11an1n64x5 FILLER_53_1103 ();
 b15zdnd00an1n02x5 FILLER_53_1167 ();
 b15zdnd00an1n01x5 FILLER_53_1169 ();
 b15zdnd11an1n64x5 FILLER_53_1173 ();
 b15zdnd11an1n64x5 FILLER_53_1237 ();
 b15zdnd11an1n32x5 FILLER_53_1301 ();
 b15zdnd11an1n16x5 FILLER_53_1333 ();
 b15zdnd11an1n08x5 FILLER_53_1349 ();
 b15zdnd11an1n64x5 FILLER_53_1360 ();
 b15zdnd11an1n64x5 FILLER_53_1424 ();
 b15zdnd11an1n64x5 FILLER_53_1488 ();
 b15zdnd11an1n64x5 FILLER_53_1552 ();
 b15zdnd11an1n64x5 FILLER_53_1616 ();
 b15zdnd11an1n32x5 FILLER_53_1680 ();
 b15zdnd11an1n08x5 FILLER_53_1712 ();
 b15zdnd11an1n04x5 FILLER_53_1720 ();
 b15zdnd00an1n02x5 FILLER_53_1724 ();
 b15zdnd00an1n01x5 FILLER_53_1726 ();
 b15zdnd11an1n64x5 FILLER_53_1735 ();
 b15zdnd11an1n32x5 FILLER_53_1799 ();
 b15zdnd11an1n08x5 FILLER_53_1831 ();
 b15zdnd11an1n04x5 FILLER_53_1839 ();
 b15zdnd00an1n02x5 FILLER_53_1843 ();
 b15zdnd00an1n01x5 FILLER_53_1845 ();
 b15zdnd11an1n64x5 FILLER_53_1849 ();
 b15zdnd11an1n64x5 FILLER_53_1913 ();
 b15zdnd11an1n64x5 FILLER_53_1977 ();
 b15zdnd11an1n64x5 FILLER_53_2041 ();
 b15zdnd11an1n64x5 FILLER_53_2105 ();
 b15zdnd11an1n64x5 FILLER_53_2169 ();
 b15zdnd11an1n32x5 FILLER_53_2233 ();
 b15zdnd11an1n16x5 FILLER_53_2265 ();
 b15zdnd00an1n02x5 FILLER_53_2281 ();
 b15zdnd00an1n01x5 FILLER_53_2283 ();
 b15zdnd11an1n64x5 FILLER_54_8 ();
 b15zdnd11an1n64x5 FILLER_54_72 ();
 b15zdnd11an1n64x5 FILLER_54_136 ();
 b15zdnd11an1n64x5 FILLER_54_200 ();
 b15zdnd11an1n64x5 FILLER_54_264 ();
 b15zdnd11an1n64x5 FILLER_54_328 ();
 b15zdnd11an1n32x5 FILLER_54_392 ();
 b15zdnd11an1n16x5 FILLER_54_424 ();
 b15zdnd11an1n32x5 FILLER_54_451 ();
 b15zdnd11an1n08x5 FILLER_54_483 ();
 b15zdnd11an1n04x5 FILLER_54_491 ();
 b15zdnd11an1n32x5 FILLER_54_535 ();
 b15zdnd11an1n08x5 FILLER_54_567 ();
 b15zdnd11an1n04x5 FILLER_54_575 ();
 b15zdnd00an1n02x5 FILLER_54_579 ();
 b15zdnd11an1n16x5 FILLER_54_623 ();
 b15zdnd11an1n08x5 FILLER_54_639 ();
 b15zdnd11an1n04x5 FILLER_54_647 ();
 b15zdnd00an1n02x5 FILLER_54_651 ();
 b15zdnd00an1n01x5 FILLER_54_653 ();
 b15zdnd11an1n16x5 FILLER_54_696 ();
 b15zdnd11an1n04x5 FILLER_54_712 ();
 b15zdnd00an1n02x5 FILLER_54_716 ();
 b15zdnd11an1n64x5 FILLER_54_726 ();
 b15zdnd11an1n04x5 FILLER_54_790 ();
 b15zdnd11an1n64x5 FILLER_54_834 ();
 b15zdnd11an1n64x5 FILLER_54_898 ();
 b15zdnd11an1n64x5 FILLER_54_962 ();
 b15zdnd11an1n64x5 FILLER_54_1026 ();
 b15zdnd11an1n64x5 FILLER_54_1090 ();
 b15zdnd11an1n16x5 FILLER_54_1154 ();
 b15zdnd00an1n02x5 FILLER_54_1170 ();
 b15zdnd11an1n64x5 FILLER_54_1186 ();
 b15zdnd11an1n64x5 FILLER_54_1250 ();
 b15zdnd11an1n16x5 FILLER_54_1314 ();
 b15zdnd11an1n08x5 FILLER_54_1330 ();
 b15zdnd11an1n64x5 FILLER_54_1382 ();
 b15zdnd11an1n64x5 FILLER_54_1446 ();
 b15zdnd11an1n64x5 FILLER_54_1510 ();
 b15zdnd11an1n64x5 FILLER_54_1574 ();
 b15zdnd11an1n64x5 FILLER_54_1638 ();
 b15zdnd11an1n64x5 FILLER_54_1702 ();
 b15zdnd11an1n64x5 FILLER_54_1766 ();
 b15zdnd11an1n32x5 FILLER_54_1830 ();
 b15zdnd11an1n08x5 FILLER_54_1862 ();
 b15zdnd11an1n04x5 FILLER_54_1870 ();
 b15zdnd00an1n02x5 FILLER_54_1874 ();
 b15zdnd00an1n01x5 FILLER_54_1876 ();
 b15zdnd11an1n32x5 FILLER_54_1886 ();
 b15zdnd11an1n08x5 FILLER_54_1918 ();
 b15zdnd11an1n04x5 FILLER_54_1926 ();
 b15zdnd00an1n02x5 FILLER_54_1930 ();
 b15zdnd11an1n64x5 FILLER_54_1941 ();
 b15zdnd11an1n32x5 FILLER_54_2005 ();
 b15zdnd11an1n08x5 FILLER_54_2037 ();
 b15zdnd11an1n04x5 FILLER_54_2045 ();
 b15zdnd00an1n01x5 FILLER_54_2049 ();
 b15zdnd11an1n64x5 FILLER_54_2054 ();
 b15zdnd11an1n32x5 FILLER_54_2118 ();
 b15zdnd11an1n04x5 FILLER_54_2150 ();
 b15zdnd11an1n64x5 FILLER_54_2162 ();
 b15zdnd11an1n32x5 FILLER_54_2226 ();
 b15zdnd11an1n16x5 FILLER_54_2258 ();
 b15zdnd00an1n02x5 FILLER_54_2274 ();
 b15zdnd11an1n64x5 FILLER_55_0 ();
 b15zdnd11an1n64x5 FILLER_55_64 ();
 b15zdnd11an1n32x5 FILLER_55_128 ();
 b15zdnd11an1n16x5 FILLER_55_160 ();
 b15zdnd11an1n08x5 FILLER_55_176 ();
 b15zdnd11an1n04x5 FILLER_55_184 ();
 b15zdnd00an1n02x5 FILLER_55_188 ();
 b15zdnd11an1n64x5 FILLER_55_194 ();
 b15zdnd11an1n64x5 FILLER_55_258 ();
 b15zdnd11an1n64x5 FILLER_55_322 ();
 b15zdnd11an1n64x5 FILLER_55_386 ();
 b15zdnd11an1n64x5 FILLER_55_450 ();
 b15zdnd11an1n08x5 FILLER_55_514 ();
 b15zdnd11an1n04x5 FILLER_55_522 ();
 b15zdnd11an1n04x5 FILLER_55_529 ();
 b15zdnd11an1n64x5 FILLER_55_536 ();
 b15zdnd11an1n64x5 FILLER_55_600 ();
 b15zdnd11an1n08x5 FILLER_55_664 ();
 b15zdnd11an1n04x5 FILLER_55_672 ();
 b15zdnd00an1n01x5 FILLER_55_676 ();
 b15zdnd11an1n64x5 FILLER_55_695 ();
 b15zdnd11an1n64x5 FILLER_55_759 ();
 b15zdnd11an1n64x5 FILLER_55_823 ();
 b15zdnd11an1n64x5 FILLER_55_887 ();
 b15zdnd11an1n64x5 FILLER_55_951 ();
 b15zdnd11an1n16x5 FILLER_55_1015 ();
 b15zdnd11an1n08x5 FILLER_55_1031 ();
 b15zdnd00an1n01x5 FILLER_55_1039 ();
 b15zdnd11an1n64x5 FILLER_55_1058 ();
 b15zdnd11an1n04x5 FILLER_55_1122 ();
 b15zdnd00an1n02x5 FILLER_55_1126 ();
 b15zdnd11an1n64x5 FILLER_55_1134 ();
 b15zdnd11an1n16x5 FILLER_55_1198 ();
 b15zdnd11an1n08x5 FILLER_55_1214 ();
 b15zdnd11an1n04x5 FILLER_55_1222 ();
 b15zdnd00an1n01x5 FILLER_55_1226 ();
 b15zdnd11an1n04x5 FILLER_55_1230 ();
 b15zdnd00an1n02x5 FILLER_55_1234 ();
 b15zdnd00an1n01x5 FILLER_55_1236 ();
 b15zdnd11an1n64x5 FILLER_55_1240 ();
 b15zdnd11an1n32x5 FILLER_55_1304 ();
 b15zdnd11an1n16x5 FILLER_55_1336 ();
 b15zdnd11an1n04x5 FILLER_55_1352 ();
 b15zdnd00an1n02x5 FILLER_55_1356 ();
 b15zdnd00an1n01x5 FILLER_55_1358 ();
 b15zdnd11an1n16x5 FILLER_55_1362 ();
 b15zdnd11an1n08x5 FILLER_55_1378 ();
 b15zdnd00an1n01x5 FILLER_55_1386 ();
 b15zdnd11an1n64x5 FILLER_55_1407 ();
 b15zdnd11an1n64x5 FILLER_55_1471 ();
 b15zdnd11an1n64x5 FILLER_55_1535 ();
 b15zdnd11an1n64x5 FILLER_55_1599 ();
 b15zdnd11an1n16x5 FILLER_55_1663 ();
 b15zdnd11an1n04x5 FILLER_55_1679 ();
 b15zdnd00an1n02x5 FILLER_55_1683 ();
 b15zdnd11an1n64x5 FILLER_55_1693 ();
 b15zdnd11an1n64x5 FILLER_55_1757 ();
 b15zdnd11an1n64x5 FILLER_55_1821 ();
 b15zdnd11an1n64x5 FILLER_55_1885 ();
 b15zdnd11an1n16x5 FILLER_55_1949 ();
 b15zdnd00an1n02x5 FILLER_55_1965 ();
 b15zdnd11an1n64x5 FILLER_55_1970 ();
 b15zdnd11an1n64x5 FILLER_55_2034 ();
 b15zdnd11an1n64x5 FILLER_55_2098 ();
 b15zdnd11an1n64x5 FILLER_55_2162 ();
 b15zdnd11an1n32x5 FILLER_55_2226 ();
 b15zdnd11an1n16x5 FILLER_55_2258 ();
 b15zdnd11an1n08x5 FILLER_55_2274 ();
 b15zdnd00an1n02x5 FILLER_55_2282 ();
 b15zdnd11an1n64x5 FILLER_56_8 ();
 b15zdnd11an1n64x5 FILLER_56_72 ();
 b15zdnd11an1n32x5 FILLER_56_136 ();
 b15zdnd11an1n16x5 FILLER_56_168 ();
 b15zdnd11an1n04x5 FILLER_56_184 ();
 b15zdnd11an1n64x5 FILLER_56_194 ();
 b15zdnd11an1n64x5 FILLER_56_258 ();
 b15zdnd11an1n64x5 FILLER_56_322 ();
 b15zdnd11an1n64x5 FILLER_56_386 ();
 b15zdnd11an1n64x5 FILLER_56_450 ();
 b15zdnd11an1n64x5 FILLER_56_514 ();
 b15zdnd11an1n64x5 FILLER_56_578 ();
 b15zdnd11an1n32x5 FILLER_56_642 ();
 b15zdnd00an1n02x5 FILLER_56_716 ();
 b15zdnd11an1n32x5 FILLER_56_726 ();
 b15zdnd11an1n16x5 FILLER_56_758 ();
 b15zdnd11an1n08x5 FILLER_56_774 ();
 b15zdnd11an1n04x5 FILLER_56_782 ();
 b15zdnd00an1n01x5 FILLER_56_786 ();
 b15zdnd11an1n64x5 FILLER_56_795 ();
 b15zdnd11an1n64x5 FILLER_56_859 ();
 b15zdnd00an1n02x5 FILLER_56_923 ();
 b15zdnd00an1n01x5 FILLER_56_925 ();
 b15zdnd11an1n08x5 FILLER_56_930 ();
 b15zdnd00an1n01x5 FILLER_56_938 ();
 b15zdnd11an1n64x5 FILLER_56_943 ();
 b15zdnd11an1n32x5 FILLER_56_1007 ();
 b15zdnd11an1n16x5 FILLER_56_1039 ();
 b15zdnd11an1n04x5 FILLER_56_1055 ();
 b15zdnd00an1n02x5 FILLER_56_1059 ();
 b15zdnd11an1n64x5 FILLER_56_1075 ();
 b15zdnd11an1n32x5 FILLER_56_1139 ();
 b15zdnd00an1n02x5 FILLER_56_1171 ();
 b15zdnd11an1n08x5 FILLER_56_1176 ();
 b15zdnd11an1n04x5 FILLER_56_1184 ();
 b15zdnd00an1n02x5 FILLER_56_1188 ();
 b15zdnd00an1n01x5 FILLER_56_1190 ();
 b15zdnd11an1n16x5 FILLER_56_1207 ();
 b15zdnd00an1n02x5 FILLER_56_1223 ();
 b15zdnd00an1n01x5 FILLER_56_1225 ();
 b15zdnd11an1n64x5 FILLER_56_1233 ();
 b15zdnd11an1n64x5 FILLER_56_1297 ();
 b15zdnd11an1n64x5 FILLER_56_1361 ();
 b15zdnd11an1n64x5 FILLER_56_1425 ();
 b15zdnd11an1n64x5 FILLER_56_1489 ();
 b15zdnd11an1n64x5 FILLER_56_1553 ();
 b15zdnd11an1n64x5 FILLER_56_1617 ();
 b15zdnd11an1n64x5 FILLER_56_1681 ();
 b15zdnd11an1n64x5 FILLER_56_1745 ();
 b15zdnd11an1n64x5 FILLER_56_1809 ();
 b15zdnd11an1n64x5 FILLER_56_1873 ();
 b15zdnd11an1n16x5 FILLER_56_1937 ();
 b15zdnd11an1n08x5 FILLER_56_1953 ();
 b15zdnd11an1n04x5 FILLER_56_1961 ();
 b15zdnd00an1n02x5 FILLER_56_1965 ();
 b15zdnd00an1n01x5 FILLER_56_1967 ();
 b15zdnd11an1n64x5 FILLER_56_1971 ();
 b15zdnd11an1n64x5 FILLER_56_2035 ();
 b15zdnd11an1n32x5 FILLER_56_2099 ();
 b15zdnd11an1n16x5 FILLER_56_2131 ();
 b15zdnd11an1n04x5 FILLER_56_2147 ();
 b15zdnd00an1n02x5 FILLER_56_2151 ();
 b15zdnd00an1n01x5 FILLER_56_2153 ();
 b15zdnd11an1n64x5 FILLER_56_2162 ();
 b15zdnd11an1n32x5 FILLER_56_2226 ();
 b15zdnd11an1n16x5 FILLER_56_2258 ();
 b15zdnd00an1n02x5 FILLER_56_2274 ();
 b15zdnd11an1n64x5 FILLER_57_0 ();
 b15zdnd11an1n64x5 FILLER_57_64 ();
 b15zdnd11an1n32x5 FILLER_57_128 ();
 b15zdnd11an1n16x5 FILLER_57_160 ();
 b15zdnd11an1n04x5 FILLER_57_176 ();
 b15zdnd00an1n02x5 FILLER_57_180 ();
 b15zdnd00an1n01x5 FILLER_57_182 ();
 b15zdnd11an1n04x5 FILLER_57_188 ();
 b15zdnd11an1n64x5 FILLER_57_195 ();
 b15zdnd11an1n64x5 FILLER_57_259 ();
 b15zdnd11an1n16x5 FILLER_57_323 ();
 b15zdnd00an1n01x5 FILLER_57_339 ();
 b15zdnd11an1n32x5 FILLER_57_344 ();
 b15zdnd11an1n16x5 FILLER_57_376 ();
 b15zdnd00an1n02x5 FILLER_57_392 ();
 b15zdnd00an1n01x5 FILLER_57_394 ();
 b15zdnd11an1n64x5 FILLER_57_406 ();
 b15zdnd11an1n64x5 FILLER_57_470 ();
 b15zdnd11an1n64x5 FILLER_57_534 ();
 b15zdnd11an1n64x5 FILLER_57_598 ();
 b15zdnd11an1n64x5 FILLER_57_662 ();
 b15zdnd11an1n64x5 FILLER_57_726 ();
 b15zdnd11an1n64x5 FILLER_57_790 ();
 b15zdnd11an1n64x5 FILLER_57_854 ();
 b15zdnd11an1n16x5 FILLER_57_918 ();
 b15zdnd00an1n02x5 FILLER_57_934 ();
 b15zdnd11an1n04x5 FILLER_57_940 ();
 b15zdnd11an1n64x5 FILLER_57_965 ();
 b15zdnd11an1n32x5 FILLER_57_1029 ();
 b15zdnd11an1n08x5 FILLER_57_1061 ();
 b15zdnd11an1n04x5 FILLER_57_1069 ();
 b15zdnd11an1n64x5 FILLER_57_1081 ();
 b15zdnd11an1n64x5 FILLER_57_1145 ();
 b15zdnd11an1n04x5 FILLER_57_1209 ();
 b15zdnd00an1n02x5 FILLER_57_1213 ();
 b15zdnd11an1n64x5 FILLER_57_1229 ();
 b15zdnd11an1n64x5 FILLER_57_1293 ();
 b15zdnd11an1n64x5 FILLER_57_1357 ();
 b15zdnd11an1n64x5 FILLER_57_1421 ();
 b15zdnd11an1n64x5 FILLER_57_1485 ();
 b15zdnd11an1n08x5 FILLER_57_1549 ();
 b15zdnd11an1n04x5 FILLER_57_1557 ();
 b15zdnd00an1n02x5 FILLER_57_1561 ();
 b15zdnd00an1n01x5 FILLER_57_1563 ();
 b15zdnd11an1n64x5 FILLER_57_1572 ();
 b15zdnd11an1n64x5 FILLER_57_1636 ();
 b15zdnd11an1n64x5 FILLER_57_1700 ();
 b15zdnd11an1n64x5 FILLER_57_1764 ();
 b15zdnd11an1n64x5 FILLER_57_1828 ();
 b15zdnd11an1n32x5 FILLER_57_1892 ();
 b15zdnd11an1n16x5 FILLER_57_1924 ();
 b15zdnd00an1n02x5 FILLER_57_1940 ();
 b15zdnd00an1n01x5 FILLER_57_1942 ();
 b15zdnd11an1n64x5 FILLER_57_1995 ();
 b15zdnd11an1n64x5 FILLER_57_2059 ();
 b15zdnd11an1n64x5 FILLER_57_2123 ();
 b15zdnd11an1n64x5 FILLER_57_2187 ();
 b15zdnd11an1n32x5 FILLER_57_2251 ();
 b15zdnd00an1n01x5 FILLER_57_2283 ();
 b15zdnd11an1n64x5 FILLER_58_8 ();
 b15zdnd11an1n64x5 FILLER_58_72 ();
 b15zdnd11an1n32x5 FILLER_58_136 ();
 b15zdnd11an1n16x5 FILLER_58_168 ();
 b15zdnd00an1n01x5 FILLER_58_184 ();
 b15zdnd11an1n64x5 FILLER_58_195 ();
 b15zdnd11an1n64x5 FILLER_58_259 ();
 b15zdnd00an1n02x5 FILLER_58_323 ();
 b15zdnd00an1n01x5 FILLER_58_325 ();
 b15zdnd11an1n32x5 FILLER_58_332 ();
 b15zdnd11an1n08x5 FILLER_58_364 ();
 b15zdnd11an1n04x5 FILLER_58_372 ();
 b15zdnd00an1n02x5 FILLER_58_376 ();
 b15zdnd00an1n01x5 FILLER_58_378 ();
 b15zdnd11an1n64x5 FILLER_58_385 ();
 b15zdnd11an1n64x5 FILLER_58_449 ();
 b15zdnd11an1n64x5 FILLER_58_513 ();
 b15zdnd11an1n64x5 FILLER_58_577 ();
 b15zdnd11an1n64x5 FILLER_58_641 ();
 b15zdnd11an1n08x5 FILLER_58_705 ();
 b15zdnd11an1n04x5 FILLER_58_713 ();
 b15zdnd00an1n01x5 FILLER_58_717 ();
 b15zdnd11an1n64x5 FILLER_58_726 ();
 b15zdnd11an1n32x5 FILLER_58_790 ();
 b15zdnd11an1n16x5 FILLER_58_822 ();
 b15zdnd00an1n01x5 FILLER_58_838 ();
 b15zdnd11an1n08x5 FILLER_58_842 ();
 b15zdnd00an1n02x5 FILLER_58_850 ();
 b15zdnd11an1n64x5 FILLER_58_868 ();
 b15zdnd11an1n64x5 FILLER_58_932 ();
 b15zdnd11an1n64x5 FILLER_58_996 ();
 b15zdnd11an1n32x5 FILLER_58_1060 ();
 b15zdnd11an1n04x5 FILLER_58_1092 ();
 b15zdnd00an1n02x5 FILLER_58_1096 ();
 b15zdnd11an1n64x5 FILLER_58_1118 ();
 b15zdnd11an1n16x5 FILLER_58_1182 ();
 b15zdnd11an1n08x5 FILLER_58_1198 ();
 b15zdnd00an1n01x5 FILLER_58_1206 ();
 b15zdnd11an1n04x5 FILLER_58_1224 ();
 b15zdnd11an1n64x5 FILLER_58_1270 ();
 b15zdnd11an1n64x5 FILLER_58_1334 ();
 b15zdnd11an1n64x5 FILLER_58_1398 ();
 b15zdnd11an1n64x5 FILLER_58_1462 ();
 b15zdnd11an1n64x5 FILLER_58_1526 ();
 b15zdnd11an1n64x5 FILLER_58_1590 ();
 b15zdnd11an1n64x5 FILLER_58_1654 ();
 b15zdnd11an1n64x5 FILLER_58_1718 ();
 b15zdnd11an1n32x5 FILLER_58_1782 ();
 b15zdnd11an1n16x5 FILLER_58_1814 ();
 b15zdnd11an1n32x5 FILLER_58_1857 ();
 b15zdnd11an1n16x5 FILLER_58_1889 ();
 b15zdnd11an1n08x5 FILLER_58_1905 ();
 b15zdnd11an1n04x5 FILLER_58_1913 ();
 b15zdnd00an1n02x5 FILLER_58_1917 ();
 b15zdnd11an1n32x5 FILLER_58_1928 ();
 b15zdnd11an1n08x5 FILLER_58_1960 ();
 b15zdnd11an1n64x5 FILLER_58_1971 ();
 b15zdnd11an1n64x5 FILLER_58_2035 ();
 b15zdnd11an1n32x5 FILLER_58_2099 ();
 b15zdnd11an1n16x5 FILLER_58_2131 ();
 b15zdnd11an1n04x5 FILLER_58_2147 ();
 b15zdnd00an1n02x5 FILLER_58_2151 ();
 b15zdnd00an1n01x5 FILLER_58_2153 ();
 b15zdnd11an1n64x5 FILLER_58_2162 ();
 b15zdnd11an1n32x5 FILLER_58_2226 ();
 b15zdnd11an1n16x5 FILLER_58_2258 ();
 b15zdnd00an1n02x5 FILLER_58_2274 ();
 b15zdnd11an1n64x5 FILLER_59_0 ();
 b15zdnd11an1n64x5 FILLER_59_64 ();
 b15zdnd11an1n32x5 FILLER_59_128 ();
 b15zdnd11an1n16x5 FILLER_59_160 ();
 b15zdnd11an1n04x5 FILLER_59_186 ();
 b15zdnd11an1n04x5 FILLER_59_201 ();
 b15zdnd11an1n32x5 FILLER_59_247 ();
 b15zdnd11an1n16x5 FILLER_59_279 ();
 b15zdnd00an1n02x5 FILLER_59_295 ();
 b15zdnd00an1n01x5 FILLER_59_297 ();
 b15zdnd11an1n16x5 FILLER_59_301 ();
 b15zdnd11an1n08x5 FILLER_59_317 ();
 b15zdnd11an1n04x5 FILLER_59_325 ();
 b15zdnd00an1n01x5 FILLER_59_329 ();
 b15zdnd11an1n64x5 FILLER_59_342 ();
 b15zdnd11an1n32x5 FILLER_59_406 ();
 b15zdnd11an1n16x5 FILLER_59_438 ();
 b15zdnd11an1n64x5 FILLER_59_457 ();
 b15zdnd11an1n64x5 FILLER_59_521 ();
 b15zdnd11an1n64x5 FILLER_59_585 ();
 b15zdnd11an1n64x5 FILLER_59_649 ();
 b15zdnd11an1n64x5 FILLER_59_713 ();
 b15zdnd11an1n32x5 FILLER_59_777 ();
 b15zdnd11an1n16x5 FILLER_59_809 ();
 b15zdnd11an1n08x5 FILLER_59_825 ();
 b15zdnd00an1n02x5 FILLER_59_833 ();
 b15zdnd00an1n01x5 FILLER_59_835 ();
 b15zdnd11an1n08x5 FILLER_59_839 ();
 b15zdnd00an1n02x5 FILLER_59_847 ();
 b15zdnd11an1n64x5 FILLER_59_852 ();
 b15zdnd11an1n64x5 FILLER_59_916 ();
 b15zdnd11an1n64x5 FILLER_59_980 ();
 b15zdnd11an1n32x5 FILLER_59_1044 ();
 b15zdnd11an1n16x5 FILLER_59_1076 ();
 b15zdnd11an1n04x5 FILLER_59_1092 ();
 b15zdnd00an1n01x5 FILLER_59_1096 ();
 b15zdnd11an1n64x5 FILLER_59_1109 ();
 b15zdnd11an1n32x5 FILLER_59_1173 ();
 b15zdnd11an1n16x5 FILLER_59_1205 ();
 b15zdnd11an1n08x5 FILLER_59_1221 ();
 b15zdnd00an1n02x5 FILLER_59_1229 ();
 b15zdnd11an1n32x5 FILLER_59_1244 ();
 b15zdnd11an1n64x5 FILLER_59_1280 ();
 b15zdnd11an1n32x5 FILLER_59_1344 ();
 b15zdnd11an1n16x5 FILLER_59_1376 ();
 b15zdnd11an1n04x5 FILLER_59_1392 ();
 b15zdnd00an1n02x5 FILLER_59_1396 ();
 b15zdnd11an1n04x5 FILLER_59_1426 ();
 b15zdnd11an1n64x5 FILLER_59_1433 ();
 b15zdnd11an1n64x5 FILLER_59_1497 ();
 b15zdnd11an1n64x5 FILLER_59_1561 ();
 b15zdnd11an1n64x5 FILLER_59_1625 ();
 b15zdnd11an1n64x5 FILLER_59_1689 ();
 b15zdnd11an1n64x5 FILLER_59_1753 ();
 b15zdnd11an1n08x5 FILLER_59_1817 ();
 b15zdnd11an1n04x5 FILLER_59_1825 ();
 b15zdnd00an1n01x5 FILLER_59_1829 ();
 b15zdnd11an1n64x5 FILLER_59_1833 ();
 b15zdnd11an1n64x5 FILLER_59_1897 ();
 b15zdnd11an1n64x5 FILLER_59_1961 ();
 b15zdnd11an1n64x5 FILLER_59_2025 ();
 b15zdnd11an1n64x5 FILLER_59_2089 ();
 b15zdnd11an1n64x5 FILLER_59_2153 ();
 b15zdnd11an1n64x5 FILLER_59_2217 ();
 b15zdnd00an1n02x5 FILLER_59_2281 ();
 b15zdnd00an1n01x5 FILLER_59_2283 ();
 b15zdnd11an1n64x5 FILLER_60_8 ();
 b15zdnd11an1n64x5 FILLER_60_72 ();
 b15zdnd11an1n32x5 FILLER_60_136 ();
 b15zdnd11an1n32x5 FILLER_60_220 ();
 b15zdnd11an1n16x5 FILLER_60_252 ();
 b15zdnd11an1n04x5 FILLER_60_268 ();
 b15zdnd00an1n02x5 FILLER_60_272 ();
 b15zdnd11an1n08x5 FILLER_60_326 ();
 b15zdnd00an1n02x5 FILLER_60_334 ();
 b15zdnd00an1n01x5 FILLER_60_336 ();
 b15zdnd11an1n04x5 FILLER_60_350 ();
 b15zdnd11an1n32x5 FILLER_60_357 ();
 b15zdnd11an1n16x5 FILLER_60_389 ();
 b15zdnd11an1n08x5 FILLER_60_405 ();
 b15zdnd11an1n04x5 FILLER_60_413 ();
 b15zdnd00an1n02x5 FILLER_60_417 ();
 b15zdnd00an1n01x5 FILLER_60_419 ();
 b15zdnd11an1n04x5 FILLER_60_423 ();
 b15zdnd11an1n64x5 FILLER_60_479 ();
 b15zdnd11an1n64x5 FILLER_60_543 ();
 b15zdnd11an1n04x5 FILLER_60_607 ();
 b15zdnd00an1n01x5 FILLER_60_611 ();
 b15zdnd11an1n64x5 FILLER_60_654 ();
 b15zdnd11an1n64x5 FILLER_60_726 ();
 b15zdnd11an1n16x5 FILLER_60_790 ();
 b15zdnd11an1n08x5 FILLER_60_806 ();
 b15zdnd00an1n01x5 FILLER_60_814 ();
 b15zdnd11an1n64x5 FILLER_60_859 ();
 b15zdnd11an1n64x5 FILLER_60_923 ();
 b15zdnd11an1n32x5 FILLER_60_987 ();
 b15zdnd11an1n04x5 FILLER_60_1019 ();
 b15zdnd00an1n02x5 FILLER_60_1023 ();
 b15zdnd00an1n01x5 FILLER_60_1025 ();
 b15zdnd11an1n64x5 FILLER_60_1030 ();
 b15zdnd11an1n64x5 FILLER_60_1094 ();
 b15zdnd11an1n32x5 FILLER_60_1158 ();
 b15zdnd00an1n02x5 FILLER_60_1190 ();
 b15zdnd11an1n32x5 FILLER_60_1199 ();
 b15zdnd11an1n08x5 FILLER_60_1231 ();
 b15zdnd00an1n01x5 FILLER_60_1239 ();
 b15zdnd11an1n64x5 FILLER_60_1254 ();
 b15zdnd11an1n64x5 FILLER_60_1318 ();
 b15zdnd11an1n08x5 FILLER_60_1382 ();
 b15zdnd11an1n04x5 FILLER_60_1390 ();
 b15zdnd00an1n02x5 FILLER_60_1394 ();
 b15zdnd11an1n32x5 FILLER_60_1438 ();
 b15zdnd11an1n16x5 FILLER_60_1470 ();
 b15zdnd11an1n08x5 FILLER_60_1486 ();
 b15zdnd00an1n01x5 FILLER_60_1494 ();
 b15zdnd11an1n64x5 FILLER_60_1499 ();
 b15zdnd11an1n64x5 FILLER_60_1563 ();
 b15zdnd11an1n64x5 FILLER_60_1627 ();
 b15zdnd11an1n64x5 FILLER_60_1691 ();
 b15zdnd11an1n64x5 FILLER_60_1755 ();
 b15zdnd11an1n64x5 FILLER_60_1819 ();
 b15zdnd11an1n64x5 FILLER_60_1883 ();
 b15zdnd11an1n64x5 FILLER_60_1947 ();
 b15zdnd11an1n64x5 FILLER_60_2011 ();
 b15zdnd11an1n64x5 FILLER_60_2075 ();
 b15zdnd11an1n08x5 FILLER_60_2139 ();
 b15zdnd11an1n04x5 FILLER_60_2147 ();
 b15zdnd00an1n02x5 FILLER_60_2151 ();
 b15zdnd00an1n01x5 FILLER_60_2153 ();
 b15zdnd11an1n64x5 FILLER_60_2162 ();
 b15zdnd11an1n32x5 FILLER_60_2226 ();
 b15zdnd11an1n16x5 FILLER_60_2258 ();
 b15zdnd00an1n02x5 FILLER_60_2274 ();
 b15zdnd11an1n64x5 FILLER_61_0 ();
 b15zdnd11an1n64x5 FILLER_61_64 ();
 b15zdnd11an1n32x5 FILLER_61_128 ();
 b15zdnd11an1n08x5 FILLER_61_160 ();
 b15zdnd11an1n04x5 FILLER_61_168 ();
 b15zdnd00an1n01x5 FILLER_61_172 ();
 b15zdnd11an1n04x5 FILLER_61_178 ();
 b15zdnd11an1n04x5 FILLER_61_185 ();
 b15zdnd11an1n64x5 FILLER_61_231 ();
 b15zdnd00an1n02x5 FILLER_61_295 ();
 b15zdnd11an1n08x5 FILLER_61_300 ();
 b15zdnd11an1n04x5 FILLER_61_308 ();
 b15zdnd00an1n02x5 FILLER_61_312 ();
 b15zdnd11an1n04x5 FILLER_61_324 ();
 b15zdnd11an1n04x5 FILLER_61_370 ();
 b15zdnd11an1n16x5 FILLER_61_381 ();
 b15zdnd11an1n04x5 FILLER_61_397 ();
 b15zdnd11an1n08x5 FILLER_61_443 ();
 b15zdnd00an1n02x5 FILLER_61_451 ();
 b15zdnd11an1n04x5 FILLER_61_456 ();
 b15zdnd11an1n64x5 FILLER_61_463 ();
 b15zdnd11an1n64x5 FILLER_61_527 ();
 b15zdnd11an1n64x5 FILLER_61_591 ();
 b15zdnd11an1n64x5 FILLER_61_655 ();
 b15zdnd00an1n01x5 FILLER_61_719 ();
 b15zdnd11an1n64x5 FILLER_61_723 ();
 b15zdnd11an1n64x5 FILLER_61_787 ();
 b15zdnd11an1n64x5 FILLER_61_851 ();
 b15zdnd11an1n64x5 FILLER_61_915 ();
 b15zdnd11an1n64x5 FILLER_61_979 ();
 b15zdnd11an1n64x5 FILLER_61_1043 ();
 b15zdnd11an1n32x5 FILLER_61_1107 ();
 b15zdnd11an1n16x5 FILLER_61_1139 ();
 b15zdnd00an1n01x5 FILLER_61_1155 ();
 b15zdnd11an1n32x5 FILLER_61_1159 ();
 b15zdnd11an1n08x5 FILLER_61_1191 ();
 b15zdnd00an1n02x5 FILLER_61_1199 ();
 b15zdnd00an1n01x5 FILLER_61_1201 ();
 b15zdnd11an1n64x5 FILLER_61_1208 ();
 b15zdnd11an1n16x5 FILLER_61_1272 ();
 b15zdnd11an1n04x5 FILLER_61_1288 ();
 b15zdnd11an1n64x5 FILLER_61_1302 ();
 b15zdnd11an1n16x5 FILLER_61_1366 ();
 b15zdnd11an1n08x5 FILLER_61_1382 ();
 b15zdnd11an1n08x5 FILLER_61_1407 ();
 b15zdnd11an1n04x5 FILLER_61_1415 ();
 b15zdnd00an1n02x5 FILLER_61_1419 ();
 b15zdnd00an1n01x5 FILLER_61_1421 ();
 b15zdnd11an1n64x5 FILLER_61_1425 ();
 b15zdnd11an1n16x5 FILLER_61_1489 ();
 b15zdnd11an1n04x5 FILLER_61_1505 ();
 b15zdnd00an1n02x5 FILLER_61_1509 ();
 b15zdnd11an1n32x5 FILLER_61_1528 ();
 b15zdnd11an1n16x5 FILLER_61_1560 ();
 b15zdnd11an1n04x5 FILLER_61_1576 ();
 b15zdnd00an1n01x5 FILLER_61_1580 ();
 b15zdnd11an1n64x5 FILLER_61_1585 ();
 b15zdnd11an1n64x5 FILLER_61_1649 ();
 b15zdnd11an1n64x5 FILLER_61_1713 ();
 b15zdnd11an1n64x5 FILLER_61_1777 ();
 b15zdnd11an1n64x5 FILLER_61_1841 ();
 b15zdnd11an1n32x5 FILLER_61_1905 ();
 b15zdnd11an1n04x5 FILLER_61_1937 ();
 b15zdnd00an1n02x5 FILLER_61_1941 ();
 b15zdnd11an1n64x5 FILLER_61_1946 ();
 b15zdnd11an1n64x5 FILLER_61_2010 ();
 b15zdnd11an1n64x5 FILLER_61_2074 ();
 b15zdnd11an1n64x5 FILLER_61_2138 ();
 b15zdnd11an1n64x5 FILLER_61_2202 ();
 b15zdnd11an1n16x5 FILLER_61_2266 ();
 b15zdnd00an1n02x5 FILLER_61_2282 ();
 b15zdnd11an1n64x5 FILLER_62_8 ();
 b15zdnd11an1n64x5 FILLER_62_72 ();
 b15zdnd11an1n32x5 FILLER_62_136 ();
 b15zdnd11an1n08x5 FILLER_62_168 ();
 b15zdnd11an1n04x5 FILLER_62_176 ();
 b15zdnd00an1n02x5 FILLER_62_180 ();
 b15zdnd11an1n08x5 FILLER_62_191 ();
 b15zdnd00an1n01x5 FILLER_62_199 ();
 b15zdnd11an1n64x5 FILLER_62_207 ();
 b15zdnd11an1n16x5 FILLER_62_271 ();
 b15zdnd11an1n08x5 FILLER_62_287 ();
 b15zdnd00an1n01x5 FILLER_62_295 ();
 b15zdnd11an1n16x5 FILLER_62_299 ();
 b15zdnd11an1n04x5 FILLER_62_315 ();
 b15zdnd00an1n02x5 FILLER_62_319 ();
 b15zdnd11an1n32x5 FILLER_62_363 ();
 b15zdnd00an1n02x5 FILLER_62_395 ();
 b15zdnd11an1n04x5 FILLER_62_449 ();
 b15zdnd11an1n64x5 FILLER_62_495 ();
 b15zdnd11an1n64x5 FILLER_62_559 ();
 b15zdnd11an1n64x5 FILLER_62_623 ();
 b15zdnd11an1n16x5 FILLER_62_687 ();
 b15zdnd11an1n08x5 FILLER_62_703 ();
 b15zdnd11an1n04x5 FILLER_62_711 ();
 b15zdnd00an1n02x5 FILLER_62_715 ();
 b15zdnd00an1n01x5 FILLER_62_717 ();
 b15zdnd11an1n64x5 FILLER_62_726 ();
 b15zdnd11an1n64x5 FILLER_62_790 ();
 b15zdnd11an1n64x5 FILLER_62_854 ();
 b15zdnd11an1n64x5 FILLER_62_918 ();
 b15zdnd11an1n64x5 FILLER_62_982 ();
 b15zdnd11an1n64x5 FILLER_62_1046 ();
 b15zdnd11an1n16x5 FILLER_62_1110 ();
 b15zdnd11an1n08x5 FILLER_62_1126 ();
 b15zdnd11an1n04x5 FILLER_62_1134 ();
 b15zdnd11an1n64x5 FILLER_62_1180 ();
 b15zdnd11an1n32x5 FILLER_62_1244 ();
 b15zdnd00an1n02x5 FILLER_62_1276 ();
 b15zdnd00an1n01x5 FILLER_62_1278 ();
 b15zdnd11an1n32x5 FILLER_62_1285 ();
 b15zdnd00an1n02x5 FILLER_62_1317 ();
 b15zdnd11an1n16x5 FILLER_62_1331 ();
 b15zdnd00an1n02x5 FILLER_62_1347 ();
 b15zdnd11an1n64x5 FILLER_62_1366 ();
 b15zdnd11an1n64x5 FILLER_62_1430 ();
 b15zdnd11an1n64x5 FILLER_62_1494 ();
 b15zdnd11an1n08x5 FILLER_62_1558 ();
 b15zdnd11an1n04x5 FILLER_62_1566 ();
 b15zdnd11an1n64x5 FILLER_62_1574 ();
 b15zdnd11an1n64x5 FILLER_62_1638 ();
 b15zdnd11an1n64x5 FILLER_62_1702 ();
 b15zdnd11an1n64x5 FILLER_62_1766 ();
 b15zdnd11an1n64x5 FILLER_62_1830 ();
 b15zdnd11an1n64x5 FILLER_62_1894 ();
 b15zdnd11an1n16x5 FILLER_62_1958 ();
 b15zdnd11an1n08x5 FILLER_62_1974 ();
 b15zdnd00an1n02x5 FILLER_62_1982 ();
 b15zdnd00an1n01x5 FILLER_62_1984 ();
 b15zdnd11an1n64x5 FILLER_62_1988 ();
 b15zdnd11an1n08x5 FILLER_62_2052 ();
 b15zdnd11an1n04x5 FILLER_62_2060 ();
 b15zdnd00an1n02x5 FILLER_62_2064 ();
 b15zdnd11an1n64x5 FILLER_62_2070 ();
 b15zdnd11an1n16x5 FILLER_62_2134 ();
 b15zdnd11an1n04x5 FILLER_62_2150 ();
 b15zdnd11an1n64x5 FILLER_62_2162 ();
 b15zdnd11an1n32x5 FILLER_62_2226 ();
 b15zdnd11an1n16x5 FILLER_62_2258 ();
 b15zdnd00an1n02x5 FILLER_62_2274 ();
 b15zdnd11an1n64x5 FILLER_63_0 ();
 b15zdnd11an1n64x5 FILLER_63_64 ();
 b15zdnd11an1n32x5 FILLER_63_128 ();
 b15zdnd11an1n16x5 FILLER_63_160 ();
 b15zdnd11an1n08x5 FILLER_63_176 ();
 b15zdnd00an1n02x5 FILLER_63_184 ();
 b15zdnd11an1n04x5 FILLER_63_189 ();
 b15zdnd11an1n64x5 FILLER_63_196 ();
 b15zdnd11an1n64x5 FILLER_63_260 ();
 b15zdnd11an1n04x5 FILLER_63_324 ();
 b15zdnd11an1n04x5 FILLER_63_337 ();
 b15zdnd11an1n64x5 FILLER_63_346 ();
 b15zdnd11an1n04x5 FILLER_63_410 ();
 b15zdnd00an1n01x5 FILLER_63_414 ();
 b15zdnd11an1n04x5 FILLER_63_418 ();
 b15zdnd11an1n64x5 FILLER_63_425 ();
 b15zdnd11an1n64x5 FILLER_63_489 ();
 b15zdnd11an1n32x5 FILLER_63_553 ();
 b15zdnd11an1n64x5 FILLER_63_616 ();
 b15zdnd11an1n64x5 FILLER_63_680 ();
 b15zdnd11an1n64x5 FILLER_63_744 ();
 b15zdnd11an1n64x5 FILLER_63_808 ();
 b15zdnd11an1n64x5 FILLER_63_872 ();
 b15zdnd11an1n64x5 FILLER_63_936 ();
 b15zdnd11an1n64x5 FILLER_63_1000 ();
 b15zdnd11an1n64x5 FILLER_63_1064 ();
 b15zdnd11an1n08x5 FILLER_63_1128 ();
 b15zdnd11an1n04x5 FILLER_63_1136 ();
 b15zdnd00an1n01x5 FILLER_63_1140 ();
 b15zdnd11an1n64x5 FILLER_63_1183 ();
 b15zdnd11an1n32x5 FILLER_63_1247 ();
 b15zdnd11an1n16x5 FILLER_63_1279 ();
 b15zdnd11an1n08x5 FILLER_63_1295 ();
 b15zdnd00an1n02x5 FILLER_63_1303 ();
 b15zdnd00an1n01x5 FILLER_63_1305 ();
 b15zdnd11an1n32x5 FILLER_63_1310 ();
 b15zdnd11an1n08x5 FILLER_63_1342 ();
 b15zdnd11an1n04x5 FILLER_63_1350 ();
 b15zdnd00an1n02x5 FILLER_63_1354 ();
 b15zdnd00an1n01x5 FILLER_63_1356 ();
 b15zdnd11an1n04x5 FILLER_63_1369 ();
 b15zdnd11an1n64x5 FILLER_63_1379 ();
 b15zdnd11an1n64x5 FILLER_63_1443 ();
 b15zdnd11an1n04x5 FILLER_63_1507 ();
 b15zdnd00an1n02x5 FILLER_63_1511 ();
 b15zdnd00an1n01x5 FILLER_63_1513 ();
 b15zdnd11an1n64x5 FILLER_63_1535 ();
 b15zdnd11an1n64x5 FILLER_63_1599 ();
 b15zdnd11an1n64x5 FILLER_63_1663 ();
 b15zdnd11an1n64x5 FILLER_63_1727 ();
 b15zdnd11an1n64x5 FILLER_63_1791 ();
 b15zdnd11an1n64x5 FILLER_63_1855 ();
 b15zdnd11an1n08x5 FILLER_63_1919 ();
 b15zdnd00an1n02x5 FILLER_63_1927 ();
 b15zdnd00an1n01x5 FILLER_63_1929 ();
 b15zdnd11an1n04x5 FILLER_63_1933 ();
 b15zdnd11an1n32x5 FILLER_63_1940 ();
 b15zdnd00an1n01x5 FILLER_63_1972 ();
 b15zdnd11an1n64x5 FILLER_63_2025 ();
 b15zdnd11an1n64x5 FILLER_63_2089 ();
 b15zdnd11an1n64x5 FILLER_63_2153 ();
 b15zdnd11an1n64x5 FILLER_63_2217 ();
 b15zdnd00an1n02x5 FILLER_63_2281 ();
 b15zdnd00an1n01x5 FILLER_63_2283 ();
 b15zdnd11an1n64x5 FILLER_64_8 ();
 b15zdnd11an1n64x5 FILLER_64_72 ();
 b15zdnd11an1n64x5 FILLER_64_136 ();
 b15zdnd11an1n32x5 FILLER_64_200 ();
 b15zdnd11an1n08x5 FILLER_64_232 ();
 b15zdnd11an1n04x5 FILLER_64_240 ();
 b15zdnd00an1n02x5 FILLER_64_244 ();
 b15zdnd11an1n64x5 FILLER_64_288 ();
 b15zdnd11an1n64x5 FILLER_64_352 ();
 b15zdnd11an1n64x5 FILLER_64_416 ();
 b15zdnd11an1n64x5 FILLER_64_480 ();
 b15zdnd11an1n32x5 FILLER_64_544 ();
 b15zdnd11an1n16x5 FILLER_64_576 ();
 b15zdnd11an1n04x5 FILLER_64_592 ();
 b15zdnd00an1n02x5 FILLER_64_596 ();
 b15zdnd00an1n01x5 FILLER_64_598 ();
 b15zdnd11an1n64x5 FILLER_64_608 ();
 b15zdnd11an1n32x5 FILLER_64_672 ();
 b15zdnd11an1n08x5 FILLER_64_704 ();
 b15zdnd11an1n04x5 FILLER_64_712 ();
 b15zdnd00an1n02x5 FILLER_64_716 ();
 b15zdnd11an1n64x5 FILLER_64_726 ();
 b15zdnd11an1n64x5 FILLER_64_790 ();
 b15zdnd11an1n64x5 FILLER_64_854 ();
 b15zdnd11an1n64x5 FILLER_64_918 ();
 b15zdnd11an1n64x5 FILLER_64_982 ();
 b15zdnd11an1n64x5 FILLER_64_1046 ();
 b15zdnd11an1n08x5 FILLER_64_1110 ();
 b15zdnd00an1n02x5 FILLER_64_1118 ();
 b15zdnd11an1n64x5 FILLER_64_1162 ();
 b15zdnd11an1n08x5 FILLER_64_1226 ();
 b15zdnd11an1n04x5 FILLER_64_1234 ();
 b15zdnd11an1n64x5 FILLER_64_1254 ();
 b15zdnd11an1n16x5 FILLER_64_1318 ();
 b15zdnd11an1n04x5 FILLER_64_1334 ();
 b15zdnd00an1n02x5 FILLER_64_1338 ();
 b15zdnd00an1n01x5 FILLER_64_1340 ();
 b15zdnd11an1n08x5 FILLER_64_1345 ();
 b15zdnd11an1n04x5 FILLER_64_1353 ();
 b15zdnd00an1n02x5 FILLER_64_1357 ();
 b15zdnd11an1n04x5 FILLER_64_1362 ();
 b15zdnd00an1n01x5 FILLER_64_1366 ();
 b15zdnd11an1n08x5 FILLER_64_1381 ();
 b15zdnd00an1n02x5 FILLER_64_1389 ();
 b15zdnd00an1n01x5 FILLER_64_1391 ();
 b15zdnd11an1n16x5 FILLER_64_1395 ();
 b15zdnd11an1n64x5 FILLER_64_1425 ();
 b15zdnd11an1n64x5 FILLER_64_1489 ();
 b15zdnd11an1n64x5 FILLER_64_1553 ();
 b15zdnd11an1n64x5 FILLER_64_1617 ();
 b15zdnd11an1n32x5 FILLER_64_1681 ();
 b15zdnd11an1n16x5 FILLER_64_1713 ();
 b15zdnd11an1n08x5 FILLER_64_1729 ();
 b15zdnd11an1n04x5 FILLER_64_1737 ();
 b15zdnd00an1n02x5 FILLER_64_1741 ();
 b15zdnd00an1n01x5 FILLER_64_1743 ();
 b15zdnd11an1n64x5 FILLER_64_1748 ();
 b15zdnd11an1n08x5 FILLER_64_1812 ();
 b15zdnd11an1n04x5 FILLER_64_1820 ();
 b15zdnd11an1n08x5 FILLER_64_1827 ();
 b15zdnd00an1n02x5 FILLER_64_1835 ();
 b15zdnd00an1n01x5 FILLER_64_1837 ();
 b15zdnd11an1n64x5 FILLER_64_1841 ();
 b15zdnd11an1n04x5 FILLER_64_1905 ();
 b15zdnd00an1n01x5 FILLER_64_1909 ();
 b15zdnd11an1n16x5 FILLER_64_1962 ();
 b15zdnd11an1n08x5 FILLER_64_1978 ();
 b15zdnd11an1n04x5 FILLER_64_1986 ();
 b15zdnd11an1n04x5 FILLER_64_1993 ();
 b15zdnd11an1n64x5 FILLER_64_2000 ();
 b15zdnd00an1n01x5 FILLER_64_2064 ();
 b15zdnd11an1n64x5 FILLER_64_2069 ();
 b15zdnd11an1n16x5 FILLER_64_2133 ();
 b15zdnd11an1n04x5 FILLER_64_2149 ();
 b15zdnd00an1n01x5 FILLER_64_2153 ();
 b15zdnd11an1n64x5 FILLER_64_2162 ();
 b15zdnd11an1n32x5 FILLER_64_2226 ();
 b15zdnd11an1n16x5 FILLER_64_2258 ();
 b15zdnd00an1n02x5 FILLER_64_2274 ();
 b15zdnd11an1n16x5 FILLER_65_0 ();
 b15zdnd11an1n08x5 FILLER_65_16 ();
 b15zdnd11an1n04x5 FILLER_65_24 ();
 b15zdnd11an1n64x5 FILLER_65_33 ();
 b15zdnd11an1n64x5 FILLER_65_97 ();
 b15zdnd11an1n64x5 FILLER_65_161 ();
 b15zdnd11an1n64x5 FILLER_65_225 ();
 b15zdnd11an1n64x5 FILLER_65_289 ();
 b15zdnd11an1n64x5 FILLER_65_353 ();
 b15zdnd11an1n64x5 FILLER_65_417 ();
 b15zdnd11an1n64x5 FILLER_65_481 ();
 b15zdnd11an1n64x5 FILLER_65_545 ();
 b15zdnd11an1n64x5 FILLER_65_609 ();
 b15zdnd11an1n64x5 FILLER_65_673 ();
 b15zdnd11an1n32x5 FILLER_65_737 ();
 b15zdnd11an1n08x5 FILLER_65_769 ();
 b15zdnd11an1n04x5 FILLER_65_777 ();
 b15zdnd00an1n01x5 FILLER_65_781 ();
 b15zdnd11an1n64x5 FILLER_65_785 ();
 b15zdnd11an1n64x5 FILLER_65_849 ();
 b15zdnd11an1n64x5 FILLER_65_913 ();
 b15zdnd11an1n64x5 FILLER_65_977 ();
 b15zdnd11an1n64x5 FILLER_65_1041 ();
 b15zdnd11an1n32x5 FILLER_65_1105 ();
 b15zdnd11an1n16x5 FILLER_65_1137 ();
 b15zdnd11an1n04x5 FILLER_65_1153 ();
 b15zdnd00an1n02x5 FILLER_65_1157 ();
 b15zdnd11an1n64x5 FILLER_65_1173 ();
 b15zdnd11an1n64x5 FILLER_65_1237 ();
 b15zdnd11an1n64x5 FILLER_65_1301 ();
 b15zdnd11an1n64x5 FILLER_65_1365 ();
 b15zdnd11an1n64x5 FILLER_65_1429 ();
 b15zdnd11an1n64x5 FILLER_65_1493 ();
 b15zdnd11an1n64x5 FILLER_65_1557 ();
 b15zdnd11an1n04x5 FILLER_65_1621 ();
 b15zdnd00an1n02x5 FILLER_65_1625 ();
 b15zdnd11an1n64x5 FILLER_65_1633 ();
 b15zdnd11an1n64x5 FILLER_65_1697 ();
 b15zdnd11an1n32x5 FILLER_65_1761 ();
 b15zdnd11an1n16x5 FILLER_65_1793 ();
 b15zdnd00an1n02x5 FILLER_65_1809 ();
 b15zdnd00an1n01x5 FILLER_65_1811 ();
 b15zdnd11an1n64x5 FILLER_65_1864 ();
 b15zdnd11an1n64x5 FILLER_65_1928 ();
 b15zdnd11an1n64x5 FILLER_65_1992 ();
 b15zdnd11an1n64x5 FILLER_65_2056 ();
 b15zdnd11an1n64x5 FILLER_65_2120 ();
 b15zdnd11an1n64x5 FILLER_65_2184 ();
 b15zdnd11an1n32x5 FILLER_65_2248 ();
 b15zdnd11an1n04x5 FILLER_65_2280 ();
 b15zdnd11an1n64x5 FILLER_66_8 ();
 b15zdnd11an1n64x5 FILLER_66_72 ();
 b15zdnd11an1n64x5 FILLER_66_136 ();
 b15zdnd11an1n64x5 FILLER_66_200 ();
 b15zdnd11an1n64x5 FILLER_66_264 ();
 b15zdnd11an1n64x5 FILLER_66_328 ();
 b15zdnd11an1n64x5 FILLER_66_392 ();
 b15zdnd11an1n64x5 FILLER_66_456 ();
 b15zdnd11an1n64x5 FILLER_66_520 ();
 b15zdnd11an1n32x5 FILLER_66_584 ();
 b15zdnd11an1n16x5 FILLER_66_616 ();
 b15zdnd11an1n08x5 FILLER_66_632 ();
 b15zdnd00an1n02x5 FILLER_66_640 ();
 b15zdnd00an1n01x5 FILLER_66_642 ();
 b15zdnd11an1n32x5 FILLER_66_661 ();
 b15zdnd11an1n04x5 FILLER_66_693 ();
 b15zdnd00an1n02x5 FILLER_66_697 ();
 b15zdnd00an1n01x5 FILLER_66_699 ();
 b15zdnd11an1n08x5 FILLER_66_706 ();
 b15zdnd11an1n04x5 FILLER_66_714 ();
 b15zdnd11an1n32x5 FILLER_66_726 ();
 b15zdnd11an1n04x5 FILLER_66_758 ();
 b15zdnd00an1n01x5 FILLER_66_762 ();
 b15zdnd11an1n64x5 FILLER_66_776 ();
 b15zdnd11an1n64x5 FILLER_66_840 ();
 b15zdnd11an1n64x5 FILLER_66_904 ();
 b15zdnd11an1n32x5 FILLER_66_968 ();
 b15zdnd11an1n16x5 FILLER_66_1000 ();
 b15zdnd11an1n08x5 FILLER_66_1016 ();
 b15zdnd11an1n04x5 FILLER_66_1027 ();
 b15zdnd11an1n64x5 FILLER_66_1034 ();
 b15zdnd11an1n64x5 FILLER_66_1098 ();
 b15zdnd11an1n64x5 FILLER_66_1162 ();
 b15zdnd11an1n64x5 FILLER_66_1226 ();
 b15zdnd00an1n02x5 FILLER_66_1290 ();
 b15zdnd00an1n01x5 FILLER_66_1292 ();
 b15zdnd11an1n32x5 FILLER_66_1304 ();
 b15zdnd11an1n08x5 FILLER_66_1336 ();
 b15zdnd00an1n02x5 FILLER_66_1344 ();
 b15zdnd00an1n01x5 FILLER_66_1346 ();
 b15zdnd11an1n64x5 FILLER_66_1361 ();
 b15zdnd11an1n64x5 FILLER_66_1425 ();
 b15zdnd11an1n64x5 FILLER_66_1489 ();
 b15zdnd11an1n32x5 FILLER_66_1553 ();
 b15zdnd11an1n16x5 FILLER_66_1585 ();
 b15zdnd11an1n04x5 FILLER_66_1601 ();
 b15zdnd11an1n64x5 FILLER_66_1609 ();
 b15zdnd11an1n32x5 FILLER_66_1673 ();
 b15zdnd00an1n02x5 FILLER_66_1705 ();
 b15zdnd00an1n01x5 FILLER_66_1707 ();
 b15zdnd11an1n64x5 FILLER_66_1712 ();
 b15zdnd11an1n16x5 FILLER_66_1776 ();
 b15zdnd11an1n08x5 FILLER_66_1792 ();
 b15zdnd00an1n02x5 FILLER_66_1800 ();
 b15zdnd11an1n64x5 FILLER_66_1854 ();
 b15zdnd11an1n64x5 FILLER_66_1918 ();
 b15zdnd11an1n64x5 FILLER_66_1982 ();
 b15zdnd11an1n64x5 FILLER_66_2046 ();
 b15zdnd11an1n32x5 FILLER_66_2110 ();
 b15zdnd11an1n08x5 FILLER_66_2142 ();
 b15zdnd11an1n04x5 FILLER_66_2150 ();
 b15zdnd11an1n64x5 FILLER_66_2162 ();
 b15zdnd11an1n32x5 FILLER_66_2226 ();
 b15zdnd11an1n16x5 FILLER_66_2258 ();
 b15zdnd00an1n02x5 FILLER_66_2274 ();
 b15zdnd11an1n64x5 FILLER_67_0 ();
 b15zdnd11an1n64x5 FILLER_67_64 ();
 b15zdnd11an1n64x5 FILLER_67_128 ();
 b15zdnd11an1n64x5 FILLER_67_192 ();
 b15zdnd11an1n64x5 FILLER_67_256 ();
 b15zdnd11an1n64x5 FILLER_67_320 ();
 b15zdnd11an1n64x5 FILLER_67_384 ();
 b15zdnd11an1n64x5 FILLER_67_448 ();
 b15zdnd11an1n64x5 FILLER_67_512 ();
 b15zdnd11an1n64x5 FILLER_67_576 ();
 b15zdnd11an1n08x5 FILLER_67_640 ();
 b15zdnd00an1n02x5 FILLER_67_648 ();
 b15zdnd11an1n16x5 FILLER_67_655 ();
 b15zdnd11an1n08x5 FILLER_67_671 ();
 b15zdnd11an1n04x5 FILLER_67_679 ();
 b15zdnd00an1n02x5 FILLER_67_683 ();
 b15zdnd11an1n04x5 FILLER_67_727 ();
 b15zdnd11an1n32x5 FILLER_67_745 ();
 b15zdnd00an1n02x5 FILLER_67_777 ();
 b15zdnd11an1n64x5 FILLER_67_793 ();
 b15zdnd11an1n64x5 FILLER_67_857 ();
 b15zdnd11an1n04x5 FILLER_67_921 ();
 b15zdnd00an1n02x5 FILLER_67_925 ();
 b15zdnd11an1n04x5 FILLER_67_930 ();
 b15zdnd11an1n64x5 FILLER_67_937 ();
 b15zdnd00an1n02x5 FILLER_67_1001 ();
 b15zdnd00an1n01x5 FILLER_67_1003 ();
 b15zdnd11an1n64x5 FILLER_67_1056 ();
 b15zdnd11an1n64x5 FILLER_67_1120 ();
 b15zdnd11an1n04x5 FILLER_67_1184 ();
 b15zdnd00an1n02x5 FILLER_67_1188 ();
 b15zdnd00an1n01x5 FILLER_67_1190 ();
 b15zdnd11an1n64x5 FILLER_67_1197 ();
 b15zdnd11an1n32x5 FILLER_67_1261 ();
 b15zdnd11an1n04x5 FILLER_67_1293 ();
 b15zdnd11an1n64x5 FILLER_67_1304 ();
 b15zdnd11an1n64x5 FILLER_67_1368 ();
 b15zdnd11an1n64x5 FILLER_67_1432 ();
 b15zdnd11an1n64x5 FILLER_67_1496 ();
 b15zdnd11an1n16x5 FILLER_67_1560 ();
 b15zdnd11an1n04x5 FILLER_67_1576 ();
 b15zdnd11an1n64x5 FILLER_67_1584 ();
 b15zdnd11an1n32x5 FILLER_67_1648 ();
 b15zdnd11an1n16x5 FILLER_67_1680 ();
 b15zdnd00an1n02x5 FILLER_67_1696 ();
 b15zdnd11an1n64x5 FILLER_67_1702 ();
 b15zdnd11an1n32x5 FILLER_67_1766 ();
 b15zdnd11an1n16x5 FILLER_67_1798 ();
 b15zdnd11an1n08x5 FILLER_67_1814 ();
 b15zdnd00an1n02x5 FILLER_67_1822 ();
 b15zdnd11an1n04x5 FILLER_67_1827 ();
 b15zdnd11an1n04x5 FILLER_67_1834 ();
 b15zdnd11an1n64x5 FILLER_67_1841 ();
 b15zdnd11an1n64x5 FILLER_67_1905 ();
 b15zdnd11an1n64x5 FILLER_67_1969 ();
 b15zdnd11an1n08x5 FILLER_67_2033 ();
 b15zdnd00an1n01x5 FILLER_67_2041 ();
 b15zdnd11an1n32x5 FILLER_67_2048 ();
 b15zdnd11an1n08x5 FILLER_67_2080 ();
 b15zdnd11an1n04x5 FILLER_67_2088 ();
 b15zdnd00an1n02x5 FILLER_67_2092 ();
 b15zdnd11an1n64x5 FILLER_67_2101 ();
 b15zdnd11an1n64x5 FILLER_67_2165 ();
 b15zdnd11an1n32x5 FILLER_67_2229 ();
 b15zdnd11an1n16x5 FILLER_67_2261 ();
 b15zdnd11an1n04x5 FILLER_67_2277 ();
 b15zdnd00an1n02x5 FILLER_67_2281 ();
 b15zdnd00an1n01x5 FILLER_67_2283 ();
 b15zdnd11an1n64x5 FILLER_68_8 ();
 b15zdnd11an1n04x5 FILLER_68_72 ();
 b15zdnd00an1n02x5 FILLER_68_76 ();
 b15zdnd00an1n01x5 FILLER_68_78 ();
 b15zdnd11an1n08x5 FILLER_68_86 ();
 b15zdnd11an1n64x5 FILLER_68_139 ();
 b15zdnd11an1n64x5 FILLER_68_203 ();
 b15zdnd11an1n64x5 FILLER_68_267 ();
 b15zdnd11an1n64x5 FILLER_68_331 ();
 b15zdnd11an1n64x5 FILLER_68_395 ();
 b15zdnd11an1n64x5 FILLER_68_459 ();
 b15zdnd11an1n64x5 FILLER_68_523 ();
 b15zdnd11an1n32x5 FILLER_68_587 ();
 b15zdnd11an1n16x5 FILLER_68_619 ();
 b15zdnd11an1n04x5 FILLER_68_635 ();
 b15zdnd11an1n04x5 FILLER_68_645 ();
 b15zdnd11an1n16x5 FILLER_68_691 ();
 b15zdnd11an1n08x5 FILLER_68_707 ();
 b15zdnd00an1n02x5 FILLER_68_715 ();
 b15zdnd00an1n01x5 FILLER_68_717 ();
 b15zdnd11an1n64x5 FILLER_68_726 ();
 b15zdnd11an1n64x5 FILLER_68_790 ();
 b15zdnd11an1n32x5 FILLER_68_854 ();
 b15zdnd11an1n16x5 FILLER_68_886 ();
 b15zdnd11an1n04x5 FILLER_68_902 ();
 b15zdnd00an1n01x5 FILLER_68_906 ();
 b15zdnd11an1n64x5 FILLER_68_959 ();
 b15zdnd00an1n02x5 FILLER_68_1023 ();
 b15zdnd11an1n16x5 FILLER_68_1028 ();
 b15zdnd11an1n08x5 FILLER_68_1044 ();
 b15zdnd11an1n04x5 FILLER_68_1052 ();
 b15zdnd00an1n02x5 FILLER_68_1056 ();
 b15zdnd00an1n01x5 FILLER_68_1058 ();
 b15zdnd11an1n64x5 FILLER_68_1062 ();
 b15zdnd11an1n16x5 FILLER_68_1126 ();
 b15zdnd11an1n04x5 FILLER_68_1142 ();
 b15zdnd00an1n01x5 FILLER_68_1146 ();
 b15zdnd11an1n64x5 FILLER_68_1164 ();
 b15zdnd11an1n64x5 FILLER_68_1228 ();
 b15zdnd11an1n32x5 FILLER_68_1292 ();
 b15zdnd11an1n04x5 FILLER_68_1324 ();
 b15zdnd11an1n32x5 FILLER_68_1348 ();
 b15zdnd11an1n08x5 FILLER_68_1380 ();
 b15zdnd00an1n02x5 FILLER_68_1388 ();
 b15zdnd00an1n01x5 FILLER_68_1390 ();
 b15zdnd11an1n32x5 FILLER_68_1398 ();
 b15zdnd11an1n08x5 FILLER_68_1430 ();
 b15zdnd11an1n04x5 FILLER_68_1438 ();
 b15zdnd00an1n01x5 FILLER_68_1442 ();
 b15zdnd11an1n04x5 FILLER_68_1450 ();
 b15zdnd11an1n32x5 FILLER_68_1485 ();
 b15zdnd11an1n08x5 FILLER_68_1517 ();
 b15zdnd11an1n04x5 FILLER_68_1525 ();
 b15zdnd00an1n02x5 FILLER_68_1529 ();
 b15zdnd00an1n01x5 FILLER_68_1531 ();
 b15zdnd11an1n64x5 FILLER_68_1538 ();
 b15zdnd11an1n64x5 FILLER_68_1602 ();
 b15zdnd11an1n32x5 FILLER_68_1666 ();
 b15zdnd11an1n04x5 FILLER_68_1698 ();
 b15zdnd11an1n16x5 FILLER_68_1706 ();
 b15zdnd11an1n08x5 FILLER_68_1722 ();
 b15zdnd00an1n02x5 FILLER_68_1730 ();
 b15zdnd11an1n64x5 FILLER_68_1736 ();
 b15zdnd11an1n16x5 FILLER_68_1800 ();
 b15zdnd11an1n04x5 FILLER_68_1816 ();
 b15zdnd11an1n04x5 FILLER_68_1832 ();
 b15zdnd11an1n64x5 FILLER_68_1839 ();
 b15zdnd11an1n64x5 FILLER_68_1903 ();
 b15zdnd11an1n64x5 FILLER_68_1967 ();
 b15zdnd11an1n64x5 FILLER_68_2031 ();
 b15zdnd11an1n32x5 FILLER_68_2095 ();
 b15zdnd11an1n16x5 FILLER_68_2127 ();
 b15zdnd11an1n08x5 FILLER_68_2143 ();
 b15zdnd00an1n02x5 FILLER_68_2151 ();
 b15zdnd00an1n01x5 FILLER_68_2153 ();
 b15zdnd11an1n64x5 FILLER_68_2162 ();
 b15zdnd11an1n32x5 FILLER_68_2226 ();
 b15zdnd11an1n04x5 FILLER_68_2258 ();
 b15zdnd00an1n02x5 FILLER_68_2262 ();
 b15zdnd11an1n04x5 FILLER_68_2272 ();
 b15zdnd11an1n64x5 FILLER_69_0 ();
 b15zdnd11an1n16x5 FILLER_69_64 ();
 b15zdnd11an1n08x5 FILLER_69_80 ();
 b15zdnd11an1n04x5 FILLER_69_88 ();
 b15zdnd11an1n64x5 FILLER_69_99 ();
 b15zdnd11an1n64x5 FILLER_69_163 ();
 b15zdnd11an1n64x5 FILLER_69_227 ();
 b15zdnd11an1n64x5 FILLER_69_291 ();
 b15zdnd11an1n64x5 FILLER_69_355 ();
 b15zdnd11an1n64x5 FILLER_69_419 ();
 b15zdnd11an1n16x5 FILLER_69_483 ();
 b15zdnd11an1n08x5 FILLER_69_499 ();
 b15zdnd00an1n01x5 FILLER_69_507 ();
 b15zdnd11an1n64x5 FILLER_69_522 ();
 b15zdnd11an1n32x5 FILLER_69_586 ();
 b15zdnd11an1n16x5 FILLER_69_618 ();
 b15zdnd11an1n08x5 FILLER_69_634 ();
 b15zdnd11an1n04x5 FILLER_69_642 ();
 b15zdnd00an1n01x5 FILLER_69_646 ();
 b15zdnd11an1n64x5 FILLER_69_668 ();
 b15zdnd11an1n64x5 FILLER_69_732 ();
 b15zdnd00an1n02x5 FILLER_69_796 ();
 b15zdnd00an1n01x5 FILLER_69_798 ();
 b15zdnd11an1n64x5 FILLER_69_802 ();
 b15zdnd11an1n32x5 FILLER_69_866 ();
 b15zdnd11an1n08x5 FILLER_69_898 ();
 b15zdnd00an1n02x5 FILLER_69_906 ();
 b15zdnd11an1n32x5 FILLER_69_960 ();
 b15zdnd11an1n16x5 FILLER_69_992 ();
 b15zdnd11an1n08x5 FILLER_69_1008 ();
 b15zdnd11an1n04x5 FILLER_69_1016 ();
 b15zdnd00an1n02x5 FILLER_69_1020 ();
 b15zdnd11an1n16x5 FILLER_69_1030 ();
 b15zdnd11an1n08x5 FILLER_69_1046 ();
 b15zdnd11an1n04x5 FILLER_69_1054 ();
 b15zdnd00an1n01x5 FILLER_69_1058 ();
 b15zdnd11an1n04x5 FILLER_69_1062 ();
 b15zdnd11an1n32x5 FILLER_69_1069 ();
 b15zdnd11an1n08x5 FILLER_69_1101 ();
 b15zdnd11an1n04x5 FILLER_69_1109 ();
 b15zdnd00an1n02x5 FILLER_69_1113 ();
 b15zdnd00an1n01x5 FILLER_69_1115 ();
 b15zdnd11an1n16x5 FILLER_69_1134 ();
 b15zdnd11an1n04x5 FILLER_69_1150 ();
 b15zdnd00an1n02x5 FILLER_69_1154 ();
 b15zdnd11an1n64x5 FILLER_69_1166 ();
 b15zdnd11an1n64x5 FILLER_69_1230 ();
 b15zdnd11an1n64x5 FILLER_69_1294 ();
 b15zdnd11an1n64x5 FILLER_69_1358 ();
 b15zdnd11an1n08x5 FILLER_69_1422 ();
 b15zdnd00an1n02x5 FILLER_69_1430 ();
 b15zdnd00an1n01x5 FILLER_69_1432 ();
 b15zdnd11an1n64x5 FILLER_69_1447 ();
 b15zdnd11an1n64x5 FILLER_69_1511 ();
 b15zdnd11an1n64x5 FILLER_69_1575 ();
 b15zdnd11an1n64x5 FILLER_69_1639 ();
 b15zdnd11an1n64x5 FILLER_69_1703 ();
 b15zdnd11an1n64x5 FILLER_69_1767 ();
 b15zdnd11an1n64x5 FILLER_69_1831 ();
 b15zdnd11an1n64x5 FILLER_69_1895 ();
 b15zdnd11an1n64x5 FILLER_69_1959 ();
 b15zdnd11an1n08x5 FILLER_69_2023 ();
 b15zdnd11an1n04x5 FILLER_69_2031 ();
 b15zdnd00an1n02x5 FILLER_69_2035 ();
 b15zdnd11an1n64x5 FILLER_69_2043 ();
 b15zdnd11an1n08x5 FILLER_69_2107 ();
 b15zdnd11an1n04x5 FILLER_69_2115 ();
 b15zdnd00an1n01x5 FILLER_69_2119 ();
 b15zdnd11an1n64x5 FILLER_69_2162 ();
 b15zdnd11an1n32x5 FILLER_69_2226 ();
 b15zdnd11an1n16x5 FILLER_69_2258 ();
 b15zdnd11an1n08x5 FILLER_69_2274 ();
 b15zdnd00an1n02x5 FILLER_69_2282 ();
 b15zdnd11an1n64x5 FILLER_70_8 ();
 b15zdnd11an1n64x5 FILLER_70_72 ();
 b15zdnd11an1n64x5 FILLER_70_136 ();
 b15zdnd11an1n64x5 FILLER_70_200 ();
 b15zdnd11an1n64x5 FILLER_70_264 ();
 b15zdnd11an1n64x5 FILLER_70_328 ();
 b15zdnd11an1n64x5 FILLER_70_392 ();
 b15zdnd11an1n32x5 FILLER_70_456 ();
 b15zdnd11an1n08x5 FILLER_70_488 ();
 b15zdnd11an1n04x5 FILLER_70_496 ();
 b15zdnd11an1n32x5 FILLER_70_542 ();
 b15zdnd11an1n16x5 FILLER_70_574 ();
 b15zdnd11an1n04x5 FILLER_70_590 ();
 b15zdnd00an1n02x5 FILLER_70_594 ();
 b15zdnd11an1n04x5 FILLER_70_599 ();
 b15zdnd11an1n08x5 FILLER_70_606 ();
 b15zdnd00an1n01x5 FILLER_70_614 ();
 b15zdnd11an1n32x5 FILLER_70_618 ();
 b15zdnd11an1n04x5 FILLER_70_650 ();
 b15zdnd00an1n01x5 FILLER_70_654 ();
 b15zdnd11an1n16x5 FILLER_70_697 ();
 b15zdnd11an1n04x5 FILLER_70_713 ();
 b15zdnd00an1n01x5 FILLER_70_717 ();
 b15zdnd11an1n32x5 FILLER_70_726 ();
 b15zdnd11an1n16x5 FILLER_70_758 ();
 b15zdnd11an1n04x5 FILLER_70_790 ();
 b15zdnd00an1n01x5 FILLER_70_794 ();
 b15zdnd11an1n04x5 FILLER_70_798 ();
 b15zdnd11an1n64x5 FILLER_70_816 ();
 b15zdnd11an1n16x5 FILLER_70_880 ();
 b15zdnd11an1n08x5 FILLER_70_896 ();
 b15zdnd11an1n04x5 FILLER_70_904 ();
 b15zdnd11an1n04x5 FILLER_70_919 ();
 b15zdnd00an1n02x5 FILLER_70_923 ();
 b15zdnd00an1n01x5 FILLER_70_925 ();
 b15zdnd11an1n04x5 FILLER_70_929 ();
 b15zdnd11an1n04x5 FILLER_70_936 ();
 b15zdnd11an1n64x5 FILLER_70_943 ();
 b15zdnd11an1n16x5 FILLER_70_1007 ();
 b15zdnd11an1n08x5 FILLER_70_1023 ();
 b15zdnd11an1n04x5 FILLER_70_1031 ();
 b15zdnd00an1n01x5 FILLER_70_1035 ();
 b15zdnd11an1n04x5 FILLER_70_1088 ();
 b15zdnd11an1n64x5 FILLER_70_1134 ();
 b15zdnd11an1n64x5 FILLER_70_1198 ();
 b15zdnd11an1n64x5 FILLER_70_1262 ();
 b15zdnd11an1n64x5 FILLER_70_1326 ();
 b15zdnd11an1n64x5 FILLER_70_1390 ();
 b15zdnd11an1n64x5 FILLER_70_1454 ();
 b15zdnd11an1n64x5 FILLER_70_1518 ();
 b15zdnd11an1n64x5 FILLER_70_1582 ();
 b15zdnd11an1n64x5 FILLER_70_1646 ();
 b15zdnd11an1n64x5 FILLER_70_1710 ();
 b15zdnd11an1n64x5 FILLER_70_1774 ();
 b15zdnd11an1n64x5 FILLER_70_1838 ();
 b15zdnd11an1n64x5 FILLER_70_1902 ();
 b15zdnd11an1n64x5 FILLER_70_1966 ();
 b15zdnd11an1n64x5 FILLER_70_2030 ();
 b15zdnd11an1n32x5 FILLER_70_2094 ();
 b15zdnd11an1n16x5 FILLER_70_2126 ();
 b15zdnd11an1n08x5 FILLER_70_2142 ();
 b15zdnd11an1n04x5 FILLER_70_2150 ();
 b15zdnd11an1n64x5 FILLER_70_2162 ();
 b15zdnd11an1n32x5 FILLER_70_2226 ();
 b15zdnd11an1n16x5 FILLER_70_2258 ();
 b15zdnd00an1n02x5 FILLER_70_2274 ();
 b15zdnd11an1n64x5 FILLER_71_0 ();
 b15zdnd11an1n64x5 FILLER_71_64 ();
 b15zdnd11an1n64x5 FILLER_71_128 ();
 b15zdnd11an1n64x5 FILLER_71_192 ();
 b15zdnd11an1n64x5 FILLER_71_256 ();
 b15zdnd11an1n64x5 FILLER_71_320 ();
 b15zdnd11an1n64x5 FILLER_71_384 ();
 b15zdnd11an1n64x5 FILLER_71_448 ();
 b15zdnd11an1n64x5 FILLER_71_512 ();
 b15zdnd11an1n08x5 FILLER_71_628 ();
 b15zdnd11an1n04x5 FILLER_71_636 ();
 b15zdnd11an1n64x5 FILLER_71_643 ();
 b15zdnd11an1n32x5 FILLER_71_749 ();
 b15zdnd11an1n08x5 FILLER_71_781 ();
 b15zdnd11an1n04x5 FILLER_71_789 ();
 b15zdnd00an1n02x5 FILLER_71_793 ();
 b15zdnd00an1n01x5 FILLER_71_795 ();
 b15zdnd11an1n16x5 FILLER_71_800 ();
 b15zdnd11an1n08x5 FILLER_71_816 ();
 b15zdnd11an1n32x5 FILLER_71_866 ();
 b15zdnd11an1n16x5 FILLER_71_898 ();
 b15zdnd11an1n08x5 FILLER_71_914 ();
 b15zdnd11an1n04x5 FILLER_71_922 ();
 b15zdnd00an1n02x5 FILLER_71_926 ();
 b15zdnd11an1n64x5 FILLER_71_931 ();
 b15zdnd11an1n64x5 FILLER_71_995 ();
 b15zdnd11an1n32x5 FILLER_71_1059 ();
 b15zdnd11an1n04x5 FILLER_71_1091 ();
 b15zdnd11an1n32x5 FILLER_71_1099 ();
 b15zdnd11an1n16x5 FILLER_71_1131 ();
 b15zdnd11an1n08x5 FILLER_71_1147 ();
 b15zdnd11an1n04x5 FILLER_71_1155 ();
 b15zdnd11an1n64x5 FILLER_71_1175 ();
 b15zdnd11an1n64x5 FILLER_71_1239 ();
 b15zdnd11an1n64x5 FILLER_71_1303 ();
 b15zdnd11an1n32x5 FILLER_71_1367 ();
 b15zdnd11an1n16x5 FILLER_71_1399 ();
 b15zdnd11an1n08x5 FILLER_71_1415 ();
 b15zdnd11an1n04x5 FILLER_71_1423 ();
 b15zdnd00an1n02x5 FILLER_71_1427 ();
 b15zdnd00an1n01x5 FILLER_71_1429 ();
 b15zdnd11an1n64x5 FILLER_71_1436 ();
 b15zdnd11an1n64x5 FILLER_71_1500 ();
 b15zdnd11an1n16x5 FILLER_71_1564 ();
 b15zdnd11an1n08x5 FILLER_71_1580 ();
 b15zdnd00an1n02x5 FILLER_71_1588 ();
 b15zdnd11an1n64x5 FILLER_71_1594 ();
 b15zdnd11an1n32x5 FILLER_71_1658 ();
 b15zdnd11an1n16x5 FILLER_71_1690 ();
 b15zdnd00an1n02x5 FILLER_71_1706 ();
 b15zdnd11an1n64x5 FILLER_71_1712 ();
 b15zdnd11an1n64x5 FILLER_71_1776 ();
 b15zdnd11an1n64x5 FILLER_71_1840 ();
 b15zdnd11an1n64x5 FILLER_71_1904 ();
 b15zdnd11an1n64x5 FILLER_71_1968 ();
 b15zdnd11an1n08x5 FILLER_71_2032 ();
 b15zdnd00an1n01x5 FILLER_71_2040 ();
 b15zdnd11an1n64x5 FILLER_71_2045 ();
 b15zdnd11an1n64x5 FILLER_71_2109 ();
 b15zdnd11an1n64x5 FILLER_71_2173 ();
 b15zdnd11an1n32x5 FILLER_71_2237 ();
 b15zdnd11an1n08x5 FILLER_71_2269 ();
 b15zdnd11an1n04x5 FILLER_71_2277 ();
 b15zdnd00an1n02x5 FILLER_71_2281 ();
 b15zdnd00an1n01x5 FILLER_71_2283 ();
 b15zdnd11an1n64x5 FILLER_72_8 ();
 b15zdnd11an1n64x5 FILLER_72_72 ();
 b15zdnd11an1n64x5 FILLER_72_136 ();
 b15zdnd11an1n64x5 FILLER_72_200 ();
 b15zdnd11an1n64x5 FILLER_72_264 ();
 b15zdnd11an1n64x5 FILLER_72_328 ();
 b15zdnd11an1n64x5 FILLER_72_392 ();
 b15zdnd11an1n64x5 FILLER_72_456 ();
 b15zdnd11an1n64x5 FILLER_72_520 ();
 b15zdnd11an1n16x5 FILLER_72_584 ();
 b15zdnd00an1n01x5 FILLER_72_600 ();
 b15zdnd11an1n32x5 FILLER_72_604 ();
 b15zdnd11an1n04x5 FILLER_72_636 ();
 b15zdnd00an1n02x5 FILLER_72_640 ();
 b15zdnd00an1n01x5 FILLER_72_642 ();
 b15zdnd11an1n32x5 FILLER_72_685 ();
 b15zdnd00an1n01x5 FILLER_72_717 ();
 b15zdnd11an1n64x5 FILLER_72_726 ();
 b15zdnd11an1n64x5 FILLER_72_794 ();
 b15zdnd11an1n64x5 FILLER_72_858 ();
 b15zdnd11an1n64x5 FILLER_72_922 ();
 b15zdnd11an1n64x5 FILLER_72_986 ();
 b15zdnd11an1n64x5 FILLER_72_1050 ();
 b15zdnd11an1n16x5 FILLER_72_1114 ();
 b15zdnd00an1n01x5 FILLER_72_1130 ();
 b15zdnd11an1n64x5 FILLER_72_1136 ();
 b15zdnd11an1n64x5 FILLER_72_1200 ();
 b15zdnd11an1n64x5 FILLER_72_1264 ();
 b15zdnd11an1n64x5 FILLER_72_1328 ();
 b15zdnd11an1n16x5 FILLER_72_1392 ();
 b15zdnd11an1n08x5 FILLER_72_1408 ();
 b15zdnd11an1n04x5 FILLER_72_1416 ();
 b15zdnd00an1n02x5 FILLER_72_1420 ();
 b15zdnd00an1n01x5 FILLER_72_1422 ();
 b15zdnd11an1n64x5 FILLER_72_1433 ();
 b15zdnd11an1n64x5 FILLER_72_1497 ();
 b15zdnd11an1n64x5 FILLER_72_1561 ();
 b15zdnd11an1n64x5 FILLER_72_1625 ();
 b15zdnd11an1n64x5 FILLER_72_1689 ();
 b15zdnd11an1n64x5 FILLER_72_1753 ();
 b15zdnd11an1n64x5 FILLER_72_1817 ();
 b15zdnd11an1n64x5 FILLER_72_1881 ();
 b15zdnd11an1n64x5 FILLER_72_1945 ();
 b15zdnd11an1n64x5 FILLER_72_2009 ();
 b15zdnd11an1n64x5 FILLER_72_2073 ();
 b15zdnd11an1n16x5 FILLER_72_2137 ();
 b15zdnd00an1n01x5 FILLER_72_2153 ();
 b15zdnd11an1n64x5 FILLER_72_2162 ();
 b15zdnd11an1n32x5 FILLER_72_2226 ();
 b15zdnd11an1n16x5 FILLER_72_2258 ();
 b15zdnd00an1n02x5 FILLER_72_2274 ();
 b15zdnd11an1n64x5 FILLER_73_0 ();
 b15zdnd11an1n64x5 FILLER_73_64 ();
 b15zdnd11an1n64x5 FILLER_73_128 ();
 b15zdnd11an1n64x5 FILLER_73_192 ();
 b15zdnd11an1n64x5 FILLER_73_256 ();
 b15zdnd11an1n64x5 FILLER_73_320 ();
 b15zdnd11an1n64x5 FILLER_73_384 ();
 b15zdnd11an1n64x5 FILLER_73_448 ();
 b15zdnd11an1n64x5 FILLER_73_512 ();
 b15zdnd11an1n64x5 FILLER_73_576 ();
 b15zdnd11an1n08x5 FILLER_73_640 ();
 b15zdnd11an1n32x5 FILLER_73_662 ();
 b15zdnd11an1n04x5 FILLER_73_694 ();
 b15zdnd00an1n02x5 FILLER_73_698 ();
 b15zdnd00an1n01x5 FILLER_73_700 ();
 b15zdnd11an1n64x5 FILLER_73_715 ();
 b15zdnd11an1n04x5 FILLER_73_779 ();
 b15zdnd11an1n04x5 FILLER_73_797 ();
 b15zdnd11an1n64x5 FILLER_73_805 ();
 b15zdnd11an1n64x5 FILLER_73_869 ();
 b15zdnd11an1n16x5 FILLER_73_933 ();
 b15zdnd11an1n08x5 FILLER_73_949 ();
 b15zdnd00an1n02x5 FILLER_73_957 ();
 b15zdnd00an1n01x5 FILLER_73_959 ();
 b15zdnd11an1n32x5 FILLER_73_969 ();
 b15zdnd11an1n08x5 FILLER_73_1001 ();
 b15zdnd11an1n04x5 FILLER_73_1009 ();
 b15zdnd00an1n02x5 FILLER_73_1013 ();
 b15zdnd00an1n01x5 FILLER_73_1015 ();
 b15zdnd11an1n64x5 FILLER_73_1025 ();
 b15zdnd11an1n64x5 FILLER_73_1089 ();
 b15zdnd11an1n64x5 FILLER_73_1153 ();
 b15zdnd11an1n64x5 FILLER_73_1217 ();
 b15zdnd11an1n64x5 FILLER_73_1281 ();
 b15zdnd11an1n64x5 FILLER_73_1345 ();
 b15zdnd11an1n08x5 FILLER_73_1409 ();
 b15zdnd11an1n04x5 FILLER_73_1417 ();
 b15zdnd11an1n64x5 FILLER_73_1437 ();
 b15zdnd11an1n64x5 FILLER_73_1501 ();
 b15zdnd11an1n32x5 FILLER_73_1565 ();
 b15zdnd00an1n02x5 FILLER_73_1597 ();
 b15zdnd11an1n64x5 FILLER_73_1630 ();
 b15zdnd11an1n64x5 FILLER_73_1694 ();
 b15zdnd11an1n64x5 FILLER_73_1758 ();
 b15zdnd11an1n04x5 FILLER_73_1822 ();
 b15zdnd11an1n64x5 FILLER_73_1854 ();
 b15zdnd11an1n64x5 FILLER_73_1918 ();
 b15zdnd11an1n64x5 FILLER_73_1982 ();
 b15zdnd11an1n64x5 FILLER_73_2046 ();
 b15zdnd11an1n64x5 FILLER_73_2110 ();
 b15zdnd11an1n64x5 FILLER_73_2174 ();
 b15zdnd11an1n32x5 FILLER_73_2238 ();
 b15zdnd11an1n08x5 FILLER_73_2270 ();
 b15zdnd11an1n04x5 FILLER_73_2278 ();
 b15zdnd00an1n02x5 FILLER_73_2282 ();
 b15zdnd11an1n64x5 FILLER_74_8 ();
 b15zdnd11an1n64x5 FILLER_74_72 ();
 b15zdnd11an1n64x5 FILLER_74_136 ();
 b15zdnd11an1n64x5 FILLER_74_200 ();
 b15zdnd11an1n64x5 FILLER_74_264 ();
 b15zdnd11an1n64x5 FILLER_74_328 ();
 b15zdnd11an1n64x5 FILLER_74_392 ();
 b15zdnd11an1n64x5 FILLER_74_456 ();
 b15zdnd11an1n64x5 FILLER_74_520 ();
 b15zdnd11an1n64x5 FILLER_74_584 ();
 b15zdnd11an1n64x5 FILLER_74_648 ();
 b15zdnd11an1n04x5 FILLER_74_712 ();
 b15zdnd00an1n02x5 FILLER_74_716 ();
 b15zdnd11an1n64x5 FILLER_74_726 ();
 b15zdnd11an1n08x5 FILLER_74_790 ();
 b15zdnd11an1n16x5 FILLER_74_814 ();
 b15zdnd11an1n08x5 FILLER_74_830 ();
 b15zdnd11an1n64x5 FILLER_74_849 ();
 b15zdnd11an1n64x5 FILLER_74_913 ();
 b15zdnd11an1n64x5 FILLER_74_977 ();
 b15zdnd11an1n32x5 FILLER_74_1041 ();
 b15zdnd11an1n16x5 FILLER_74_1073 ();
 b15zdnd11an1n04x5 FILLER_74_1089 ();
 b15zdnd00an1n02x5 FILLER_74_1093 ();
 b15zdnd11an1n64x5 FILLER_74_1099 ();
 b15zdnd11an1n64x5 FILLER_74_1163 ();
 b15zdnd11an1n64x5 FILLER_74_1227 ();
 b15zdnd11an1n64x5 FILLER_74_1291 ();
 b15zdnd11an1n64x5 FILLER_74_1355 ();
 b15zdnd11an1n64x5 FILLER_74_1419 ();
 b15zdnd11an1n64x5 FILLER_74_1483 ();
 b15zdnd11an1n64x5 FILLER_74_1547 ();
 b15zdnd11an1n64x5 FILLER_74_1611 ();
 b15zdnd11an1n64x5 FILLER_74_1675 ();
 b15zdnd11an1n64x5 FILLER_74_1739 ();
 b15zdnd11an1n64x5 FILLER_74_1803 ();
 b15zdnd11an1n16x5 FILLER_74_1867 ();
 b15zdnd00an1n02x5 FILLER_74_1883 ();
 b15zdnd00an1n01x5 FILLER_74_1885 ();
 b15zdnd11an1n32x5 FILLER_74_1900 ();
 b15zdnd00an1n01x5 FILLER_74_1932 ();
 b15zdnd11an1n16x5 FILLER_74_1937 ();
 b15zdnd11an1n08x5 FILLER_74_1953 ();
 b15zdnd11an1n04x5 FILLER_74_1961 ();
 b15zdnd00an1n02x5 FILLER_74_1965 ();
 b15zdnd11an1n64x5 FILLER_74_1998 ();
 b15zdnd11an1n64x5 FILLER_74_2062 ();
 b15zdnd11an1n16x5 FILLER_74_2126 ();
 b15zdnd11an1n08x5 FILLER_74_2142 ();
 b15zdnd11an1n04x5 FILLER_74_2150 ();
 b15zdnd11an1n64x5 FILLER_74_2162 ();
 b15zdnd11an1n32x5 FILLER_74_2226 ();
 b15zdnd11an1n16x5 FILLER_74_2258 ();
 b15zdnd00an1n02x5 FILLER_74_2274 ();
 b15zdnd11an1n64x5 FILLER_75_0 ();
 b15zdnd11an1n64x5 FILLER_75_64 ();
 b15zdnd11an1n32x5 FILLER_75_128 ();
 b15zdnd11an1n08x5 FILLER_75_160 ();
 b15zdnd00an1n02x5 FILLER_75_168 ();
 b15zdnd11an1n64x5 FILLER_75_222 ();
 b15zdnd11an1n64x5 FILLER_75_286 ();
 b15zdnd11an1n64x5 FILLER_75_350 ();
 b15zdnd11an1n16x5 FILLER_75_414 ();
 b15zdnd00an1n02x5 FILLER_75_430 ();
 b15zdnd00an1n01x5 FILLER_75_432 ();
 b15zdnd11an1n04x5 FILLER_75_438 ();
 b15zdnd11an1n32x5 FILLER_75_446 ();
 b15zdnd11an1n16x5 FILLER_75_478 ();
 b15zdnd00an1n01x5 FILLER_75_494 ();
 b15zdnd11an1n64x5 FILLER_75_498 ();
 b15zdnd11an1n64x5 FILLER_75_562 ();
 b15zdnd11an1n32x5 FILLER_75_626 ();
 b15zdnd11an1n16x5 FILLER_75_658 ();
 b15zdnd11an1n04x5 FILLER_75_684 ();
 b15zdnd11an1n64x5 FILLER_75_702 ();
 b15zdnd11an1n64x5 FILLER_75_766 ();
 b15zdnd11an1n08x5 FILLER_75_830 ();
 b15zdnd11an1n04x5 FILLER_75_838 ();
 b15zdnd00an1n02x5 FILLER_75_842 ();
 b15zdnd00an1n01x5 FILLER_75_844 ();
 b15zdnd11an1n64x5 FILLER_75_865 ();
 b15zdnd11an1n64x5 FILLER_75_929 ();
 b15zdnd11an1n64x5 FILLER_75_993 ();
 b15zdnd11an1n64x5 FILLER_75_1057 ();
 b15zdnd11an1n64x5 FILLER_75_1121 ();
 b15zdnd11an1n64x5 FILLER_75_1185 ();
 b15zdnd11an1n64x5 FILLER_75_1249 ();
 b15zdnd11an1n64x5 FILLER_75_1313 ();
 b15zdnd11an1n64x5 FILLER_75_1377 ();
 b15zdnd11an1n04x5 FILLER_75_1441 ();
 b15zdnd11an1n32x5 FILLER_75_1476 ();
 b15zdnd11an1n16x5 FILLER_75_1508 ();
 b15zdnd11an1n08x5 FILLER_75_1524 ();
 b15zdnd11an1n04x5 FILLER_75_1532 ();
 b15zdnd00an1n02x5 FILLER_75_1536 ();
 b15zdnd11an1n08x5 FILLER_75_1546 ();
 b15zdnd00an1n01x5 FILLER_75_1554 ();
 b15zdnd11an1n64x5 FILLER_75_1599 ();
 b15zdnd11an1n16x5 FILLER_75_1663 ();
 b15zdnd11an1n04x5 FILLER_75_1679 ();
 b15zdnd00an1n02x5 FILLER_75_1683 ();
 b15zdnd00an1n01x5 FILLER_75_1685 ();
 b15zdnd11an1n04x5 FILLER_75_1689 ();
 b15zdnd11an1n64x5 FILLER_75_1696 ();
 b15zdnd11an1n64x5 FILLER_75_1760 ();
 b15zdnd11an1n64x5 FILLER_75_1824 ();
 b15zdnd11an1n64x5 FILLER_75_1888 ();
 b15zdnd11an1n64x5 FILLER_75_1952 ();
 b15zdnd11an1n64x5 FILLER_75_2016 ();
 b15zdnd11an1n64x5 FILLER_75_2080 ();
 b15zdnd11an1n64x5 FILLER_75_2144 ();
 b15zdnd11an1n64x5 FILLER_75_2208 ();
 b15zdnd11an1n08x5 FILLER_75_2272 ();
 b15zdnd11an1n04x5 FILLER_75_2280 ();
 b15zdnd11an1n64x5 FILLER_76_8 ();
 b15zdnd11an1n64x5 FILLER_76_72 ();
 b15zdnd11an1n32x5 FILLER_76_136 ();
 b15zdnd11an1n16x5 FILLER_76_168 ();
 b15zdnd00an1n02x5 FILLER_76_184 ();
 b15zdnd11an1n64x5 FILLER_76_228 ();
 b15zdnd11an1n64x5 FILLER_76_292 ();
 b15zdnd11an1n08x5 FILLER_76_356 ();
 b15zdnd11an1n32x5 FILLER_76_375 ();
 b15zdnd11an1n16x5 FILLER_76_407 ();
 b15zdnd11an1n08x5 FILLER_76_423 ();
 b15zdnd11an1n16x5 FILLER_76_440 ();
 b15zdnd11an1n08x5 FILLER_76_456 ();
 b15zdnd11an1n04x5 FILLER_76_464 ();
 b15zdnd11an1n64x5 FILLER_76_520 ();
 b15zdnd11an1n64x5 FILLER_76_584 ();
 b15zdnd11an1n32x5 FILLER_76_648 ();
 b15zdnd00an1n01x5 FILLER_76_680 ();
 b15zdnd11an1n04x5 FILLER_76_695 ();
 b15zdnd00an1n02x5 FILLER_76_716 ();
 b15zdnd11an1n64x5 FILLER_76_726 ();
 b15zdnd11an1n32x5 FILLER_76_790 ();
 b15zdnd11an1n08x5 FILLER_76_822 ();
 b15zdnd00an1n01x5 FILLER_76_830 ();
 b15zdnd11an1n04x5 FILLER_76_857 ();
 b15zdnd11an1n64x5 FILLER_76_869 ();
 b15zdnd11an1n64x5 FILLER_76_933 ();
 b15zdnd11an1n08x5 FILLER_76_997 ();
 b15zdnd00an1n02x5 FILLER_76_1005 ();
 b15zdnd00an1n01x5 FILLER_76_1007 ();
 b15zdnd11an1n04x5 FILLER_76_1011 ();
 b15zdnd11an1n64x5 FILLER_76_1042 ();
 b15zdnd11an1n32x5 FILLER_76_1106 ();
 b15zdnd11an1n04x5 FILLER_76_1138 ();
 b15zdnd00an1n02x5 FILLER_76_1142 ();
 b15zdnd11an1n04x5 FILLER_76_1158 ();
 b15zdnd11an1n64x5 FILLER_76_1173 ();
 b15zdnd11an1n64x5 FILLER_76_1237 ();
 b15zdnd11an1n64x5 FILLER_76_1301 ();
 b15zdnd11an1n64x5 FILLER_76_1365 ();
 b15zdnd11an1n64x5 FILLER_76_1429 ();
 b15zdnd11an1n64x5 FILLER_76_1493 ();
 b15zdnd11an1n08x5 FILLER_76_1557 ();
 b15zdnd11an1n04x5 FILLER_76_1565 ();
 b15zdnd00an1n01x5 FILLER_76_1569 ();
 b15zdnd11an1n04x5 FILLER_76_1573 ();
 b15zdnd11an1n64x5 FILLER_76_1580 ();
 b15zdnd11an1n16x5 FILLER_76_1644 ();
 b15zdnd11an1n04x5 FILLER_76_1660 ();
 b15zdnd11an1n64x5 FILLER_76_1708 ();
 b15zdnd11an1n64x5 FILLER_76_1772 ();
 b15zdnd11an1n64x5 FILLER_76_1836 ();
 b15zdnd11an1n64x5 FILLER_76_1900 ();
 b15zdnd11an1n64x5 FILLER_76_1964 ();
 b15zdnd11an1n64x5 FILLER_76_2028 ();
 b15zdnd11an1n32x5 FILLER_76_2092 ();
 b15zdnd11an1n16x5 FILLER_76_2124 ();
 b15zdnd11an1n08x5 FILLER_76_2140 ();
 b15zdnd11an1n04x5 FILLER_76_2148 ();
 b15zdnd00an1n02x5 FILLER_76_2152 ();
 b15zdnd11an1n64x5 FILLER_76_2162 ();
 b15zdnd11an1n32x5 FILLER_76_2226 ();
 b15zdnd11an1n16x5 FILLER_76_2258 ();
 b15zdnd00an1n02x5 FILLER_76_2274 ();
 b15zdnd11an1n64x5 FILLER_77_0 ();
 b15zdnd11an1n64x5 FILLER_77_64 ();
 b15zdnd11an1n32x5 FILLER_77_128 ();
 b15zdnd11an1n16x5 FILLER_77_160 ();
 b15zdnd11an1n08x5 FILLER_77_176 ();
 b15zdnd11an1n04x5 FILLER_77_184 ();
 b15zdnd00an1n02x5 FILLER_77_188 ();
 b15zdnd11an1n04x5 FILLER_77_193 ();
 b15zdnd11an1n04x5 FILLER_77_200 ();
 b15zdnd11an1n64x5 FILLER_77_207 ();
 b15zdnd11an1n64x5 FILLER_77_271 ();
 b15zdnd11an1n64x5 FILLER_77_335 ();
 b15zdnd11an1n32x5 FILLER_77_399 ();
 b15zdnd00an1n02x5 FILLER_77_431 ();
 b15zdnd11an1n08x5 FILLER_77_442 ();
 b15zdnd11an1n04x5 FILLER_77_450 ();
 b15zdnd00an1n01x5 FILLER_77_454 ();
 b15zdnd11an1n04x5 FILLER_77_497 ();
 b15zdnd11an1n64x5 FILLER_77_504 ();
 b15zdnd11an1n32x5 FILLER_77_568 ();
 b15zdnd11an1n08x5 FILLER_77_600 ();
 b15zdnd11an1n04x5 FILLER_77_608 ();
 b15zdnd00an1n02x5 FILLER_77_612 ();
 b15zdnd00an1n01x5 FILLER_77_614 ();
 b15zdnd11an1n16x5 FILLER_77_626 ();
 b15zdnd11an1n08x5 FILLER_77_642 ();
 b15zdnd00an1n02x5 FILLER_77_650 ();
 b15zdnd00an1n01x5 FILLER_77_652 ();
 b15zdnd11an1n32x5 FILLER_77_661 ();
 b15zdnd11an1n16x5 FILLER_77_693 ();
 b15zdnd11an1n04x5 FILLER_77_709 ();
 b15zdnd00an1n02x5 FILLER_77_713 ();
 b15zdnd00an1n01x5 FILLER_77_715 ();
 b15zdnd11an1n64x5 FILLER_77_723 ();
 b15zdnd11an1n04x5 FILLER_77_787 ();
 b15zdnd00an1n02x5 FILLER_77_791 ();
 b15zdnd00an1n01x5 FILLER_77_793 ();
 b15zdnd11an1n64x5 FILLER_77_806 ();
 b15zdnd11an1n64x5 FILLER_77_870 ();
 b15zdnd11an1n32x5 FILLER_77_934 ();
 b15zdnd11an1n16x5 FILLER_77_966 ();
 b15zdnd11an1n08x5 FILLER_77_982 ();
 b15zdnd00an1n02x5 FILLER_77_990 ();
 b15zdnd00an1n01x5 FILLER_77_992 ();
 b15zdnd11an1n64x5 FILLER_77_1002 ();
 b15zdnd11an1n64x5 FILLER_77_1066 ();
 b15zdnd11an1n64x5 FILLER_77_1130 ();
 b15zdnd11an1n64x5 FILLER_77_1194 ();
 b15zdnd11an1n64x5 FILLER_77_1258 ();
 b15zdnd11an1n64x5 FILLER_77_1322 ();
 b15zdnd11an1n64x5 FILLER_77_1386 ();
 b15zdnd11an1n64x5 FILLER_77_1450 ();
 b15zdnd11an1n32x5 FILLER_77_1514 ();
 b15zdnd11an1n16x5 FILLER_77_1546 ();
 b15zdnd11an1n04x5 FILLER_77_1562 ();
 b15zdnd00an1n02x5 FILLER_77_1566 ();
 b15zdnd11an1n04x5 FILLER_77_1574 ();
 b15zdnd11an1n64x5 FILLER_77_1581 ();
 b15zdnd11an1n32x5 FILLER_77_1645 ();
 b15zdnd11an1n08x5 FILLER_77_1677 ();
 b15zdnd00an1n02x5 FILLER_77_1685 ();
 b15zdnd11an1n64x5 FILLER_77_1690 ();
 b15zdnd11an1n08x5 FILLER_77_1754 ();
 b15zdnd00an1n02x5 FILLER_77_1762 ();
 b15zdnd11an1n64x5 FILLER_77_1772 ();
 b15zdnd11an1n64x5 FILLER_77_1836 ();
 b15zdnd11an1n64x5 FILLER_77_1900 ();
 b15zdnd11an1n64x5 FILLER_77_1964 ();
 b15zdnd11an1n64x5 FILLER_77_2028 ();
 b15zdnd11an1n64x5 FILLER_77_2092 ();
 b15zdnd11an1n64x5 FILLER_77_2156 ();
 b15zdnd11an1n64x5 FILLER_77_2220 ();
 b15zdnd11an1n64x5 FILLER_78_8 ();
 b15zdnd11an1n64x5 FILLER_78_72 ();
 b15zdnd11an1n64x5 FILLER_78_136 ();
 b15zdnd11an1n64x5 FILLER_78_200 ();
 b15zdnd11an1n64x5 FILLER_78_264 ();
 b15zdnd11an1n64x5 FILLER_78_328 ();
 b15zdnd11an1n08x5 FILLER_78_392 ();
 b15zdnd11an1n08x5 FILLER_78_405 ();
 b15zdnd11an1n04x5 FILLER_78_413 ();
 b15zdnd00an1n02x5 FILLER_78_417 ();
 b15zdnd00an1n01x5 FILLER_78_419 ();
 b15zdnd11an1n04x5 FILLER_78_431 ();
 b15zdnd00an1n02x5 FILLER_78_435 ();
 b15zdnd00an1n01x5 FILLER_78_437 ();
 b15zdnd11an1n32x5 FILLER_78_443 ();
 b15zdnd11an1n08x5 FILLER_78_475 ();
 b15zdnd00an1n02x5 FILLER_78_483 ();
 b15zdnd00an1n01x5 FILLER_78_485 ();
 b15zdnd11an1n64x5 FILLER_78_489 ();
 b15zdnd11an1n64x5 FILLER_78_553 ();
 b15zdnd11an1n32x5 FILLER_78_617 ();
 b15zdnd11an1n08x5 FILLER_78_649 ();
 b15zdnd11an1n04x5 FILLER_78_657 ();
 b15zdnd00an1n02x5 FILLER_78_661 ();
 b15zdnd11an1n16x5 FILLER_78_669 ();
 b15zdnd11an1n04x5 FILLER_78_685 ();
 b15zdnd00an1n01x5 FILLER_78_689 ();
 b15zdnd11an1n16x5 FILLER_78_697 ();
 b15zdnd11an1n04x5 FILLER_78_713 ();
 b15zdnd00an1n01x5 FILLER_78_717 ();
 b15zdnd11an1n64x5 FILLER_78_726 ();
 b15zdnd11an1n64x5 FILLER_78_790 ();
 b15zdnd11an1n64x5 FILLER_78_854 ();
 b15zdnd11an1n64x5 FILLER_78_918 ();
 b15zdnd11an1n64x5 FILLER_78_982 ();
 b15zdnd11an1n64x5 FILLER_78_1046 ();
 b15zdnd11an1n64x5 FILLER_78_1110 ();
 b15zdnd11an1n64x5 FILLER_78_1174 ();
 b15zdnd11an1n64x5 FILLER_78_1238 ();
 b15zdnd11an1n64x5 FILLER_78_1302 ();
 b15zdnd11an1n64x5 FILLER_78_1366 ();
 b15zdnd11an1n64x5 FILLER_78_1430 ();
 b15zdnd11an1n64x5 FILLER_78_1494 ();
 b15zdnd11an1n32x5 FILLER_78_1558 ();
 b15zdnd11an1n16x5 FILLER_78_1590 ();
 b15zdnd00an1n02x5 FILLER_78_1606 ();
 b15zdnd00an1n01x5 FILLER_78_1608 ();
 b15zdnd11an1n64x5 FILLER_78_1612 ();
 b15zdnd11an1n64x5 FILLER_78_1676 ();
 b15zdnd11an1n64x5 FILLER_78_1740 ();
 b15zdnd11an1n32x5 FILLER_78_1810 ();
 b15zdnd11an1n16x5 FILLER_78_1842 ();
 b15zdnd11an1n08x5 FILLER_78_1858 ();
 b15zdnd00an1n02x5 FILLER_78_1866 ();
 b15zdnd00an1n01x5 FILLER_78_1868 ();
 b15zdnd11an1n64x5 FILLER_78_1889 ();
 b15zdnd11an1n64x5 FILLER_78_1953 ();
 b15zdnd11an1n64x5 FILLER_78_2017 ();
 b15zdnd11an1n64x5 FILLER_78_2081 ();
 b15zdnd11an1n08x5 FILLER_78_2145 ();
 b15zdnd00an1n01x5 FILLER_78_2153 ();
 b15zdnd11an1n64x5 FILLER_78_2162 ();
 b15zdnd11an1n32x5 FILLER_78_2226 ();
 b15zdnd11an1n16x5 FILLER_78_2258 ();
 b15zdnd00an1n02x5 FILLER_78_2274 ();
 b15zdnd11an1n64x5 FILLER_79_0 ();
 b15zdnd11an1n64x5 FILLER_79_64 ();
 b15zdnd11an1n64x5 FILLER_79_128 ();
 b15zdnd11an1n64x5 FILLER_79_192 ();
 b15zdnd11an1n64x5 FILLER_79_256 ();
 b15zdnd11an1n64x5 FILLER_79_320 ();
 b15zdnd11an1n64x5 FILLER_79_384 ();
 b15zdnd11an1n64x5 FILLER_79_448 ();
 b15zdnd11an1n64x5 FILLER_79_512 ();
 b15zdnd11an1n64x5 FILLER_79_576 ();
 b15zdnd11an1n64x5 FILLER_79_640 ();
 b15zdnd11an1n64x5 FILLER_79_704 ();
 b15zdnd11an1n64x5 FILLER_79_768 ();
 b15zdnd11an1n64x5 FILLER_79_832 ();
 b15zdnd11an1n64x5 FILLER_79_896 ();
 b15zdnd11an1n64x5 FILLER_79_960 ();
 b15zdnd11an1n64x5 FILLER_79_1024 ();
 b15zdnd11an1n64x5 FILLER_79_1088 ();
 b15zdnd11an1n08x5 FILLER_79_1152 ();
 b15zdnd11an1n04x5 FILLER_79_1160 ();
 b15zdnd11an1n16x5 FILLER_79_1167 ();
 b15zdnd11an1n08x5 FILLER_79_1183 ();
 b15zdnd00an1n02x5 FILLER_79_1191 ();
 b15zdnd11an1n64x5 FILLER_79_1207 ();
 b15zdnd11an1n64x5 FILLER_79_1271 ();
 b15zdnd11an1n64x5 FILLER_79_1335 ();
 b15zdnd11an1n32x5 FILLER_79_1399 ();
 b15zdnd11an1n16x5 FILLER_79_1431 ();
 b15zdnd11an1n08x5 FILLER_79_1447 ();
 b15zdnd11an1n04x5 FILLER_79_1455 ();
 b15zdnd00an1n01x5 FILLER_79_1459 ();
 b15zdnd11an1n64x5 FILLER_79_1473 ();
 b15zdnd11an1n32x5 FILLER_79_1537 ();
 b15zdnd00an1n01x5 FILLER_79_1569 ();
 b15zdnd11an1n16x5 FILLER_79_1576 ();
 b15zdnd11an1n04x5 FILLER_79_1592 ();
 b15zdnd00an1n02x5 FILLER_79_1596 ();
 b15zdnd00an1n01x5 FILLER_79_1598 ();
 b15zdnd11an1n64x5 FILLER_79_1612 ();
 b15zdnd11an1n32x5 FILLER_79_1676 ();
 b15zdnd00an1n02x5 FILLER_79_1708 ();
 b15zdnd00an1n01x5 FILLER_79_1710 ();
 b15zdnd11an1n16x5 FILLER_79_1735 ();
 b15zdnd00an1n02x5 FILLER_79_1751 ();
 b15zdnd11an1n64x5 FILLER_79_1757 ();
 b15zdnd11an1n64x5 FILLER_79_1821 ();
 b15zdnd11an1n16x5 FILLER_79_1885 ();
 b15zdnd11an1n04x5 FILLER_79_1901 ();
 b15zdnd00an1n02x5 FILLER_79_1905 ();
 b15zdnd11an1n64x5 FILLER_79_1915 ();
 b15zdnd11an1n64x5 FILLER_79_1979 ();
 b15zdnd11an1n64x5 FILLER_79_2043 ();
 b15zdnd11an1n64x5 FILLER_79_2107 ();
 b15zdnd11an1n64x5 FILLER_79_2171 ();
 b15zdnd11an1n32x5 FILLER_79_2235 ();
 b15zdnd11an1n16x5 FILLER_79_2267 ();
 b15zdnd00an1n01x5 FILLER_79_2283 ();
 b15zdnd11an1n64x5 FILLER_80_8 ();
 b15zdnd11an1n64x5 FILLER_80_72 ();
 b15zdnd11an1n64x5 FILLER_80_136 ();
 b15zdnd11an1n64x5 FILLER_80_200 ();
 b15zdnd11an1n64x5 FILLER_80_264 ();
 b15zdnd11an1n32x5 FILLER_80_328 ();
 b15zdnd11an1n08x5 FILLER_80_360 ();
 b15zdnd11an1n04x5 FILLER_80_368 ();
 b15zdnd00an1n02x5 FILLER_80_372 ();
 b15zdnd00an1n01x5 FILLER_80_374 ();
 b15zdnd11an1n64x5 FILLER_80_378 ();
 b15zdnd11an1n64x5 FILLER_80_442 ();
 b15zdnd11an1n64x5 FILLER_80_506 ();
 b15zdnd11an1n64x5 FILLER_80_570 ();
 b15zdnd11an1n32x5 FILLER_80_634 ();
 b15zdnd11an1n08x5 FILLER_80_666 ();
 b15zdnd11an1n04x5 FILLER_80_674 ();
 b15zdnd00an1n02x5 FILLER_80_678 ();
 b15zdnd00an1n01x5 FILLER_80_680 ();
 b15zdnd11an1n04x5 FILLER_80_702 ();
 b15zdnd00an1n01x5 FILLER_80_706 ();
 b15zdnd11an1n04x5 FILLER_80_714 ();
 b15zdnd11an1n16x5 FILLER_80_726 ();
 b15zdnd11an1n08x5 FILLER_80_742 ();
 b15zdnd11an1n04x5 FILLER_80_750 ();
 b15zdnd00an1n02x5 FILLER_80_754 ();
 b15zdnd00an1n01x5 FILLER_80_756 ();
 b15zdnd11an1n64x5 FILLER_80_799 ();
 b15zdnd11an1n64x5 FILLER_80_863 ();
 b15zdnd11an1n64x5 FILLER_80_927 ();
 b15zdnd11an1n64x5 FILLER_80_991 ();
 b15zdnd11an1n64x5 FILLER_80_1055 ();
 b15zdnd11an1n64x5 FILLER_80_1119 ();
 b15zdnd11an1n64x5 FILLER_80_1183 ();
 b15zdnd11an1n32x5 FILLER_80_1247 ();
 b15zdnd11an1n08x5 FILLER_80_1279 ();
 b15zdnd11an1n64x5 FILLER_80_1290 ();
 b15zdnd11an1n16x5 FILLER_80_1354 ();
 b15zdnd11an1n08x5 FILLER_80_1370 ();
 b15zdnd00an1n02x5 FILLER_80_1378 ();
 b15zdnd11an1n32x5 FILLER_80_1416 ();
 b15zdnd11an1n16x5 FILLER_80_1448 ();
 b15zdnd11an1n08x5 FILLER_80_1464 ();
 b15zdnd11an1n64x5 FILLER_80_1475 ();
 b15zdnd11an1n64x5 FILLER_80_1539 ();
 b15zdnd11an1n64x5 FILLER_80_1603 ();
 b15zdnd11an1n32x5 FILLER_80_1667 ();
 b15zdnd11an1n16x5 FILLER_80_1699 ();
 b15zdnd00an1n01x5 FILLER_80_1715 ();
 b15zdnd11an1n08x5 FILLER_80_1724 ();
 b15zdnd11an1n04x5 FILLER_80_1732 ();
 b15zdnd11an1n04x5 FILLER_80_1742 ();
 b15zdnd11an1n64x5 FILLER_80_1751 ();
 b15zdnd11an1n64x5 FILLER_80_1815 ();
 b15zdnd11an1n64x5 FILLER_80_1879 ();
 b15zdnd11an1n64x5 FILLER_80_1943 ();
 b15zdnd11an1n64x5 FILLER_80_2007 ();
 b15zdnd11an1n64x5 FILLER_80_2071 ();
 b15zdnd11an1n16x5 FILLER_80_2135 ();
 b15zdnd00an1n02x5 FILLER_80_2151 ();
 b15zdnd00an1n01x5 FILLER_80_2153 ();
 b15zdnd11an1n64x5 FILLER_80_2162 ();
 b15zdnd11an1n32x5 FILLER_80_2226 ();
 b15zdnd11an1n16x5 FILLER_80_2258 ();
 b15zdnd00an1n02x5 FILLER_80_2274 ();
 b15zdnd11an1n64x5 FILLER_81_0 ();
 b15zdnd11an1n64x5 FILLER_81_64 ();
 b15zdnd11an1n64x5 FILLER_81_128 ();
 b15zdnd11an1n64x5 FILLER_81_192 ();
 b15zdnd11an1n64x5 FILLER_81_256 ();
 b15zdnd11an1n32x5 FILLER_81_320 ();
 b15zdnd11an1n16x5 FILLER_81_352 ();
 b15zdnd11an1n04x5 FILLER_81_368 ();
 b15zdnd00an1n01x5 FILLER_81_372 ();
 b15zdnd11an1n64x5 FILLER_81_380 ();
 b15zdnd11an1n64x5 FILLER_81_444 ();
 b15zdnd11an1n64x5 FILLER_81_508 ();
 b15zdnd11an1n64x5 FILLER_81_572 ();
 b15zdnd11an1n64x5 FILLER_81_636 ();
 b15zdnd11an1n64x5 FILLER_81_700 ();
 b15zdnd11an1n64x5 FILLER_81_764 ();
 b15zdnd11an1n64x5 FILLER_81_828 ();
 b15zdnd11an1n64x5 FILLER_81_892 ();
 b15zdnd11an1n64x5 FILLER_81_956 ();
 b15zdnd11an1n64x5 FILLER_81_1020 ();
 b15zdnd11an1n64x5 FILLER_81_1084 ();
 b15zdnd11an1n64x5 FILLER_81_1148 ();
 b15zdnd11an1n32x5 FILLER_81_1212 ();
 b15zdnd11an1n16x5 FILLER_81_1244 ();
 b15zdnd11an1n08x5 FILLER_81_1260 ();
 b15zdnd11an1n04x5 FILLER_81_1268 ();
 b15zdnd11an1n04x5 FILLER_81_1275 ();
 b15zdnd11an1n04x5 FILLER_81_1282 ();
 b15zdnd11an1n04x5 FILLER_81_1289 ();
 b15zdnd11an1n64x5 FILLER_81_1296 ();
 b15zdnd11an1n64x5 FILLER_81_1360 ();
 b15zdnd11an1n64x5 FILLER_81_1424 ();
 b15zdnd11an1n64x5 FILLER_81_1488 ();
 b15zdnd11an1n32x5 FILLER_81_1552 ();
 b15zdnd11an1n08x5 FILLER_81_1584 ();
 b15zdnd11an1n04x5 FILLER_81_1592 ();
 b15zdnd11an1n64x5 FILLER_81_1599 ();
 b15zdnd11an1n32x5 FILLER_81_1663 ();
 b15zdnd11an1n16x5 FILLER_81_1695 ();
 b15zdnd11an1n08x5 FILLER_81_1711 ();
 b15zdnd11an1n04x5 FILLER_81_1719 ();
 b15zdnd00an1n02x5 FILLER_81_1723 ();
 b15zdnd00an1n01x5 FILLER_81_1725 ();
 b15zdnd11an1n64x5 FILLER_81_1740 ();
 b15zdnd11an1n64x5 FILLER_81_1804 ();
 b15zdnd11an1n64x5 FILLER_81_1868 ();
 b15zdnd11an1n64x5 FILLER_81_1932 ();
 b15zdnd11an1n64x5 FILLER_81_1996 ();
 b15zdnd11an1n64x5 FILLER_81_2060 ();
 b15zdnd11an1n64x5 FILLER_81_2124 ();
 b15zdnd11an1n64x5 FILLER_81_2188 ();
 b15zdnd11an1n32x5 FILLER_81_2252 ();
 b15zdnd11an1n64x5 FILLER_82_8 ();
 b15zdnd11an1n64x5 FILLER_82_72 ();
 b15zdnd11an1n64x5 FILLER_82_136 ();
 b15zdnd11an1n64x5 FILLER_82_200 ();
 b15zdnd11an1n64x5 FILLER_82_264 ();
 b15zdnd11an1n32x5 FILLER_82_328 ();
 b15zdnd11an1n16x5 FILLER_82_360 ();
 b15zdnd00an1n02x5 FILLER_82_376 ();
 b15zdnd11an1n64x5 FILLER_82_383 ();
 b15zdnd11an1n64x5 FILLER_82_447 ();
 b15zdnd11an1n64x5 FILLER_82_511 ();
 b15zdnd11an1n64x5 FILLER_82_575 ();
 b15zdnd11an1n64x5 FILLER_82_639 ();
 b15zdnd11an1n08x5 FILLER_82_703 ();
 b15zdnd11an1n04x5 FILLER_82_711 ();
 b15zdnd00an1n02x5 FILLER_82_715 ();
 b15zdnd00an1n01x5 FILLER_82_717 ();
 b15zdnd11an1n64x5 FILLER_82_726 ();
 b15zdnd11an1n64x5 FILLER_82_790 ();
 b15zdnd11an1n64x5 FILLER_82_854 ();
 b15zdnd11an1n64x5 FILLER_82_918 ();
 b15zdnd11an1n64x5 FILLER_82_982 ();
 b15zdnd11an1n64x5 FILLER_82_1046 ();
 b15zdnd11an1n32x5 FILLER_82_1110 ();
 b15zdnd11an1n16x5 FILLER_82_1142 ();
 b15zdnd11an1n04x5 FILLER_82_1158 ();
 b15zdnd00an1n02x5 FILLER_82_1162 ();
 b15zdnd11an1n64x5 FILLER_82_1178 ();
 b15zdnd11an1n16x5 FILLER_82_1242 ();
 b15zdnd11an1n04x5 FILLER_82_1258 ();
 b15zdnd11an1n64x5 FILLER_82_1314 ();
 b15zdnd11an1n32x5 FILLER_82_1378 ();
 b15zdnd11an1n04x5 FILLER_82_1410 ();
 b15zdnd11an1n04x5 FILLER_82_1434 ();
 b15zdnd11an1n08x5 FILLER_82_1452 ();
 b15zdnd00an1n02x5 FILLER_82_1460 ();
 b15zdnd00an1n01x5 FILLER_82_1462 ();
 b15zdnd11an1n16x5 FILLER_82_1466 ();
 b15zdnd11an1n04x5 FILLER_82_1482 ();
 b15zdnd00an1n02x5 FILLER_82_1486 ();
 b15zdnd00an1n01x5 FILLER_82_1488 ();
 b15zdnd11an1n64x5 FILLER_82_1497 ();
 b15zdnd11an1n64x5 FILLER_82_1561 ();
 b15zdnd11an1n64x5 FILLER_82_1625 ();
 b15zdnd11an1n32x5 FILLER_82_1689 ();
 b15zdnd11an1n04x5 FILLER_82_1721 ();
 b15zdnd00an1n02x5 FILLER_82_1725 ();
 b15zdnd00an1n01x5 FILLER_82_1727 ();
 b15zdnd11an1n04x5 FILLER_82_1735 ();
 b15zdnd11an1n04x5 FILLER_82_1748 ();
 b15zdnd00an1n01x5 FILLER_82_1752 ();
 b15zdnd11an1n64x5 FILLER_82_1757 ();
 b15zdnd11an1n16x5 FILLER_82_1821 ();
 b15zdnd11an1n08x5 FILLER_82_1837 ();
 b15zdnd11an1n64x5 FILLER_82_1853 ();
 b15zdnd11an1n64x5 FILLER_82_1917 ();
 b15zdnd11an1n64x5 FILLER_82_1981 ();
 b15zdnd11an1n32x5 FILLER_82_2045 ();
 b15zdnd11an1n08x5 FILLER_82_2077 ();
 b15zdnd00an1n01x5 FILLER_82_2085 ();
 b15zdnd11an1n64x5 FILLER_82_2090 ();
 b15zdnd11an1n64x5 FILLER_82_2162 ();
 b15zdnd11an1n32x5 FILLER_82_2226 ();
 b15zdnd11an1n16x5 FILLER_82_2258 ();
 b15zdnd00an1n02x5 FILLER_82_2274 ();
 b15zdnd11an1n64x5 FILLER_83_0 ();
 b15zdnd11an1n64x5 FILLER_83_64 ();
 b15zdnd11an1n64x5 FILLER_83_128 ();
 b15zdnd11an1n64x5 FILLER_83_192 ();
 b15zdnd11an1n64x5 FILLER_83_256 ();
 b15zdnd11an1n64x5 FILLER_83_320 ();
 b15zdnd11an1n32x5 FILLER_83_384 ();
 b15zdnd11an1n16x5 FILLER_83_416 ();
 b15zdnd11an1n08x5 FILLER_83_432 ();
 b15zdnd11an1n64x5 FILLER_83_444 ();
 b15zdnd11an1n64x5 FILLER_83_508 ();
 b15zdnd11an1n64x5 FILLER_83_572 ();
 b15zdnd11an1n64x5 FILLER_83_636 ();
 b15zdnd11an1n64x5 FILLER_83_700 ();
 b15zdnd11an1n64x5 FILLER_83_764 ();
 b15zdnd11an1n64x5 FILLER_83_828 ();
 b15zdnd11an1n32x5 FILLER_83_892 ();
 b15zdnd11an1n08x5 FILLER_83_924 ();
 b15zdnd11an1n04x5 FILLER_83_932 ();
 b15zdnd00an1n01x5 FILLER_83_936 ();
 b15zdnd11an1n64x5 FILLER_83_940 ();
 b15zdnd11an1n16x5 FILLER_83_1004 ();
 b15zdnd00an1n01x5 FILLER_83_1020 ();
 b15zdnd11an1n04x5 FILLER_83_1024 ();
 b15zdnd11an1n04x5 FILLER_83_1031 ();
 b15zdnd11an1n64x5 FILLER_83_1038 ();
 b15zdnd11an1n32x5 FILLER_83_1102 ();
 b15zdnd11an1n16x5 FILLER_83_1134 ();
 b15zdnd00an1n02x5 FILLER_83_1150 ();
 b15zdnd00an1n01x5 FILLER_83_1152 ();
 b15zdnd11an1n32x5 FILLER_83_1195 ();
 b15zdnd11an1n16x5 FILLER_83_1227 ();
 b15zdnd11an1n08x5 FILLER_83_1243 ();
 b15zdnd00an1n02x5 FILLER_83_1251 ();
 b15zdnd11an1n04x5 FILLER_83_1305 ();
 b15zdnd11an1n04x5 FILLER_83_1312 ();
 b15zdnd11an1n04x5 FILLER_83_1319 ();
 b15zdnd11an1n64x5 FILLER_83_1326 ();
 b15zdnd11an1n32x5 FILLER_83_1390 ();
 b15zdnd11an1n08x5 FILLER_83_1422 ();
 b15zdnd00an1n01x5 FILLER_83_1430 ();
 b15zdnd11an1n64x5 FILLER_83_1446 ();
 b15zdnd11an1n64x5 FILLER_83_1510 ();
 b15zdnd11an1n64x5 FILLER_83_1574 ();
 b15zdnd11an1n64x5 FILLER_83_1638 ();
 b15zdnd11an1n16x5 FILLER_83_1702 ();
 b15zdnd11an1n04x5 FILLER_83_1718 ();
 b15zdnd11an1n64x5 FILLER_83_1738 ();
 b15zdnd11an1n64x5 FILLER_83_1802 ();
 b15zdnd11an1n64x5 FILLER_83_1866 ();
 b15zdnd11an1n64x5 FILLER_83_1930 ();
 b15zdnd11an1n64x5 FILLER_83_1994 ();
 b15zdnd11an1n64x5 FILLER_83_2058 ();
 b15zdnd11an1n64x5 FILLER_83_2122 ();
 b15zdnd11an1n64x5 FILLER_83_2186 ();
 b15zdnd11an1n32x5 FILLER_83_2250 ();
 b15zdnd00an1n02x5 FILLER_83_2282 ();
 b15zdnd11an1n64x5 FILLER_84_8 ();
 b15zdnd11an1n64x5 FILLER_84_72 ();
 b15zdnd11an1n64x5 FILLER_84_136 ();
 b15zdnd11an1n16x5 FILLER_84_200 ();
 b15zdnd11an1n04x5 FILLER_84_216 ();
 b15zdnd00an1n02x5 FILLER_84_220 ();
 b15zdnd00an1n01x5 FILLER_84_222 ();
 b15zdnd11an1n64x5 FILLER_84_226 ();
 b15zdnd11an1n64x5 FILLER_84_290 ();
 b15zdnd11an1n16x5 FILLER_84_354 ();
 b15zdnd11an1n08x5 FILLER_84_370 ();
 b15zdnd00an1n02x5 FILLER_84_378 ();
 b15zdnd00an1n01x5 FILLER_84_380 ();
 b15zdnd11an1n08x5 FILLER_84_385 ();
 b15zdnd11an1n04x5 FILLER_84_393 ();
 b15zdnd00an1n01x5 FILLER_84_397 ();
 b15zdnd11an1n64x5 FILLER_84_406 ();
 b15zdnd11an1n64x5 FILLER_84_470 ();
 b15zdnd11an1n64x5 FILLER_84_534 ();
 b15zdnd11an1n16x5 FILLER_84_598 ();
 b15zdnd00an1n02x5 FILLER_84_614 ();
 b15zdnd11an1n64x5 FILLER_84_619 ();
 b15zdnd11an1n32x5 FILLER_84_683 ();
 b15zdnd00an1n02x5 FILLER_84_715 ();
 b15zdnd00an1n01x5 FILLER_84_717 ();
 b15zdnd11an1n64x5 FILLER_84_726 ();
 b15zdnd11an1n64x5 FILLER_84_790 ();
 b15zdnd11an1n32x5 FILLER_84_854 ();
 b15zdnd11an1n16x5 FILLER_84_886 ();
 b15zdnd11an1n08x5 FILLER_84_902 ();
 b15zdnd11an1n32x5 FILLER_84_962 ();
 b15zdnd11an1n08x5 FILLER_84_994 ();
 b15zdnd11an1n64x5 FILLER_84_1054 ();
 b15zdnd11an1n64x5 FILLER_84_1118 ();
 b15zdnd11an1n64x5 FILLER_84_1182 ();
 b15zdnd11an1n16x5 FILLER_84_1246 ();
 b15zdnd11an1n08x5 FILLER_84_1262 ();
 b15zdnd00an1n02x5 FILLER_84_1270 ();
 b15zdnd00an1n01x5 FILLER_84_1272 ();
 b15zdnd11an1n04x5 FILLER_84_1276 ();
 b15zdnd11an1n64x5 FILLER_84_1332 ();
 b15zdnd11an1n64x5 FILLER_84_1396 ();
 b15zdnd11an1n64x5 FILLER_84_1460 ();
 b15zdnd11an1n32x5 FILLER_84_1524 ();
 b15zdnd11an1n08x5 FILLER_84_1556 ();
 b15zdnd11an1n64x5 FILLER_84_1575 ();
 b15zdnd11an1n64x5 FILLER_84_1639 ();
 b15zdnd11an1n64x5 FILLER_84_1703 ();
 b15zdnd11an1n64x5 FILLER_84_1767 ();
 b15zdnd11an1n64x5 FILLER_84_1831 ();
 b15zdnd11an1n64x5 FILLER_84_1895 ();
 b15zdnd11an1n64x5 FILLER_84_1959 ();
 b15zdnd11an1n64x5 FILLER_84_2023 ();
 b15zdnd11an1n08x5 FILLER_84_2087 ();
 b15zdnd00an1n02x5 FILLER_84_2095 ();
 b15zdnd11an1n32x5 FILLER_84_2101 ();
 b15zdnd11an1n16x5 FILLER_84_2133 ();
 b15zdnd11an1n04x5 FILLER_84_2149 ();
 b15zdnd00an1n01x5 FILLER_84_2153 ();
 b15zdnd11an1n64x5 FILLER_84_2162 ();
 b15zdnd11an1n32x5 FILLER_84_2226 ();
 b15zdnd11an1n16x5 FILLER_84_2258 ();
 b15zdnd00an1n02x5 FILLER_84_2274 ();
 b15zdnd11an1n64x5 FILLER_85_0 ();
 b15zdnd11an1n64x5 FILLER_85_64 ();
 b15zdnd11an1n32x5 FILLER_85_128 ();
 b15zdnd11an1n16x5 FILLER_85_160 ();
 b15zdnd11an1n08x5 FILLER_85_176 ();
 b15zdnd00an1n02x5 FILLER_85_184 ();
 b15zdnd11an1n04x5 FILLER_85_226 ();
 b15zdnd11an1n64x5 FILLER_85_233 ();
 b15zdnd11an1n32x5 FILLER_85_297 ();
 b15zdnd11an1n16x5 FILLER_85_329 ();
 b15zdnd11an1n08x5 FILLER_85_345 ();
 b15zdnd11an1n04x5 FILLER_85_353 ();
 b15zdnd00an1n02x5 FILLER_85_357 ();
 b15zdnd11an1n16x5 FILLER_85_362 ();
 b15zdnd11an1n04x5 FILLER_85_378 ();
 b15zdnd11an1n64x5 FILLER_85_424 ();
 b15zdnd11an1n64x5 FILLER_85_488 ();
 b15zdnd11an1n32x5 FILLER_85_552 ();
 b15zdnd11an1n04x5 FILLER_85_584 ();
 b15zdnd00an1n01x5 FILLER_85_588 ();
 b15zdnd11an1n64x5 FILLER_85_641 ();
 b15zdnd11an1n64x5 FILLER_85_705 ();
 b15zdnd11an1n64x5 FILLER_85_769 ();
 b15zdnd11an1n64x5 FILLER_85_833 ();
 b15zdnd11an1n08x5 FILLER_85_897 ();
 b15zdnd00an1n02x5 FILLER_85_905 ();
 b15zdnd00an1n01x5 FILLER_85_907 ();
 b15zdnd11an1n32x5 FILLER_85_960 ();
 b15zdnd00an1n02x5 FILLER_85_992 ();
 b15zdnd00an1n01x5 FILLER_85_994 ();
 b15zdnd11an1n64x5 FILLER_85_1047 ();
 b15zdnd11an1n64x5 FILLER_85_1111 ();
 b15zdnd11an1n64x5 FILLER_85_1175 ();
 b15zdnd11an1n32x5 FILLER_85_1239 ();
 b15zdnd11an1n08x5 FILLER_85_1271 ();
 b15zdnd11an1n08x5 FILLER_85_1282 ();
 b15zdnd00an1n02x5 FILLER_85_1290 ();
 b15zdnd00an1n01x5 FILLER_85_1292 ();
 b15zdnd11an1n64x5 FILLER_85_1345 ();
 b15zdnd11an1n64x5 FILLER_85_1409 ();
 b15zdnd11an1n64x5 FILLER_85_1473 ();
 b15zdnd11an1n64x5 FILLER_85_1537 ();
 b15zdnd11an1n64x5 FILLER_85_1601 ();
 b15zdnd11an1n64x5 FILLER_85_1665 ();
 b15zdnd11an1n64x5 FILLER_85_1729 ();
 b15zdnd11an1n64x5 FILLER_85_1793 ();
 b15zdnd11an1n64x5 FILLER_85_1857 ();
 b15zdnd11an1n64x5 FILLER_85_1921 ();
 b15zdnd11an1n64x5 FILLER_85_1985 ();
 b15zdnd11an1n64x5 FILLER_85_2049 ();
 b15zdnd11an1n32x5 FILLER_85_2113 ();
 b15zdnd00an1n02x5 FILLER_85_2145 ();
 b15zdnd11an1n64x5 FILLER_85_2170 ();
 b15zdnd11an1n32x5 FILLER_85_2234 ();
 b15zdnd11an1n16x5 FILLER_85_2266 ();
 b15zdnd00an1n02x5 FILLER_85_2282 ();
 b15zdnd11an1n16x5 FILLER_86_8 ();
 b15zdnd11an1n08x5 FILLER_86_24 ();
 b15zdnd11an1n04x5 FILLER_86_32 ();
 b15zdnd11an1n64x5 FILLER_86_40 ();
 b15zdnd11an1n64x5 FILLER_86_104 ();
 b15zdnd11an1n64x5 FILLER_86_168 ();
 b15zdnd11an1n32x5 FILLER_86_232 ();
 b15zdnd00an1n01x5 FILLER_86_264 ();
 b15zdnd11an1n32x5 FILLER_86_269 ();
 b15zdnd11an1n16x5 FILLER_86_301 ();
 b15zdnd11an1n08x5 FILLER_86_317 ();
 b15zdnd11an1n04x5 FILLER_86_325 ();
 b15zdnd00an1n02x5 FILLER_86_329 ();
 b15zdnd00an1n01x5 FILLER_86_331 ();
 b15zdnd11an1n64x5 FILLER_86_384 ();
 b15zdnd11an1n64x5 FILLER_86_448 ();
 b15zdnd11an1n64x5 FILLER_86_512 ();
 b15zdnd11an1n32x5 FILLER_86_576 ();
 b15zdnd11an1n04x5 FILLER_86_611 ();
 b15zdnd11an1n64x5 FILLER_86_618 ();
 b15zdnd11an1n32x5 FILLER_86_682 ();
 b15zdnd11an1n04x5 FILLER_86_714 ();
 b15zdnd11an1n04x5 FILLER_86_726 ();
 b15zdnd11an1n64x5 FILLER_86_734 ();
 b15zdnd11an1n64x5 FILLER_86_798 ();
 b15zdnd11an1n64x5 FILLER_86_862 ();
 b15zdnd00an1n02x5 FILLER_86_926 ();
 b15zdnd11an1n04x5 FILLER_86_931 ();
 b15zdnd11an1n04x5 FILLER_86_938 ();
 b15zdnd11an1n64x5 FILLER_86_945 ();
 b15zdnd11an1n08x5 FILLER_86_1009 ();
 b15zdnd00an1n02x5 FILLER_86_1017 ();
 b15zdnd00an1n01x5 FILLER_86_1019 ();
 b15zdnd11an1n04x5 FILLER_86_1023 ();
 b15zdnd11an1n64x5 FILLER_86_1030 ();
 b15zdnd00an1n01x5 FILLER_86_1094 ();
 b15zdnd11an1n64x5 FILLER_86_1099 ();
 b15zdnd11an1n64x5 FILLER_86_1163 ();
 b15zdnd11an1n32x5 FILLER_86_1227 ();
 b15zdnd11an1n16x5 FILLER_86_1259 ();
 b15zdnd00an1n02x5 FILLER_86_1275 ();
 b15zdnd00an1n01x5 FILLER_86_1277 ();
 b15zdnd11an1n04x5 FILLER_86_1305 ();
 b15zdnd00an1n02x5 FILLER_86_1309 ();
 b15zdnd00an1n01x5 FILLER_86_1311 ();
 b15zdnd11an1n04x5 FILLER_86_1315 ();
 b15zdnd11an1n64x5 FILLER_86_1322 ();
 b15zdnd11an1n64x5 FILLER_86_1386 ();
 b15zdnd11an1n08x5 FILLER_86_1450 ();
 b15zdnd11an1n04x5 FILLER_86_1458 ();
 b15zdnd00an1n02x5 FILLER_86_1462 ();
 b15zdnd11an1n32x5 FILLER_86_1474 ();
 b15zdnd11an1n16x5 FILLER_86_1506 ();
 b15zdnd11an1n08x5 FILLER_86_1522 ();
 b15zdnd11an1n04x5 FILLER_86_1530 ();
 b15zdnd00an1n02x5 FILLER_86_1534 ();
 b15zdnd00an1n01x5 FILLER_86_1536 ();
 b15zdnd11an1n64x5 FILLER_86_1540 ();
 b15zdnd11an1n64x5 FILLER_86_1604 ();
 b15zdnd11an1n64x5 FILLER_86_1668 ();
 b15zdnd11an1n64x5 FILLER_86_1732 ();
 b15zdnd11an1n16x5 FILLER_86_1796 ();
 b15zdnd11an1n08x5 FILLER_86_1812 ();
 b15zdnd11an1n04x5 FILLER_86_1820 ();
 b15zdnd00an1n01x5 FILLER_86_1824 ();
 b15zdnd11an1n64x5 FILLER_86_1829 ();
 b15zdnd11an1n64x5 FILLER_86_1893 ();
 b15zdnd11an1n64x5 FILLER_86_1957 ();
 b15zdnd11an1n04x5 FILLER_86_2021 ();
 b15zdnd00an1n02x5 FILLER_86_2025 ();
 b15zdnd11an1n64x5 FILLER_86_2030 ();
 b15zdnd11an1n08x5 FILLER_86_2094 ();
 b15zdnd11an1n32x5 FILLER_86_2108 ();
 b15zdnd11an1n08x5 FILLER_86_2140 ();
 b15zdnd11an1n04x5 FILLER_86_2148 ();
 b15zdnd00an1n02x5 FILLER_86_2152 ();
 b15zdnd11an1n64x5 FILLER_86_2162 ();
 b15zdnd11an1n32x5 FILLER_86_2226 ();
 b15zdnd11an1n16x5 FILLER_86_2258 ();
 b15zdnd00an1n02x5 FILLER_86_2274 ();
 b15zdnd11an1n08x5 FILLER_87_0 ();
 b15zdnd11an1n04x5 FILLER_87_8 ();
 b15zdnd00an1n02x5 FILLER_87_12 ();
 b15zdnd11an1n64x5 FILLER_87_56 ();
 b15zdnd11an1n64x5 FILLER_87_120 ();
 b15zdnd11an1n32x5 FILLER_87_184 ();
 b15zdnd11an1n16x5 FILLER_87_216 ();
 b15zdnd11an1n08x5 FILLER_87_232 ();
 b15zdnd11an1n64x5 FILLER_87_282 ();
 b15zdnd00an1n02x5 FILLER_87_346 ();
 b15zdnd11an1n04x5 FILLER_87_351 ();
 b15zdnd00an1n02x5 FILLER_87_355 ();
 b15zdnd00an1n01x5 FILLER_87_357 ();
 b15zdnd11an1n64x5 FILLER_87_361 ();
 b15zdnd11an1n64x5 FILLER_87_425 ();
 b15zdnd11an1n64x5 FILLER_87_489 ();
 b15zdnd11an1n64x5 FILLER_87_553 ();
 b15zdnd11an1n32x5 FILLER_87_617 ();
 b15zdnd11an1n16x5 FILLER_87_649 ();
 b15zdnd11an1n04x5 FILLER_87_665 ();
 b15zdnd00an1n02x5 FILLER_87_669 ();
 b15zdnd00an1n01x5 FILLER_87_671 ();
 b15zdnd11an1n64x5 FILLER_87_682 ();
 b15zdnd11an1n64x5 FILLER_87_746 ();
 b15zdnd11an1n64x5 FILLER_87_810 ();
 b15zdnd11an1n32x5 FILLER_87_874 ();
 b15zdnd11an1n16x5 FILLER_87_906 ();
 b15zdnd11an1n04x5 FILLER_87_922 ();
 b15zdnd00an1n02x5 FILLER_87_926 ();
 b15zdnd11an1n08x5 FILLER_87_931 ();
 b15zdnd00an1n01x5 FILLER_87_939 ();
 b15zdnd11an1n64x5 FILLER_87_943 ();
 b15zdnd11an1n08x5 FILLER_87_1007 ();
 b15zdnd11an1n04x5 FILLER_87_1015 ();
 b15zdnd00an1n01x5 FILLER_87_1019 ();
 b15zdnd11an1n64x5 FILLER_87_1023 ();
 b15zdnd11an1n08x5 FILLER_87_1087 ();
 b15zdnd00an1n01x5 FILLER_87_1095 ();
 b15zdnd11an1n64x5 FILLER_87_1102 ();
 b15zdnd11an1n64x5 FILLER_87_1166 ();
 b15zdnd11an1n64x5 FILLER_87_1230 ();
 b15zdnd11an1n08x5 FILLER_87_1303 ();
 b15zdnd11an1n04x5 FILLER_87_1311 ();
 b15zdnd00an1n02x5 FILLER_87_1315 ();
 b15zdnd00an1n01x5 FILLER_87_1317 ();
 b15zdnd11an1n64x5 FILLER_87_1321 ();
 b15zdnd11an1n64x5 FILLER_87_1385 ();
 b15zdnd11an1n08x5 FILLER_87_1449 ();
 b15zdnd00an1n01x5 FILLER_87_1457 ();
 b15zdnd11an1n64x5 FILLER_87_1474 ();
 b15zdnd11an1n16x5 FILLER_87_1552 ();
 b15zdnd11an1n08x5 FILLER_87_1568 ();
 b15zdnd00an1n02x5 FILLER_87_1576 ();
 b15zdnd00an1n01x5 FILLER_87_1578 ();
 b15zdnd11an1n04x5 FILLER_87_1593 ();
 b15zdnd11an1n64x5 FILLER_87_1610 ();
 b15zdnd11an1n64x5 FILLER_87_1674 ();
 b15zdnd11an1n64x5 FILLER_87_1738 ();
 b15zdnd11an1n64x5 FILLER_87_1802 ();
 b15zdnd11an1n64x5 FILLER_87_1866 ();
 b15zdnd11an1n64x5 FILLER_87_1930 ();
 b15zdnd11an1n32x5 FILLER_87_2046 ();
 b15zdnd11an1n16x5 FILLER_87_2078 ();
 b15zdnd11an1n08x5 FILLER_87_2094 ();
 b15zdnd11an1n04x5 FILLER_87_2102 ();
 b15zdnd11an1n64x5 FILLER_87_2110 ();
 b15zdnd11an1n64x5 FILLER_87_2174 ();
 b15zdnd11an1n32x5 FILLER_87_2238 ();
 b15zdnd11an1n08x5 FILLER_87_2270 ();
 b15zdnd11an1n04x5 FILLER_87_2278 ();
 b15zdnd00an1n02x5 FILLER_87_2282 ();
 b15zdnd11an1n64x5 FILLER_88_8 ();
 b15zdnd11an1n64x5 FILLER_88_72 ();
 b15zdnd11an1n64x5 FILLER_88_136 ();
 b15zdnd11an1n64x5 FILLER_88_200 ();
 b15zdnd11an1n16x5 FILLER_88_264 ();
 b15zdnd11an1n04x5 FILLER_88_280 ();
 b15zdnd00an1n01x5 FILLER_88_284 ();
 b15zdnd11an1n64x5 FILLER_88_293 ();
 b15zdnd11an1n64x5 FILLER_88_357 ();
 b15zdnd11an1n32x5 FILLER_88_421 ();
 b15zdnd11an1n64x5 FILLER_88_456 ();
 b15zdnd11an1n64x5 FILLER_88_520 ();
 b15zdnd11an1n64x5 FILLER_88_584 ();
 b15zdnd11an1n32x5 FILLER_88_648 ();
 b15zdnd11an1n16x5 FILLER_88_680 ();
 b15zdnd11an1n08x5 FILLER_88_696 ();
 b15zdnd11an1n04x5 FILLER_88_704 ();
 b15zdnd00an1n01x5 FILLER_88_708 ();
 b15zdnd11an1n04x5 FILLER_88_713 ();
 b15zdnd00an1n01x5 FILLER_88_717 ();
 b15zdnd11an1n64x5 FILLER_88_726 ();
 b15zdnd11an1n64x5 FILLER_88_790 ();
 b15zdnd11an1n64x5 FILLER_88_854 ();
 b15zdnd11an1n64x5 FILLER_88_918 ();
 b15zdnd11an1n64x5 FILLER_88_982 ();
 b15zdnd11an1n64x5 FILLER_88_1046 ();
 b15zdnd11an1n64x5 FILLER_88_1110 ();
 b15zdnd11an1n64x5 FILLER_88_1174 ();
 b15zdnd11an1n64x5 FILLER_88_1238 ();
 b15zdnd11an1n64x5 FILLER_88_1302 ();
 b15zdnd11an1n64x5 FILLER_88_1366 ();
 b15zdnd11an1n64x5 FILLER_88_1430 ();
 b15zdnd11an1n64x5 FILLER_88_1494 ();
 b15zdnd11an1n64x5 FILLER_88_1558 ();
 b15zdnd11an1n64x5 FILLER_88_1622 ();
 b15zdnd11an1n64x5 FILLER_88_1686 ();
 b15zdnd11an1n16x5 FILLER_88_1750 ();
 b15zdnd11an1n08x5 FILLER_88_1766 ();
 b15zdnd00an1n02x5 FILLER_88_1774 ();
 b15zdnd11an1n32x5 FILLER_88_1821 ();
 b15zdnd11an1n08x5 FILLER_88_1853 ();
 b15zdnd11an1n04x5 FILLER_88_1864 ();
 b15zdnd11an1n64x5 FILLER_88_1871 ();
 b15zdnd11an1n64x5 FILLER_88_1935 ();
 b15zdnd00an1n02x5 FILLER_88_1999 ();
 b15zdnd11an1n64x5 FILLER_88_2053 ();
 b15zdnd11an1n32x5 FILLER_88_2117 ();
 b15zdnd11an1n04x5 FILLER_88_2149 ();
 b15zdnd00an1n01x5 FILLER_88_2153 ();
 b15zdnd11an1n64x5 FILLER_88_2162 ();
 b15zdnd11an1n32x5 FILLER_88_2226 ();
 b15zdnd11an1n16x5 FILLER_88_2258 ();
 b15zdnd00an1n02x5 FILLER_88_2274 ();
 b15zdnd11an1n64x5 FILLER_89_0 ();
 b15zdnd11an1n64x5 FILLER_89_64 ();
 b15zdnd11an1n64x5 FILLER_89_128 ();
 b15zdnd11an1n64x5 FILLER_89_192 ();
 b15zdnd11an1n04x5 FILLER_89_256 ();
 b15zdnd00an1n02x5 FILLER_89_260 ();
 b15zdnd11an1n64x5 FILLER_89_301 ();
 b15zdnd11an1n32x5 FILLER_89_365 ();
 b15zdnd11an1n16x5 FILLER_89_397 ();
 b15zdnd11an1n04x5 FILLER_89_413 ();
 b15zdnd11an1n04x5 FILLER_89_457 ();
 b15zdnd11an1n64x5 FILLER_89_464 ();
 b15zdnd11an1n64x5 FILLER_89_528 ();
 b15zdnd11an1n64x5 FILLER_89_592 ();
 b15zdnd11an1n64x5 FILLER_89_656 ();
 b15zdnd11an1n64x5 FILLER_89_720 ();
 b15zdnd11an1n04x5 FILLER_89_784 ();
 b15zdnd00an1n01x5 FILLER_89_788 ();
 b15zdnd11an1n16x5 FILLER_89_792 ();
 b15zdnd11an1n64x5 FILLER_89_811 ();
 b15zdnd11an1n32x5 FILLER_89_875 ();
 b15zdnd11an1n16x5 FILLER_89_907 ();
 b15zdnd11an1n08x5 FILLER_89_923 ();
 b15zdnd11an1n04x5 FILLER_89_931 ();
 b15zdnd00an1n02x5 FILLER_89_935 ();
 b15zdnd00an1n01x5 FILLER_89_937 ();
 b15zdnd11an1n64x5 FILLER_89_942 ();
 b15zdnd11an1n64x5 FILLER_89_1006 ();
 b15zdnd11an1n64x5 FILLER_89_1070 ();
 b15zdnd11an1n64x5 FILLER_89_1134 ();
 b15zdnd11an1n64x5 FILLER_89_1198 ();
 b15zdnd11an1n64x5 FILLER_89_1262 ();
 b15zdnd11an1n64x5 FILLER_89_1326 ();
 b15zdnd11an1n64x5 FILLER_89_1390 ();
 b15zdnd11an1n64x5 FILLER_89_1454 ();
 b15zdnd11an1n08x5 FILLER_89_1518 ();
 b15zdnd00an1n02x5 FILLER_89_1526 ();
 b15zdnd00an1n01x5 FILLER_89_1528 ();
 b15zdnd11an1n64x5 FILLER_89_1543 ();
 b15zdnd11an1n64x5 FILLER_89_1607 ();
 b15zdnd11an1n64x5 FILLER_89_1671 ();
 b15zdnd11an1n64x5 FILLER_89_1735 ();
 b15zdnd11an1n32x5 FILLER_89_1799 ();
 b15zdnd11an1n08x5 FILLER_89_1831 ();
 b15zdnd11an1n04x5 FILLER_89_1839 ();
 b15zdnd11an1n04x5 FILLER_89_1895 ();
 b15zdnd11an1n64x5 FILLER_89_1902 ();
 b15zdnd11an1n32x5 FILLER_89_1966 ();
 b15zdnd11an1n08x5 FILLER_89_1998 ();
 b15zdnd11an1n04x5 FILLER_89_2006 ();
 b15zdnd00an1n02x5 FILLER_89_2010 ();
 b15zdnd11an1n04x5 FILLER_89_2015 ();
 b15zdnd11an1n04x5 FILLER_89_2022 ();
 b15zdnd11an1n32x5 FILLER_89_2029 ();
 b15zdnd11an1n08x5 FILLER_89_2061 ();
 b15zdnd00an1n02x5 FILLER_89_2069 ();
 b15zdnd00an1n01x5 FILLER_89_2071 ();
 b15zdnd11an1n64x5 FILLER_89_2083 ();
 b15zdnd11an1n64x5 FILLER_89_2147 ();
 b15zdnd11an1n64x5 FILLER_89_2211 ();
 b15zdnd11an1n08x5 FILLER_89_2275 ();
 b15zdnd00an1n01x5 FILLER_89_2283 ();
 b15zdnd11an1n64x5 FILLER_90_8 ();
 b15zdnd11an1n64x5 FILLER_90_72 ();
 b15zdnd11an1n64x5 FILLER_90_136 ();
 b15zdnd11an1n32x5 FILLER_90_200 ();
 b15zdnd11an1n08x5 FILLER_90_232 ();
 b15zdnd11an1n04x5 FILLER_90_240 ();
 b15zdnd00an1n02x5 FILLER_90_244 ();
 b15zdnd00an1n01x5 FILLER_90_246 ();
 b15zdnd11an1n64x5 FILLER_90_289 ();
 b15zdnd11an1n64x5 FILLER_90_353 ();
 b15zdnd11an1n64x5 FILLER_90_417 ();
 b15zdnd11an1n64x5 FILLER_90_481 ();
 b15zdnd11an1n04x5 FILLER_90_545 ();
 b15zdnd00an1n02x5 FILLER_90_549 ();
 b15zdnd11an1n04x5 FILLER_90_569 ();
 b15zdnd11an1n08x5 FILLER_90_604 ();
 b15zdnd11an1n16x5 FILLER_90_622 ();
 b15zdnd00an1n02x5 FILLER_90_638 ();
 b15zdnd00an1n01x5 FILLER_90_640 ();
 b15zdnd11an1n04x5 FILLER_90_648 ();
 b15zdnd11an1n32x5 FILLER_90_663 ();
 b15zdnd11an1n16x5 FILLER_90_695 ();
 b15zdnd11an1n04x5 FILLER_90_711 ();
 b15zdnd00an1n02x5 FILLER_90_715 ();
 b15zdnd00an1n01x5 FILLER_90_717 ();
 b15zdnd11an1n08x5 FILLER_90_726 ();
 b15zdnd11an1n04x5 FILLER_90_734 ();
 b15zdnd00an1n01x5 FILLER_90_738 ();
 b15zdnd11an1n04x5 FILLER_90_760 ();
 b15zdnd11an1n16x5 FILLER_90_767 ();
 b15zdnd11an1n04x5 FILLER_90_783 ();
 b15zdnd00an1n01x5 FILLER_90_787 ();
 b15zdnd11an1n64x5 FILLER_90_840 ();
 b15zdnd11an1n64x5 FILLER_90_904 ();
 b15zdnd11an1n64x5 FILLER_90_968 ();
 b15zdnd11an1n64x5 FILLER_90_1032 ();
 b15zdnd11an1n32x5 FILLER_90_1096 ();
 b15zdnd11an1n08x5 FILLER_90_1128 ();
 b15zdnd11an1n04x5 FILLER_90_1136 ();
 b15zdnd11an1n64x5 FILLER_90_1160 ();
 b15zdnd11an1n64x5 FILLER_90_1224 ();
 b15zdnd11an1n64x5 FILLER_90_1288 ();
 b15zdnd11an1n32x5 FILLER_90_1352 ();
 b15zdnd11an1n08x5 FILLER_90_1384 ();
 b15zdnd11an1n04x5 FILLER_90_1392 ();
 b15zdnd00an1n02x5 FILLER_90_1396 ();
 b15zdnd00an1n01x5 FILLER_90_1398 ();
 b15zdnd11an1n64x5 FILLER_90_1403 ();
 b15zdnd11an1n64x5 FILLER_90_1467 ();
 b15zdnd11an1n32x5 FILLER_90_1531 ();
 b15zdnd11an1n16x5 FILLER_90_1563 ();
 b15zdnd11an1n08x5 FILLER_90_1579 ();
 b15zdnd11an1n04x5 FILLER_90_1587 ();
 b15zdnd00an1n01x5 FILLER_90_1591 ();
 b15zdnd11an1n64x5 FILLER_90_1608 ();
 b15zdnd11an1n64x5 FILLER_90_1672 ();
 b15zdnd11an1n64x5 FILLER_90_1736 ();
 b15zdnd11an1n32x5 FILLER_90_1800 ();
 b15zdnd11an1n16x5 FILLER_90_1832 ();
 b15zdnd11an1n08x5 FILLER_90_1848 ();
 b15zdnd11an1n04x5 FILLER_90_1856 ();
 b15zdnd11an1n04x5 FILLER_90_1863 ();
 b15zdnd11an1n64x5 FILLER_90_1919 ();
 b15zdnd11an1n16x5 FILLER_90_1983 ();
 b15zdnd11an1n04x5 FILLER_90_1999 ();
 b15zdnd00an1n01x5 FILLER_90_2003 ();
 b15zdnd11an1n04x5 FILLER_90_2011 ();
 b15zdnd11an1n08x5 FILLER_90_2018 ();
 b15zdnd11an1n64x5 FILLER_90_2029 ();
 b15zdnd11an1n32x5 FILLER_90_2093 ();
 b15zdnd11an1n16x5 FILLER_90_2125 ();
 b15zdnd11an1n08x5 FILLER_90_2141 ();
 b15zdnd11an1n04x5 FILLER_90_2149 ();
 b15zdnd00an1n01x5 FILLER_90_2153 ();
 b15zdnd11an1n64x5 FILLER_90_2162 ();
 b15zdnd11an1n32x5 FILLER_90_2226 ();
 b15zdnd11an1n16x5 FILLER_90_2258 ();
 b15zdnd00an1n02x5 FILLER_90_2274 ();
 b15zdnd11an1n64x5 FILLER_91_0 ();
 b15zdnd11an1n64x5 FILLER_91_64 ();
 b15zdnd11an1n64x5 FILLER_91_128 ();
 b15zdnd11an1n64x5 FILLER_91_192 ();
 b15zdnd11an1n64x5 FILLER_91_256 ();
 b15zdnd11an1n64x5 FILLER_91_320 ();
 b15zdnd11an1n64x5 FILLER_91_384 ();
 b15zdnd11an1n64x5 FILLER_91_448 ();
 b15zdnd11an1n32x5 FILLER_91_512 ();
 b15zdnd11an1n08x5 FILLER_91_544 ();
 b15zdnd11an1n04x5 FILLER_91_552 ();
 b15zdnd00an1n01x5 FILLER_91_556 ();
 b15zdnd11an1n64x5 FILLER_91_567 ();
 b15zdnd11an1n64x5 FILLER_91_631 ();
 b15zdnd11an1n32x5 FILLER_91_695 ();
 b15zdnd11an1n16x5 FILLER_91_727 ();
 b15zdnd11an1n08x5 FILLER_91_743 ();
 b15zdnd11an1n04x5 FILLER_91_754 ();
 b15zdnd11an1n04x5 FILLER_91_761 ();
 b15zdnd11an1n04x5 FILLER_91_817 ();
 b15zdnd11an1n64x5 FILLER_91_824 ();
 b15zdnd11an1n32x5 FILLER_91_888 ();
 b15zdnd11an1n08x5 FILLER_91_920 ();
 b15zdnd11an1n04x5 FILLER_91_928 ();
 b15zdnd00an1n01x5 FILLER_91_932 ();
 b15zdnd11an1n64x5 FILLER_91_937 ();
 b15zdnd11an1n64x5 FILLER_91_1001 ();
 b15zdnd11an1n64x5 FILLER_91_1065 ();
 b15zdnd11an1n04x5 FILLER_91_1129 ();
 b15zdnd11an1n64x5 FILLER_91_1145 ();
 b15zdnd11an1n64x5 FILLER_91_1209 ();
 b15zdnd11an1n64x5 FILLER_91_1273 ();
 b15zdnd11an1n64x5 FILLER_91_1337 ();
 b15zdnd11an1n64x5 FILLER_91_1401 ();
 b15zdnd11an1n16x5 FILLER_91_1465 ();
 b15zdnd11an1n04x5 FILLER_91_1481 ();
 b15zdnd11an1n64x5 FILLER_91_1499 ();
 b15zdnd11an1n64x5 FILLER_91_1563 ();
 b15zdnd11an1n64x5 FILLER_91_1627 ();
 b15zdnd11an1n16x5 FILLER_91_1691 ();
 b15zdnd11an1n08x5 FILLER_91_1707 ();
 b15zdnd11an1n64x5 FILLER_91_1723 ();
 b15zdnd11an1n64x5 FILLER_91_1787 ();
 b15zdnd11an1n32x5 FILLER_91_1851 ();
 b15zdnd00an1n02x5 FILLER_91_1883 ();
 b15zdnd00an1n01x5 FILLER_91_1885 ();
 b15zdnd11an1n04x5 FILLER_91_1889 ();
 b15zdnd11an1n64x5 FILLER_91_1896 ();
 b15zdnd11an1n64x5 FILLER_91_1960 ();
 b15zdnd11an1n64x5 FILLER_91_2024 ();
 b15zdnd11an1n64x5 FILLER_91_2088 ();
 b15zdnd11an1n64x5 FILLER_91_2152 ();
 b15zdnd11an1n64x5 FILLER_91_2216 ();
 b15zdnd11an1n04x5 FILLER_91_2280 ();
 b15zdnd11an1n64x5 FILLER_92_8 ();
 b15zdnd11an1n64x5 FILLER_92_72 ();
 b15zdnd11an1n64x5 FILLER_92_136 ();
 b15zdnd11an1n64x5 FILLER_92_200 ();
 b15zdnd11an1n64x5 FILLER_92_264 ();
 b15zdnd11an1n16x5 FILLER_92_328 ();
 b15zdnd11an1n08x5 FILLER_92_344 ();
 b15zdnd11an1n32x5 FILLER_92_394 ();
 b15zdnd11an1n16x5 FILLER_92_426 ();
 b15zdnd11an1n08x5 FILLER_92_442 ();
 b15zdnd00an1n02x5 FILLER_92_450 ();
 b15zdnd00an1n01x5 FILLER_92_452 ();
 b15zdnd11an1n16x5 FILLER_92_505 ();
 b15zdnd11an1n64x5 FILLER_92_552 ();
 b15zdnd11an1n64x5 FILLER_92_616 ();
 b15zdnd11an1n32x5 FILLER_92_680 ();
 b15zdnd11an1n04x5 FILLER_92_712 ();
 b15zdnd00an1n02x5 FILLER_92_716 ();
 b15zdnd11an1n08x5 FILLER_92_726 ();
 b15zdnd11an1n04x5 FILLER_92_734 ();
 b15zdnd11an1n04x5 FILLER_92_790 ();
 b15zdnd11an1n08x5 FILLER_92_797 ();
 b15zdnd00an1n02x5 FILLER_92_805 ();
 b15zdnd00an1n01x5 FILLER_92_807 ();
 b15zdnd11an1n64x5 FILLER_92_811 ();
 b15zdnd11an1n32x5 FILLER_92_875 ();
 b15zdnd11an1n08x5 FILLER_92_907 ();
 b15zdnd11an1n32x5 FILLER_92_919 ();
 b15zdnd11an1n08x5 FILLER_92_951 ();
 b15zdnd11an1n64x5 FILLER_92_1001 ();
 b15zdnd11an1n32x5 FILLER_92_1065 ();
 b15zdnd11an1n16x5 FILLER_92_1097 ();
 b15zdnd11an1n08x5 FILLER_92_1113 ();
 b15zdnd00an1n02x5 FILLER_92_1121 ();
 b15zdnd00an1n01x5 FILLER_92_1123 ();
 b15zdnd11an1n32x5 FILLER_92_1144 ();
 b15zdnd11an1n64x5 FILLER_92_1179 ();
 b15zdnd11an1n64x5 FILLER_92_1243 ();
 b15zdnd11an1n64x5 FILLER_92_1307 ();
 b15zdnd11an1n64x5 FILLER_92_1371 ();
 b15zdnd11an1n32x5 FILLER_92_1435 ();
 b15zdnd11an1n08x5 FILLER_92_1467 ();
 b15zdnd00an1n02x5 FILLER_92_1475 ();
 b15zdnd00an1n01x5 FILLER_92_1477 ();
 b15zdnd11an1n64x5 FILLER_92_1506 ();
 b15zdnd11an1n16x5 FILLER_92_1570 ();
 b15zdnd00an1n01x5 FILLER_92_1586 ();
 b15zdnd11an1n04x5 FILLER_92_1595 ();
 b15zdnd11an1n32x5 FILLER_92_1608 ();
 b15zdnd11an1n16x5 FILLER_92_1640 ();
 b15zdnd00an1n02x5 FILLER_92_1656 ();
 b15zdnd00an1n01x5 FILLER_92_1658 ();
 b15zdnd11an1n64x5 FILLER_92_1683 ();
 b15zdnd11an1n64x5 FILLER_92_1747 ();
 b15zdnd11an1n16x5 FILLER_92_1811 ();
 b15zdnd11an1n08x5 FILLER_92_1827 ();
 b15zdnd11an1n04x5 FILLER_92_1835 ();
 b15zdnd00an1n02x5 FILLER_92_1839 ();
 b15zdnd00an1n01x5 FILLER_92_1841 ();
 b15zdnd11an1n32x5 FILLER_92_1845 ();
 b15zdnd11an1n16x5 FILLER_92_1877 ();
 b15zdnd11an1n08x5 FILLER_92_1893 ();
 b15zdnd11an1n04x5 FILLER_92_1901 ();
 b15zdnd11an1n32x5 FILLER_92_1914 ();
 b15zdnd11an1n08x5 FILLER_92_1946 ();
 b15zdnd11an1n04x5 FILLER_92_1954 ();
 b15zdnd00an1n02x5 FILLER_92_1958 ();
 b15zdnd11an1n64x5 FILLER_92_1969 ();
 b15zdnd11an1n64x5 FILLER_92_2033 ();
 b15zdnd11an1n32x5 FILLER_92_2097 ();
 b15zdnd11an1n16x5 FILLER_92_2129 ();
 b15zdnd11an1n08x5 FILLER_92_2145 ();
 b15zdnd00an1n01x5 FILLER_92_2153 ();
 b15zdnd11an1n64x5 FILLER_92_2162 ();
 b15zdnd11an1n32x5 FILLER_92_2226 ();
 b15zdnd11an1n16x5 FILLER_92_2258 ();
 b15zdnd00an1n02x5 FILLER_92_2274 ();
 b15zdnd11an1n64x5 FILLER_93_0 ();
 b15zdnd11an1n64x5 FILLER_93_64 ();
 b15zdnd11an1n64x5 FILLER_93_128 ();
 b15zdnd11an1n64x5 FILLER_93_192 ();
 b15zdnd11an1n64x5 FILLER_93_256 ();
 b15zdnd11an1n64x5 FILLER_93_320 ();
 b15zdnd11an1n64x5 FILLER_93_384 ();
 b15zdnd11an1n16x5 FILLER_93_448 ();
 b15zdnd11an1n08x5 FILLER_93_464 ();
 b15zdnd11an1n04x5 FILLER_93_472 ();
 b15zdnd11an1n04x5 FILLER_93_479 ();
 b15zdnd11an1n64x5 FILLER_93_486 ();
 b15zdnd11an1n04x5 FILLER_93_550 ();
 b15zdnd00an1n01x5 FILLER_93_554 ();
 b15zdnd11an1n64x5 FILLER_93_561 ();
 b15zdnd11an1n64x5 FILLER_93_625 ();
 b15zdnd11an1n32x5 FILLER_93_689 ();
 b15zdnd11an1n16x5 FILLER_93_721 ();
 b15zdnd11an1n08x5 FILLER_93_737 ();
 b15zdnd00an1n02x5 FILLER_93_745 ();
 b15zdnd00an1n01x5 FILLER_93_747 ();
 b15zdnd11an1n32x5 FILLER_93_754 ();
 b15zdnd11an1n04x5 FILLER_93_786 ();
 b15zdnd00an1n01x5 FILLER_93_790 ();
 b15zdnd11an1n64x5 FILLER_93_794 ();
 b15zdnd11an1n64x5 FILLER_93_858 ();
 b15zdnd11an1n64x5 FILLER_93_922 ();
 b15zdnd11an1n64x5 FILLER_93_986 ();
 b15zdnd11an1n64x5 FILLER_93_1050 ();
 b15zdnd11an1n32x5 FILLER_93_1114 ();
 b15zdnd11an1n08x5 FILLER_93_1149 ();
 b15zdnd11an1n04x5 FILLER_93_1157 ();
 b15zdnd00an1n02x5 FILLER_93_1161 ();
 b15zdnd00an1n01x5 FILLER_93_1163 ();
 b15zdnd11an1n64x5 FILLER_93_1178 ();
 b15zdnd11an1n64x5 FILLER_93_1242 ();
 b15zdnd11an1n64x5 FILLER_93_1306 ();
 b15zdnd11an1n64x5 FILLER_93_1370 ();
 b15zdnd11an1n32x5 FILLER_93_1434 ();
 b15zdnd11an1n04x5 FILLER_93_1490 ();
 b15zdnd11an1n32x5 FILLER_93_1501 ();
 b15zdnd11an1n04x5 FILLER_93_1533 ();
 b15zdnd00an1n01x5 FILLER_93_1537 ();
 b15zdnd11an1n64x5 FILLER_93_1551 ();
 b15zdnd11an1n64x5 FILLER_93_1615 ();
 b15zdnd11an1n64x5 FILLER_93_1679 ();
 b15zdnd11an1n64x5 FILLER_93_1743 ();
 b15zdnd11an1n32x5 FILLER_93_1807 ();
 b15zdnd00an1n02x5 FILLER_93_1839 ();
 b15zdnd00an1n01x5 FILLER_93_1841 ();
 b15zdnd11an1n64x5 FILLER_93_1869 ();
 b15zdnd11an1n08x5 FILLER_93_1933 ();
 b15zdnd00an1n02x5 FILLER_93_1941 ();
 b15zdnd11an1n64x5 FILLER_93_1952 ();
 b15zdnd11an1n64x5 FILLER_93_2016 ();
 b15zdnd11an1n64x5 FILLER_93_2080 ();
 b15zdnd11an1n64x5 FILLER_93_2144 ();
 b15zdnd11an1n64x5 FILLER_93_2208 ();
 b15zdnd11an1n08x5 FILLER_93_2272 ();
 b15zdnd11an1n04x5 FILLER_93_2280 ();
 b15zdnd11an1n64x5 FILLER_94_8 ();
 b15zdnd11an1n64x5 FILLER_94_72 ();
 b15zdnd11an1n64x5 FILLER_94_136 ();
 b15zdnd11an1n64x5 FILLER_94_200 ();
 b15zdnd11an1n64x5 FILLER_94_264 ();
 b15zdnd11an1n64x5 FILLER_94_328 ();
 b15zdnd11an1n64x5 FILLER_94_392 ();
 b15zdnd11an1n16x5 FILLER_94_456 ();
 b15zdnd00an1n02x5 FILLER_94_472 ();
 b15zdnd00an1n01x5 FILLER_94_474 ();
 b15zdnd11an1n64x5 FILLER_94_478 ();
 b15zdnd11an1n64x5 FILLER_94_542 ();
 b15zdnd11an1n64x5 FILLER_94_606 ();
 b15zdnd11an1n32x5 FILLER_94_670 ();
 b15zdnd11an1n16x5 FILLER_94_702 ();
 b15zdnd11an1n64x5 FILLER_94_726 ();
 b15zdnd11an1n64x5 FILLER_94_790 ();
 b15zdnd11an1n64x5 FILLER_94_854 ();
 b15zdnd11an1n64x5 FILLER_94_918 ();
 b15zdnd11an1n64x5 FILLER_94_982 ();
 b15zdnd11an1n64x5 FILLER_94_1046 ();
 b15zdnd11an1n16x5 FILLER_94_1110 ();
 b15zdnd11an1n08x5 FILLER_94_1126 ();
 b15zdnd00an1n01x5 FILLER_94_1134 ();
 b15zdnd11an1n64x5 FILLER_94_1149 ();
 b15zdnd11an1n64x5 FILLER_94_1213 ();
 b15zdnd11an1n32x5 FILLER_94_1277 ();
 b15zdnd11an1n04x5 FILLER_94_1309 ();
 b15zdnd00an1n01x5 FILLER_94_1313 ();
 b15zdnd11an1n64x5 FILLER_94_1323 ();
 b15zdnd11an1n64x5 FILLER_94_1387 ();
 b15zdnd11an1n64x5 FILLER_94_1451 ();
 b15zdnd11an1n32x5 FILLER_94_1515 ();
 b15zdnd00an1n01x5 FILLER_94_1547 ();
 b15zdnd11an1n64x5 FILLER_94_1551 ();
 b15zdnd11an1n16x5 FILLER_94_1615 ();
 b15zdnd11an1n08x5 FILLER_94_1631 ();
 b15zdnd11an1n04x5 FILLER_94_1639 ();
 b15zdnd00an1n02x5 FILLER_94_1643 ();
 b15zdnd11an1n16x5 FILLER_94_1676 ();
 b15zdnd11an1n04x5 FILLER_94_1692 ();
 b15zdnd00an1n02x5 FILLER_94_1696 ();
 b15zdnd11an1n16x5 FILLER_94_1704 ();
 b15zdnd11an1n08x5 FILLER_94_1720 ();
 b15zdnd11an1n64x5 FILLER_94_1734 ();
 b15zdnd11an1n64x5 FILLER_94_1798 ();
 b15zdnd11an1n08x5 FILLER_94_1862 ();
 b15zdnd00an1n01x5 FILLER_94_1870 ();
 b15zdnd11an1n64x5 FILLER_94_1874 ();
 b15zdnd11an1n64x5 FILLER_94_1938 ();
 b15zdnd11an1n64x5 FILLER_94_2002 ();
 b15zdnd11an1n64x5 FILLER_94_2066 ();
 b15zdnd11an1n16x5 FILLER_94_2130 ();
 b15zdnd11an1n08x5 FILLER_94_2146 ();
 b15zdnd11an1n64x5 FILLER_94_2162 ();
 b15zdnd11an1n32x5 FILLER_94_2226 ();
 b15zdnd11an1n16x5 FILLER_94_2258 ();
 b15zdnd00an1n02x5 FILLER_94_2274 ();
 b15zdnd11an1n64x5 FILLER_95_0 ();
 b15zdnd11an1n64x5 FILLER_95_64 ();
 b15zdnd11an1n64x5 FILLER_95_128 ();
 b15zdnd11an1n64x5 FILLER_95_192 ();
 b15zdnd11an1n32x5 FILLER_95_256 ();
 b15zdnd11an1n08x5 FILLER_95_288 ();
 b15zdnd11an1n64x5 FILLER_95_302 ();
 b15zdnd11an1n64x5 FILLER_95_366 ();
 b15zdnd11an1n64x5 FILLER_95_430 ();
 b15zdnd11an1n64x5 FILLER_95_494 ();
 b15zdnd11an1n64x5 FILLER_95_558 ();
 b15zdnd11an1n64x5 FILLER_95_622 ();
 b15zdnd11an1n64x5 FILLER_95_686 ();
 b15zdnd11an1n64x5 FILLER_95_750 ();
 b15zdnd11an1n64x5 FILLER_95_814 ();
 b15zdnd11an1n64x5 FILLER_95_878 ();
 b15zdnd11an1n64x5 FILLER_95_942 ();
 b15zdnd11an1n64x5 FILLER_95_1006 ();
 b15zdnd11an1n32x5 FILLER_95_1070 ();
 b15zdnd11an1n16x5 FILLER_95_1102 ();
 b15zdnd11an1n08x5 FILLER_95_1118 ();
 b15zdnd11an1n04x5 FILLER_95_1126 ();
 b15zdnd00an1n02x5 FILLER_95_1130 ();
 b15zdnd00an1n01x5 FILLER_95_1132 ();
 b15zdnd11an1n64x5 FILLER_95_1150 ();
 b15zdnd11an1n64x5 FILLER_95_1214 ();
 b15zdnd11an1n64x5 FILLER_95_1278 ();
 b15zdnd11an1n64x5 FILLER_95_1342 ();
 b15zdnd11an1n64x5 FILLER_95_1406 ();
 b15zdnd11an1n64x5 FILLER_95_1470 ();
 b15zdnd11an1n64x5 FILLER_95_1534 ();
 b15zdnd11an1n64x5 FILLER_95_1598 ();
 b15zdnd11an1n64x5 FILLER_95_1674 ();
 b15zdnd11an1n64x5 FILLER_95_1738 ();
 b15zdnd11an1n32x5 FILLER_95_1802 ();
 b15zdnd11an1n08x5 FILLER_95_1834 ();
 b15zdnd11an1n04x5 FILLER_95_1842 ();
 b15zdnd00an1n02x5 FILLER_95_1846 ();
 b15zdnd00an1n01x5 FILLER_95_1848 ();
 b15zdnd11an1n08x5 FILLER_95_1852 ();
 b15zdnd11an1n04x5 FILLER_95_1860 ();
 b15zdnd11an1n04x5 FILLER_95_1867 ();
 b15zdnd11an1n64x5 FILLER_95_1874 ();
 b15zdnd11an1n64x5 FILLER_95_1938 ();
 b15zdnd11an1n08x5 FILLER_95_2002 ();
 b15zdnd00an1n02x5 FILLER_95_2010 ();
 b15zdnd11an1n04x5 FILLER_95_2015 ();
 b15zdnd11an1n64x5 FILLER_95_2022 ();
 b15zdnd11an1n64x5 FILLER_95_2086 ();
 b15zdnd11an1n64x5 FILLER_95_2150 ();
 b15zdnd11an1n64x5 FILLER_95_2214 ();
 b15zdnd11an1n04x5 FILLER_95_2278 ();
 b15zdnd00an1n02x5 FILLER_95_2282 ();
 b15zdnd11an1n64x5 FILLER_96_8 ();
 b15zdnd11an1n64x5 FILLER_96_72 ();
 b15zdnd11an1n64x5 FILLER_96_136 ();
 b15zdnd11an1n64x5 FILLER_96_200 ();
 b15zdnd11an1n64x5 FILLER_96_264 ();
 b15zdnd11an1n64x5 FILLER_96_328 ();
 b15zdnd11an1n64x5 FILLER_96_392 ();
 b15zdnd11an1n64x5 FILLER_96_456 ();
 b15zdnd11an1n64x5 FILLER_96_520 ();
 b15zdnd11an1n64x5 FILLER_96_584 ();
 b15zdnd11an1n64x5 FILLER_96_648 ();
 b15zdnd11an1n04x5 FILLER_96_712 ();
 b15zdnd00an1n02x5 FILLER_96_716 ();
 b15zdnd11an1n64x5 FILLER_96_726 ();
 b15zdnd11an1n64x5 FILLER_96_790 ();
 b15zdnd11an1n64x5 FILLER_96_854 ();
 b15zdnd11an1n64x5 FILLER_96_918 ();
 b15zdnd11an1n64x5 FILLER_96_982 ();
 b15zdnd11an1n64x5 FILLER_96_1046 ();
 b15zdnd11an1n32x5 FILLER_96_1110 ();
 b15zdnd11an1n16x5 FILLER_96_1142 ();
 b15zdnd11an1n08x5 FILLER_96_1158 ();
 b15zdnd11an1n04x5 FILLER_96_1166 ();
 b15zdnd00an1n02x5 FILLER_96_1170 ();
 b15zdnd11an1n64x5 FILLER_96_1190 ();
 b15zdnd11an1n64x5 FILLER_96_1254 ();
 b15zdnd11an1n64x5 FILLER_96_1318 ();
 b15zdnd11an1n64x5 FILLER_96_1382 ();
 b15zdnd11an1n64x5 FILLER_96_1446 ();
 b15zdnd11an1n64x5 FILLER_96_1510 ();
 b15zdnd11an1n64x5 FILLER_96_1574 ();
 b15zdnd11an1n04x5 FILLER_96_1638 ();
 b15zdnd00an1n02x5 FILLER_96_1642 ();
 b15zdnd11an1n04x5 FILLER_96_1661 ();
 b15zdnd00an1n01x5 FILLER_96_1665 ();
 b15zdnd11an1n16x5 FILLER_96_1708 ();
 b15zdnd11an1n04x5 FILLER_96_1724 ();
 b15zdnd00an1n01x5 FILLER_96_1728 ();
 b15zdnd11an1n64x5 FILLER_96_1735 ();
 b15zdnd11an1n32x5 FILLER_96_1799 ();
 b15zdnd11an1n08x5 FILLER_96_1831 ();
 b15zdnd11an1n04x5 FILLER_96_1839 ();
 b15zdnd00an1n02x5 FILLER_96_1843 ();
 b15zdnd00an1n01x5 FILLER_96_1845 ();
 b15zdnd11an1n32x5 FILLER_96_1898 ();
 b15zdnd11an1n08x5 FILLER_96_1930 ();
 b15zdnd11an1n04x5 FILLER_96_1938 ();
 b15zdnd11an1n32x5 FILLER_96_1951 ();
 b15zdnd11an1n08x5 FILLER_96_1983 ();
 b15zdnd00an1n02x5 FILLER_96_1991 ();
 b15zdnd00an1n01x5 FILLER_96_1993 ();
 b15zdnd11an1n64x5 FILLER_96_2046 ();
 b15zdnd11an1n32x5 FILLER_96_2110 ();
 b15zdnd11an1n08x5 FILLER_96_2142 ();
 b15zdnd11an1n04x5 FILLER_96_2150 ();
 b15zdnd11an1n64x5 FILLER_96_2162 ();
 b15zdnd11an1n32x5 FILLER_96_2226 ();
 b15zdnd11an1n16x5 FILLER_96_2258 ();
 b15zdnd00an1n02x5 FILLER_96_2274 ();
 b15zdnd11an1n64x5 FILLER_97_0 ();
 b15zdnd11an1n64x5 FILLER_97_64 ();
 b15zdnd11an1n64x5 FILLER_97_128 ();
 b15zdnd11an1n64x5 FILLER_97_192 ();
 b15zdnd11an1n64x5 FILLER_97_256 ();
 b15zdnd11an1n64x5 FILLER_97_320 ();
 b15zdnd11an1n64x5 FILLER_97_384 ();
 b15zdnd11an1n32x5 FILLER_97_448 ();
 b15zdnd11an1n16x5 FILLER_97_480 ();
 b15zdnd11an1n08x5 FILLER_97_496 ();
 b15zdnd11an1n04x5 FILLER_97_504 ();
 b15zdnd00an1n01x5 FILLER_97_508 ();
 b15zdnd11an1n64x5 FILLER_97_518 ();
 b15zdnd11an1n64x5 FILLER_97_582 ();
 b15zdnd11an1n64x5 FILLER_97_646 ();
 b15zdnd11an1n64x5 FILLER_97_710 ();
 b15zdnd11an1n64x5 FILLER_97_774 ();
 b15zdnd11an1n64x5 FILLER_97_838 ();
 b15zdnd11an1n64x5 FILLER_97_902 ();
 b15zdnd11an1n64x5 FILLER_97_966 ();
 b15zdnd11an1n64x5 FILLER_97_1030 ();
 b15zdnd11an1n64x5 FILLER_97_1094 ();
 b15zdnd11an1n64x5 FILLER_97_1158 ();
 b15zdnd11an1n64x5 FILLER_97_1222 ();
 b15zdnd11an1n08x5 FILLER_97_1286 ();
 b15zdnd11an1n64x5 FILLER_97_1303 ();
 b15zdnd11an1n64x5 FILLER_97_1367 ();
 b15zdnd11an1n64x5 FILLER_97_1431 ();
 b15zdnd11an1n64x5 FILLER_97_1495 ();
 b15zdnd11an1n64x5 FILLER_97_1559 ();
 b15zdnd11an1n64x5 FILLER_97_1623 ();
 b15zdnd11an1n64x5 FILLER_97_1687 ();
 b15zdnd11an1n64x5 FILLER_97_1751 ();
 b15zdnd11an1n16x5 FILLER_97_1815 ();
 b15zdnd11an1n08x5 FILLER_97_1831 ();
 b15zdnd11an1n04x5 FILLER_97_1839 ();
 b15zdnd00an1n01x5 FILLER_97_1843 ();
 b15zdnd11an1n32x5 FILLER_97_1847 ();
 b15zdnd11an1n08x5 FILLER_97_1879 ();
 b15zdnd11an1n04x5 FILLER_97_1887 ();
 b15zdnd11an1n64x5 FILLER_97_1898 ();
 b15zdnd11an1n16x5 FILLER_97_1962 ();
 b15zdnd11an1n08x5 FILLER_97_1978 ();
 b15zdnd11an1n04x5 FILLER_97_1986 ();
 b15zdnd11an1n64x5 FILLER_97_2042 ();
 b15zdnd11an1n64x5 FILLER_97_2106 ();
 b15zdnd11an1n64x5 FILLER_97_2170 ();
 b15zdnd11an1n32x5 FILLER_97_2234 ();
 b15zdnd11an1n16x5 FILLER_97_2266 ();
 b15zdnd00an1n02x5 FILLER_97_2282 ();
 b15zdnd11an1n64x5 FILLER_98_8 ();
 b15zdnd11an1n64x5 FILLER_98_72 ();
 b15zdnd11an1n64x5 FILLER_98_136 ();
 b15zdnd11an1n64x5 FILLER_98_200 ();
 b15zdnd11an1n64x5 FILLER_98_264 ();
 b15zdnd11an1n64x5 FILLER_98_328 ();
 b15zdnd11an1n64x5 FILLER_98_392 ();
 b15zdnd11an1n64x5 FILLER_98_456 ();
 b15zdnd11an1n64x5 FILLER_98_520 ();
 b15zdnd11an1n64x5 FILLER_98_584 ();
 b15zdnd11an1n64x5 FILLER_98_648 ();
 b15zdnd11an1n04x5 FILLER_98_712 ();
 b15zdnd00an1n02x5 FILLER_98_716 ();
 b15zdnd11an1n64x5 FILLER_98_726 ();
 b15zdnd11an1n32x5 FILLER_98_842 ();
 b15zdnd11an1n16x5 FILLER_98_874 ();
 b15zdnd00an1n02x5 FILLER_98_890 ();
 b15zdnd00an1n01x5 FILLER_98_892 ();
 b15zdnd11an1n64x5 FILLER_98_897 ();
 b15zdnd11an1n64x5 FILLER_98_961 ();
 b15zdnd11an1n64x5 FILLER_98_1025 ();
 b15zdnd11an1n64x5 FILLER_98_1089 ();
 b15zdnd11an1n64x5 FILLER_98_1153 ();
 b15zdnd11an1n64x5 FILLER_98_1217 ();
 b15zdnd11an1n64x5 FILLER_98_1281 ();
 b15zdnd11an1n64x5 FILLER_98_1345 ();
 b15zdnd11an1n32x5 FILLER_98_1409 ();
 b15zdnd11an1n16x5 FILLER_98_1441 ();
 b15zdnd11an1n32x5 FILLER_98_1473 ();
 b15zdnd11an1n16x5 FILLER_98_1505 ();
 b15zdnd11an1n08x5 FILLER_98_1521 ();
 b15zdnd11an1n04x5 FILLER_98_1529 ();
 b15zdnd00an1n01x5 FILLER_98_1533 ();
 b15zdnd11an1n64x5 FILLER_98_1550 ();
 b15zdnd11an1n64x5 FILLER_98_1614 ();
 b15zdnd11an1n32x5 FILLER_98_1678 ();
 b15zdnd00an1n02x5 FILLER_98_1710 ();
 b15zdnd11an1n04x5 FILLER_98_1715 ();
 b15zdnd11an1n08x5 FILLER_98_1722 ();
 b15zdnd00an1n01x5 FILLER_98_1730 ();
 b15zdnd11an1n64x5 FILLER_98_1737 ();
 b15zdnd11an1n16x5 FILLER_98_1801 ();
 b15zdnd11an1n04x5 FILLER_98_1817 ();
 b15zdnd11an1n32x5 FILLER_98_1873 ();
 b15zdnd11an1n04x5 FILLER_98_1905 ();
 b15zdnd00an1n02x5 FILLER_98_1909 ();
 b15zdnd11an1n64x5 FILLER_98_1919 ();
 b15zdnd11an1n16x5 FILLER_98_1983 ();
 b15zdnd11an1n08x5 FILLER_98_1999 ();
 b15zdnd11an1n04x5 FILLER_98_2007 ();
 b15zdnd00an1n02x5 FILLER_98_2011 ();
 b15zdnd11an1n04x5 FILLER_98_2016 ();
 b15zdnd11an1n04x5 FILLER_98_2023 ();
 b15zdnd11an1n64x5 FILLER_98_2030 ();
 b15zdnd11an1n32x5 FILLER_98_2094 ();
 b15zdnd11an1n16x5 FILLER_98_2126 ();
 b15zdnd11an1n08x5 FILLER_98_2142 ();
 b15zdnd11an1n04x5 FILLER_98_2150 ();
 b15zdnd11an1n64x5 FILLER_98_2162 ();
 b15zdnd11an1n32x5 FILLER_98_2226 ();
 b15zdnd11an1n16x5 FILLER_98_2258 ();
 b15zdnd00an1n02x5 FILLER_98_2274 ();
 b15zdnd11an1n64x5 FILLER_99_0 ();
 b15zdnd11an1n64x5 FILLER_99_64 ();
 b15zdnd11an1n64x5 FILLER_99_128 ();
 b15zdnd11an1n32x5 FILLER_99_192 ();
 b15zdnd11an1n16x5 FILLER_99_224 ();
 b15zdnd00an1n02x5 FILLER_99_240 ();
 b15zdnd00an1n01x5 FILLER_99_242 ();
 b15zdnd11an1n64x5 FILLER_99_254 ();
 b15zdnd11an1n64x5 FILLER_99_318 ();
 b15zdnd11an1n64x5 FILLER_99_382 ();
 b15zdnd11an1n64x5 FILLER_99_446 ();
 b15zdnd11an1n64x5 FILLER_99_510 ();
 b15zdnd11an1n32x5 FILLER_99_574 ();
 b15zdnd11an1n16x5 FILLER_99_606 ();
 b15zdnd00an1n02x5 FILLER_99_622 ();
 b15zdnd00an1n01x5 FILLER_99_624 ();
 b15zdnd11an1n64x5 FILLER_99_633 ();
 b15zdnd11an1n64x5 FILLER_99_697 ();
 b15zdnd11an1n16x5 FILLER_99_761 ();
 b15zdnd00an1n01x5 FILLER_99_777 ();
 b15zdnd11an1n04x5 FILLER_99_805 ();
 b15zdnd11an1n04x5 FILLER_99_812 ();
 b15zdnd11an1n04x5 FILLER_99_819 ();
 b15zdnd00an1n02x5 FILLER_99_823 ();
 b15zdnd11an1n16x5 FILLER_99_856 ();
 b15zdnd11an1n04x5 FILLER_99_872 ();
 b15zdnd00an1n02x5 FILLER_99_876 ();
 b15zdnd00an1n01x5 FILLER_99_878 ();
 b15zdnd11an1n64x5 FILLER_99_883 ();
 b15zdnd11an1n16x5 FILLER_99_947 ();
 b15zdnd11an1n08x5 FILLER_99_963 ();
 b15zdnd11an1n04x5 FILLER_99_971 ();
 b15zdnd00an1n01x5 FILLER_99_975 ();
 b15zdnd11an1n64x5 FILLER_99_985 ();
 b15zdnd11an1n64x5 FILLER_99_1049 ();
 b15zdnd11an1n64x5 FILLER_99_1113 ();
 b15zdnd11an1n64x5 FILLER_99_1177 ();
 b15zdnd11an1n64x5 FILLER_99_1241 ();
 b15zdnd11an1n64x5 FILLER_99_1305 ();
 b15zdnd11an1n64x5 FILLER_99_1369 ();
 b15zdnd11an1n16x5 FILLER_99_1433 ();
 b15zdnd11an1n08x5 FILLER_99_1449 ();
 b15zdnd00an1n02x5 FILLER_99_1457 ();
 b15zdnd00an1n01x5 FILLER_99_1459 ();
 b15zdnd11an1n16x5 FILLER_99_1473 ();
 b15zdnd11an1n04x5 FILLER_99_1489 ();
 b15zdnd00an1n02x5 FILLER_99_1493 ();
 b15zdnd00an1n01x5 FILLER_99_1495 ();
 b15zdnd11an1n64x5 FILLER_99_1516 ();
 b15zdnd11an1n64x5 FILLER_99_1580 ();
 b15zdnd11an1n32x5 FILLER_99_1644 ();
 b15zdnd11an1n16x5 FILLER_99_1676 ();
 b15zdnd00an1n02x5 FILLER_99_1692 ();
 b15zdnd11an1n64x5 FILLER_99_1746 ();
 b15zdnd11an1n32x5 FILLER_99_1810 ();
 b15zdnd11an1n08x5 FILLER_99_1842 ();
 b15zdnd11an1n04x5 FILLER_99_1850 ();
 b15zdnd00an1n01x5 FILLER_99_1854 ();
 b15zdnd11an1n64x5 FILLER_99_1858 ();
 b15zdnd11an1n32x5 FILLER_99_1922 ();
 b15zdnd11an1n16x5 FILLER_99_1954 ();
 b15zdnd11an1n16x5 FILLER_99_1987 ();
 b15zdnd11an1n08x5 FILLER_99_2003 ();
 b15zdnd00an1n02x5 FILLER_99_2011 ();
 b15zdnd11an1n64x5 FILLER_99_2016 ();
 b15zdnd11an1n08x5 FILLER_99_2080 ();
 b15zdnd11an1n04x5 FILLER_99_2094 ();
 b15zdnd00an1n02x5 FILLER_99_2098 ();
 b15zdnd00an1n01x5 FILLER_99_2100 ();
 b15zdnd11an1n64x5 FILLER_99_2107 ();
 b15zdnd11an1n64x5 FILLER_99_2171 ();
 b15zdnd11an1n32x5 FILLER_99_2235 ();
 b15zdnd11an1n16x5 FILLER_99_2267 ();
 b15zdnd00an1n01x5 FILLER_99_2283 ();
 b15zdnd11an1n64x5 FILLER_100_8 ();
 b15zdnd11an1n64x5 FILLER_100_72 ();
 b15zdnd11an1n64x5 FILLER_100_136 ();
 b15zdnd11an1n64x5 FILLER_100_200 ();
 b15zdnd11an1n64x5 FILLER_100_264 ();
 b15zdnd11an1n64x5 FILLER_100_328 ();
 b15zdnd11an1n64x5 FILLER_100_392 ();
 b15zdnd11an1n64x5 FILLER_100_456 ();
 b15zdnd11an1n64x5 FILLER_100_520 ();
 b15zdnd11an1n64x5 FILLER_100_584 ();
 b15zdnd11an1n64x5 FILLER_100_648 ();
 b15zdnd11an1n04x5 FILLER_100_712 ();
 b15zdnd00an1n02x5 FILLER_100_716 ();
 b15zdnd11an1n32x5 FILLER_100_726 ();
 b15zdnd11an1n16x5 FILLER_100_758 ();
 b15zdnd00an1n02x5 FILLER_100_774 ();
 b15zdnd11an1n32x5 FILLER_100_779 ();
 b15zdnd00an1n02x5 FILLER_100_811 ();
 b15zdnd11an1n64x5 FILLER_100_816 ();
 b15zdnd11an1n32x5 FILLER_100_880 ();
 b15zdnd11an1n16x5 FILLER_100_912 ();
 b15zdnd11an1n08x5 FILLER_100_928 ();
 b15zdnd00an1n01x5 FILLER_100_936 ();
 b15zdnd11an1n64x5 FILLER_100_941 ();
 b15zdnd11an1n32x5 FILLER_100_1005 ();
 b15zdnd11an1n08x5 FILLER_100_1037 ();
 b15zdnd11an1n04x5 FILLER_100_1045 ();
 b15zdnd00an1n02x5 FILLER_100_1049 ();
 b15zdnd11an1n04x5 FILLER_100_1059 ();
 b15zdnd11an1n64x5 FILLER_100_1066 ();
 b15zdnd11an1n64x5 FILLER_100_1130 ();
 b15zdnd11an1n64x5 FILLER_100_1194 ();
 b15zdnd11an1n64x5 FILLER_100_1258 ();
 b15zdnd11an1n64x5 FILLER_100_1322 ();
 b15zdnd11an1n16x5 FILLER_100_1386 ();
 b15zdnd11an1n08x5 FILLER_100_1402 ();
 b15zdnd11an1n04x5 FILLER_100_1410 ();
 b15zdnd00an1n02x5 FILLER_100_1414 ();
 b15zdnd11an1n04x5 FILLER_100_1452 ();
 b15zdnd11an1n08x5 FILLER_100_1459 ();
 b15zdnd00an1n02x5 FILLER_100_1467 ();
 b15zdnd11an1n04x5 FILLER_100_1479 ();
 b15zdnd11an1n64x5 FILLER_100_1507 ();
 b15zdnd11an1n64x5 FILLER_100_1571 ();
 b15zdnd11an1n64x5 FILLER_100_1635 ();
 b15zdnd11an1n16x5 FILLER_100_1699 ();
 b15zdnd11an1n04x5 FILLER_100_1715 ();
 b15zdnd11an1n64x5 FILLER_100_1722 ();
 b15zdnd11an1n64x5 FILLER_100_1786 ();
 b15zdnd11an1n64x5 FILLER_100_1850 ();
 b15zdnd11an1n64x5 FILLER_100_1914 ();
 b15zdnd11an1n64x5 FILLER_100_1978 ();
 b15zdnd11an1n32x5 FILLER_100_2042 ();
 b15zdnd11an1n16x5 FILLER_100_2074 ();
 b15zdnd11an1n08x5 FILLER_100_2090 ();
 b15zdnd00an1n02x5 FILLER_100_2098 ();
 b15zdnd11an1n16x5 FILLER_100_2124 ();
 b15zdnd11an1n08x5 FILLER_100_2140 ();
 b15zdnd11an1n04x5 FILLER_100_2148 ();
 b15zdnd00an1n02x5 FILLER_100_2152 ();
 b15zdnd11an1n64x5 FILLER_100_2162 ();
 b15zdnd11an1n32x5 FILLER_100_2226 ();
 b15zdnd11an1n16x5 FILLER_100_2258 ();
 b15zdnd00an1n02x5 FILLER_100_2274 ();
 b15zdnd11an1n64x5 FILLER_101_0 ();
 b15zdnd11an1n64x5 FILLER_101_64 ();
 b15zdnd11an1n64x5 FILLER_101_128 ();
 b15zdnd11an1n64x5 FILLER_101_192 ();
 b15zdnd11an1n64x5 FILLER_101_256 ();
 b15zdnd11an1n64x5 FILLER_101_320 ();
 b15zdnd11an1n64x5 FILLER_101_384 ();
 b15zdnd11an1n32x5 FILLER_101_448 ();
 b15zdnd11an1n16x5 FILLER_101_480 ();
 b15zdnd11an1n04x5 FILLER_101_496 ();
 b15zdnd00an1n01x5 FILLER_101_500 ();
 b15zdnd11an1n32x5 FILLER_101_519 ();
 b15zdnd11an1n64x5 FILLER_101_554 ();
 b15zdnd11an1n32x5 FILLER_101_618 ();
 b15zdnd11an1n16x5 FILLER_101_650 ();
 b15zdnd00an1n02x5 FILLER_101_666 ();
 b15zdnd11an1n64x5 FILLER_101_689 ();
 b15zdnd11an1n32x5 FILLER_101_753 ();
 b15zdnd11an1n04x5 FILLER_101_785 ();
 b15zdnd11an1n64x5 FILLER_101_796 ();
 b15zdnd11an1n32x5 FILLER_101_860 ();
 b15zdnd11an1n64x5 FILLER_101_903 ();
 b15zdnd11an1n64x5 FILLER_101_967 ();
 b15zdnd11an1n16x5 FILLER_101_1031 ();
 b15zdnd11an1n08x5 FILLER_101_1047 ();
 b15zdnd11an1n04x5 FILLER_101_1055 ();
 b15zdnd11an1n64x5 FILLER_101_1062 ();
 b15zdnd11an1n08x5 FILLER_101_1126 ();
 b15zdnd11an1n04x5 FILLER_101_1134 ();
 b15zdnd11an1n64x5 FILLER_101_1147 ();
 b15zdnd11an1n64x5 FILLER_101_1211 ();
 b15zdnd11an1n64x5 FILLER_101_1275 ();
 b15zdnd11an1n64x5 FILLER_101_1339 ();
 b15zdnd11an1n64x5 FILLER_101_1403 ();
 b15zdnd11an1n04x5 FILLER_101_1467 ();
 b15zdnd00an1n02x5 FILLER_101_1471 ();
 b15zdnd11an1n64x5 FILLER_101_1476 ();
 b15zdnd11an1n64x5 FILLER_101_1540 ();
 b15zdnd11an1n64x5 FILLER_101_1604 ();
 b15zdnd11an1n64x5 FILLER_101_1668 ();
 b15zdnd11an1n64x5 FILLER_101_1732 ();
 b15zdnd11an1n64x5 FILLER_101_1796 ();
 b15zdnd11an1n64x5 FILLER_101_1860 ();
 b15zdnd11an1n64x5 FILLER_101_1924 ();
 b15zdnd11an1n64x5 FILLER_101_1988 ();
 b15zdnd11an1n64x5 FILLER_101_2052 ();
 b15zdnd11an1n64x5 FILLER_101_2116 ();
 b15zdnd11an1n16x5 FILLER_101_2180 ();
 b15zdnd11an1n08x5 FILLER_101_2196 ();
 b15zdnd11an1n04x5 FILLER_101_2204 ();
 b15zdnd00an1n01x5 FILLER_101_2208 ();
 b15zdnd11an1n64x5 FILLER_101_2217 ();
 b15zdnd00an1n02x5 FILLER_101_2281 ();
 b15zdnd00an1n01x5 FILLER_101_2283 ();
 b15zdnd11an1n64x5 FILLER_102_8 ();
 b15zdnd11an1n64x5 FILLER_102_72 ();
 b15zdnd11an1n64x5 FILLER_102_136 ();
 b15zdnd11an1n64x5 FILLER_102_200 ();
 b15zdnd11an1n64x5 FILLER_102_264 ();
 b15zdnd11an1n64x5 FILLER_102_328 ();
 b15zdnd11an1n64x5 FILLER_102_392 ();
 b15zdnd11an1n64x5 FILLER_102_456 ();
 b15zdnd11an1n64x5 FILLER_102_520 ();
 b15zdnd11an1n16x5 FILLER_102_584 ();
 b15zdnd11an1n08x5 FILLER_102_600 ();
 b15zdnd00an1n02x5 FILLER_102_608 ();
 b15zdnd11an1n64x5 FILLER_102_614 ();
 b15zdnd11an1n32x5 FILLER_102_678 ();
 b15zdnd11an1n08x5 FILLER_102_710 ();
 b15zdnd11an1n32x5 FILLER_102_726 ();
 b15zdnd11an1n08x5 FILLER_102_758 ();
 b15zdnd11an1n64x5 FILLER_102_775 ();
 b15zdnd11an1n64x5 FILLER_102_839 ();
 b15zdnd11an1n64x5 FILLER_102_903 ();
 b15zdnd11an1n32x5 FILLER_102_967 ();
 b15zdnd11an1n16x5 FILLER_102_999 ();
 b15zdnd00an1n01x5 FILLER_102_1015 ();
 b15zdnd11an1n08x5 FILLER_102_1025 ();
 b15zdnd11an1n04x5 FILLER_102_1033 ();
 b15zdnd00an1n02x5 FILLER_102_1037 ();
 b15zdnd11an1n64x5 FILLER_102_1083 ();
 b15zdnd11an1n64x5 FILLER_102_1147 ();
 b15zdnd11an1n64x5 FILLER_102_1211 ();
 b15zdnd11an1n64x5 FILLER_102_1275 ();
 b15zdnd11an1n64x5 FILLER_102_1339 ();
 b15zdnd11an1n64x5 FILLER_102_1403 ();
 b15zdnd11an1n64x5 FILLER_102_1467 ();
 b15zdnd11an1n64x5 FILLER_102_1531 ();
 b15zdnd11an1n64x5 FILLER_102_1595 ();
 b15zdnd11an1n64x5 FILLER_102_1659 ();
 b15zdnd11an1n64x5 FILLER_102_1723 ();
 b15zdnd11an1n64x5 FILLER_102_1787 ();
 b15zdnd11an1n64x5 FILLER_102_1851 ();
 b15zdnd11an1n64x5 FILLER_102_1915 ();
 b15zdnd11an1n64x5 FILLER_102_1979 ();
 b15zdnd11an1n64x5 FILLER_102_2043 ();
 b15zdnd11an1n32x5 FILLER_102_2107 ();
 b15zdnd11an1n08x5 FILLER_102_2139 ();
 b15zdnd11an1n04x5 FILLER_102_2147 ();
 b15zdnd00an1n02x5 FILLER_102_2151 ();
 b15zdnd00an1n01x5 FILLER_102_2153 ();
 b15zdnd11an1n64x5 FILLER_102_2162 ();
 b15zdnd11an1n32x5 FILLER_102_2226 ();
 b15zdnd11an1n16x5 FILLER_102_2258 ();
 b15zdnd00an1n02x5 FILLER_102_2274 ();
 b15zdnd11an1n64x5 FILLER_103_0 ();
 b15zdnd11an1n64x5 FILLER_103_64 ();
 b15zdnd11an1n64x5 FILLER_103_128 ();
 b15zdnd11an1n64x5 FILLER_103_192 ();
 b15zdnd11an1n64x5 FILLER_103_256 ();
 b15zdnd11an1n64x5 FILLER_103_320 ();
 b15zdnd11an1n64x5 FILLER_103_384 ();
 b15zdnd11an1n64x5 FILLER_103_448 ();
 b15zdnd11an1n64x5 FILLER_103_512 ();
 b15zdnd11an1n32x5 FILLER_103_576 ();
 b15zdnd11an1n16x5 FILLER_103_608 ();
 b15zdnd11an1n08x5 FILLER_103_624 ();
 b15zdnd00an1n01x5 FILLER_103_632 ();
 b15zdnd11an1n16x5 FILLER_103_659 ();
 b15zdnd11an1n04x5 FILLER_103_675 ();
 b15zdnd11an1n64x5 FILLER_103_682 ();
 b15zdnd11an1n64x5 FILLER_103_746 ();
 b15zdnd11an1n64x5 FILLER_103_810 ();
 b15zdnd11an1n64x5 FILLER_103_874 ();
 b15zdnd11an1n64x5 FILLER_103_938 ();
 b15zdnd11an1n32x5 FILLER_103_1002 ();
 b15zdnd11an1n16x5 FILLER_103_1034 ();
 b15zdnd11an1n08x5 FILLER_103_1050 ();
 b15zdnd00an1n01x5 FILLER_103_1058 ();
 b15zdnd11an1n64x5 FILLER_103_1062 ();
 b15zdnd11an1n64x5 FILLER_103_1126 ();
 b15zdnd11an1n64x5 FILLER_103_1190 ();
 b15zdnd11an1n16x5 FILLER_103_1254 ();
 b15zdnd11an1n04x5 FILLER_103_1270 ();
 b15zdnd00an1n02x5 FILLER_103_1274 ();
 b15zdnd00an1n01x5 FILLER_103_1276 ();
 b15zdnd11an1n04x5 FILLER_103_1280 ();
 b15zdnd11an1n04x5 FILLER_103_1287 ();
 b15zdnd11an1n16x5 FILLER_103_1294 ();
 b15zdnd00an1n01x5 FILLER_103_1310 ();
 b15zdnd11an1n64x5 FILLER_103_1363 ();
 b15zdnd11an1n04x5 FILLER_103_1427 ();
 b15zdnd11an1n64x5 FILLER_103_1435 ();
 b15zdnd11an1n64x5 FILLER_103_1499 ();
 b15zdnd11an1n64x5 FILLER_103_1563 ();
 b15zdnd11an1n64x5 FILLER_103_1627 ();
 b15zdnd11an1n32x5 FILLER_103_1691 ();
 b15zdnd00an1n01x5 FILLER_103_1723 ();
 b15zdnd11an1n64x5 FILLER_103_1766 ();
 b15zdnd11an1n16x5 FILLER_103_1830 ();
 b15zdnd00an1n02x5 FILLER_103_1846 ();
 b15zdnd11an1n64x5 FILLER_103_1859 ();
 b15zdnd11an1n64x5 FILLER_103_1923 ();
 b15zdnd11an1n64x5 FILLER_103_1987 ();
 b15zdnd11an1n32x5 FILLER_103_2051 ();
 b15zdnd11an1n64x5 FILLER_103_2093 ();
 b15zdnd11an1n64x5 FILLER_103_2157 ();
 b15zdnd11an1n32x5 FILLER_103_2221 ();
 b15zdnd11an1n16x5 FILLER_103_2253 ();
 b15zdnd11an1n08x5 FILLER_103_2269 ();
 b15zdnd11an1n04x5 FILLER_103_2277 ();
 b15zdnd00an1n02x5 FILLER_103_2281 ();
 b15zdnd00an1n01x5 FILLER_103_2283 ();
 b15zdnd11an1n64x5 FILLER_104_8 ();
 b15zdnd11an1n64x5 FILLER_104_72 ();
 b15zdnd11an1n64x5 FILLER_104_136 ();
 b15zdnd11an1n64x5 FILLER_104_200 ();
 b15zdnd11an1n64x5 FILLER_104_264 ();
 b15zdnd11an1n64x5 FILLER_104_328 ();
 b15zdnd11an1n64x5 FILLER_104_392 ();
 b15zdnd11an1n64x5 FILLER_104_456 ();
 b15zdnd11an1n64x5 FILLER_104_520 ();
 b15zdnd11an1n64x5 FILLER_104_584 ();
 b15zdnd11an1n08x5 FILLER_104_648 ();
 b15zdnd11an1n04x5 FILLER_104_656 ();
 b15zdnd00an1n01x5 FILLER_104_660 ();
 b15zdnd11an1n04x5 FILLER_104_689 ();
 b15zdnd11an1n16x5 FILLER_104_696 ();
 b15zdnd11an1n04x5 FILLER_104_712 ();
 b15zdnd00an1n02x5 FILLER_104_716 ();
 b15zdnd11an1n64x5 FILLER_104_726 ();
 b15zdnd11an1n64x5 FILLER_104_790 ();
 b15zdnd11an1n64x5 FILLER_104_854 ();
 b15zdnd11an1n64x5 FILLER_104_918 ();
 b15zdnd11an1n32x5 FILLER_104_982 ();
 b15zdnd11an1n08x5 FILLER_104_1014 ();
 b15zdnd11an1n04x5 FILLER_104_1022 ();
 b15zdnd00an1n02x5 FILLER_104_1026 ();
 b15zdnd11an1n64x5 FILLER_104_1031 ();
 b15zdnd11an1n64x5 FILLER_104_1095 ();
 b15zdnd11an1n64x5 FILLER_104_1159 ();
 b15zdnd11an1n32x5 FILLER_104_1223 ();
 b15zdnd11an1n08x5 FILLER_104_1255 ();
 b15zdnd11an1n04x5 FILLER_104_1263 ();
 b15zdnd00an1n02x5 FILLER_104_1267 ();
 b15zdnd11an1n04x5 FILLER_104_1321 ();
 b15zdnd11an1n04x5 FILLER_104_1328 ();
 b15zdnd00an1n02x5 FILLER_104_1332 ();
 b15zdnd11an1n04x5 FILLER_104_1337 ();
 b15zdnd11an1n64x5 FILLER_104_1344 ();
 b15zdnd11an1n64x5 FILLER_104_1408 ();
 b15zdnd11an1n64x5 FILLER_104_1472 ();
 b15zdnd11an1n64x5 FILLER_104_1536 ();
 b15zdnd11an1n64x5 FILLER_104_1600 ();
 b15zdnd11an1n64x5 FILLER_104_1664 ();
 b15zdnd00an1n02x5 FILLER_104_1728 ();
 b15zdnd00an1n01x5 FILLER_104_1730 ();
 b15zdnd11an1n08x5 FILLER_104_1737 ();
 b15zdnd00an1n01x5 FILLER_104_1745 ();
 b15zdnd11an1n64x5 FILLER_104_1777 ();
 b15zdnd11an1n64x5 FILLER_104_1841 ();
 b15zdnd11an1n64x5 FILLER_104_1905 ();
 b15zdnd11an1n64x5 FILLER_104_1969 ();
 b15zdnd11an1n64x5 FILLER_104_2033 ();
 b15zdnd11an1n32x5 FILLER_104_2097 ();
 b15zdnd11an1n16x5 FILLER_104_2129 ();
 b15zdnd11an1n08x5 FILLER_104_2145 ();
 b15zdnd00an1n01x5 FILLER_104_2153 ();
 b15zdnd11an1n64x5 FILLER_104_2162 ();
 b15zdnd11an1n32x5 FILLER_104_2226 ();
 b15zdnd11an1n16x5 FILLER_104_2258 ();
 b15zdnd00an1n02x5 FILLER_104_2274 ();
 b15zdnd11an1n64x5 FILLER_105_0 ();
 b15zdnd11an1n64x5 FILLER_105_64 ();
 b15zdnd11an1n64x5 FILLER_105_128 ();
 b15zdnd11an1n64x5 FILLER_105_192 ();
 b15zdnd11an1n64x5 FILLER_105_256 ();
 b15zdnd11an1n64x5 FILLER_105_320 ();
 b15zdnd11an1n32x5 FILLER_105_384 ();
 b15zdnd11an1n08x5 FILLER_105_416 ();
 b15zdnd11an1n16x5 FILLER_105_435 ();
 b15zdnd11an1n08x5 FILLER_105_454 ();
 b15zdnd00an1n02x5 FILLER_105_462 ();
 b15zdnd11an1n64x5 FILLER_105_467 ();
 b15zdnd11an1n16x5 FILLER_105_531 ();
 b15zdnd00an1n02x5 FILLER_105_547 ();
 b15zdnd00an1n01x5 FILLER_105_549 ();
 b15zdnd11an1n64x5 FILLER_105_571 ();
 b15zdnd11an1n32x5 FILLER_105_635 ();
 b15zdnd11an1n04x5 FILLER_105_667 ();
 b15zdnd11an1n64x5 FILLER_105_691 ();
 b15zdnd11an1n64x5 FILLER_105_755 ();
 b15zdnd11an1n64x5 FILLER_105_819 ();
 b15zdnd11an1n64x5 FILLER_105_883 ();
 b15zdnd11an1n64x5 FILLER_105_947 ();
 b15zdnd11an1n08x5 FILLER_105_1011 ();
 b15zdnd11an1n04x5 FILLER_105_1019 ();
 b15zdnd00an1n02x5 FILLER_105_1023 ();
 b15zdnd11an1n64x5 FILLER_105_1039 ();
 b15zdnd11an1n16x5 FILLER_105_1103 ();
 b15zdnd00an1n01x5 FILLER_105_1119 ();
 b15zdnd11an1n64x5 FILLER_105_1130 ();
 b15zdnd11an1n64x5 FILLER_105_1194 ();
 b15zdnd11an1n04x5 FILLER_105_1310 ();
 b15zdnd11an1n04x5 FILLER_105_1317 ();
 b15zdnd11an1n04x5 FILLER_105_1324 ();
 b15zdnd11an1n04x5 FILLER_105_1331 ();
 b15zdnd11an1n64x5 FILLER_105_1338 ();
 b15zdnd11an1n32x5 FILLER_105_1402 ();
 b15zdnd11an1n04x5 FILLER_105_1434 ();
 b15zdnd11an1n64x5 FILLER_105_1449 ();
 b15zdnd11an1n64x5 FILLER_105_1513 ();
 b15zdnd11an1n08x5 FILLER_105_1577 ();
 b15zdnd11an1n04x5 FILLER_105_1585 ();
 b15zdnd00an1n02x5 FILLER_105_1589 ();
 b15zdnd11an1n04x5 FILLER_105_1594 ();
 b15zdnd11an1n64x5 FILLER_105_1601 ();
 b15zdnd11an1n64x5 FILLER_105_1665 ();
 b15zdnd00an1n02x5 FILLER_105_1729 ();
 b15zdnd00an1n01x5 FILLER_105_1731 ();
 b15zdnd11an1n64x5 FILLER_105_1746 ();
 b15zdnd11an1n64x5 FILLER_105_1810 ();
 b15zdnd11an1n64x5 FILLER_105_1874 ();
 b15zdnd11an1n64x5 FILLER_105_1938 ();
 b15zdnd11an1n64x5 FILLER_105_2002 ();
 b15zdnd11an1n64x5 FILLER_105_2066 ();
 b15zdnd11an1n64x5 FILLER_105_2130 ();
 b15zdnd11an1n64x5 FILLER_105_2194 ();
 b15zdnd11an1n16x5 FILLER_105_2258 ();
 b15zdnd11an1n08x5 FILLER_105_2274 ();
 b15zdnd00an1n02x5 FILLER_105_2282 ();
 b15zdnd11an1n64x5 FILLER_106_8 ();
 b15zdnd11an1n64x5 FILLER_106_72 ();
 b15zdnd11an1n32x5 FILLER_106_136 ();
 b15zdnd11an1n16x5 FILLER_106_168 ();
 b15zdnd11an1n04x5 FILLER_106_184 ();
 b15zdnd00an1n01x5 FILLER_106_188 ();
 b15zdnd11an1n64x5 FILLER_106_220 ();
 b15zdnd11an1n32x5 FILLER_106_284 ();
 b15zdnd11an1n16x5 FILLER_106_316 ();
 b15zdnd11an1n04x5 FILLER_106_335 ();
 b15zdnd11an1n04x5 FILLER_106_344 ();
 b15zdnd11an1n32x5 FILLER_106_390 ();
 b15zdnd11an1n08x5 FILLER_106_422 ();
 b15zdnd00an1n02x5 FILLER_106_430 ();
 b15zdnd00an1n01x5 FILLER_106_432 ();
 b15zdnd11an1n04x5 FILLER_106_475 ();
 b15zdnd11an1n64x5 FILLER_106_482 ();
 b15zdnd11an1n16x5 FILLER_106_546 ();
 b15zdnd11an1n04x5 FILLER_106_562 ();
 b15zdnd00an1n02x5 FILLER_106_566 ();
 b15zdnd00an1n01x5 FILLER_106_568 ();
 b15zdnd11an1n64x5 FILLER_106_573 ();
 b15zdnd11an1n64x5 FILLER_106_637 ();
 b15zdnd11an1n16x5 FILLER_106_701 ();
 b15zdnd00an1n01x5 FILLER_106_717 ();
 b15zdnd11an1n32x5 FILLER_106_726 ();
 b15zdnd11an1n16x5 FILLER_106_758 ();
 b15zdnd11an1n08x5 FILLER_106_774 ();
 b15zdnd11an1n04x5 FILLER_106_782 ();
 b15zdnd11an1n64x5 FILLER_106_795 ();
 b15zdnd11an1n64x5 FILLER_106_859 ();
 b15zdnd11an1n32x5 FILLER_106_923 ();
 b15zdnd11an1n16x5 FILLER_106_955 ();
 b15zdnd11an1n08x5 FILLER_106_971 ();
 b15zdnd11an1n04x5 FILLER_106_979 ();
 b15zdnd11an1n64x5 FILLER_106_997 ();
 b15zdnd11an1n16x5 FILLER_106_1061 ();
 b15zdnd11an1n04x5 FILLER_106_1077 ();
 b15zdnd11an1n64x5 FILLER_106_1087 ();
 b15zdnd11an1n64x5 FILLER_106_1151 ();
 b15zdnd11an1n32x5 FILLER_106_1215 ();
 b15zdnd11an1n16x5 FILLER_106_1247 ();
 b15zdnd11an1n08x5 FILLER_106_1263 ();
 b15zdnd11an1n04x5 FILLER_106_1271 ();
 b15zdnd00an1n01x5 FILLER_106_1275 ();
 b15zdnd11an1n04x5 FILLER_106_1279 ();
 b15zdnd11an1n64x5 FILLER_106_1335 ();
 b15zdnd11an1n64x5 FILLER_106_1399 ();
 b15zdnd11an1n64x5 FILLER_106_1463 ();
 b15zdnd11an1n32x5 FILLER_106_1527 ();
 b15zdnd11an1n16x5 FILLER_106_1559 ();
 b15zdnd11an1n64x5 FILLER_106_1617 ();
 b15zdnd11an1n64x5 FILLER_106_1681 ();
 b15zdnd11an1n64x5 FILLER_106_1745 ();
 b15zdnd11an1n64x5 FILLER_106_1809 ();
 b15zdnd11an1n64x5 FILLER_106_1873 ();
 b15zdnd11an1n64x5 FILLER_106_1937 ();
 b15zdnd11an1n64x5 FILLER_106_2001 ();
 b15zdnd11an1n64x5 FILLER_106_2065 ();
 b15zdnd11an1n16x5 FILLER_106_2129 ();
 b15zdnd11an1n08x5 FILLER_106_2145 ();
 b15zdnd00an1n01x5 FILLER_106_2153 ();
 b15zdnd11an1n64x5 FILLER_106_2162 ();
 b15zdnd11an1n32x5 FILLER_106_2226 ();
 b15zdnd11an1n16x5 FILLER_106_2258 ();
 b15zdnd00an1n02x5 FILLER_106_2274 ();
 b15zdnd11an1n08x5 FILLER_107_0 ();
 b15zdnd11an1n04x5 FILLER_107_8 ();
 b15zdnd00an1n02x5 FILLER_107_12 ();
 b15zdnd11an1n64x5 FILLER_107_18 ();
 b15zdnd11an1n64x5 FILLER_107_82 ();
 b15zdnd11an1n64x5 FILLER_107_146 ();
 b15zdnd11an1n64x5 FILLER_107_210 ();
 b15zdnd11an1n16x5 FILLER_107_274 ();
 b15zdnd11an1n08x5 FILLER_107_290 ();
 b15zdnd11an1n04x5 FILLER_107_298 ();
 b15zdnd00an1n01x5 FILLER_107_302 ();
 b15zdnd11an1n04x5 FILLER_107_355 ();
 b15zdnd11an1n04x5 FILLER_107_365 ();
 b15zdnd00an1n02x5 FILLER_107_369 ();
 b15zdnd00an1n01x5 FILLER_107_371 ();
 b15zdnd11an1n04x5 FILLER_107_379 ();
 b15zdnd00an1n02x5 FILLER_107_383 ();
 b15zdnd00an1n01x5 FILLER_107_385 ();
 b15zdnd11an1n16x5 FILLER_107_396 ();
 b15zdnd11an1n08x5 FILLER_107_417 ();
 b15zdnd11an1n04x5 FILLER_107_425 ();
 b15zdnd00an1n01x5 FILLER_107_429 ();
 b15zdnd11an1n64x5 FILLER_107_482 ();
 b15zdnd11an1n64x5 FILLER_107_546 ();
 b15zdnd11an1n64x5 FILLER_107_610 ();
 b15zdnd11an1n64x5 FILLER_107_674 ();
 b15zdnd11an1n16x5 FILLER_107_738 ();
 b15zdnd11an1n08x5 FILLER_107_754 ();
 b15zdnd11an1n04x5 FILLER_107_762 ();
 b15zdnd11an1n64x5 FILLER_107_775 ();
 b15zdnd11an1n64x5 FILLER_107_839 ();
 b15zdnd11an1n08x5 FILLER_107_903 ();
 b15zdnd11an1n64x5 FILLER_107_935 ();
 b15zdnd11an1n08x5 FILLER_107_999 ();
 b15zdnd11an1n04x5 FILLER_107_1007 ();
 b15zdnd00an1n01x5 FILLER_107_1011 ();
 b15zdnd11an1n04x5 FILLER_107_1032 ();
 b15zdnd11an1n04x5 FILLER_107_1050 ();
 b15zdnd00an1n02x5 FILLER_107_1054 ();
 b15zdnd00an1n01x5 FILLER_107_1056 ();
 b15zdnd11an1n64x5 FILLER_107_1099 ();
 b15zdnd11an1n04x5 FILLER_107_1163 ();
 b15zdnd00an1n02x5 FILLER_107_1167 ();
 b15zdnd00an1n01x5 FILLER_107_1169 ();
 b15zdnd11an1n04x5 FILLER_107_1186 ();
 b15zdnd11an1n64x5 FILLER_107_1211 ();
 b15zdnd11an1n32x5 FILLER_107_1275 ();
 b15zdnd11an1n64x5 FILLER_107_1310 ();
 b15zdnd11an1n64x5 FILLER_107_1374 ();
 b15zdnd11an1n64x5 FILLER_107_1438 ();
 b15zdnd11an1n64x5 FILLER_107_1502 ();
 b15zdnd11an1n04x5 FILLER_107_1566 ();
 b15zdnd00an1n02x5 FILLER_107_1570 ();
 b15zdnd00an1n01x5 FILLER_107_1572 ();
 b15zdnd11an1n64x5 FILLER_107_1625 ();
 b15zdnd11an1n08x5 FILLER_107_1689 ();
 b15zdnd11an1n04x5 FILLER_107_1697 ();
 b15zdnd00an1n02x5 FILLER_107_1701 ();
 b15zdnd00an1n01x5 FILLER_107_1703 ();
 b15zdnd11an1n16x5 FILLER_107_1725 ();
 b15zdnd11an1n08x5 FILLER_107_1741 ();
 b15zdnd00an1n01x5 FILLER_107_1749 ();
 b15zdnd11an1n64x5 FILLER_107_1756 ();
 b15zdnd11an1n64x5 FILLER_107_1820 ();
 b15zdnd11an1n64x5 FILLER_107_1884 ();
 b15zdnd11an1n64x5 FILLER_107_1948 ();
 b15zdnd11an1n64x5 FILLER_107_2012 ();
 b15zdnd11an1n64x5 FILLER_107_2076 ();
 b15zdnd11an1n64x5 FILLER_107_2140 ();
 b15zdnd11an1n64x5 FILLER_107_2204 ();
 b15zdnd11an1n16x5 FILLER_107_2268 ();
 b15zdnd11an1n32x5 FILLER_108_8 ();
 b15zdnd11an1n16x5 FILLER_108_40 ();
 b15zdnd11an1n08x5 FILLER_108_56 ();
 b15zdnd11an1n04x5 FILLER_108_64 ();
 b15zdnd00an1n01x5 FILLER_108_68 ();
 b15zdnd11an1n64x5 FILLER_108_73 ();
 b15zdnd11an1n32x5 FILLER_108_137 ();
 b15zdnd11an1n16x5 FILLER_108_169 ();
 b15zdnd11an1n08x5 FILLER_108_185 ();
 b15zdnd11an1n04x5 FILLER_108_193 ();
 b15zdnd00an1n02x5 FILLER_108_197 ();
 b15zdnd11an1n64x5 FILLER_108_202 ();
 b15zdnd11an1n32x5 FILLER_108_266 ();
 b15zdnd11an1n08x5 FILLER_108_298 ();
 b15zdnd11an1n04x5 FILLER_108_306 ();
 b15zdnd00an1n01x5 FILLER_108_310 ();
 b15zdnd11an1n04x5 FILLER_108_314 ();
 b15zdnd11an1n04x5 FILLER_108_321 ();
 b15zdnd11an1n04x5 FILLER_108_367 ();
 b15zdnd11an1n08x5 FILLER_108_413 ();
 b15zdnd00an1n02x5 FILLER_108_421 ();
 b15zdnd00an1n01x5 FILLER_108_423 ();
 b15zdnd11an1n64x5 FILLER_108_466 ();
 b15zdnd11an1n64x5 FILLER_108_530 ();
 b15zdnd11an1n64x5 FILLER_108_594 ();
 b15zdnd11an1n32x5 FILLER_108_658 ();
 b15zdnd11an1n16x5 FILLER_108_690 ();
 b15zdnd11an1n08x5 FILLER_108_706 ();
 b15zdnd11an1n04x5 FILLER_108_714 ();
 b15zdnd11an1n64x5 FILLER_108_726 ();
 b15zdnd11an1n64x5 FILLER_108_790 ();
 b15zdnd11an1n64x5 FILLER_108_854 ();
 b15zdnd11an1n64x5 FILLER_108_918 ();
 b15zdnd11an1n32x5 FILLER_108_982 ();
 b15zdnd11an1n16x5 FILLER_108_1014 ();
 b15zdnd00an1n01x5 FILLER_108_1030 ();
 b15zdnd11an1n04x5 FILLER_108_1034 ();
 b15zdnd11an1n08x5 FILLER_108_1080 ();
 b15zdnd11an1n04x5 FILLER_108_1088 ();
 b15zdnd00an1n01x5 FILLER_108_1092 ();
 b15zdnd11an1n64x5 FILLER_108_1100 ();
 b15zdnd11an1n16x5 FILLER_108_1164 ();
 b15zdnd11an1n04x5 FILLER_108_1180 ();
 b15zdnd00an1n02x5 FILLER_108_1184 ();
 b15zdnd00an1n01x5 FILLER_108_1186 ();
 b15zdnd11an1n64x5 FILLER_108_1201 ();
 b15zdnd00an1n02x5 FILLER_108_1265 ();
 b15zdnd11an1n64x5 FILLER_108_1293 ();
 b15zdnd11an1n32x5 FILLER_108_1357 ();
 b15zdnd11an1n16x5 FILLER_108_1389 ();
 b15zdnd11an1n08x5 FILLER_108_1405 ();
 b15zdnd11an1n04x5 FILLER_108_1413 ();
 b15zdnd11an1n32x5 FILLER_108_1425 ();
 b15zdnd11an1n08x5 FILLER_108_1457 ();
 b15zdnd00an1n02x5 FILLER_108_1465 ();
 b15zdnd11an1n32x5 FILLER_108_1489 ();
 b15zdnd11an1n08x5 FILLER_108_1521 ();
 b15zdnd00an1n02x5 FILLER_108_1529 ();
 b15zdnd11an1n16x5 FILLER_108_1542 ();
 b15zdnd11an1n08x5 FILLER_108_1558 ();
 b15zdnd11an1n04x5 FILLER_108_1566 ();
 b15zdnd00an1n02x5 FILLER_108_1570 ();
 b15zdnd11an1n04x5 FILLER_108_1579 ();
 b15zdnd11an1n64x5 FILLER_108_1625 ();
 b15zdnd11an1n64x5 FILLER_108_1689 ();
 b15zdnd11an1n64x5 FILLER_108_1753 ();
 b15zdnd11an1n64x5 FILLER_108_1817 ();
 b15zdnd11an1n64x5 FILLER_108_1881 ();
 b15zdnd11an1n64x5 FILLER_108_1945 ();
 b15zdnd11an1n64x5 FILLER_108_2009 ();
 b15zdnd11an1n16x5 FILLER_108_2073 ();
 b15zdnd11an1n04x5 FILLER_108_2089 ();
 b15zdnd00an1n01x5 FILLER_108_2093 ();
 b15zdnd11an1n04x5 FILLER_108_2108 ();
 b15zdnd11an1n16x5 FILLER_108_2132 ();
 b15zdnd11an1n04x5 FILLER_108_2148 ();
 b15zdnd00an1n02x5 FILLER_108_2152 ();
 b15zdnd11an1n32x5 FILLER_108_2162 ();
 b15zdnd11an1n16x5 FILLER_108_2194 ();
 b15zdnd11an1n32x5 FILLER_108_2227 ();
 b15zdnd11an1n16x5 FILLER_108_2259 ();
 b15zdnd00an1n01x5 FILLER_108_2275 ();
 b15zdnd11an1n64x5 FILLER_109_0 ();
 b15zdnd11an1n04x5 FILLER_109_64 ();
 b15zdnd00an1n02x5 FILLER_109_68 ();
 b15zdnd11an1n64x5 FILLER_109_82 ();
 b15zdnd11an1n32x5 FILLER_109_146 ();
 b15zdnd11an1n16x5 FILLER_109_178 ();
 b15zdnd11an1n04x5 FILLER_109_194 ();
 b15zdnd11an1n64x5 FILLER_109_201 ();
 b15zdnd11an1n32x5 FILLER_109_265 ();
 b15zdnd11an1n16x5 FILLER_109_297 ();
 b15zdnd11an1n08x5 FILLER_109_313 ();
 b15zdnd00an1n02x5 FILLER_109_321 ();
 b15zdnd11an1n04x5 FILLER_109_326 ();
 b15zdnd11an1n04x5 FILLER_109_335 ();
 b15zdnd11an1n04x5 FILLER_109_345 ();
 b15zdnd00an1n02x5 FILLER_109_349 ();
 b15zdnd00an1n01x5 FILLER_109_351 ();
 b15zdnd11an1n04x5 FILLER_109_394 ();
 b15zdnd11an1n16x5 FILLER_109_401 ();
 b15zdnd11an1n04x5 FILLER_109_417 ();
 b15zdnd00an1n02x5 FILLER_109_421 ();
 b15zdnd11an1n64x5 FILLER_109_465 ();
 b15zdnd11an1n32x5 FILLER_109_529 ();
 b15zdnd11an1n04x5 FILLER_109_561 ();
 b15zdnd00an1n02x5 FILLER_109_565 ();
 b15zdnd00an1n01x5 FILLER_109_567 ();
 b15zdnd11an1n64x5 FILLER_109_575 ();
 b15zdnd11an1n64x5 FILLER_109_639 ();
 b15zdnd11an1n64x5 FILLER_109_703 ();
 b15zdnd11an1n64x5 FILLER_109_767 ();
 b15zdnd11an1n64x5 FILLER_109_831 ();
 b15zdnd11an1n64x5 FILLER_109_895 ();
 b15zdnd11an1n64x5 FILLER_109_959 ();
 b15zdnd11an1n08x5 FILLER_109_1023 ();
 b15zdnd11an1n04x5 FILLER_109_1045 ();
 b15zdnd11an1n64x5 FILLER_109_1052 ();
 b15zdnd11an1n64x5 FILLER_109_1116 ();
 b15zdnd11an1n64x5 FILLER_109_1180 ();
 b15zdnd11an1n64x5 FILLER_109_1244 ();
 b15zdnd11an1n64x5 FILLER_109_1308 ();
 b15zdnd11an1n64x5 FILLER_109_1372 ();
 b15zdnd11an1n08x5 FILLER_109_1436 ();
 b15zdnd11an1n04x5 FILLER_109_1444 ();
 b15zdnd00an1n02x5 FILLER_109_1448 ();
 b15zdnd00an1n01x5 FILLER_109_1450 ();
 b15zdnd11an1n16x5 FILLER_109_1495 ();
 b15zdnd11an1n04x5 FILLER_109_1511 ();
 b15zdnd00an1n02x5 FILLER_109_1515 ();
 b15zdnd11an1n04x5 FILLER_109_1548 ();
 b15zdnd11an1n04x5 FILLER_109_1564 ();
 b15zdnd11an1n32x5 FILLER_109_1610 ();
 b15zdnd11an1n16x5 FILLER_109_1642 ();
 b15zdnd11an1n04x5 FILLER_109_1658 ();
 b15zdnd00an1n02x5 FILLER_109_1662 ();
 b15zdnd11an1n04x5 FILLER_109_1667 ();
 b15zdnd11an1n64x5 FILLER_109_1684 ();
 b15zdnd11an1n64x5 FILLER_109_1748 ();
 b15zdnd11an1n64x5 FILLER_109_1812 ();
 b15zdnd11an1n64x5 FILLER_109_1876 ();
 b15zdnd11an1n64x5 FILLER_109_1940 ();
 b15zdnd11an1n64x5 FILLER_109_2004 ();
 b15zdnd11an1n64x5 FILLER_109_2068 ();
 b15zdnd11an1n64x5 FILLER_109_2132 ();
 b15zdnd11an1n64x5 FILLER_109_2196 ();
 b15zdnd11an1n16x5 FILLER_109_2260 ();
 b15zdnd11an1n08x5 FILLER_109_2276 ();
 b15zdnd11an1n64x5 FILLER_110_8 ();
 b15zdnd11an1n64x5 FILLER_110_72 ();
 b15zdnd11an1n32x5 FILLER_110_136 ();
 b15zdnd11an1n04x5 FILLER_110_168 ();
 b15zdnd00an1n02x5 FILLER_110_172 ();
 b15zdnd00an1n01x5 FILLER_110_174 ();
 b15zdnd11an1n64x5 FILLER_110_227 ();
 b15zdnd11an1n32x5 FILLER_110_291 ();
 b15zdnd11an1n04x5 FILLER_110_323 ();
 b15zdnd00an1n02x5 FILLER_110_327 ();
 b15zdnd00an1n01x5 FILLER_110_329 ();
 b15zdnd11an1n04x5 FILLER_110_333 ();
 b15zdnd00an1n01x5 FILLER_110_337 ();
 b15zdnd11an1n04x5 FILLER_110_342 ();
 b15zdnd00an1n02x5 FILLER_110_346 ();
 b15zdnd00an1n01x5 FILLER_110_348 ();
 b15zdnd11an1n04x5 FILLER_110_353 ();
 b15zdnd00an1n02x5 FILLER_110_357 ();
 b15zdnd11an1n16x5 FILLER_110_363 ();
 b15zdnd11an1n08x5 FILLER_110_379 ();
 b15zdnd11an1n64x5 FILLER_110_402 ();
 b15zdnd11an1n64x5 FILLER_110_466 ();
 b15zdnd11an1n64x5 FILLER_110_530 ();
 b15zdnd11an1n64x5 FILLER_110_594 ();
 b15zdnd11an1n32x5 FILLER_110_658 ();
 b15zdnd11an1n16x5 FILLER_110_690 ();
 b15zdnd11an1n08x5 FILLER_110_706 ();
 b15zdnd11an1n04x5 FILLER_110_714 ();
 b15zdnd11an1n64x5 FILLER_110_726 ();
 b15zdnd11an1n64x5 FILLER_110_790 ();
 b15zdnd11an1n16x5 FILLER_110_854 ();
 b15zdnd11an1n08x5 FILLER_110_870 ();
 b15zdnd00an1n01x5 FILLER_110_878 ();
 b15zdnd11an1n04x5 FILLER_110_885 ();
 b15zdnd11an1n32x5 FILLER_110_909 ();
 b15zdnd00an1n02x5 FILLER_110_941 ();
 b15zdnd11an1n08x5 FILLER_110_957 ();
 b15zdnd00an1n02x5 FILLER_110_965 ();
 b15zdnd11an1n16x5 FILLER_110_975 ();
 b15zdnd11an1n08x5 FILLER_110_991 ();
 b15zdnd00an1n02x5 FILLER_110_999 ();
 b15zdnd00an1n01x5 FILLER_110_1001 ();
 b15zdnd11an1n04x5 FILLER_110_1044 ();
 b15zdnd11an1n64x5 FILLER_110_1061 ();
 b15zdnd11an1n64x5 FILLER_110_1125 ();
 b15zdnd11an1n64x5 FILLER_110_1189 ();
 b15zdnd11an1n64x5 FILLER_110_1253 ();
 b15zdnd11an1n64x5 FILLER_110_1317 ();
 b15zdnd11an1n64x5 FILLER_110_1381 ();
 b15zdnd11an1n16x5 FILLER_110_1445 ();
 b15zdnd00an1n02x5 FILLER_110_1461 ();
 b15zdnd00an1n01x5 FILLER_110_1463 ();
 b15zdnd11an1n04x5 FILLER_110_1467 ();
 b15zdnd11an1n04x5 FILLER_110_1474 ();
 b15zdnd11an1n16x5 FILLER_110_1481 ();
 b15zdnd11an1n08x5 FILLER_110_1497 ();
 b15zdnd11an1n04x5 FILLER_110_1505 ();
 b15zdnd00an1n01x5 FILLER_110_1509 ();
 b15zdnd11an1n04x5 FILLER_110_1513 ();
 b15zdnd11an1n64x5 FILLER_110_1527 ();
 b15zdnd11an1n04x5 FILLER_110_1591 ();
 b15zdnd00an1n02x5 FILLER_110_1595 ();
 b15zdnd00an1n01x5 FILLER_110_1597 ();
 b15zdnd11an1n64x5 FILLER_110_1601 ();
 b15zdnd11an1n16x5 FILLER_110_1665 ();
 b15zdnd00an1n01x5 FILLER_110_1681 ();
 b15zdnd11an1n64x5 FILLER_110_1685 ();
 b15zdnd11an1n04x5 FILLER_110_1749 ();
 b15zdnd00an1n02x5 FILLER_110_1753 ();
 b15zdnd11an1n64x5 FILLER_110_1761 ();
 b15zdnd11an1n64x5 FILLER_110_1825 ();
 b15zdnd11an1n08x5 FILLER_110_1889 ();
 b15zdnd00an1n02x5 FILLER_110_1897 ();
 b15zdnd00an1n01x5 FILLER_110_1899 ();
 b15zdnd11an1n64x5 FILLER_110_1904 ();
 b15zdnd11an1n64x5 FILLER_110_1968 ();
 b15zdnd11an1n64x5 FILLER_110_2032 ();
 b15zdnd11an1n32x5 FILLER_110_2096 ();
 b15zdnd11an1n16x5 FILLER_110_2128 ();
 b15zdnd11an1n08x5 FILLER_110_2144 ();
 b15zdnd00an1n02x5 FILLER_110_2152 ();
 b15zdnd11an1n64x5 FILLER_110_2162 ();
 b15zdnd11an1n32x5 FILLER_110_2226 ();
 b15zdnd11an1n16x5 FILLER_110_2258 ();
 b15zdnd00an1n02x5 FILLER_110_2274 ();
 b15zdnd11an1n64x5 FILLER_111_0 ();
 b15zdnd11an1n64x5 FILLER_111_64 ();
 b15zdnd11an1n32x5 FILLER_111_128 ();
 b15zdnd11an1n04x5 FILLER_111_160 ();
 b15zdnd00an1n02x5 FILLER_111_164 ();
 b15zdnd11an1n04x5 FILLER_111_169 ();
 b15zdnd11an1n64x5 FILLER_111_225 ();
 b15zdnd11an1n16x5 FILLER_111_289 ();
 b15zdnd11an1n08x5 FILLER_111_305 ();
 b15zdnd11an1n04x5 FILLER_111_313 ();
 b15zdnd11an1n64x5 FILLER_111_342 ();
 b15zdnd11an1n64x5 FILLER_111_406 ();
 b15zdnd11an1n64x5 FILLER_111_470 ();
 b15zdnd11an1n64x5 FILLER_111_534 ();
 b15zdnd11an1n64x5 FILLER_111_598 ();
 b15zdnd11an1n08x5 FILLER_111_662 ();
 b15zdnd11an1n04x5 FILLER_111_670 ();
 b15zdnd00an1n02x5 FILLER_111_674 ();
 b15zdnd11an1n64x5 FILLER_111_696 ();
 b15zdnd11an1n64x5 FILLER_111_760 ();
 b15zdnd11an1n64x5 FILLER_111_824 ();
 b15zdnd11an1n32x5 FILLER_111_888 ();
 b15zdnd11an1n16x5 FILLER_111_920 ();
 b15zdnd00an1n01x5 FILLER_111_936 ();
 b15zdnd11an1n32x5 FILLER_111_979 ();
 b15zdnd11an1n16x5 FILLER_111_1011 ();
 b15zdnd00an1n02x5 FILLER_111_1027 ();
 b15zdnd11an1n64x5 FILLER_111_1045 ();
 b15zdnd11an1n64x5 FILLER_111_1109 ();
 b15zdnd11an1n64x5 FILLER_111_1173 ();
 b15zdnd11an1n16x5 FILLER_111_1237 ();
 b15zdnd11an1n04x5 FILLER_111_1253 ();
 b15zdnd00an1n02x5 FILLER_111_1257 ();
 b15zdnd00an1n01x5 FILLER_111_1259 ();
 b15zdnd11an1n64x5 FILLER_111_1268 ();
 b15zdnd11an1n64x5 FILLER_111_1332 ();
 b15zdnd11an1n32x5 FILLER_111_1396 ();
 b15zdnd11an1n16x5 FILLER_111_1428 ();
 b15zdnd11an1n08x5 FILLER_111_1444 ();
 b15zdnd00an1n02x5 FILLER_111_1452 ();
 b15zdnd11an1n04x5 FILLER_111_1474 ();
 b15zdnd11an1n08x5 FILLER_111_1498 ();
 b15zdnd11an1n04x5 FILLER_111_1506 ();
 b15zdnd00an1n02x5 FILLER_111_1510 ();
 b15zdnd11an1n16x5 FILLER_111_1522 ();
 b15zdnd11an1n04x5 FILLER_111_1538 ();
 b15zdnd11an1n64x5 FILLER_111_1550 ();
 b15zdnd11an1n64x5 FILLER_111_1614 ();
 b15zdnd11an1n64x5 FILLER_111_1678 ();
 b15zdnd11an1n64x5 FILLER_111_1742 ();
 b15zdnd11an1n64x5 FILLER_111_1806 ();
 b15zdnd11an1n16x5 FILLER_111_1870 ();
 b15zdnd11an1n08x5 FILLER_111_1886 ();
 b15zdnd00an1n01x5 FILLER_111_1894 ();
 b15zdnd11an1n64x5 FILLER_111_1899 ();
 b15zdnd11an1n04x5 FILLER_111_1963 ();
 b15zdnd00an1n02x5 FILLER_111_1967 ();
 b15zdnd00an1n01x5 FILLER_111_1969 ();
 b15zdnd11an1n32x5 FILLER_111_1978 ();
 b15zdnd00an1n02x5 FILLER_111_2010 ();
 b15zdnd11an1n16x5 FILLER_111_2016 ();
 b15zdnd11an1n08x5 FILLER_111_2032 ();
 b15zdnd00an1n01x5 FILLER_111_2040 ();
 b15zdnd11an1n16x5 FILLER_111_2061 ();
 b15zdnd11an1n04x5 FILLER_111_2088 ();
 b15zdnd11an1n64x5 FILLER_111_2102 ();
 b15zdnd11an1n64x5 FILLER_111_2166 ();
 b15zdnd11an1n16x5 FILLER_111_2230 ();
 b15zdnd11an1n08x5 FILLER_111_2246 ();
 b15zdnd11an1n04x5 FILLER_111_2254 ();
 b15zdnd11an1n04x5 FILLER_111_2262 ();
 b15zdnd00an1n02x5 FILLER_111_2266 ();
 b15zdnd11an1n08x5 FILLER_111_2272 ();
 b15zdnd11an1n04x5 FILLER_111_2280 ();
 b15zdnd11an1n64x5 FILLER_112_8 ();
 b15zdnd11an1n64x5 FILLER_112_72 ();
 b15zdnd11an1n32x5 FILLER_112_136 ();
 b15zdnd11an1n16x5 FILLER_112_168 ();
 b15zdnd00an1n02x5 FILLER_112_184 ();
 b15zdnd00an1n01x5 FILLER_112_186 ();
 b15zdnd11an1n04x5 FILLER_112_190 ();
 b15zdnd11an1n04x5 FILLER_112_197 ();
 b15zdnd00an1n02x5 FILLER_112_201 ();
 b15zdnd11an1n04x5 FILLER_112_206 ();
 b15zdnd11an1n64x5 FILLER_112_224 ();
 b15zdnd11an1n64x5 FILLER_112_288 ();
 b15zdnd11an1n64x5 FILLER_112_352 ();
 b15zdnd11an1n64x5 FILLER_112_416 ();
 b15zdnd11an1n64x5 FILLER_112_480 ();
 b15zdnd11an1n64x5 FILLER_112_544 ();
 b15zdnd11an1n16x5 FILLER_112_608 ();
 b15zdnd00an1n02x5 FILLER_112_624 ();
 b15zdnd11an1n64x5 FILLER_112_629 ();
 b15zdnd11an1n16x5 FILLER_112_693 ();
 b15zdnd11an1n08x5 FILLER_112_709 ();
 b15zdnd00an1n01x5 FILLER_112_717 ();
 b15zdnd11an1n64x5 FILLER_112_726 ();
 b15zdnd11an1n64x5 FILLER_112_790 ();
 b15zdnd11an1n64x5 FILLER_112_854 ();
 b15zdnd11an1n08x5 FILLER_112_918 ();
 b15zdnd11an1n64x5 FILLER_112_978 ();
 b15zdnd11an1n64x5 FILLER_112_1042 ();
 b15zdnd11an1n64x5 FILLER_112_1106 ();
 b15zdnd11an1n64x5 FILLER_112_1170 ();
 b15zdnd11an1n64x5 FILLER_112_1234 ();
 b15zdnd11an1n64x5 FILLER_112_1298 ();
 b15zdnd11an1n64x5 FILLER_112_1362 ();
 b15zdnd11an1n64x5 FILLER_112_1426 ();
 b15zdnd11an1n16x5 FILLER_112_1490 ();
 b15zdnd00an1n02x5 FILLER_112_1506 ();
 b15zdnd00an1n01x5 FILLER_112_1508 ();
 b15zdnd11an1n04x5 FILLER_112_1515 ();
 b15zdnd00an1n02x5 FILLER_112_1519 ();
 b15zdnd11an1n64x5 FILLER_112_1524 ();
 b15zdnd11an1n64x5 FILLER_112_1588 ();
 b15zdnd11an1n08x5 FILLER_112_1652 ();
 b15zdnd00an1n02x5 FILLER_112_1660 ();
 b15zdnd00an1n01x5 FILLER_112_1662 ();
 b15zdnd11an1n64x5 FILLER_112_1672 ();
 b15zdnd11an1n64x5 FILLER_112_1736 ();
 b15zdnd11an1n64x5 FILLER_112_1800 ();
 b15zdnd11an1n64x5 FILLER_112_1864 ();
 b15zdnd11an1n64x5 FILLER_112_1928 ();
 b15zdnd11an1n16x5 FILLER_112_1992 ();
 b15zdnd11an1n64x5 FILLER_112_2012 ();
 b15zdnd11an1n64x5 FILLER_112_2076 ();
 b15zdnd11an1n08x5 FILLER_112_2140 ();
 b15zdnd11an1n04x5 FILLER_112_2148 ();
 b15zdnd00an1n02x5 FILLER_112_2152 ();
 b15zdnd11an1n64x5 FILLER_112_2162 ();
 b15zdnd11an1n16x5 FILLER_112_2226 ();
 b15zdnd11an1n08x5 FILLER_112_2242 ();
 b15zdnd00an1n02x5 FILLER_112_2250 ();
 b15zdnd11an1n04x5 FILLER_112_2256 ();
 b15zdnd11an1n04x5 FILLER_112_2264 ();
 b15zdnd11an1n04x5 FILLER_112_2272 ();
 b15zdnd11an1n64x5 FILLER_113_0 ();
 b15zdnd11an1n64x5 FILLER_113_64 ();
 b15zdnd11an1n64x5 FILLER_113_128 ();
 b15zdnd11an1n08x5 FILLER_113_192 ();
 b15zdnd11an1n04x5 FILLER_113_200 ();
 b15zdnd00an1n02x5 FILLER_113_204 ();
 b15zdnd11an1n64x5 FILLER_113_226 ();
 b15zdnd11an1n16x5 FILLER_113_290 ();
 b15zdnd11an1n08x5 FILLER_113_306 ();
 b15zdnd00an1n02x5 FILLER_113_314 ();
 b15zdnd11an1n64x5 FILLER_113_327 ();
 b15zdnd11an1n64x5 FILLER_113_391 ();
 b15zdnd11an1n64x5 FILLER_113_455 ();
 b15zdnd11an1n64x5 FILLER_113_519 ();
 b15zdnd11an1n32x5 FILLER_113_583 ();
 b15zdnd11an1n08x5 FILLER_113_615 ();
 b15zdnd00an1n02x5 FILLER_113_623 ();
 b15zdnd11an1n32x5 FILLER_113_652 ();
 b15zdnd11an1n64x5 FILLER_113_726 ();
 b15zdnd11an1n64x5 FILLER_113_790 ();
 b15zdnd11an1n64x5 FILLER_113_854 ();
 b15zdnd11an1n16x5 FILLER_113_918 ();
 b15zdnd11an1n08x5 FILLER_113_934 ();
 b15zdnd11an1n04x5 FILLER_113_942 ();
 b15zdnd11an1n04x5 FILLER_113_949 ();
 b15zdnd11an1n04x5 FILLER_113_956 ();
 b15zdnd11an1n32x5 FILLER_113_963 ();
 b15zdnd11an1n16x5 FILLER_113_995 ();
 b15zdnd11an1n08x5 FILLER_113_1011 ();
 b15zdnd11an1n04x5 FILLER_113_1019 ();
 b15zdnd11an1n04x5 FILLER_113_1029 ();
 b15zdnd00an1n02x5 FILLER_113_1033 ();
 b15zdnd11an1n64x5 FILLER_113_1049 ();
 b15zdnd11an1n32x5 FILLER_113_1113 ();
 b15zdnd11an1n16x5 FILLER_113_1145 ();
 b15zdnd00an1n02x5 FILLER_113_1161 ();
 b15zdnd00an1n01x5 FILLER_113_1163 ();
 b15zdnd11an1n64x5 FILLER_113_1180 ();
 b15zdnd11an1n64x5 FILLER_113_1244 ();
 b15zdnd11an1n64x5 FILLER_113_1308 ();
 b15zdnd11an1n64x5 FILLER_113_1372 ();
 b15zdnd11an1n64x5 FILLER_113_1436 ();
 b15zdnd11an1n64x5 FILLER_113_1500 ();
 b15zdnd11an1n64x5 FILLER_113_1564 ();
 b15zdnd11an1n64x5 FILLER_113_1628 ();
 b15zdnd11an1n64x5 FILLER_113_1692 ();
 b15zdnd11an1n64x5 FILLER_113_1756 ();
 b15zdnd11an1n32x5 FILLER_113_1820 ();
 b15zdnd11an1n16x5 FILLER_113_1852 ();
 b15zdnd11an1n04x5 FILLER_113_1868 ();
 b15zdnd00an1n01x5 FILLER_113_1872 ();
 b15zdnd11an1n32x5 FILLER_113_1877 ();
 b15zdnd11an1n16x5 FILLER_113_1909 ();
 b15zdnd11an1n04x5 FILLER_113_1925 ();
 b15zdnd00an1n02x5 FILLER_113_1929 ();
 b15zdnd00an1n01x5 FILLER_113_1931 ();
 b15zdnd11an1n64x5 FILLER_113_1938 ();
 b15zdnd11an1n64x5 FILLER_113_2002 ();
 b15zdnd11an1n64x5 FILLER_113_2066 ();
 b15zdnd11an1n32x5 FILLER_113_2130 ();
 b15zdnd11an1n16x5 FILLER_113_2162 ();
 b15zdnd11an1n08x5 FILLER_113_2178 ();
 b15zdnd11an1n04x5 FILLER_113_2186 ();
 b15zdnd11an1n32x5 FILLER_113_2202 ();
 b15zdnd11an1n04x5 FILLER_113_2234 ();
 b15zdnd00an1n02x5 FILLER_113_2238 ();
 b15zdnd00an1n02x5 FILLER_113_2282 ();
 b15zdnd11an1n64x5 FILLER_114_8 ();
 b15zdnd11an1n64x5 FILLER_114_72 ();
 b15zdnd11an1n64x5 FILLER_114_136 ();
 b15zdnd11an1n32x5 FILLER_114_200 ();
 b15zdnd00an1n02x5 FILLER_114_232 ();
 b15zdnd00an1n01x5 FILLER_114_234 ();
 b15zdnd11an1n64x5 FILLER_114_277 ();
 b15zdnd11an1n64x5 FILLER_114_341 ();
 b15zdnd11an1n04x5 FILLER_114_405 ();
 b15zdnd00an1n01x5 FILLER_114_409 ();
 b15zdnd11an1n64x5 FILLER_114_441 ();
 b15zdnd11an1n64x5 FILLER_114_505 ();
 b15zdnd11an1n16x5 FILLER_114_569 ();
 b15zdnd11an1n04x5 FILLER_114_585 ();
 b15zdnd00an1n02x5 FILLER_114_589 ();
 b15zdnd11an1n64x5 FILLER_114_594 ();
 b15zdnd11an1n32x5 FILLER_114_658 ();
 b15zdnd11an1n16x5 FILLER_114_690 ();
 b15zdnd11an1n08x5 FILLER_114_706 ();
 b15zdnd11an1n04x5 FILLER_114_714 ();
 b15zdnd11an1n64x5 FILLER_114_726 ();
 b15zdnd11an1n64x5 FILLER_114_790 ();
 b15zdnd11an1n64x5 FILLER_114_854 ();
 b15zdnd11an1n32x5 FILLER_114_918 ();
 b15zdnd00an1n01x5 FILLER_114_950 ();
 b15zdnd11an1n64x5 FILLER_114_993 ();
 b15zdnd11an1n64x5 FILLER_114_1057 ();
 b15zdnd11an1n64x5 FILLER_114_1121 ();
 b15zdnd11an1n64x5 FILLER_114_1185 ();
 b15zdnd11an1n64x5 FILLER_114_1249 ();
 b15zdnd11an1n64x5 FILLER_114_1313 ();
 b15zdnd11an1n64x5 FILLER_114_1377 ();
 b15zdnd11an1n64x5 FILLER_114_1441 ();
 b15zdnd11an1n64x5 FILLER_114_1505 ();
 b15zdnd11an1n64x5 FILLER_114_1569 ();
 b15zdnd11an1n16x5 FILLER_114_1633 ();
 b15zdnd11an1n08x5 FILLER_114_1649 ();
 b15zdnd11an1n64x5 FILLER_114_1671 ();
 b15zdnd11an1n64x5 FILLER_114_1735 ();
 b15zdnd11an1n64x5 FILLER_114_1799 ();
 b15zdnd11an1n64x5 FILLER_114_1863 ();
 b15zdnd11an1n64x5 FILLER_114_1927 ();
 b15zdnd11an1n64x5 FILLER_114_1991 ();
 b15zdnd11an1n64x5 FILLER_114_2055 ();
 b15zdnd11an1n32x5 FILLER_114_2119 ();
 b15zdnd00an1n02x5 FILLER_114_2151 ();
 b15zdnd00an1n01x5 FILLER_114_2153 ();
 b15zdnd11an1n64x5 FILLER_114_2162 ();
 b15zdnd11an1n04x5 FILLER_114_2226 ();
 b15zdnd00an1n02x5 FILLER_114_2230 ();
 b15zdnd00an1n02x5 FILLER_114_2274 ();
 b15zdnd11an1n64x5 FILLER_115_0 ();
 b15zdnd11an1n64x5 FILLER_115_64 ();
 b15zdnd11an1n64x5 FILLER_115_128 ();
 b15zdnd11an1n16x5 FILLER_115_192 ();
 b15zdnd11an1n08x5 FILLER_115_208 ();
 b15zdnd00an1n01x5 FILLER_115_216 ();
 b15zdnd11an1n64x5 FILLER_115_259 ();
 b15zdnd11an1n64x5 FILLER_115_323 ();
 b15zdnd11an1n64x5 FILLER_115_387 ();
 b15zdnd11an1n64x5 FILLER_115_451 ();
 b15zdnd11an1n32x5 FILLER_115_515 ();
 b15zdnd11an1n16x5 FILLER_115_547 ();
 b15zdnd11an1n08x5 FILLER_115_563 ();
 b15zdnd00an1n02x5 FILLER_115_571 ();
 b15zdnd11an1n64x5 FILLER_115_601 ();
 b15zdnd11an1n64x5 FILLER_115_665 ();
 b15zdnd11an1n64x5 FILLER_115_729 ();
 b15zdnd11an1n64x5 FILLER_115_793 ();
 b15zdnd11an1n64x5 FILLER_115_857 ();
 b15zdnd11an1n64x5 FILLER_115_921 ();
 b15zdnd11an1n32x5 FILLER_115_985 ();
 b15zdnd11an1n16x5 FILLER_115_1017 ();
 b15zdnd11an1n08x5 FILLER_115_1033 ();
 b15zdnd11an1n04x5 FILLER_115_1041 ();
 b15zdnd11an1n64x5 FILLER_115_1048 ();
 b15zdnd11an1n64x5 FILLER_115_1112 ();
 b15zdnd11an1n64x5 FILLER_115_1186 ();
 b15zdnd11an1n64x5 FILLER_115_1250 ();
 b15zdnd11an1n64x5 FILLER_115_1314 ();
 b15zdnd11an1n64x5 FILLER_115_1378 ();
 b15zdnd11an1n64x5 FILLER_115_1442 ();
 b15zdnd11an1n64x5 FILLER_115_1522 ();
 b15zdnd11an1n64x5 FILLER_115_1586 ();
 b15zdnd11an1n32x5 FILLER_115_1650 ();
 b15zdnd11an1n04x5 FILLER_115_1682 ();
 b15zdnd00an1n02x5 FILLER_115_1686 ();
 b15zdnd11an1n32x5 FILLER_115_1699 ();
 b15zdnd11an1n08x5 FILLER_115_1731 ();
 b15zdnd11an1n04x5 FILLER_115_1739 ();
 b15zdnd00an1n02x5 FILLER_115_1743 ();
 b15zdnd11an1n64x5 FILLER_115_1762 ();
 b15zdnd11an1n64x5 FILLER_115_1826 ();
 b15zdnd11an1n64x5 FILLER_115_1890 ();
 b15zdnd11an1n64x5 FILLER_115_1954 ();
 b15zdnd11an1n32x5 FILLER_115_2018 ();
 b15zdnd11an1n04x5 FILLER_115_2050 ();
 b15zdnd00an1n02x5 FILLER_115_2054 ();
 b15zdnd00an1n01x5 FILLER_115_2056 ();
 b15zdnd11an1n04x5 FILLER_115_2060 ();
 b15zdnd11an1n64x5 FILLER_115_2067 ();
 b15zdnd11an1n64x5 FILLER_115_2131 ();
 b15zdnd11an1n32x5 FILLER_115_2195 ();
 b15zdnd11an1n04x5 FILLER_115_2227 ();
 b15zdnd00an1n01x5 FILLER_115_2231 ();
 b15zdnd11an1n04x5 FILLER_115_2236 ();
 b15zdnd00an1n02x5 FILLER_115_2282 ();
 b15zdnd11an1n64x5 FILLER_116_8 ();
 b15zdnd11an1n64x5 FILLER_116_72 ();
 b15zdnd11an1n64x5 FILLER_116_136 ();
 b15zdnd11an1n16x5 FILLER_116_200 ();
 b15zdnd11an1n08x5 FILLER_116_216 ();
 b15zdnd00an1n02x5 FILLER_116_224 ();
 b15zdnd00an1n01x5 FILLER_116_226 ();
 b15zdnd11an1n08x5 FILLER_116_233 ();
 b15zdnd11an1n04x5 FILLER_116_241 ();
 b15zdnd00an1n01x5 FILLER_116_245 ();
 b15zdnd11an1n64x5 FILLER_116_249 ();
 b15zdnd00an1n02x5 FILLER_116_313 ();
 b15zdnd00an1n01x5 FILLER_116_315 ();
 b15zdnd11an1n64x5 FILLER_116_325 ();
 b15zdnd11an1n64x5 FILLER_116_389 ();
 b15zdnd11an1n64x5 FILLER_116_453 ();
 b15zdnd11an1n64x5 FILLER_116_517 ();
 b15zdnd11an1n08x5 FILLER_116_581 ();
 b15zdnd11an1n04x5 FILLER_116_589 ();
 b15zdnd00an1n02x5 FILLER_116_593 ();
 b15zdnd11an1n64x5 FILLER_116_598 ();
 b15zdnd11an1n32x5 FILLER_116_662 ();
 b15zdnd11an1n16x5 FILLER_116_694 ();
 b15zdnd11an1n08x5 FILLER_116_710 ();
 b15zdnd11an1n64x5 FILLER_116_726 ();
 b15zdnd11an1n64x5 FILLER_116_790 ();
 b15zdnd11an1n64x5 FILLER_116_854 ();
 b15zdnd11an1n16x5 FILLER_116_918 ();
 b15zdnd11an1n08x5 FILLER_116_934 ();
 b15zdnd00an1n02x5 FILLER_116_942 ();
 b15zdnd11an1n04x5 FILLER_116_964 ();
 b15zdnd00an1n02x5 FILLER_116_968 ();
 b15zdnd00an1n01x5 FILLER_116_970 ();
 b15zdnd11an1n32x5 FILLER_116_985 ();
 b15zdnd11an1n16x5 FILLER_116_1017 ();
 b15zdnd11an1n08x5 FILLER_116_1033 ();
 b15zdnd00an1n01x5 FILLER_116_1041 ();
 b15zdnd11an1n64x5 FILLER_116_1058 ();
 b15zdnd11an1n64x5 FILLER_116_1122 ();
 b15zdnd11an1n08x5 FILLER_116_1186 ();
 b15zdnd00an1n02x5 FILLER_116_1194 ();
 b15zdnd00an1n01x5 FILLER_116_1196 ();
 b15zdnd11an1n64x5 FILLER_116_1201 ();
 b15zdnd11an1n64x5 FILLER_116_1265 ();
 b15zdnd11an1n64x5 FILLER_116_1329 ();
 b15zdnd11an1n64x5 FILLER_116_1393 ();
 b15zdnd11an1n64x5 FILLER_116_1457 ();
 b15zdnd11an1n32x5 FILLER_116_1521 ();
 b15zdnd11an1n32x5 FILLER_116_1565 ();
 b15zdnd00an1n01x5 FILLER_116_1597 ();
 b15zdnd11an1n64x5 FILLER_116_1618 ();
 b15zdnd11an1n64x5 FILLER_116_1682 ();
 b15zdnd11an1n32x5 FILLER_116_1746 ();
 b15zdnd11an1n08x5 FILLER_116_1778 ();
 b15zdnd11an1n04x5 FILLER_116_1786 ();
 b15zdnd00an1n02x5 FILLER_116_1790 ();
 b15zdnd00an1n01x5 FILLER_116_1792 ();
 b15zdnd11an1n04x5 FILLER_116_1811 ();
 b15zdnd11an1n64x5 FILLER_116_1829 ();
 b15zdnd11an1n64x5 FILLER_116_1893 ();
 b15zdnd11an1n64x5 FILLER_116_1957 ();
 b15zdnd11an1n16x5 FILLER_116_2021 ();
 b15zdnd00an1n02x5 FILLER_116_2037 ();
 b15zdnd11an1n32x5 FILLER_116_2091 ();
 b15zdnd11an1n16x5 FILLER_116_2123 ();
 b15zdnd11an1n08x5 FILLER_116_2139 ();
 b15zdnd11an1n04x5 FILLER_116_2147 ();
 b15zdnd00an1n02x5 FILLER_116_2151 ();
 b15zdnd00an1n01x5 FILLER_116_2153 ();
 b15zdnd00an1n02x5 FILLER_116_2162 ();
 b15zdnd11an1n16x5 FILLER_116_2206 ();
 b15zdnd11an1n08x5 FILLER_116_2222 ();
 b15zdnd00an1n02x5 FILLER_116_2230 ();
 b15zdnd00an1n02x5 FILLER_116_2274 ();
 b15zdnd11an1n64x5 FILLER_117_0 ();
 b15zdnd11an1n64x5 FILLER_117_64 ();
 b15zdnd11an1n64x5 FILLER_117_128 ();
 b15zdnd11an1n64x5 FILLER_117_192 ();
 b15zdnd11an1n64x5 FILLER_117_256 ();
 b15zdnd11an1n64x5 FILLER_117_320 ();
 b15zdnd11an1n64x5 FILLER_117_384 ();
 b15zdnd11an1n16x5 FILLER_117_448 ();
 b15zdnd00an1n01x5 FILLER_117_464 ();
 b15zdnd11an1n64x5 FILLER_117_468 ();
 b15zdnd11an1n32x5 FILLER_117_532 ();
 b15zdnd11an1n04x5 FILLER_117_564 ();
 b15zdnd00an1n02x5 FILLER_117_568 ();
 b15zdnd00an1n01x5 FILLER_117_570 ();
 b15zdnd11an1n64x5 FILLER_117_611 ();
 b15zdnd11an1n64x5 FILLER_117_675 ();
 b15zdnd11an1n64x5 FILLER_117_739 ();
 b15zdnd11an1n64x5 FILLER_117_803 ();
 b15zdnd11an1n64x5 FILLER_117_867 ();
 b15zdnd11an1n64x5 FILLER_117_931 ();
 b15zdnd11an1n64x5 FILLER_117_995 ();
 b15zdnd11an1n32x5 FILLER_117_1059 ();
 b15zdnd11an1n16x5 FILLER_117_1091 ();
 b15zdnd00an1n02x5 FILLER_117_1107 ();
 b15zdnd00an1n01x5 FILLER_117_1109 ();
 b15zdnd11an1n32x5 FILLER_117_1131 ();
 b15zdnd11an1n16x5 FILLER_117_1163 ();
 b15zdnd11an1n04x5 FILLER_117_1179 ();
 b15zdnd00an1n01x5 FILLER_117_1183 ();
 b15zdnd11an1n64x5 FILLER_117_1188 ();
 b15zdnd11an1n64x5 FILLER_117_1252 ();
 b15zdnd11an1n64x5 FILLER_117_1316 ();
 b15zdnd11an1n64x5 FILLER_117_1380 ();
 b15zdnd11an1n64x5 FILLER_117_1444 ();
 b15zdnd11an1n64x5 FILLER_117_1508 ();
 b15zdnd11an1n64x5 FILLER_117_1572 ();
 b15zdnd11an1n32x5 FILLER_117_1636 ();
 b15zdnd11an1n16x5 FILLER_117_1668 ();
 b15zdnd11an1n08x5 FILLER_117_1684 ();
 b15zdnd11an1n04x5 FILLER_117_1692 ();
 b15zdnd00an1n01x5 FILLER_117_1696 ();
 b15zdnd11an1n16x5 FILLER_117_1705 ();
 b15zdnd11an1n04x5 FILLER_117_1721 ();
 b15zdnd11an1n64x5 FILLER_117_1728 ();
 b15zdnd11an1n32x5 FILLER_117_1792 ();
 b15zdnd11an1n16x5 FILLER_117_1824 ();
 b15zdnd11an1n08x5 FILLER_117_1840 ();
 b15zdnd11an1n04x5 FILLER_117_1848 ();
 b15zdnd00an1n01x5 FILLER_117_1852 ();
 b15zdnd11an1n04x5 FILLER_117_1856 ();
 b15zdnd11an1n64x5 FILLER_117_1863 ();
 b15zdnd11an1n64x5 FILLER_117_1927 ();
 b15zdnd11an1n16x5 FILLER_117_1991 ();
 b15zdnd11an1n04x5 FILLER_117_2007 ();
 b15zdnd11an1n08x5 FILLER_117_2053 ();
 b15zdnd00an1n02x5 FILLER_117_2061 ();
 b15zdnd00an1n01x5 FILLER_117_2063 ();
 b15zdnd11an1n32x5 FILLER_117_2067 ();
 b15zdnd00an1n01x5 FILLER_117_2099 ();
 b15zdnd11an1n04x5 FILLER_117_2142 ();
 b15zdnd11an1n32x5 FILLER_117_2188 ();
 b15zdnd11an1n08x5 FILLER_117_2220 ();
 b15zdnd00an1n02x5 FILLER_117_2228 ();
 b15zdnd00an1n01x5 FILLER_117_2230 ();
 b15zdnd11an1n04x5 FILLER_117_2273 ();
 b15zdnd00an1n02x5 FILLER_117_2281 ();
 b15zdnd00an1n01x5 FILLER_117_2283 ();
 b15zdnd11an1n64x5 FILLER_118_8 ();
 b15zdnd11an1n64x5 FILLER_118_72 ();
 b15zdnd11an1n64x5 FILLER_118_136 ();
 b15zdnd11an1n32x5 FILLER_118_200 ();
 b15zdnd11an1n04x5 FILLER_118_232 ();
 b15zdnd00an1n01x5 FILLER_118_236 ();
 b15zdnd11an1n64x5 FILLER_118_252 ();
 b15zdnd11an1n64x5 FILLER_118_316 ();
 b15zdnd11an1n32x5 FILLER_118_380 ();
 b15zdnd11an1n16x5 FILLER_118_412 ();
 b15zdnd00an1n01x5 FILLER_118_428 ();
 b15zdnd11an1n04x5 FILLER_118_469 ();
 b15zdnd11an1n08x5 FILLER_118_476 ();
 b15zdnd11an1n64x5 FILLER_118_491 ();
 b15zdnd11an1n04x5 FILLER_118_555 ();
 b15zdnd11an1n08x5 FILLER_118_601 ();
 b15zdnd11an1n04x5 FILLER_118_609 ();
 b15zdnd00an1n02x5 FILLER_118_613 ();
 b15zdnd11an1n64x5 FILLER_118_618 ();
 b15zdnd11an1n32x5 FILLER_118_682 ();
 b15zdnd11an1n04x5 FILLER_118_714 ();
 b15zdnd11an1n32x5 FILLER_118_726 ();
 b15zdnd11an1n16x5 FILLER_118_758 ();
 b15zdnd11an1n08x5 FILLER_118_774 ();
 b15zdnd11an1n64x5 FILLER_118_785 ();
 b15zdnd11an1n64x5 FILLER_118_849 ();
 b15zdnd11an1n64x5 FILLER_118_913 ();
 b15zdnd11an1n64x5 FILLER_118_977 ();
 b15zdnd11an1n32x5 FILLER_118_1041 ();
 b15zdnd11an1n04x5 FILLER_118_1073 ();
 b15zdnd00an1n01x5 FILLER_118_1077 ();
 b15zdnd11an1n16x5 FILLER_118_1084 ();
 b15zdnd11an1n08x5 FILLER_118_1100 ();
 b15zdnd11an1n04x5 FILLER_118_1108 ();
 b15zdnd00an1n02x5 FILLER_118_1112 ();
 b15zdnd11an1n64x5 FILLER_118_1118 ();
 b15zdnd11an1n64x5 FILLER_118_1182 ();
 b15zdnd11an1n16x5 FILLER_118_1246 ();
 b15zdnd11an1n04x5 FILLER_118_1262 ();
 b15zdnd00an1n02x5 FILLER_118_1266 ();
 b15zdnd11an1n64x5 FILLER_118_1276 ();
 b15zdnd11an1n64x5 FILLER_118_1340 ();
 b15zdnd11an1n64x5 FILLER_118_1404 ();
 b15zdnd11an1n64x5 FILLER_118_1468 ();
 b15zdnd11an1n64x5 FILLER_118_1532 ();
 b15zdnd11an1n16x5 FILLER_118_1596 ();
 b15zdnd11an1n08x5 FILLER_118_1612 ();
 b15zdnd11an1n04x5 FILLER_118_1620 ();
 b15zdnd11an1n32x5 FILLER_118_1635 ();
 b15zdnd11an1n08x5 FILLER_118_1667 ();
 b15zdnd11an1n04x5 FILLER_118_1675 ();
 b15zdnd00an1n01x5 FILLER_118_1679 ();
 b15zdnd11an1n08x5 FILLER_118_1693 ();
 b15zdnd11an1n04x5 FILLER_118_1701 ();
 b15zdnd00an1n01x5 FILLER_118_1705 ();
 b15zdnd11an1n08x5 FILLER_118_1709 ();
 b15zdnd00an1n02x5 FILLER_118_1717 ();
 b15zdnd00an1n01x5 FILLER_118_1719 ();
 b15zdnd11an1n04x5 FILLER_118_1723 ();
 b15zdnd11an1n64x5 FILLER_118_1730 ();
 b15zdnd11an1n32x5 FILLER_118_1794 ();
 b15zdnd11an1n08x5 FILLER_118_1826 ();
 b15zdnd11an1n04x5 FILLER_118_1834 ();
 b15zdnd11an1n04x5 FILLER_118_1882 ();
 b15zdnd00an1n02x5 FILLER_118_1886 ();
 b15zdnd00an1n01x5 FILLER_118_1888 ();
 b15zdnd11an1n64x5 FILLER_118_1892 ();
 b15zdnd11an1n16x5 FILLER_118_1956 ();
 b15zdnd11an1n04x5 FILLER_118_1972 ();
 b15zdnd11an1n64x5 FILLER_118_2018 ();
 b15zdnd11an1n64x5 FILLER_118_2082 ();
 b15zdnd11an1n08x5 FILLER_118_2146 ();
 b15zdnd11an1n08x5 FILLER_118_2162 ();
 b15zdnd11an1n04x5 FILLER_118_2170 ();
 b15zdnd11an1n16x5 FILLER_118_2216 ();
 b15zdnd00an1n02x5 FILLER_118_2274 ();
 b15zdnd11an1n64x5 FILLER_119_0 ();
 b15zdnd11an1n64x5 FILLER_119_64 ();
 b15zdnd11an1n64x5 FILLER_119_128 ();
 b15zdnd11an1n64x5 FILLER_119_192 ();
 b15zdnd11an1n64x5 FILLER_119_256 ();
 b15zdnd11an1n64x5 FILLER_119_320 ();
 b15zdnd11an1n64x5 FILLER_119_384 ();
 b15zdnd11an1n64x5 FILLER_119_448 ();
 b15zdnd11an1n64x5 FILLER_119_512 ();
 b15zdnd11an1n16x5 FILLER_119_576 ();
 b15zdnd11an1n08x5 FILLER_119_592 ();
 b15zdnd00an1n02x5 FILLER_119_600 ();
 b15zdnd00an1n01x5 FILLER_119_602 ();
 b15zdnd11an1n64x5 FILLER_119_606 ();
 b15zdnd11an1n64x5 FILLER_119_670 ();
 b15zdnd00an1n02x5 FILLER_119_734 ();
 b15zdnd00an1n01x5 FILLER_119_736 ();
 b15zdnd11an1n04x5 FILLER_119_789 ();
 b15zdnd00an1n02x5 FILLER_119_793 ();
 b15zdnd00an1n01x5 FILLER_119_795 ();
 b15zdnd11an1n04x5 FILLER_119_799 ();
 b15zdnd11an1n04x5 FILLER_119_806 ();
 b15zdnd11an1n64x5 FILLER_119_813 ();
 b15zdnd11an1n64x5 FILLER_119_877 ();
 b15zdnd11an1n32x5 FILLER_119_941 ();
 b15zdnd11an1n04x5 FILLER_119_973 ();
 b15zdnd00an1n02x5 FILLER_119_977 ();
 b15zdnd11an1n64x5 FILLER_119_1011 ();
 b15zdnd11an1n16x5 FILLER_119_1075 ();
 b15zdnd11an1n08x5 FILLER_119_1091 ();
 b15zdnd00an1n02x5 FILLER_119_1099 ();
 b15zdnd00an1n01x5 FILLER_119_1101 ();
 b15zdnd11an1n64x5 FILLER_119_1109 ();
 b15zdnd11an1n64x5 FILLER_119_1173 ();
 b15zdnd11an1n64x5 FILLER_119_1237 ();
 b15zdnd11an1n64x5 FILLER_119_1301 ();
 b15zdnd11an1n64x5 FILLER_119_1365 ();
 b15zdnd11an1n16x5 FILLER_119_1429 ();
 b15zdnd11an1n64x5 FILLER_119_1455 ();
 b15zdnd11an1n64x5 FILLER_119_1519 ();
 b15zdnd11an1n32x5 FILLER_119_1583 ();
 b15zdnd11an1n04x5 FILLER_119_1615 ();
 b15zdnd11an1n64x5 FILLER_119_1624 ();
 b15zdnd11an1n08x5 FILLER_119_1688 ();
 b15zdnd11an1n04x5 FILLER_119_1696 ();
 b15zdnd00an1n01x5 FILLER_119_1700 ();
 b15zdnd11an1n64x5 FILLER_119_1753 ();
 b15zdnd11an1n16x5 FILLER_119_1817 ();
 b15zdnd11an1n08x5 FILLER_119_1833 ();
 b15zdnd11an1n04x5 FILLER_119_1883 ();
 b15zdnd11an1n04x5 FILLER_119_1929 ();
 b15zdnd11an1n64x5 FILLER_119_1940 ();
 b15zdnd11an1n32x5 FILLER_119_2004 ();
 b15zdnd11an1n16x5 FILLER_119_2036 ();
 b15zdnd11an1n08x5 FILLER_119_2052 ();
 b15zdnd11an1n04x5 FILLER_119_2060 ();
 b15zdnd00an1n02x5 FILLER_119_2064 ();
 b15zdnd11an1n16x5 FILLER_119_2080 ();
 b15zdnd11an1n08x5 FILLER_119_2096 ();
 b15zdnd11an1n04x5 FILLER_119_2104 ();
 b15zdnd00an1n01x5 FILLER_119_2108 ();
 b15zdnd11an1n64x5 FILLER_119_2116 ();
 b15zdnd11an1n64x5 FILLER_119_2180 ();
 b15zdnd00an1n02x5 FILLER_119_2244 ();
 b15zdnd00an1n01x5 FILLER_119_2246 ();
 b15zdnd11an1n04x5 FILLER_119_2254 ();
 b15zdnd11an1n16x5 FILLER_119_2262 ();
 b15zdnd11an1n04x5 FILLER_119_2278 ();
 b15zdnd00an1n02x5 FILLER_119_2282 ();
 b15zdnd11an1n64x5 FILLER_120_8 ();
 b15zdnd11an1n64x5 FILLER_120_72 ();
 b15zdnd11an1n64x5 FILLER_120_136 ();
 b15zdnd11an1n64x5 FILLER_120_200 ();
 b15zdnd11an1n08x5 FILLER_120_264 ();
 b15zdnd00an1n01x5 FILLER_120_272 ();
 b15zdnd11an1n32x5 FILLER_120_277 ();
 b15zdnd11an1n16x5 FILLER_120_309 ();
 b15zdnd00an1n02x5 FILLER_120_325 ();
 b15zdnd00an1n01x5 FILLER_120_327 ();
 b15zdnd11an1n64x5 FILLER_120_336 ();
 b15zdnd11an1n64x5 FILLER_120_400 ();
 b15zdnd11an1n64x5 FILLER_120_464 ();
 b15zdnd11an1n08x5 FILLER_120_528 ();
 b15zdnd11an1n04x5 FILLER_120_536 ();
 b15zdnd00an1n01x5 FILLER_120_540 ();
 b15zdnd11an1n64x5 FILLER_120_559 ();
 b15zdnd11an1n64x5 FILLER_120_623 ();
 b15zdnd11an1n16x5 FILLER_120_687 ();
 b15zdnd11an1n08x5 FILLER_120_703 ();
 b15zdnd11an1n04x5 FILLER_120_711 ();
 b15zdnd00an1n02x5 FILLER_120_715 ();
 b15zdnd00an1n01x5 FILLER_120_717 ();
 b15zdnd11an1n32x5 FILLER_120_726 ();
 b15zdnd00an1n02x5 FILLER_120_758 ();
 b15zdnd11an1n04x5 FILLER_120_763 ();
 b15zdnd11an1n32x5 FILLER_120_819 ();
 b15zdnd11an1n16x5 FILLER_120_851 ();
 b15zdnd11an1n04x5 FILLER_120_867 ();
 b15zdnd00an1n02x5 FILLER_120_871 ();
 b15zdnd00an1n01x5 FILLER_120_873 ();
 b15zdnd11an1n64x5 FILLER_120_878 ();
 b15zdnd11an1n32x5 FILLER_120_953 ();
 b15zdnd11an1n08x5 FILLER_120_985 ();
 b15zdnd11an1n04x5 FILLER_120_993 ();
 b15zdnd00an1n01x5 FILLER_120_997 ();
 b15zdnd11an1n64x5 FILLER_120_1019 ();
 b15zdnd11an1n64x5 FILLER_120_1083 ();
 b15zdnd11an1n32x5 FILLER_120_1147 ();
 b15zdnd11an1n08x5 FILLER_120_1179 ();
 b15zdnd00an1n01x5 FILLER_120_1187 ();
 b15zdnd11an1n64x5 FILLER_120_1192 ();
 b15zdnd11an1n64x5 FILLER_120_1256 ();
 b15zdnd11an1n64x5 FILLER_120_1320 ();
 b15zdnd11an1n16x5 FILLER_120_1384 ();
 b15zdnd11an1n04x5 FILLER_120_1400 ();
 b15zdnd00an1n01x5 FILLER_120_1404 ();
 b15zdnd11an1n64x5 FILLER_120_1413 ();
 b15zdnd11an1n64x5 FILLER_120_1477 ();
 b15zdnd11an1n08x5 FILLER_120_1541 ();
 b15zdnd00an1n01x5 FILLER_120_1549 ();
 b15zdnd11an1n64x5 FILLER_120_1560 ();
 b15zdnd11an1n16x5 FILLER_120_1624 ();
 b15zdnd11an1n08x5 FILLER_120_1640 ();
 b15zdnd11an1n04x5 FILLER_120_1648 ();
 b15zdnd00an1n02x5 FILLER_120_1652 ();
 b15zdnd00an1n01x5 FILLER_120_1654 ();
 b15zdnd11an1n64x5 FILLER_120_1671 ();
 b15zdnd11an1n64x5 FILLER_120_1735 ();
 b15zdnd11an1n32x5 FILLER_120_1799 ();
 b15zdnd11an1n16x5 FILLER_120_1831 ();
 b15zdnd11an1n08x5 FILLER_120_1847 ();
 b15zdnd00an1n02x5 FILLER_120_1855 ();
 b15zdnd11an1n04x5 FILLER_120_1860 ();
 b15zdnd11an1n04x5 FILLER_120_1874 ();
 b15zdnd00an1n02x5 FILLER_120_1878 ();
 b15zdnd11an1n04x5 FILLER_120_1893 ();
 b15zdnd11an1n64x5 FILLER_120_1900 ();
 b15zdnd11an1n64x5 FILLER_120_1964 ();
 b15zdnd11an1n32x5 FILLER_120_2028 ();
 b15zdnd11an1n16x5 FILLER_120_2060 ();
 b15zdnd11an1n04x5 FILLER_120_2076 ();
 b15zdnd11an1n04x5 FILLER_120_2084 ();
 b15zdnd11an1n32x5 FILLER_120_2099 ();
 b15zdnd11an1n16x5 FILLER_120_2131 ();
 b15zdnd11an1n04x5 FILLER_120_2147 ();
 b15zdnd00an1n02x5 FILLER_120_2151 ();
 b15zdnd00an1n01x5 FILLER_120_2153 ();
 b15zdnd11an1n64x5 FILLER_120_2162 ();
 b15zdnd11an1n32x5 FILLER_120_2226 ();
 b15zdnd11an1n16x5 FILLER_120_2258 ();
 b15zdnd00an1n02x5 FILLER_120_2274 ();
 b15zdnd11an1n64x5 FILLER_121_0 ();
 b15zdnd11an1n64x5 FILLER_121_64 ();
 b15zdnd11an1n64x5 FILLER_121_128 ();
 b15zdnd11an1n64x5 FILLER_121_192 ();
 b15zdnd11an1n64x5 FILLER_121_256 ();
 b15zdnd11an1n32x5 FILLER_121_320 ();
 b15zdnd11an1n16x5 FILLER_121_352 ();
 b15zdnd11an1n08x5 FILLER_121_368 ();
 b15zdnd00an1n01x5 FILLER_121_376 ();
 b15zdnd11an1n64x5 FILLER_121_386 ();
 b15zdnd11an1n64x5 FILLER_121_450 ();
 b15zdnd11an1n64x5 FILLER_121_514 ();
 b15zdnd11an1n64x5 FILLER_121_578 ();
 b15zdnd11an1n32x5 FILLER_121_642 ();
 b15zdnd11an1n08x5 FILLER_121_674 ();
 b15zdnd11an1n04x5 FILLER_121_682 ();
 b15zdnd00an1n02x5 FILLER_121_686 ();
 b15zdnd00an1n01x5 FILLER_121_688 ();
 b15zdnd11an1n32x5 FILLER_121_709 ();
 b15zdnd11an1n16x5 FILLER_121_741 ();
 b15zdnd11an1n04x5 FILLER_121_757 ();
 b15zdnd00an1n01x5 FILLER_121_761 ();
 b15zdnd11an1n04x5 FILLER_121_765 ();
 b15zdnd11an1n08x5 FILLER_121_772 ();
 b15zdnd00an1n01x5 FILLER_121_780 ();
 b15zdnd11an1n32x5 FILLER_121_833 ();
 b15zdnd11an1n16x5 FILLER_121_865 ();
 b15zdnd00an1n02x5 FILLER_121_881 ();
 b15zdnd00an1n01x5 FILLER_121_883 ();
 b15zdnd11an1n64x5 FILLER_121_888 ();
 b15zdnd11an1n64x5 FILLER_121_952 ();
 b15zdnd11an1n64x5 FILLER_121_1016 ();
 b15zdnd11an1n32x5 FILLER_121_1080 ();
 b15zdnd11an1n16x5 FILLER_121_1112 ();
 b15zdnd11an1n04x5 FILLER_121_1128 ();
 b15zdnd00an1n02x5 FILLER_121_1132 ();
 b15zdnd11an1n64x5 FILLER_121_1143 ();
 b15zdnd11an1n16x5 FILLER_121_1207 ();
 b15zdnd00an1n02x5 FILLER_121_1223 ();
 b15zdnd00an1n01x5 FILLER_121_1225 ();
 b15zdnd11an1n32x5 FILLER_121_1235 ();
 b15zdnd11an1n16x5 FILLER_121_1267 ();
 b15zdnd00an1n02x5 FILLER_121_1283 ();
 b15zdnd11an1n04x5 FILLER_121_1289 ();
 b15zdnd00an1n02x5 FILLER_121_1293 ();
 b15zdnd11an1n16x5 FILLER_121_1299 ();
 b15zdnd11an1n08x5 FILLER_121_1315 ();
 b15zdnd11an1n04x5 FILLER_121_1323 ();
 b15zdnd00an1n01x5 FILLER_121_1327 ();
 b15zdnd11an1n64x5 FILLER_121_1334 ();
 b15zdnd11an1n32x5 FILLER_121_1398 ();
 b15zdnd11an1n04x5 FILLER_121_1430 ();
 b15zdnd00an1n02x5 FILLER_121_1434 ();
 b15zdnd00an1n01x5 FILLER_121_1436 ();
 b15zdnd11an1n04x5 FILLER_121_1453 ();
 b15zdnd11an1n64x5 FILLER_121_1467 ();
 b15zdnd11an1n16x5 FILLER_121_1531 ();
 b15zdnd11an1n04x5 FILLER_121_1547 ();
 b15zdnd00an1n01x5 FILLER_121_1551 ();
 b15zdnd11an1n04x5 FILLER_121_1561 ();
 b15zdnd11an1n64x5 FILLER_121_1586 ();
 b15zdnd11an1n64x5 FILLER_121_1650 ();
 b15zdnd11an1n08x5 FILLER_121_1714 ();
 b15zdnd00an1n02x5 FILLER_121_1722 ();
 b15zdnd11an1n64x5 FILLER_121_1750 ();
 b15zdnd11an1n32x5 FILLER_121_1814 ();
 b15zdnd11an1n08x5 FILLER_121_1846 ();
 b15zdnd00an1n02x5 FILLER_121_1854 ();
 b15zdnd11an1n08x5 FILLER_121_1872 ();
 b15zdnd11an1n04x5 FILLER_121_1880 ();
 b15zdnd00an1n02x5 FILLER_121_1884 ();
 b15zdnd11an1n04x5 FILLER_121_1910 ();
 b15zdnd11an1n64x5 FILLER_121_1934 ();
 b15zdnd11an1n64x5 FILLER_121_1998 ();
 b15zdnd11an1n32x5 FILLER_121_2062 ();
 b15zdnd11an1n04x5 FILLER_121_2094 ();
 b15zdnd00an1n01x5 FILLER_121_2098 ();
 b15zdnd11an1n16x5 FILLER_121_2119 ();
 b15zdnd11an1n04x5 FILLER_121_2135 ();
 b15zdnd11an1n64x5 FILLER_121_2165 ();
 b15zdnd11an1n32x5 FILLER_121_2229 ();
 b15zdnd11an1n16x5 FILLER_121_2261 ();
 b15zdnd11an1n04x5 FILLER_121_2277 ();
 b15zdnd00an1n02x5 FILLER_121_2281 ();
 b15zdnd00an1n01x5 FILLER_121_2283 ();
 b15zdnd11an1n64x5 FILLER_122_8 ();
 b15zdnd11an1n64x5 FILLER_122_72 ();
 b15zdnd11an1n64x5 FILLER_122_136 ();
 b15zdnd11an1n64x5 FILLER_122_200 ();
 b15zdnd11an1n04x5 FILLER_122_264 ();
 b15zdnd11an1n64x5 FILLER_122_280 ();
 b15zdnd11an1n64x5 FILLER_122_344 ();
 b15zdnd11an1n64x5 FILLER_122_408 ();
 b15zdnd11an1n64x5 FILLER_122_472 ();
 b15zdnd11an1n32x5 FILLER_122_536 ();
 b15zdnd11an1n04x5 FILLER_122_568 ();
 b15zdnd00an1n02x5 FILLER_122_572 ();
 b15zdnd00an1n01x5 FILLER_122_574 ();
 b15zdnd11an1n04x5 FILLER_122_578 ();
 b15zdnd11an1n64x5 FILLER_122_585 ();
 b15zdnd11an1n64x5 FILLER_122_649 ();
 b15zdnd11an1n04x5 FILLER_122_713 ();
 b15zdnd00an1n01x5 FILLER_122_717 ();
 b15zdnd11an1n16x5 FILLER_122_726 ();
 b15zdnd11an1n08x5 FILLER_122_742 ();
 b15zdnd11an1n04x5 FILLER_122_750 ();
 b15zdnd00an1n02x5 FILLER_122_754 ();
 b15zdnd00an1n01x5 FILLER_122_756 ();
 b15zdnd11an1n04x5 FILLER_122_809 ();
 b15zdnd11an1n64x5 FILLER_122_816 ();
 b15zdnd11an1n64x5 FILLER_122_880 ();
 b15zdnd11an1n64x5 FILLER_122_944 ();
 b15zdnd11an1n04x5 FILLER_122_1008 ();
 b15zdnd00an1n01x5 FILLER_122_1012 ();
 b15zdnd11an1n64x5 FILLER_122_1021 ();
 b15zdnd11an1n32x5 FILLER_122_1127 ();
 b15zdnd11an1n16x5 FILLER_122_1159 ();
 b15zdnd11an1n08x5 FILLER_122_1175 ();
 b15zdnd11an1n04x5 FILLER_122_1204 ();
 b15zdnd11an1n04x5 FILLER_122_1217 ();
 b15zdnd11an1n04x5 FILLER_122_1230 ();
 b15zdnd11an1n08x5 FILLER_122_1242 ();
 b15zdnd11an1n04x5 FILLER_122_1250 ();
 b15zdnd00an1n02x5 FILLER_122_1254 ();
 b15zdnd11an1n64x5 FILLER_122_1265 ();
 b15zdnd11an1n04x5 FILLER_122_1329 ();
 b15zdnd00an1n02x5 FILLER_122_1333 ();
 b15zdnd11an1n64x5 FILLER_122_1341 ();
 b15zdnd11an1n64x5 FILLER_122_1405 ();
 b15zdnd11an1n64x5 FILLER_122_1469 ();
 b15zdnd11an1n64x5 FILLER_122_1533 ();
 b15zdnd11an1n64x5 FILLER_122_1597 ();
 b15zdnd11an1n16x5 FILLER_122_1661 ();
 b15zdnd11an1n08x5 FILLER_122_1677 ();
 b15zdnd11an1n04x5 FILLER_122_1685 ();
 b15zdnd11an1n64x5 FILLER_122_1700 ();
 b15zdnd11an1n64x5 FILLER_122_1764 ();
 b15zdnd11an1n64x5 FILLER_122_1828 ();
 b15zdnd11an1n64x5 FILLER_122_1892 ();
 b15zdnd11an1n16x5 FILLER_122_1956 ();
 b15zdnd11an1n04x5 FILLER_122_1972 ();
 b15zdnd00an1n02x5 FILLER_122_1976 ();
 b15zdnd11an1n32x5 FILLER_122_2002 ();
 b15zdnd11an1n64x5 FILLER_122_2040 ();
 b15zdnd11an1n08x5 FILLER_122_2104 ();
 b15zdnd11an1n04x5 FILLER_122_2115 ();
 b15zdnd00an1n02x5 FILLER_122_2119 ();
 b15zdnd00an1n02x5 FILLER_122_2152 ();
 b15zdnd11an1n32x5 FILLER_122_2162 ();
 b15zdnd11an1n08x5 FILLER_122_2194 ();
 b15zdnd11an1n04x5 FILLER_122_2202 ();
 b15zdnd00an1n01x5 FILLER_122_2206 ();
 b15zdnd11an1n32x5 FILLER_122_2225 ();
 b15zdnd11an1n16x5 FILLER_122_2257 ();
 b15zdnd00an1n02x5 FILLER_122_2273 ();
 b15zdnd00an1n01x5 FILLER_122_2275 ();
 b15zdnd11an1n64x5 FILLER_123_0 ();
 b15zdnd11an1n64x5 FILLER_123_64 ();
 b15zdnd11an1n64x5 FILLER_123_128 ();
 b15zdnd11an1n64x5 FILLER_123_192 ();
 b15zdnd11an1n08x5 FILLER_123_256 ();
 b15zdnd11an1n04x5 FILLER_123_264 ();
 b15zdnd00an1n01x5 FILLER_123_268 ();
 b15zdnd11an1n64x5 FILLER_123_276 ();
 b15zdnd11an1n64x5 FILLER_123_340 ();
 b15zdnd11an1n08x5 FILLER_123_404 ();
 b15zdnd11an1n04x5 FILLER_123_412 ();
 b15zdnd00an1n02x5 FILLER_123_416 ();
 b15zdnd11an1n32x5 FILLER_123_436 ();
 b15zdnd11an1n04x5 FILLER_123_468 ();
 b15zdnd00an1n01x5 FILLER_123_472 ();
 b15zdnd11an1n64x5 FILLER_123_476 ();
 b15zdnd11an1n16x5 FILLER_123_540 ();
 b15zdnd00an1n02x5 FILLER_123_556 ();
 b15zdnd11an1n32x5 FILLER_123_586 ();
 b15zdnd11an1n16x5 FILLER_123_618 ();
 b15zdnd11an1n04x5 FILLER_123_634 ();
 b15zdnd00an1n02x5 FILLER_123_638 ();
 b15zdnd00an1n01x5 FILLER_123_640 ();
 b15zdnd11an1n04x5 FILLER_123_683 ();
 b15zdnd00an1n02x5 FILLER_123_687 ();
 b15zdnd11an1n16x5 FILLER_123_731 ();
 b15zdnd11an1n08x5 FILLER_123_747 ();
 b15zdnd11an1n04x5 FILLER_123_755 ();
 b15zdnd00an1n02x5 FILLER_123_759 ();
 b15zdnd00an1n01x5 FILLER_123_761 ();
 b15zdnd11an1n08x5 FILLER_123_765 ();
 b15zdnd11an1n04x5 FILLER_123_773 ();
 b15zdnd00an1n02x5 FILLER_123_777 ();
 b15zdnd00an1n01x5 FILLER_123_779 ();
 b15zdnd11an1n04x5 FILLER_123_783 ();
 b15zdnd11an1n04x5 FILLER_123_790 ();
 b15zdnd11an1n64x5 FILLER_123_797 ();
 b15zdnd11an1n04x5 FILLER_123_861 ();
 b15zdnd00an1n02x5 FILLER_123_865 ();
 b15zdnd11an1n64x5 FILLER_123_871 ();
 b15zdnd11an1n64x5 FILLER_123_935 ();
 b15zdnd11an1n64x5 FILLER_123_999 ();
 b15zdnd00an1n01x5 FILLER_123_1063 ();
 b15zdnd11an1n16x5 FILLER_123_1081 ();
 b15zdnd11an1n08x5 FILLER_123_1097 ();
 b15zdnd11an1n04x5 FILLER_123_1105 ();
 b15zdnd00an1n02x5 FILLER_123_1109 ();
 b15zdnd11an1n64x5 FILLER_123_1143 ();
 b15zdnd11an1n64x5 FILLER_123_1207 ();
 b15zdnd11an1n08x5 FILLER_123_1271 ();
 b15zdnd11an1n04x5 FILLER_123_1279 ();
 b15zdnd00an1n02x5 FILLER_123_1283 ();
 b15zdnd00an1n01x5 FILLER_123_1285 ();
 b15zdnd11an1n64x5 FILLER_123_1294 ();
 b15zdnd11an1n64x5 FILLER_123_1358 ();
 b15zdnd11an1n64x5 FILLER_123_1422 ();
 b15zdnd11an1n32x5 FILLER_123_1486 ();
 b15zdnd11an1n04x5 FILLER_123_1518 ();
 b15zdnd11an1n64x5 FILLER_123_1531 ();
 b15zdnd11an1n64x5 FILLER_123_1595 ();
 b15zdnd11an1n08x5 FILLER_123_1659 ();
 b15zdnd11an1n04x5 FILLER_123_1667 ();
 b15zdnd11an1n64x5 FILLER_123_1676 ();
 b15zdnd11an1n32x5 FILLER_123_1740 ();
 b15zdnd11an1n04x5 FILLER_123_1772 ();
 b15zdnd00an1n02x5 FILLER_123_1776 ();
 b15zdnd00an1n01x5 FILLER_123_1778 ();
 b15zdnd11an1n64x5 FILLER_123_1815 ();
 b15zdnd11an1n64x5 FILLER_123_1879 ();
 b15zdnd11an1n64x5 FILLER_123_1943 ();
 b15zdnd11an1n64x5 FILLER_123_2007 ();
 b15zdnd11an1n64x5 FILLER_123_2071 ();
 b15zdnd11an1n64x5 FILLER_123_2135 ();
 b15zdnd11an1n64x5 FILLER_123_2199 ();
 b15zdnd11an1n16x5 FILLER_123_2263 ();
 b15zdnd11an1n04x5 FILLER_123_2279 ();
 b15zdnd00an1n01x5 FILLER_123_2283 ();
 b15zdnd11an1n64x5 FILLER_124_8 ();
 b15zdnd11an1n64x5 FILLER_124_72 ();
 b15zdnd11an1n64x5 FILLER_124_136 ();
 b15zdnd11an1n64x5 FILLER_124_200 ();
 b15zdnd11an1n32x5 FILLER_124_264 ();
 b15zdnd11an1n08x5 FILLER_124_296 ();
 b15zdnd00an1n02x5 FILLER_124_304 ();
 b15zdnd11an1n64x5 FILLER_124_312 ();
 b15zdnd11an1n32x5 FILLER_124_376 ();
 b15zdnd11an1n16x5 FILLER_124_408 ();
 b15zdnd11an1n08x5 FILLER_124_424 ();
 b15zdnd11an1n04x5 FILLER_124_432 ();
 b15zdnd00an1n01x5 FILLER_124_436 ();
 b15zdnd11an1n04x5 FILLER_124_477 ();
 b15zdnd11an1n64x5 FILLER_124_484 ();
 b15zdnd11an1n64x5 FILLER_124_548 ();
 b15zdnd11an1n64x5 FILLER_124_612 ();
 b15zdnd11an1n32x5 FILLER_124_676 ();
 b15zdnd11an1n08x5 FILLER_124_708 ();
 b15zdnd00an1n02x5 FILLER_124_716 ();
 b15zdnd11an1n64x5 FILLER_124_726 ();
 b15zdnd11an1n64x5 FILLER_124_790 ();
 b15zdnd11an1n64x5 FILLER_124_854 ();
 b15zdnd11an1n64x5 FILLER_124_918 ();
 b15zdnd11an1n64x5 FILLER_124_982 ();
 b15zdnd11an1n64x5 FILLER_124_1046 ();
 b15zdnd11an1n64x5 FILLER_124_1110 ();
 b15zdnd11an1n64x5 FILLER_124_1174 ();
 b15zdnd11an1n64x5 FILLER_124_1238 ();
 b15zdnd11an1n16x5 FILLER_124_1302 ();
 b15zdnd11an1n04x5 FILLER_124_1318 ();
 b15zdnd00an1n02x5 FILLER_124_1322 ();
 b15zdnd00an1n01x5 FILLER_124_1324 ();
 b15zdnd11an1n04x5 FILLER_124_1328 ();
 b15zdnd11an1n64x5 FILLER_124_1335 ();
 b15zdnd11an1n64x5 FILLER_124_1399 ();
 b15zdnd11an1n64x5 FILLER_124_1463 ();
 b15zdnd11an1n64x5 FILLER_124_1527 ();
 b15zdnd11an1n64x5 FILLER_124_1591 ();
 b15zdnd11an1n64x5 FILLER_124_1655 ();
 b15zdnd11an1n64x5 FILLER_124_1719 ();
 b15zdnd11an1n64x5 FILLER_124_1783 ();
 b15zdnd11an1n64x5 FILLER_124_1847 ();
 b15zdnd11an1n64x5 FILLER_124_1911 ();
 b15zdnd11an1n64x5 FILLER_124_1975 ();
 b15zdnd11an1n64x5 FILLER_124_2039 ();
 b15zdnd11an1n32x5 FILLER_124_2103 ();
 b15zdnd11an1n16x5 FILLER_124_2135 ();
 b15zdnd00an1n02x5 FILLER_124_2151 ();
 b15zdnd00an1n01x5 FILLER_124_2153 ();
 b15zdnd11an1n64x5 FILLER_124_2162 ();
 b15zdnd11an1n32x5 FILLER_124_2226 ();
 b15zdnd11an1n16x5 FILLER_124_2258 ();
 b15zdnd00an1n02x5 FILLER_124_2274 ();
 b15zdnd11an1n64x5 FILLER_125_0 ();
 b15zdnd11an1n64x5 FILLER_125_64 ();
 b15zdnd11an1n64x5 FILLER_125_128 ();
 b15zdnd11an1n64x5 FILLER_125_192 ();
 b15zdnd11an1n64x5 FILLER_125_256 ();
 b15zdnd11an1n64x5 FILLER_125_320 ();
 b15zdnd11an1n64x5 FILLER_125_384 ();
 b15zdnd11an1n64x5 FILLER_125_448 ();
 b15zdnd11an1n64x5 FILLER_125_512 ();
 b15zdnd11an1n64x5 FILLER_125_576 ();
 b15zdnd11an1n64x5 FILLER_125_640 ();
 b15zdnd11an1n64x5 FILLER_125_704 ();
 b15zdnd11an1n64x5 FILLER_125_768 ();
 b15zdnd11an1n64x5 FILLER_125_832 ();
 b15zdnd11an1n32x5 FILLER_125_896 ();
 b15zdnd11an1n16x5 FILLER_125_928 ();
 b15zdnd00an1n02x5 FILLER_125_944 ();
 b15zdnd11an1n64x5 FILLER_125_963 ();
 b15zdnd11an1n16x5 FILLER_125_1027 ();
 b15zdnd11an1n08x5 FILLER_125_1043 ();
 b15zdnd11an1n04x5 FILLER_125_1051 ();
 b15zdnd00an1n01x5 FILLER_125_1055 ();
 b15zdnd11an1n32x5 FILLER_125_1065 ();
 b15zdnd11an1n16x5 FILLER_125_1097 ();
 b15zdnd11an1n04x5 FILLER_125_1113 ();
 b15zdnd00an1n01x5 FILLER_125_1117 ();
 b15zdnd11an1n64x5 FILLER_125_1129 ();
 b15zdnd11an1n64x5 FILLER_125_1193 ();
 b15zdnd11an1n16x5 FILLER_125_1257 ();
 b15zdnd11an1n08x5 FILLER_125_1273 ();
 b15zdnd11an1n04x5 FILLER_125_1281 ();
 b15zdnd00an1n02x5 FILLER_125_1285 ();
 b15zdnd00an1n01x5 FILLER_125_1287 ();
 b15zdnd11an1n04x5 FILLER_125_1292 ();
 b15zdnd11an1n04x5 FILLER_125_1302 ();
 b15zdnd11an1n64x5 FILLER_125_1358 ();
 b15zdnd11an1n32x5 FILLER_125_1422 ();
 b15zdnd11an1n04x5 FILLER_125_1454 ();
 b15zdnd00an1n02x5 FILLER_125_1458 ();
 b15zdnd11an1n64x5 FILLER_125_1480 ();
 b15zdnd11an1n64x5 FILLER_125_1544 ();
 b15zdnd11an1n64x5 FILLER_125_1608 ();
 b15zdnd11an1n64x5 FILLER_125_1672 ();
 b15zdnd11an1n64x5 FILLER_125_1736 ();
 b15zdnd11an1n64x5 FILLER_125_1800 ();
 b15zdnd11an1n64x5 FILLER_125_1864 ();
 b15zdnd11an1n64x5 FILLER_125_1928 ();
 b15zdnd11an1n64x5 FILLER_125_1992 ();
 b15zdnd11an1n64x5 FILLER_125_2056 ();
 b15zdnd11an1n64x5 FILLER_125_2120 ();
 b15zdnd11an1n64x5 FILLER_125_2184 ();
 b15zdnd11an1n32x5 FILLER_125_2248 ();
 b15zdnd11an1n04x5 FILLER_125_2280 ();
 b15zdnd11an1n64x5 FILLER_126_8 ();
 b15zdnd11an1n64x5 FILLER_126_72 ();
 b15zdnd11an1n64x5 FILLER_126_136 ();
 b15zdnd11an1n64x5 FILLER_126_200 ();
 b15zdnd11an1n16x5 FILLER_126_264 ();
 b15zdnd11an1n64x5 FILLER_126_284 ();
 b15zdnd11an1n64x5 FILLER_126_348 ();
 b15zdnd11an1n64x5 FILLER_126_412 ();
 b15zdnd11an1n64x5 FILLER_126_476 ();
 b15zdnd11an1n64x5 FILLER_126_540 ();
 b15zdnd11an1n64x5 FILLER_126_604 ();
 b15zdnd11an1n32x5 FILLER_126_668 ();
 b15zdnd11an1n16x5 FILLER_126_700 ();
 b15zdnd00an1n02x5 FILLER_126_716 ();
 b15zdnd11an1n64x5 FILLER_126_726 ();
 b15zdnd11an1n64x5 FILLER_126_790 ();
 b15zdnd11an1n04x5 FILLER_126_854 ();
 b15zdnd00an1n02x5 FILLER_126_858 ();
 b15zdnd00an1n01x5 FILLER_126_860 ();
 b15zdnd11an1n64x5 FILLER_126_865 ();
 b15zdnd11an1n64x5 FILLER_126_929 ();
 b15zdnd11an1n64x5 FILLER_126_993 ();
 b15zdnd11an1n32x5 FILLER_126_1057 ();
 b15zdnd11an1n16x5 FILLER_126_1089 ();
 b15zdnd11an1n04x5 FILLER_126_1105 ();
 b15zdnd00an1n02x5 FILLER_126_1109 ();
 b15zdnd11an1n16x5 FILLER_126_1142 ();
 b15zdnd11an1n04x5 FILLER_126_1158 ();
 b15zdnd00an1n02x5 FILLER_126_1162 ();
 b15zdnd00an1n01x5 FILLER_126_1164 ();
 b15zdnd11an1n16x5 FILLER_126_1176 ();
 b15zdnd11an1n08x5 FILLER_126_1192 ();
 b15zdnd00an1n02x5 FILLER_126_1200 ();
 b15zdnd11an1n64x5 FILLER_126_1212 ();
 b15zdnd11an1n16x5 FILLER_126_1276 ();
 b15zdnd11an1n04x5 FILLER_126_1292 ();
 b15zdnd00an1n01x5 FILLER_126_1296 ();
 b15zdnd11an1n08x5 FILLER_126_1311 ();
 b15zdnd00an1n02x5 FILLER_126_1319 ();
 b15zdnd11an1n04x5 FILLER_126_1327 ();
 b15zdnd11an1n64x5 FILLER_126_1334 ();
 b15zdnd11an1n32x5 FILLER_126_1398 ();
 b15zdnd11an1n16x5 FILLER_126_1430 ();
 b15zdnd11an1n08x5 FILLER_126_1446 ();
 b15zdnd11an1n04x5 FILLER_126_1454 ();
 b15zdnd00an1n02x5 FILLER_126_1458 ();
 b15zdnd11an1n64x5 FILLER_126_1474 ();
 b15zdnd11an1n64x5 FILLER_126_1538 ();
 b15zdnd11an1n32x5 FILLER_126_1602 ();
 b15zdnd11an1n16x5 FILLER_126_1634 ();
 b15zdnd11an1n08x5 FILLER_126_1650 ();
 b15zdnd11an1n04x5 FILLER_126_1658 ();
 b15zdnd00an1n02x5 FILLER_126_1662 ();
 b15zdnd11an1n64x5 FILLER_126_1684 ();
 b15zdnd11an1n64x5 FILLER_126_1748 ();
 b15zdnd11an1n16x5 FILLER_126_1812 ();
 b15zdnd11an1n04x5 FILLER_126_1828 ();
 b15zdnd00an1n01x5 FILLER_126_1832 ();
 b15zdnd11an1n64x5 FILLER_126_1850 ();
 b15zdnd11an1n04x5 FILLER_126_1914 ();
 b15zdnd11an1n64x5 FILLER_126_1932 ();
 b15zdnd11an1n64x5 FILLER_126_1996 ();
 b15zdnd11an1n64x5 FILLER_126_2060 ();
 b15zdnd11an1n16x5 FILLER_126_2124 ();
 b15zdnd11an1n08x5 FILLER_126_2140 ();
 b15zdnd11an1n04x5 FILLER_126_2148 ();
 b15zdnd00an1n02x5 FILLER_126_2152 ();
 b15zdnd11an1n64x5 FILLER_126_2162 ();
 b15zdnd11an1n32x5 FILLER_126_2226 ();
 b15zdnd11an1n16x5 FILLER_126_2258 ();
 b15zdnd00an1n02x5 FILLER_126_2274 ();
 b15zdnd11an1n64x5 FILLER_127_0 ();
 b15zdnd11an1n64x5 FILLER_127_64 ();
 b15zdnd11an1n64x5 FILLER_127_128 ();
 b15zdnd11an1n64x5 FILLER_127_192 ();
 b15zdnd11an1n16x5 FILLER_127_256 ();
 b15zdnd11an1n08x5 FILLER_127_272 ();
 b15zdnd00an1n02x5 FILLER_127_280 ();
 b15zdnd11an1n64x5 FILLER_127_292 ();
 b15zdnd11an1n64x5 FILLER_127_356 ();
 b15zdnd11an1n64x5 FILLER_127_420 ();
 b15zdnd11an1n64x5 FILLER_127_484 ();
 b15zdnd11an1n64x5 FILLER_127_548 ();
 b15zdnd11an1n64x5 FILLER_127_612 ();
 b15zdnd11an1n64x5 FILLER_127_676 ();
 b15zdnd11an1n64x5 FILLER_127_740 ();
 b15zdnd11an1n32x5 FILLER_127_804 ();
 b15zdnd11an1n08x5 FILLER_127_836 ();
 b15zdnd00an1n01x5 FILLER_127_844 ();
 b15zdnd11an1n64x5 FILLER_127_853 ();
 b15zdnd11an1n64x5 FILLER_127_923 ();
 b15zdnd11an1n64x5 FILLER_127_987 ();
 b15zdnd11an1n32x5 FILLER_127_1051 ();
 b15zdnd11an1n16x5 FILLER_127_1083 ();
 b15zdnd11an1n08x5 FILLER_127_1099 ();
 b15zdnd11an1n04x5 FILLER_127_1107 ();
 b15zdnd00an1n02x5 FILLER_127_1111 ();
 b15zdnd11an1n64x5 FILLER_127_1122 ();
 b15zdnd11an1n64x5 FILLER_127_1186 ();
 b15zdnd11an1n16x5 FILLER_127_1250 ();
 b15zdnd11an1n08x5 FILLER_127_1266 ();
 b15zdnd11an1n04x5 FILLER_127_1274 ();
 b15zdnd00an1n02x5 FILLER_127_1278 ();
 b15zdnd11an1n64x5 FILLER_127_1284 ();
 b15zdnd11an1n08x5 FILLER_127_1348 ();
 b15zdnd00an1n01x5 FILLER_127_1356 ();
 b15zdnd11an1n32x5 FILLER_127_1369 ();
 b15zdnd00an1n01x5 FILLER_127_1401 ();
 b15zdnd11an1n64x5 FILLER_127_1416 ();
 b15zdnd11an1n64x5 FILLER_127_1480 ();
 b15zdnd11an1n64x5 FILLER_127_1544 ();
 b15zdnd11an1n64x5 FILLER_127_1608 ();
 b15zdnd11an1n64x5 FILLER_127_1672 ();
 b15zdnd11an1n64x5 FILLER_127_1736 ();
 b15zdnd11an1n64x5 FILLER_127_1800 ();
 b15zdnd11an1n64x5 FILLER_127_1864 ();
 b15zdnd11an1n64x5 FILLER_127_1928 ();
 b15zdnd11an1n32x5 FILLER_127_1992 ();
 b15zdnd11an1n08x5 FILLER_127_2024 ();
 b15zdnd11an1n04x5 FILLER_127_2032 ();
 b15zdnd00an1n01x5 FILLER_127_2036 ();
 b15zdnd11an1n64x5 FILLER_127_2081 ();
 b15zdnd11an1n64x5 FILLER_127_2145 ();
 b15zdnd11an1n64x5 FILLER_127_2209 ();
 b15zdnd11an1n08x5 FILLER_127_2273 ();
 b15zdnd00an1n02x5 FILLER_127_2281 ();
 b15zdnd00an1n01x5 FILLER_127_2283 ();
 b15zdnd11an1n64x5 FILLER_128_8 ();
 b15zdnd00an1n02x5 FILLER_128_72 ();
 b15zdnd00an1n01x5 FILLER_128_74 ();
 b15zdnd11an1n64x5 FILLER_128_80 ();
 b15zdnd11an1n64x5 FILLER_128_144 ();
 b15zdnd11an1n16x5 FILLER_128_208 ();
 b15zdnd11an1n08x5 FILLER_128_224 ();
 b15zdnd00an1n02x5 FILLER_128_232 ();
 b15zdnd00an1n01x5 FILLER_128_234 ();
 b15zdnd11an1n16x5 FILLER_128_246 ();
 b15zdnd11an1n08x5 FILLER_128_262 ();
 b15zdnd11an1n04x5 FILLER_128_270 ();
 b15zdnd11an1n64x5 FILLER_128_284 ();
 b15zdnd11an1n64x5 FILLER_128_348 ();
 b15zdnd11an1n16x5 FILLER_128_412 ();
 b15zdnd11an1n64x5 FILLER_128_435 ();
 b15zdnd11an1n64x5 FILLER_128_499 ();
 b15zdnd11an1n64x5 FILLER_128_563 ();
 b15zdnd11an1n64x5 FILLER_128_627 ();
 b15zdnd11an1n16x5 FILLER_128_691 ();
 b15zdnd11an1n08x5 FILLER_128_707 ();
 b15zdnd00an1n02x5 FILLER_128_715 ();
 b15zdnd00an1n01x5 FILLER_128_717 ();
 b15zdnd11an1n64x5 FILLER_128_726 ();
 b15zdnd11an1n16x5 FILLER_128_790 ();
 b15zdnd11an1n08x5 FILLER_128_806 ();
 b15zdnd11an1n64x5 FILLER_128_822 ();
 b15zdnd11an1n32x5 FILLER_128_886 ();
 b15zdnd11an1n16x5 FILLER_128_918 ();
 b15zdnd11an1n08x5 FILLER_128_934 ();
 b15zdnd11an1n04x5 FILLER_128_942 ();
 b15zdnd00an1n02x5 FILLER_128_946 ();
 b15zdnd00an1n01x5 FILLER_128_948 ();
 b15zdnd11an1n64x5 FILLER_128_960 ();
 b15zdnd11an1n64x5 FILLER_128_1024 ();
 b15zdnd11an1n64x5 FILLER_128_1088 ();
 b15zdnd11an1n64x5 FILLER_128_1152 ();
 b15zdnd11an1n64x5 FILLER_128_1216 ();
 b15zdnd11an1n64x5 FILLER_128_1280 ();
 b15zdnd11an1n64x5 FILLER_128_1344 ();
 b15zdnd11an1n64x5 FILLER_128_1408 ();
 b15zdnd11an1n64x5 FILLER_128_1472 ();
 b15zdnd11an1n16x5 FILLER_128_1536 ();
 b15zdnd11an1n04x5 FILLER_128_1552 ();
 b15zdnd00an1n02x5 FILLER_128_1556 ();
 b15zdnd11an1n64x5 FILLER_128_1567 ();
 b15zdnd11an1n64x5 FILLER_128_1631 ();
 b15zdnd11an1n64x5 FILLER_128_1695 ();
 b15zdnd11an1n64x5 FILLER_128_1759 ();
 b15zdnd11an1n64x5 FILLER_128_1823 ();
 b15zdnd11an1n64x5 FILLER_128_1887 ();
 b15zdnd11an1n32x5 FILLER_128_1951 ();
 b15zdnd11an1n16x5 FILLER_128_1983 ();
 b15zdnd11an1n08x5 FILLER_128_1999 ();
 b15zdnd00an1n02x5 FILLER_128_2007 ();
 b15zdnd00an1n01x5 FILLER_128_2009 ();
 b15zdnd11an1n08x5 FILLER_128_2024 ();
 b15zdnd11an1n04x5 FILLER_128_2032 ();
 b15zdnd11an1n16x5 FILLER_128_2042 ();
 b15zdnd11an1n16x5 FILLER_128_2061 ();
 b15zdnd11an1n64x5 FILLER_128_2080 ();
 b15zdnd11an1n08x5 FILLER_128_2144 ();
 b15zdnd00an1n02x5 FILLER_128_2152 ();
 b15zdnd11an1n64x5 FILLER_128_2162 ();
 b15zdnd11an1n32x5 FILLER_128_2226 ();
 b15zdnd11an1n16x5 FILLER_128_2258 ();
 b15zdnd00an1n02x5 FILLER_128_2274 ();
 b15zdnd11an1n64x5 FILLER_129_0 ();
 b15zdnd11an1n08x5 FILLER_129_64 ();
 b15zdnd00an1n02x5 FILLER_129_72 ();
 b15zdnd11an1n64x5 FILLER_129_81 ();
 b15zdnd11an1n64x5 FILLER_129_145 ();
 b15zdnd11an1n64x5 FILLER_129_209 ();
 b15zdnd11an1n08x5 FILLER_129_273 ();
 b15zdnd00an1n01x5 FILLER_129_281 ();
 b15zdnd11an1n04x5 FILLER_129_292 ();
 b15zdnd11an1n64x5 FILLER_129_304 ();
 b15zdnd11an1n32x5 FILLER_129_368 ();
 b15zdnd11an1n16x5 FILLER_129_400 ();
 b15zdnd11an1n08x5 FILLER_129_416 ();
 b15zdnd11an1n04x5 FILLER_129_424 ();
 b15zdnd00an1n01x5 FILLER_129_428 ();
 b15zdnd11an1n16x5 FILLER_129_436 ();
 b15zdnd11an1n64x5 FILLER_129_494 ();
 b15zdnd11an1n64x5 FILLER_129_558 ();
 b15zdnd11an1n64x5 FILLER_129_622 ();
 b15zdnd11an1n08x5 FILLER_129_686 ();
 b15zdnd11an1n04x5 FILLER_129_694 ();
 b15zdnd00an1n02x5 FILLER_129_698 ();
 b15zdnd11an1n64x5 FILLER_129_742 ();
 b15zdnd11an1n64x5 FILLER_129_806 ();
 b15zdnd11an1n64x5 FILLER_129_870 ();
 b15zdnd11an1n64x5 FILLER_129_934 ();
 b15zdnd11an1n08x5 FILLER_129_998 ();
 b15zdnd11an1n04x5 FILLER_129_1006 ();
 b15zdnd00an1n02x5 FILLER_129_1010 ();
 b15zdnd11an1n64x5 FILLER_129_1019 ();
 b15zdnd11an1n64x5 FILLER_129_1083 ();
 b15zdnd11an1n64x5 FILLER_129_1147 ();
 b15zdnd11an1n64x5 FILLER_129_1211 ();
 b15zdnd11an1n16x5 FILLER_129_1275 ();
 b15zdnd11an1n08x5 FILLER_129_1291 ();
 b15zdnd00an1n02x5 FILLER_129_1299 ();
 b15zdnd11an1n64x5 FILLER_129_1307 ();
 b15zdnd11an1n64x5 FILLER_129_1371 ();
 b15zdnd11an1n64x5 FILLER_129_1447 ();
 b15zdnd11an1n32x5 FILLER_129_1511 ();
 b15zdnd11an1n16x5 FILLER_129_1543 ();
 b15zdnd11an1n08x5 FILLER_129_1559 ();
 b15zdnd00an1n02x5 FILLER_129_1567 ();
 b15zdnd11an1n64x5 FILLER_129_1578 ();
 b15zdnd11an1n64x5 FILLER_129_1642 ();
 b15zdnd11an1n64x5 FILLER_129_1706 ();
 b15zdnd11an1n64x5 FILLER_129_1770 ();
 b15zdnd11an1n64x5 FILLER_129_1834 ();
 b15zdnd11an1n64x5 FILLER_129_1898 ();
 b15zdnd11an1n32x5 FILLER_129_1962 ();
 b15zdnd11an1n16x5 FILLER_129_1994 ();
 b15zdnd00an1n02x5 FILLER_129_2010 ();
 b15zdnd11an1n04x5 FILLER_129_2057 ();
 b15zdnd11an1n64x5 FILLER_129_2064 ();
 b15zdnd11an1n64x5 FILLER_129_2128 ();
 b15zdnd11an1n64x5 FILLER_129_2192 ();
 b15zdnd11an1n16x5 FILLER_129_2256 ();
 b15zdnd11an1n08x5 FILLER_129_2272 ();
 b15zdnd11an1n04x5 FILLER_129_2280 ();
 b15zdnd11an1n64x5 FILLER_130_8 ();
 b15zdnd11an1n64x5 FILLER_130_72 ();
 b15zdnd11an1n64x5 FILLER_130_136 ();
 b15zdnd11an1n32x5 FILLER_130_200 ();
 b15zdnd11an1n16x5 FILLER_130_232 ();
 b15zdnd11an1n08x5 FILLER_130_248 ();
 b15zdnd11an1n04x5 FILLER_130_256 ();
 b15zdnd11an1n32x5 FILLER_130_302 ();
 b15zdnd11an1n04x5 FILLER_130_334 ();
 b15zdnd11an1n64x5 FILLER_130_352 ();
 b15zdnd11an1n64x5 FILLER_130_416 ();
 b15zdnd11an1n64x5 FILLER_130_480 ();
 b15zdnd11an1n64x5 FILLER_130_544 ();
 b15zdnd11an1n64x5 FILLER_130_608 ();
 b15zdnd11an1n32x5 FILLER_130_672 ();
 b15zdnd11an1n08x5 FILLER_130_704 ();
 b15zdnd11an1n04x5 FILLER_130_712 ();
 b15zdnd00an1n02x5 FILLER_130_716 ();
 b15zdnd11an1n64x5 FILLER_130_726 ();
 b15zdnd11an1n64x5 FILLER_130_790 ();
 b15zdnd11an1n64x5 FILLER_130_854 ();
 b15zdnd11an1n64x5 FILLER_130_918 ();
 b15zdnd11an1n32x5 FILLER_130_982 ();
 b15zdnd00an1n02x5 FILLER_130_1014 ();
 b15zdnd11an1n08x5 FILLER_130_1025 ();
 b15zdnd11an1n04x5 FILLER_130_1033 ();
 b15zdnd11an1n64x5 FILLER_130_1040 ();
 b15zdnd11an1n64x5 FILLER_130_1104 ();
 b15zdnd11an1n64x5 FILLER_130_1168 ();
 b15zdnd11an1n64x5 FILLER_130_1232 ();
 b15zdnd11an1n64x5 FILLER_130_1296 ();
 b15zdnd11an1n64x5 FILLER_130_1360 ();
 b15zdnd11an1n64x5 FILLER_130_1424 ();
 b15zdnd11an1n64x5 FILLER_130_1488 ();
 b15zdnd11an1n64x5 FILLER_130_1552 ();
 b15zdnd11an1n32x5 FILLER_130_1616 ();
 b15zdnd11an1n16x5 FILLER_130_1648 ();
 b15zdnd00an1n02x5 FILLER_130_1664 ();
 b15zdnd11an1n08x5 FILLER_130_1674 ();
 b15zdnd11an1n32x5 FILLER_130_1690 ();
 b15zdnd11an1n16x5 FILLER_130_1722 ();
 b15zdnd11an1n64x5 FILLER_130_1747 ();
 b15zdnd11an1n08x5 FILLER_130_1811 ();
 b15zdnd11an1n04x5 FILLER_130_1819 ();
 b15zdnd11an1n64x5 FILLER_130_1826 ();
 b15zdnd11an1n64x5 FILLER_130_1890 ();
 b15zdnd11an1n64x5 FILLER_130_1954 ();
 b15zdnd11an1n32x5 FILLER_130_2018 ();
 b15zdnd00an1n02x5 FILLER_130_2050 ();
 b15zdnd11an1n64x5 FILLER_130_2058 ();
 b15zdnd11an1n32x5 FILLER_130_2122 ();
 b15zdnd11an1n64x5 FILLER_130_2162 ();
 b15zdnd11an1n32x5 FILLER_130_2226 ();
 b15zdnd11an1n16x5 FILLER_130_2258 ();
 b15zdnd00an1n02x5 FILLER_130_2274 ();
 b15zdnd11an1n64x5 FILLER_131_0 ();
 b15zdnd11an1n64x5 FILLER_131_64 ();
 b15zdnd11an1n64x5 FILLER_131_128 ();
 b15zdnd11an1n64x5 FILLER_131_192 ();
 b15zdnd11an1n32x5 FILLER_131_256 ();
 b15zdnd11an1n64x5 FILLER_131_330 ();
 b15zdnd11an1n64x5 FILLER_131_394 ();
 b15zdnd11an1n64x5 FILLER_131_458 ();
 b15zdnd11an1n64x5 FILLER_131_522 ();
 b15zdnd11an1n64x5 FILLER_131_586 ();
 b15zdnd11an1n64x5 FILLER_131_650 ();
 b15zdnd11an1n64x5 FILLER_131_714 ();
 b15zdnd11an1n64x5 FILLER_131_778 ();
 b15zdnd11an1n32x5 FILLER_131_842 ();
 b15zdnd11an1n64x5 FILLER_131_888 ();
 b15zdnd11an1n32x5 FILLER_131_952 ();
 b15zdnd11an1n16x5 FILLER_131_984 ();
 b15zdnd11an1n08x5 FILLER_131_1000 ();
 b15zdnd00an1n02x5 FILLER_131_1008 ();
 b15zdnd11an1n32x5 FILLER_131_1062 ();
 b15zdnd11an1n16x5 FILLER_131_1094 ();
 b15zdnd11an1n04x5 FILLER_131_1110 ();
 b15zdnd00an1n01x5 FILLER_131_1114 ();
 b15zdnd11an1n64x5 FILLER_131_1124 ();
 b15zdnd11an1n64x5 FILLER_131_1188 ();
 b15zdnd11an1n64x5 FILLER_131_1252 ();
 b15zdnd11an1n64x5 FILLER_131_1316 ();
 b15zdnd11an1n08x5 FILLER_131_1380 ();
 b15zdnd00an1n02x5 FILLER_131_1388 ();
 b15zdnd00an1n01x5 FILLER_131_1390 ();
 b15zdnd11an1n64x5 FILLER_131_1412 ();
 b15zdnd11an1n64x5 FILLER_131_1476 ();
 b15zdnd11an1n64x5 FILLER_131_1540 ();
 b15zdnd11an1n64x5 FILLER_131_1604 ();
 b15zdnd11an1n64x5 FILLER_131_1668 ();
 b15zdnd11an1n64x5 FILLER_131_1732 ();
 b15zdnd11an1n64x5 FILLER_131_1796 ();
 b15zdnd11an1n64x5 FILLER_131_1860 ();
 b15zdnd11an1n64x5 FILLER_131_1924 ();
 b15zdnd11an1n64x5 FILLER_131_1988 ();
 b15zdnd11an1n64x5 FILLER_131_2052 ();
 b15zdnd11an1n64x5 FILLER_131_2116 ();
 b15zdnd11an1n64x5 FILLER_131_2180 ();
 b15zdnd11an1n32x5 FILLER_131_2244 ();
 b15zdnd11an1n08x5 FILLER_131_2276 ();
 b15zdnd11an1n08x5 FILLER_132_8 ();
 b15zdnd11an1n04x5 FILLER_132_16 ();
 b15zdnd00an1n01x5 FILLER_132_20 ();
 b15zdnd11an1n64x5 FILLER_132_25 ();
 b15zdnd11an1n64x5 FILLER_132_89 ();
 b15zdnd11an1n64x5 FILLER_132_153 ();
 b15zdnd11an1n32x5 FILLER_132_217 ();
 b15zdnd11an1n16x5 FILLER_132_249 ();
 b15zdnd11an1n08x5 FILLER_132_265 ();
 b15zdnd11an1n04x5 FILLER_132_273 ();
 b15zdnd00an1n02x5 FILLER_132_277 ();
 b15zdnd00an1n01x5 FILLER_132_279 ();
 b15zdnd11an1n64x5 FILLER_132_322 ();
 b15zdnd11an1n64x5 FILLER_132_386 ();
 b15zdnd11an1n64x5 FILLER_132_450 ();
 b15zdnd11an1n64x5 FILLER_132_514 ();
 b15zdnd11an1n64x5 FILLER_132_578 ();
 b15zdnd11an1n08x5 FILLER_132_642 ();
 b15zdnd00an1n02x5 FILLER_132_650 ();
 b15zdnd00an1n01x5 FILLER_132_652 ();
 b15zdnd11an1n32x5 FILLER_132_661 ();
 b15zdnd11an1n16x5 FILLER_132_693 ();
 b15zdnd11an1n08x5 FILLER_132_709 ();
 b15zdnd00an1n01x5 FILLER_132_717 ();
 b15zdnd11an1n64x5 FILLER_132_726 ();
 b15zdnd11an1n64x5 FILLER_132_790 ();
 b15zdnd00an1n01x5 FILLER_132_854 ();
 b15zdnd11an1n64x5 FILLER_132_859 ();
 b15zdnd11an1n64x5 FILLER_132_923 ();
 b15zdnd11an1n32x5 FILLER_132_987 ();
 b15zdnd11an1n08x5 FILLER_132_1019 ();
 b15zdnd00an1n02x5 FILLER_132_1027 ();
 b15zdnd11an1n04x5 FILLER_132_1032 ();
 b15zdnd11an1n64x5 FILLER_132_1039 ();
 b15zdnd11an1n64x5 FILLER_132_1103 ();
 b15zdnd11an1n64x5 FILLER_132_1167 ();
 b15zdnd11an1n64x5 FILLER_132_1231 ();
 b15zdnd11an1n08x5 FILLER_132_1295 ();
 b15zdnd11an1n04x5 FILLER_132_1303 ();
 b15zdnd00an1n02x5 FILLER_132_1307 ();
 b15zdnd11an1n64x5 FILLER_132_1325 ();
 b15zdnd11an1n16x5 FILLER_132_1389 ();
 b15zdnd11an1n08x5 FILLER_132_1405 ();
 b15zdnd11an1n04x5 FILLER_132_1413 ();
 b15zdnd00an1n02x5 FILLER_132_1417 ();
 b15zdnd11an1n64x5 FILLER_132_1428 ();
 b15zdnd11an1n64x5 FILLER_132_1492 ();
 b15zdnd11an1n64x5 FILLER_132_1556 ();
 b15zdnd11an1n32x5 FILLER_132_1620 ();
 b15zdnd11an1n08x5 FILLER_132_1652 ();
 b15zdnd11an1n04x5 FILLER_132_1660 ();
 b15zdnd11an1n32x5 FILLER_132_1668 ();
 b15zdnd11an1n04x5 FILLER_132_1700 ();
 b15zdnd00an1n01x5 FILLER_132_1704 ();
 b15zdnd11an1n64x5 FILLER_132_1716 ();
 b15zdnd11an1n64x5 FILLER_132_1780 ();
 b15zdnd11an1n64x5 FILLER_132_1844 ();
 b15zdnd11an1n32x5 FILLER_132_1908 ();
 b15zdnd11an1n16x5 FILLER_132_1940 ();
 b15zdnd00an1n02x5 FILLER_132_1956 ();
 b15zdnd11an1n64x5 FILLER_132_1961 ();
 b15zdnd11an1n64x5 FILLER_132_2025 ();
 b15zdnd11an1n64x5 FILLER_132_2089 ();
 b15zdnd00an1n01x5 FILLER_132_2153 ();
 b15zdnd11an1n64x5 FILLER_132_2162 ();
 b15zdnd11an1n32x5 FILLER_132_2226 ();
 b15zdnd11an1n16x5 FILLER_132_2258 ();
 b15zdnd00an1n02x5 FILLER_132_2274 ();
 b15zdnd11an1n04x5 FILLER_133_0 ();
 b15zdnd00an1n02x5 FILLER_133_4 ();
 b15zdnd11an1n64x5 FILLER_133_48 ();
 b15zdnd11an1n08x5 FILLER_133_112 ();
 b15zdnd11an1n04x5 FILLER_133_120 ();
 b15zdnd00an1n01x5 FILLER_133_124 ();
 b15zdnd11an1n08x5 FILLER_133_156 ();
 b15zdnd11an1n04x5 FILLER_133_164 ();
 b15zdnd00an1n02x5 FILLER_133_168 ();
 b15zdnd00an1n01x5 FILLER_133_170 ();
 b15zdnd11an1n64x5 FILLER_133_174 ();
 b15zdnd00an1n02x5 FILLER_133_238 ();
 b15zdnd11an1n64x5 FILLER_133_292 ();
 b15zdnd11an1n64x5 FILLER_133_356 ();
 b15zdnd11an1n32x5 FILLER_133_420 ();
 b15zdnd11an1n08x5 FILLER_133_452 ();
 b15zdnd00an1n02x5 FILLER_133_460 ();
 b15zdnd11an1n64x5 FILLER_133_466 ();
 b15zdnd11an1n64x5 FILLER_133_530 ();
 b15zdnd11an1n64x5 FILLER_133_594 ();
 b15zdnd11an1n16x5 FILLER_133_658 ();
 b15zdnd11an1n04x5 FILLER_133_674 ();
 b15zdnd11an1n64x5 FILLER_133_695 ();
 b15zdnd11an1n64x5 FILLER_133_759 ();
 b15zdnd11an1n64x5 FILLER_133_823 ();
 b15zdnd11an1n64x5 FILLER_133_887 ();
 b15zdnd11an1n64x5 FILLER_133_951 ();
 b15zdnd00an1n02x5 FILLER_133_1015 ();
 b15zdnd00an1n01x5 FILLER_133_1017 ();
 b15zdnd11an1n64x5 FILLER_133_1027 ();
 b15zdnd11an1n64x5 FILLER_133_1091 ();
 b15zdnd11an1n64x5 FILLER_133_1155 ();
 b15zdnd11an1n64x5 FILLER_133_1219 ();
 b15zdnd11an1n16x5 FILLER_133_1283 ();
 b15zdnd11an1n08x5 FILLER_133_1299 ();
 b15zdnd00an1n01x5 FILLER_133_1307 ();
 b15zdnd11an1n64x5 FILLER_133_1328 ();
 b15zdnd11an1n64x5 FILLER_133_1392 ();
 b15zdnd11an1n64x5 FILLER_133_1456 ();
 b15zdnd11an1n64x5 FILLER_133_1520 ();
 b15zdnd11an1n64x5 FILLER_133_1584 ();
 b15zdnd11an1n64x5 FILLER_133_1648 ();
 b15zdnd11an1n64x5 FILLER_133_1712 ();
 b15zdnd11an1n64x5 FILLER_133_1776 ();
 b15zdnd11an1n64x5 FILLER_133_1844 ();
 b15zdnd11an1n32x5 FILLER_133_1908 ();
 b15zdnd11an1n16x5 FILLER_133_1940 ();
 b15zdnd00an1n01x5 FILLER_133_1956 ();
 b15zdnd11an1n64x5 FILLER_133_1971 ();
 b15zdnd11an1n64x5 FILLER_133_2035 ();
 b15zdnd11an1n64x5 FILLER_133_2099 ();
 b15zdnd11an1n64x5 FILLER_133_2163 ();
 b15zdnd11an1n32x5 FILLER_133_2227 ();
 b15zdnd11an1n16x5 FILLER_133_2259 ();
 b15zdnd11an1n08x5 FILLER_133_2275 ();
 b15zdnd00an1n01x5 FILLER_133_2283 ();
 b15zdnd11an1n64x5 FILLER_134_8 ();
 b15zdnd11an1n64x5 FILLER_134_72 ();
 b15zdnd11an1n08x5 FILLER_134_136 ();
 b15zdnd00an1n01x5 FILLER_134_144 ();
 b15zdnd11an1n64x5 FILLER_134_187 ();
 b15zdnd11an1n04x5 FILLER_134_251 ();
 b15zdnd00an1n01x5 FILLER_134_255 ();
 b15zdnd11an1n04x5 FILLER_134_259 ();
 b15zdnd11an1n04x5 FILLER_134_266 ();
 b15zdnd11an1n64x5 FILLER_134_273 ();
 b15zdnd11an1n64x5 FILLER_134_337 ();
 b15zdnd11an1n32x5 FILLER_134_401 ();
 b15zdnd11an1n16x5 FILLER_134_433 ();
 b15zdnd00an1n02x5 FILLER_134_449 ();
 b15zdnd00an1n01x5 FILLER_134_451 ();
 b15zdnd11an1n04x5 FILLER_134_455 ();
 b15zdnd11an1n64x5 FILLER_134_474 ();
 b15zdnd11an1n64x5 FILLER_134_538 ();
 b15zdnd11an1n08x5 FILLER_134_602 ();
 b15zdnd00an1n02x5 FILLER_134_610 ();
 b15zdnd00an1n01x5 FILLER_134_612 ();
 b15zdnd11an1n64x5 FILLER_134_616 ();
 b15zdnd11an1n08x5 FILLER_134_680 ();
 b15zdnd11an1n04x5 FILLER_134_688 ();
 b15zdnd11an1n04x5 FILLER_134_712 ();
 b15zdnd00an1n02x5 FILLER_134_716 ();
 b15zdnd11an1n04x5 FILLER_134_726 ();
 b15zdnd00an1n02x5 FILLER_134_730 ();
 b15zdnd00an1n01x5 FILLER_134_732 ();
 b15zdnd11an1n64x5 FILLER_134_737 ();
 b15zdnd11an1n64x5 FILLER_134_801 ();
 b15zdnd00an1n02x5 FILLER_134_865 ();
 b15zdnd11an1n16x5 FILLER_134_870 ();
 b15zdnd11an1n04x5 FILLER_134_886 ();
 b15zdnd11an1n64x5 FILLER_134_914 ();
 b15zdnd11an1n16x5 FILLER_134_978 ();
 b15zdnd11an1n08x5 FILLER_134_994 ();
 b15zdnd11an1n16x5 FILLER_134_1018 ();
 b15zdnd11an1n08x5 FILLER_134_1034 ();
 b15zdnd11an1n04x5 FILLER_134_1042 ();
 b15zdnd11an1n64x5 FILLER_134_1057 ();
 b15zdnd11an1n32x5 FILLER_134_1121 ();
 b15zdnd11an1n04x5 FILLER_134_1153 ();
 b15zdnd00an1n02x5 FILLER_134_1157 ();
 b15zdnd11an1n32x5 FILLER_134_1167 ();
 b15zdnd11an1n16x5 FILLER_134_1199 ();
 b15zdnd11an1n08x5 FILLER_134_1215 ();
 b15zdnd11an1n64x5 FILLER_134_1265 ();
 b15zdnd11an1n64x5 FILLER_134_1329 ();
 b15zdnd11an1n64x5 FILLER_134_1393 ();
 b15zdnd11an1n64x5 FILLER_134_1457 ();
 b15zdnd11an1n64x5 FILLER_134_1521 ();
 b15zdnd11an1n64x5 FILLER_134_1585 ();
 b15zdnd11an1n64x5 FILLER_134_1649 ();
 b15zdnd11an1n64x5 FILLER_134_1713 ();
 b15zdnd11an1n64x5 FILLER_134_1777 ();
 b15zdnd11an1n64x5 FILLER_134_1841 ();
 b15zdnd11an1n32x5 FILLER_134_1905 ();
 b15zdnd11an1n08x5 FILLER_134_1937 ();
 b15zdnd00an1n02x5 FILLER_134_1945 ();
 b15zdnd11an1n64x5 FILLER_134_1950 ();
 b15zdnd11an1n64x5 FILLER_134_2014 ();
 b15zdnd11an1n64x5 FILLER_134_2078 ();
 b15zdnd11an1n08x5 FILLER_134_2142 ();
 b15zdnd11an1n04x5 FILLER_134_2150 ();
 b15zdnd11an1n64x5 FILLER_134_2162 ();
 b15zdnd11an1n32x5 FILLER_134_2226 ();
 b15zdnd11an1n16x5 FILLER_134_2258 ();
 b15zdnd00an1n02x5 FILLER_134_2274 ();
 b15zdnd11an1n64x5 FILLER_135_0 ();
 b15zdnd11an1n64x5 FILLER_135_64 ();
 b15zdnd11an1n16x5 FILLER_135_128 ();
 b15zdnd11an1n64x5 FILLER_135_196 ();
 b15zdnd11an1n64x5 FILLER_135_260 ();
 b15zdnd11an1n64x5 FILLER_135_324 ();
 b15zdnd11an1n64x5 FILLER_135_388 ();
 b15zdnd11an1n64x5 FILLER_135_467 ();
 b15zdnd11an1n32x5 FILLER_135_531 ();
 b15zdnd11an1n16x5 FILLER_135_563 ();
 b15zdnd11an1n04x5 FILLER_135_579 ();
 b15zdnd00an1n02x5 FILLER_135_583 ();
 b15zdnd00an1n01x5 FILLER_135_585 ();
 b15zdnd11an1n04x5 FILLER_135_638 ();
 b15zdnd11an1n08x5 FILLER_135_648 ();
 b15zdnd00an1n02x5 FILLER_135_656 ();
 b15zdnd11an1n64x5 FILLER_135_700 ();
 b15zdnd11an1n64x5 FILLER_135_764 ();
 b15zdnd11an1n64x5 FILLER_135_828 ();
 b15zdnd11an1n64x5 FILLER_135_892 ();
 b15zdnd11an1n64x5 FILLER_135_956 ();
 b15zdnd11an1n64x5 FILLER_135_1020 ();
 b15zdnd11an1n64x5 FILLER_135_1084 ();
 b15zdnd11an1n64x5 FILLER_135_1148 ();
 b15zdnd11an1n64x5 FILLER_135_1212 ();
 b15zdnd11an1n64x5 FILLER_135_1276 ();
 b15zdnd11an1n64x5 FILLER_135_1340 ();
 b15zdnd11an1n64x5 FILLER_135_1404 ();
 b15zdnd11an1n64x5 FILLER_135_1468 ();
 b15zdnd11an1n64x5 FILLER_135_1532 ();
 b15zdnd11an1n64x5 FILLER_135_1596 ();
 b15zdnd11an1n64x5 FILLER_135_1660 ();
 b15zdnd11an1n64x5 FILLER_135_1724 ();
 b15zdnd11an1n64x5 FILLER_135_1788 ();
 b15zdnd11an1n64x5 FILLER_135_1852 ();
 b15zdnd11an1n64x5 FILLER_135_1916 ();
 b15zdnd11an1n64x5 FILLER_135_1980 ();
 b15zdnd11an1n64x5 FILLER_135_2044 ();
 b15zdnd11an1n32x5 FILLER_135_2108 ();
 b15zdnd11an1n16x5 FILLER_135_2140 ();
 b15zdnd00an1n02x5 FILLER_135_2156 ();
 b15zdnd00an1n01x5 FILLER_135_2158 ();
 b15zdnd11an1n64x5 FILLER_135_2162 ();
 b15zdnd11an1n32x5 FILLER_135_2226 ();
 b15zdnd11an1n04x5 FILLER_135_2258 ();
 b15zdnd00an1n02x5 FILLER_135_2262 ();
 b15zdnd11an1n16x5 FILLER_135_2268 ();
 b15zdnd11an1n16x5 FILLER_136_8 ();
 b15zdnd11an1n04x5 FILLER_136_24 ();
 b15zdnd00an1n01x5 FILLER_136_28 ();
 b15zdnd11an1n64x5 FILLER_136_33 ();
 b15zdnd11an1n64x5 FILLER_136_97 ();
 b15zdnd00an1n01x5 FILLER_136_161 ();
 b15zdnd11an1n04x5 FILLER_136_165 ();
 b15zdnd11an1n64x5 FILLER_136_172 ();
 b15zdnd11an1n64x5 FILLER_136_236 ();
 b15zdnd11an1n64x5 FILLER_136_300 ();
 b15zdnd11an1n16x5 FILLER_136_364 ();
 b15zdnd11an1n08x5 FILLER_136_380 ();
 b15zdnd00an1n02x5 FILLER_136_388 ();
 b15zdnd11an1n64x5 FILLER_136_393 ();
 b15zdnd11an1n64x5 FILLER_136_457 ();
 b15zdnd11an1n64x5 FILLER_136_521 ();
 b15zdnd11an1n16x5 FILLER_136_585 ();
 b15zdnd00an1n02x5 FILLER_136_601 ();
 b15zdnd00an1n01x5 FILLER_136_603 ();
 b15zdnd11an1n04x5 FILLER_136_607 ();
 b15zdnd00an1n01x5 FILLER_136_611 ();
 b15zdnd11an1n32x5 FILLER_136_615 ();
 b15zdnd11an1n08x5 FILLER_136_647 ();
 b15zdnd11an1n04x5 FILLER_136_655 ();
 b15zdnd00an1n02x5 FILLER_136_659 ();
 b15zdnd11an1n04x5 FILLER_136_692 ();
 b15zdnd00an1n02x5 FILLER_136_716 ();
 b15zdnd11an1n64x5 FILLER_136_726 ();
 b15zdnd11an1n64x5 FILLER_136_790 ();
 b15zdnd11an1n64x5 FILLER_136_854 ();
 b15zdnd11an1n64x5 FILLER_136_918 ();
 b15zdnd11an1n64x5 FILLER_136_982 ();
 b15zdnd11an1n64x5 FILLER_136_1046 ();
 b15zdnd11an1n64x5 FILLER_136_1110 ();
 b15zdnd11an1n64x5 FILLER_136_1174 ();
 b15zdnd11an1n64x5 FILLER_136_1238 ();
 b15zdnd11an1n64x5 FILLER_136_1302 ();
 b15zdnd11an1n64x5 FILLER_136_1366 ();
 b15zdnd11an1n64x5 FILLER_136_1430 ();
 b15zdnd11an1n64x5 FILLER_136_1494 ();
 b15zdnd11an1n64x5 FILLER_136_1558 ();
 b15zdnd11an1n64x5 FILLER_136_1622 ();
 b15zdnd11an1n64x5 FILLER_136_1686 ();
 b15zdnd11an1n64x5 FILLER_136_1750 ();
 b15zdnd11an1n64x5 FILLER_136_1814 ();
 b15zdnd11an1n64x5 FILLER_136_1878 ();
 b15zdnd11an1n64x5 FILLER_136_1942 ();
 b15zdnd11an1n64x5 FILLER_136_2006 ();
 b15zdnd11an1n64x5 FILLER_136_2070 ();
 b15zdnd11an1n16x5 FILLER_136_2134 ();
 b15zdnd11an1n04x5 FILLER_136_2150 ();
 b15zdnd11an1n08x5 FILLER_136_2162 ();
 b15zdnd11an1n04x5 FILLER_136_2170 ();
 b15zdnd00an1n02x5 FILLER_136_2174 ();
 b15zdnd11an1n32x5 FILLER_136_2184 ();
 b15zdnd00an1n01x5 FILLER_136_2216 ();
 b15zdnd11an1n32x5 FILLER_136_2225 ();
 b15zdnd11an1n08x5 FILLER_136_2257 ();
 b15zdnd11an1n04x5 FILLER_136_2265 ();
 b15zdnd00an1n01x5 FILLER_136_2269 ();
 b15zdnd00an1n02x5 FILLER_136_2274 ();
 b15zdnd11an1n64x5 FILLER_137_0 ();
 b15zdnd11an1n64x5 FILLER_137_64 ();
 b15zdnd11an1n32x5 FILLER_137_128 ();
 b15zdnd11an1n16x5 FILLER_137_160 ();
 b15zdnd00an1n01x5 FILLER_137_176 ();
 b15zdnd11an1n04x5 FILLER_137_180 ();
 b15zdnd11an1n64x5 FILLER_137_226 ();
 b15zdnd11an1n64x5 FILLER_137_290 ();
 b15zdnd11an1n08x5 FILLER_137_354 ();
 b15zdnd00an1n01x5 FILLER_137_362 ();
 b15zdnd11an1n32x5 FILLER_137_415 ();
 b15zdnd11an1n08x5 FILLER_137_447 ();
 b15zdnd11an1n04x5 FILLER_137_455 ();
 b15zdnd00an1n01x5 FILLER_137_459 ();
 b15zdnd11an1n64x5 FILLER_137_502 ();
 b15zdnd11an1n64x5 FILLER_137_566 ();
 b15zdnd11an1n64x5 FILLER_137_630 ();
 b15zdnd11an1n64x5 FILLER_137_694 ();
 b15zdnd11an1n64x5 FILLER_137_758 ();
 b15zdnd11an1n64x5 FILLER_137_822 ();
 b15zdnd11an1n32x5 FILLER_137_886 ();
 b15zdnd11an1n08x5 FILLER_137_918 ();
 b15zdnd11an1n04x5 FILLER_137_926 ();
 b15zdnd00an1n01x5 FILLER_137_930 ();
 b15zdnd11an1n32x5 FILLER_137_947 ();
 b15zdnd11an1n16x5 FILLER_137_979 ();
 b15zdnd00an1n02x5 FILLER_137_995 ();
 b15zdnd00an1n01x5 FILLER_137_997 ();
 b15zdnd11an1n64x5 FILLER_137_1013 ();
 b15zdnd11an1n64x5 FILLER_137_1077 ();
 b15zdnd11an1n64x5 FILLER_137_1141 ();
 b15zdnd11an1n64x5 FILLER_137_1205 ();
 b15zdnd11an1n64x5 FILLER_137_1269 ();
 b15zdnd11an1n64x5 FILLER_137_1333 ();
 b15zdnd11an1n64x5 FILLER_137_1397 ();
 b15zdnd11an1n64x5 FILLER_137_1461 ();
 b15zdnd11an1n64x5 FILLER_137_1525 ();
 b15zdnd11an1n64x5 FILLER_137_1589 ();
 b15zdnd11an1n64x5 FILLER_137_1653 ();
 b15zdnd11an1n64x5 FILLER_137_1717 ();
 b15zdnd11an1n64x5 FILLER_137_1781 ();
 b15zdnd11an1n64x5 FILLER_137_1845 ();
 b15zdnd11an1n64x5 FILLER_137_1909 ();
 b15zdnd11an1n32x5 FILLER_137_1973 ();
 b15zdnd11an1n16x5 FILLER_137_2005 ();
 b15zdnd11an1n08x5 FILLER_137_2021 ();
 b15zdnd00an1n02x5 FILLER_137_2029 ();
 b15zdnd11an1n64x5 FILLER_137_2083 ();
 b15zdnd11an1n16x5 FILLER_137_2147 ();
 b15zdnd00an1n02x5 FILLER_137_2163 ();
 b15zdnd00an1n01x5 FILLER_137_2165 ();
 b15zdnd11an1n64x5 FILLER_137_2181 ();
 b15zdnd11an1n32x5 FILLER_137_2245 ();
 b15zdnd11an1n04x5 FILLER_137_2277 ();
 b15zdnd00an1n02x5 FILLER_137_2281 ();
 b15zdnd00an1n01x5 FILLER_137_2283 ();
 b15zdnd11an1n64x5 FILLER_138_8 ();
 b15zdnd11an1n64x5 FILLER_138_72 ();
 b15zdnd11an1n16x5 FILLER_138_136 ();
 b15zdnd00an1n02x5 FILLER_138_152 ();
 b15zdnd11an1n64x5 FILLER_138_206 ();
 b15zdnd11an1n64x5 FILLER_138_270 ();
 b15zdnd11an1n32x5 FILLER_138_334 ();
 b15zdnd11an1n16x5 FILLER_138_366 ();
 b15zdnd00an1n02x5 FILLER_138_382 ();
 b15zdnd11an1n04x5 FILLER_138_387 ();
 b15zdnd00an1n01x5 FILLER_138_391 ();
 b15zdnd11an1n32x5 FILLER_138_395 ();
 b15zdnd00an1n02x5 FILLER_138_427 ();
 b15zdnd00an1n01x5 FILLER_138_429 ();
 b15zdnd11an1n04x5 FILLER_138_436 ();
 b15zdnd11an1n04x5 FILLER_138_444 ();
 b15zdnd11an1n04x5 FILLER_138_490 ();
 b15zdnd11an1n16x5 FILLER_138_503 ();
 b15zdnd11an1n04x5 FILLER_138_519 ();
 b15zdnd00an1n02x5 FILLER_138_523 ();
 b15zdnd00an1n01x5 FILLER_138_525 ();
 b15zdnd11an1n64x5 FILLER_138_529 ();
 b15zdnd11an1n64x5 FILLER_138_593 ();
 b15zdnd11an1n32x5 FILLER_138_657 ();
 b15zdnd11an1n16x5 FILLER_138_689 ();
 b15zdnd11an1n04x5 FILLER_138_705 ();
 b15zdnd00an1n01x5 FILLER_138_709 ();
 b15zdnd00an1n02x5 FILLER_138_716 ();
 b15zdnd11an1n64x5 FILLER_138_726 ();
 b15zdnd11an1n64x5 FILLER_138_790 ();
 b15zdnd11an1n08x5 FILLER_138_854 ();
 b15zdnd00an1n02x5 FILLER_138_862 ();
 b15zdnd11an1n16x5 FILLER_138_878 ();
 b15zdnd11an1n08x5 FILLER_138_894 ();
 b15zdnd11an1n04x5 FILLER_138_902 ();
 b15zdnd11an1n64x5 FILLER_138_922 ();
 b15zdnd11an1n16x5 FILLER_138_986 ();
 b15zdnd11an1n08x5 FILLER_138_1002 ();
 b15zdnd11an1n04x5 FILLER_138_1010 ();
 b15zdnd00an1n02x5 FILLER_138_1014 ();
 b15zdnd11an1n64x5 FILLER_138_1026 ();
 b15zdnd11an1n64x5 FILLER_138_1090 ();
 b15zdnd11an1n64x5 FILLER_138_1154 ();
 b15zdnd11an1n64x5 FILLER_138_1218 ();
 b15zdnd11an1n64x5 FILLER_138_1282 ();
 b15zdnd11an1n64x5 FILLER_138_1346 ();
 b15zdnd11an1n64x5 FILLER_138_1410 ();
 b15zdnd11an1n64x5 FILLER_138_1474 ();
 b15zdnd11an1n64x5 FILLER_138_1538 ();
 b15zdnd11an1n64x5 FILLER_138_1602 ();
 b15zdnd11an1n16x5 FILLER_138_1666 ();
 b15zdnd11an1n04x5 FILLER_138_1682 ();
 b15zdnd11an1n64x5 FILLER_138_1697 ();
 b15zdnd11an1n64x5 FILLER_138_1761 ();
 b15zdnd11an1n64x5 FILLER_138_1825 ();
 b15zdnd11an1n64x5 FILLER_138_1889 ();
 b15zdnd11an1n64x5 FILLER_138_1953 ();
 b15zdnd11an1n32x5 FILLER_138_2017 ();
 b15zdnd11an1n04x5 FILLER_138_2052 ();
 b15zdnd11an1n04x5 FILLER_138_2059 ();
 b15zdnd11an1n64x5 FILLER_138_2066 ();
 b15zdnd11an1n16x5 FILLER_138_2130 ();
 b15zdnd11an1n08x5 FILLER_138_2146 ();
 b15zdnd11an1n08x5 FILLER_138_2162 ();
 b15zdnd00an1n01x5 FILLER_138_2170 ();
 b15zdnd11an1n32x5 FILLER_138_2182 ();
 b15zdnd11an1n16x5 FILLER_138_2214 ();
 b15zdnd11an1n08x5 FILLER_138_2230 ();
 b15zdnd11an1n04x5 FILLER_138_2238 ();
 b15zdnd11an1n16x5 FILLER_138_2246 ();
 b15zdnd11an1n08x5 FILLER_138_2262 ();
 b15zdnd11an1n04x5 FILLER_138_2270 ();
 b15zdnd00an1n02x5 FILLER_138_2274 ();
 b15zdnd11an1n64x5 FILLER_139_0 ();
 b15zdnd11an1n64x5 FILLER_139_64 ();
 b15zdnd11an1n32x5 FILLER_139_128 ();
 b15zdnd11an1n08x5 FILLER_139_160 ();
 b15zdnd11an1n04x5 FILLER_139_168 ();
 b15zdnd00an1n01x5 FILLER_139_172 ();
 b15zdnd11an1n04x5 FILLER_139_176 ();
 b15zdnd11an1n64x5 FILLER_139_183 ();
 b15zdnd11an1n64x5 FILLER_139_247 ();
 b15zdnd11an1n64x5 FILLER_139_311 ();
 b15zdnd11an1n32x5 FILLER_139_375 ();
 b15zdnd11an1n08x5 FILLER_139_407 ();
 b15zdnd11an1n04x5 FILLER_139_415 ();
 b15zdnd00an1n02x5 FILLER_139_419 ();
 b15zdnd00an1n01x5 FILLER_139_421 ();
 b15zdnd11an1n16x5 FILLER_139_464 ();
 b15zdnd00an1n02x5 FILLER_139_480 ();
 b15zdnd00an1n01x5 FILLER_139_482 ();
 b15zdnd11an1n08x5 FILLER_139_525 ();
 b15zdnd11an1n64x5 FILLER_139_536 ();
 b15zdnd11an1n64x5 FILLER_139_600 ();
 b15zdnd11an1n16x5 FILLER_139_664 ();
 b15zdnd11an1n08x5 FILLER_139_680 ();
 b15zdnd00an1n02x5 FILLER_139_688 ();
 b15zdnd00an1n01x5 FILLER_139_690 ();
 b15zdnd11an1n64x5 FILLER_139_703 ();
 b15zdnd11an1n64x5 FILLER_139_767 ();
 b15zdnd11an1n64x5 FILLER_139_831 ();
 b15zdnd11an1n16x5 FILLER_139_895 ();
 b15zdnd11an1n08x5 FILLER_139_911 ();
 b15zdnd11an1n04x5 FILLER_139_919 ();
 b15zdnd00an1n02x5 FILLER_139_923 ();
 b15zdnd11an1n04x5 FILLER_139_939 ();
 b15zdnd11an1n32x5 FILLER_139_946 ();
 b15zdnd11an1n16x5 FILLER_139_978 ();
 b15zdnd11an1n04x5 FILLER_139_994 ();
 b15zdnd00an1n02x5 FILLER_139_998 ();
 b15zdnd00an1n01x5 FILLER_139_1000 ();
 b15zdnd11an1n16x5 FILLER_139_1007 ();
 b15zdnd11an1n04x5 FILLER_139_1023 ();
 b15zdnd11an1n64x5 FILLER_139_1031 ();
 b15zdnd11an1n64x5 FILLER_139_1095 ();
 b15zdnd11an1n64x5 FILLER_139_1159 ();
 b15zdnd11an1n64x5 FILLER_139_1223 ();
 b15zdnd11an1n64x5 FILLER_139_1287 ();
 b15zdnd11an1n64x5 FILLER_139_1351 ();
 b15zdnd11an1n64x5 FILLER_139_1415 ();
 b15zdnd11an1n64x5 FILLER_139_1479 ();
 b15zdnd11an1n64x5 FILLER_139_1543 ();
 b15zdnd11an1n64x5 FILLER_139_1607 ();
 b15zdnd11an1n32x5 FILLER_139_1671 ();
 b15zdnd11an1n16x5 FILLER_139_1703 ();
 b15zdnd11an1n04x5 FILLER_139_1719 ();
 b15zdnd11an1n04x5 FILLER_139_1726 ();
 b15zdnd11an1n32x5 FILLER_139_1733 ();
 b15zdnd11an1n16x5 FILLER_139_1765 ();
 b15zdnd11an1n04x5 FILLER_139_1784 ();
 b15zdnd11an1n32x5 FILLER_139_1791 ();
 b15zdnd11an1n16x5 FILLER_139_1823 ();
 b15zdnd11an1n08x5 FILLER_139_1839 ();
 b15zdnd11an1n04x5 FILLER_139_1847 ();
 b15zdnd00an1n02x5 FILLER_139_1851 ();
 b15zdnd00an1n01x5 FILLER_139_1853 ();
 b15zdnd11an1n64x5 FILLER_139_1874 ();
 b15zdnd11an1n64x5 FILLER_139_1938 ();
 b15zdnd11an1n64x5 FILLER_139_2002 ();
 b15zdnd11an1n32x5 FILLER_139_2066 ();
 b15zdnd11an1n16x5 FILLER_139_2098 ();
 b15zdnd11an1n08x5 FILLER_139_2114 ();
 b15zdnd11an1n04x5 FILLER_139_2122 ();
 b15zdnd00an1n02x5 FILLER_139_2126 ();
 b15zdnd00an1n01x5 FILLER_139_2128 ();
 b15zdnd11an1n08x5 FILLER_139_2171 ();
 b15zdnd00an1n01x5 FILLER_139_2179 ();
 b15zdnd11an1n64x5 FILLER_139_2194 ();
 b15zdnd11an1n16x5 FILLER_139_2258 ();
 b15zdnd11an1n08x5 FILLER_139_2274 ();
 b15zdnd00an1n02x5 FILLER_139_2282 ();
 b15zdnd11an1n64x5 FILLER_140_8 ();
 b15zdnd11an1n64x5 FILLER_140_72 ();
 b15zdnd11an1n64x5 FILLER_140_136 ();
 b15zdnd11an1n64x5 FILLER_140_200 ();
 b15zdnd11an1n64x5 FILLER_140_264 ();
 b15zdnd11an1n64x5 FILLER_140_328 ();
 b15zdnd11an1n16x5 FILLER_140_392 ();
 b15zdnd11an1n04x5 FILLER_140_408 ();
 b15zdnd00an1n01x5 FILLER_140_412 ();
 b15zdnd11an1n04x5 FILLER_140_455 ();
 b15zdnd11an1n04x5 FILLER_140_468 ();
 b15zdnd11an1n04x5 FILLER_140_479 ();
 b15zdnd11an1n08x5 FILLER_140_488 ();
 b15zdnd11an1n04x5 FILLER_140_496 ();
 b15zdnd00an1n02x5 FILLER_140_500 ();
 b15zdnd00an1n01x5 FILLER_140_502 ();
 b15zdnd11an1n64x5 FILLER_140_555 ();
 b15zdnd11an1n64x5 FILLER_140_619 ();
 b15zdnd11an1n32x5 FILLER_140_683 ();
 b15zdnd00an1n02x5 FILLER_140_715 ();
 b15zdnd00an1n01x5 FILLER_140_717 ();
 b15zdnd11an1n64x5 FILLER_140_726 ();
 b15zdnd11an1n64x5 FILLER_140_790 ();
 b15zdnd11an1n64x5 FILLER_140_854 ();
 b15zdnd11an1n04x5 FILLER_140_918 ();
 b15zdnd00an1n02x5 FILLER_140_922 ();
 b15zdnd00an1n01x5 FILLER_140_924 ();
 b15zdnd11an1n04x5 FILLER_140_928 ();
 b15zdnd00an1n02x5 FILLER_140_932 ();
 b15zdnd11an1n16x5 FILLER_140_944 ();
 b15zdnd11an1n04x5 FILLER_140_960 ();
 b15zdnd00an1n02x5 FILLER_140_964 ();
 b15zdnd00an1n01x5 FILLER_140_966 ();
 b15zdnd11an1n08x5 FILLER_140_993 ();
 b15zdnd11an1n64x5 FILLER_140_1021 ();
 b15zdnd11an1n64x5 FILLER_140_1085 ();
 b15zdnd11an1n64x5 FILLER_140_1149 ();
 b15zdnd11an1n64x5 FILLER_140_1213 ();
 b15zdnd11an1n64x5 FILLER_140_1277 ();
 b15zdnd11an1n64x5 FILLER_140_1341 ();
 b15zdnd11an1n16x5 FILLER_140_1405 ();
 b15zdnd11an1n04x5 FILLER_140_1421 ();
 b15zdnd11an1n16x5 FILLER_140_1477 ();
 b15zdnd11an1n04x5 FILLER_140_1493 ();
 b15zdnd00an1n01x5 FILLER_140_1497 ();
 b15zdnd11an1n64x5 FILLER_140_1505 ();
 b15zdnd11an1n32x5 FILLER_140_1569 ();
 b15zdnd11an1n16x5 FILLER_140_1601 ();
 b15zdnd00an1n02x5 FILLER_140_1617 ();
 b15zdnd00an1n01x5 FILLER_140_1619 ();
 b15zdnd11an1n32x5 FILLER_140_1634 ();
 b15zdnd00an1n01x5 FILLER_140_1666 ();
 b15zdnd11an1n16x5 FILLER_140_1671 ();
 b15zdnd11an1n08x5 FILLER_140_1687 ();
 b15zdnd00an1n01x5 FILLER_140_1695 ();
 b15zdnd11an1n16x5 FILLER_140_1748 ();
 b15zdnd11an1n04x5 FILLER_140_1764 ();
 b15zdnd11an1n16x5 FILLER_140_1820 ();
 b15zdnd11an1n08x5 FILLER_140_1836 ();
 b15zdnd11an1n04x5 FILLER_140_1844 ();
 b15zdnd00an1n01x5 FILLER_140_1848 ();
 b15zdnd11an1n08x5 FILLER_140_1853 ();
 b15zdnd11an1n04x5 FILLER_140_1861 ();
 b15zdnd11an1n64x5 FILLER_140_1885 ();
 b15zdnd11an1n64x5 FILLER_140_1949 ();
 b15zdnd11an1n64x5 FILLER_140_2013 ();
 b15zdnd11an1n08x5 FILLER_140_2077 ();
 b15zdnd11an1n04x5 FILLER_140_2085 ();
 b15zdnd11an1n16x5 FILLER_140_2131 ();
 b15zdnd11an1n04x5 FILLER_140_2147 ();
 b15zdnd00an1n02x5 FILLER_140_2151 ();
 b15zdnd00an1n01x5 FILLER_140_2153 ();
 b15zdnd00an1n02x5 FILLER_140_2162 ();
 b15zdnd11an1n32x5 FILLER_140_2206 ();
 b15zdnd11an1n16x5 FILLER_140_2238 ();
 b15zdnd11an1n08x5 FILLER_140_2254 ();
 b15zdnd11an1n04x5 FILLER_140_2262 ();
 b15zdnd00an1n02x5 FILLER_140_2274 ();
 b15zdnd11an1n64x5 FILLER_141_0 ();
 b15zdnd11an1n64x5 FILLER_141_64 ();
 b15zdnd11an1n64x5 FILLER_141_128 ();
 b15zdnd11an1n64x5 FILLER_141_192 ();
 b15zdnd11an1n64x5 FILLER_141_256 ();
 b15zdnd11an1n64x5 FILLER_141_320 ();
 b15zdnd11an1n08x5 FILLER_141_384 ();
 b15zdnd11an1n04x5 FILLER_141_392 ();
 b15zdnd00an1n02x5 FILLER_141_396 ();
 b15zdnd00an1n01x5 FILLER_141_398 ();
 b15zdnd11an1n08x5 FILLER_141_441 ();
 b15zdnd11an1n04x5 FILLER_141_449 ();
 b15zdnd00an1n01x5 FILLER_141_453 ();
 b15zdnd11an1n08x5 FILLER_141_457 ();
 b15zdnd11an1n04x5 FILLER_141_465 ();
 b15zdnd11an1n04x5 FILLER_141_474 ();
 b15zdnd00an1n02x5 FILLER_141_478 ();
 b15zdnd00an1n01x5 FILLER_141_480 ();
 b15zdnd11an1n08x5 FILLER_141_485 ();
 b15zdnd11an1n04x5 FILLER_141_493 ();
 b15zdnd00an1n02x5 FILLER_141_497 ();
 b15zdnd00an1n01x5 FILLER_141_499 ();
 b15zdnd11an1n04x5 FILLER_141_507 ();
 b15zdnd11an1n04x5 FILLER_141_514 ();
 b15zdnd00an1n02x5 FILLER_141_518 ();
 b15zdnd11an1n04x5 FILLER_141_526 ();
 b15zdnd11an1n04x5 FILLER_141_533 ();
 b15zdnd11an1n64x5 FILLER_141_579 ();
 b15zdnd11an1n64x5 FILLER_141_643 ();
 b15zdnd11an1n08x5 FILLER_141_707 ();
 b15zdnd11an1n04x5 FILLER_141_715 ();
 b15zdnd00an1n01x5 FILLER_141_719 ();
 b15zdnd11an1n64x5 FILLER_141_740 ();
 b15zdnd11an1n16x5 FILLER_141_804 ();
 b15zdnd11an1n04x5 FILLER_141_820 ();
 b15zdnd00an1n01x5 FILLER_141_824 ();
 b15zdnd11an1n64x5 FILLER_141_828 ();
 b15zdnd11an1n64x5 FILLER_141_892 ();
 b15zdnd11an1n16x5 FILLER_141_956 ();
 b15zdnd11an1n08x5 FILLER_141_972 ();
 b15zdnd11an1n04x5 FILLER_141_980 ();
 b15zdnd00an1n01x5 FILLER_141_984 ();
 b15zdnd11an1n32x5 FILLER_141_1016 ();
 b15zdnd11an1n08x5 FILLER_141_1048 ();
 b15zdnd11an1n04x5 FILLER_141_1056 ();
 b15zdnd11an1n64x5 FILLER_141_1069 ();
 b15zdnd11an1n16x5 FILLER_141_1133 ();
 b15zdnd00an1n02x5 FILLER_141_1149 ();
 b15zdnd11an1n64x5 FILLER_141_1159 ();
 b15zdnd11an1n64x5 FILLER_141_1223 ();
 b15zdnd11an1n64x5 FILLER_141_1287 ();
 b15zdnd11an1n64x5 FILLER_141_1351 ();
 b15zdnd11an1n16x5 FILLER_141_1415 ();
 b15zdnd11an1n08x5 FILLER_141_1431 ();
 b15zdnd11an1n04x5 FILLER_141_1439 ();
 b15zdnd00an1n01x5 FILLER_141_1443 ();
 b15zdnd11an1n04x5 FILLER_141_1447 ();
 b15zdnd11an1n04x5 FILLER_141_1454 ();
 b15zdnd11an1n64x5 FILLER_141_1461 ();
 b15zdnd11an1n64x5 FILLER_141_1525 ();
 b15zdnd11an1n64x5 FILLER_141_1589 ();
 b15zdnd11an1n08x5 FILLER_141_1653 ();
 b15zdnd11an1n04x5 FILLER_141_1665 ();
 b15zdnd11an1n16x5 FILLER_141_1673 ();
 b15zdnd11an1n08x5 FILLER_141_1689 ();
 b15zdnd11an1n04x5 FILLER_141_1697 ();
 b15zdnd00an1n02x5 FILLER_141_1701 ();
 b15zdnd11an1n04x5 FILLER_141_1755 ();
 b15zdnd11an1n64x5 FILLER_141_1811 ();
 b15zdnd11an1n32x5 FILLER_141_1875 ();
 b15zdnd11an1n16x5 FILLER_141_1907 ();
 b15zdnd11an1n04x5 FILLER_141_1923 ();
 b15zdnd00an1n02x5 FILLER_141_1927 ();
 b15zdnd11an1n64x5 FILLER_141_1942 ();
 b15zdnd11an1n64x5 FILLER_141_2006 ();
 b15zdnd11an1n64x5 FILLER_141_2070 ();
 b15zdnd11an1n08x5 FILLER_141_2134 ();
 b15zdnd00an1n02x5 FILLER_141_2142 ();
 b15zdnd11an1n04x5 FILLER_141_2186 ();
 b15zdnd11an1n32x5 FILLER_141_2232 ();
 b15zdnd11an1n16x5 FILLER_141_2264 ();
 b15zdnd11an1n04x5 FILLER_141_2280 ();
 b15zdnd11an1n64x5 FILLER_142_8 ();
 b15zdnd11an1n64x5 FILLER_142_72 ();
 b15zdnd11an1n64x5 FILLER_142_136 ();
 b15zdnd11an1n64x5 FILLER_142_200 ();
 b15zdnd11an1n64x5 FILLER_142_264 ();
 b15zdnd11an1n64x5 FILLER_142_328 ();
 b15zdnd11an1n32x5 FILLER_142_392 ();
 b15zdnd11an1n08x5 FILLER_142_424 ();
 b15zdnd11an1n64x5 FILLER_142_436 ();
 b15zdnd11an1n08x5 FILLER_142_500 ();
 b15zdnd11an1n04x5 FILLER_142_508 ();
 b15zdnd11an1n04x5 FILLER_142_554 ();
 b15zdnd11an1n32x5 FILLER_142_565 ();
 b15zdnd11an1n16x5 FILLER_142_597 ();
 b15zdnd11an1n04x5 FILLER_142_613 ();
 b15zdnd11an1n16x5 FILLER_142_659 ();
 b15zdnd00an1n02x5 FILLER_142_675 ();
 b15zdnd11an1n16x5 FILLER_142_698 ();
 b15zdnd11an1n04x5 FILLER_142_714 ();
 b15zdnd11an1n64x5 FILLER_142_726 ();
 b15zdnd11an1n08x5 FILLER_142_790 ();
 b15zdnd00an1n02x5 FILLER_142_798 ();
 b15zdnd00an1n01x5 FILLER_142_800 ();
 b15zdnd11an1n64x5 FILLER_142_845 ();
 b15zdnd11an1n64x5 FILLER_142_909 ();
 b15zdnd11an1n64x5 FILLER_142_973 ();
 b15zdnd11an1n64x5 FILLER_142_1037 ();
 b15zdnd11an1n08x5 FILLER_142_1101 ();
 b15zdnd00an1n02x5 FILLER_142_1109 ();
 b15zdnd00an1n01x5 FILLER_142_1111 ();
 b15zdnd11an1n04x5 FILLER_142_1164 ();
 b15zdnd00an1n02x5 FILLER_142_1168 ();
 b15zdnd00an1n01x5 FILLER_142_1170 ();
 b15zdnd11an1n64x5 FILLER_142_1179 ();
 b15zdnd11an1n16x5 FILLER_142_1243 ();
 b15zdnd00an1n02x5 FILLER_142_1259 ();
 b15zdnd11an1n64x5 FILLER_142_1269 ();
 b15zdnd11an1n64x5 FILLER_142_1333 ();
 b15zdnd11an1n16x5 FILLER_142_1397 ();
 b15zdnd00an1n01x5 FILLER_142_1413 ();
 b15zdnd11an1n08x5 FILLER_142_1423 ();
 b15zdnd11an1n04x5 FILLER_142_1431 ();
 b15zdnd00an1n02x5 FILLER_142_1435 ();
 b15zdnd11an1n64x5 FILLER_142_1479 ();
 b15zdnd11an1n64x5 FILLER_142_1543 ();
 b15zdnd11an1n64x5 FILLER_142_1607 ();
 b15zdnd11an1n08x5 FILLER_142_1671 ();
 b15zdnd00an1n01x5 FILLER_142_1679 ();
 b15zdnd11an1n16x5 FILLER_142_1688 ();
 b15zdnd11an1n08x5 FILLER_142_1704 ();
 b15zdnd00an1n02x5 FILLER_142_1712 ();
 b15zdnd11an1n04x5 FILLER_142_1717 ();
 b15zdnd11an1n04x5 FILLER_142_1724 ();
 b15zdnd11an1n04x5 FILLER_142_1731 ();
 b15zdnd11an1n32x5 FILLER_142_1738 ();
 b15zdnd11an1n08x5 FILLER_142_1770 ();
 b15zdnd00an1n01x5 FILLER_142_1778 ();
 b15zdnd11an1n04x5 FILLER_142_1782 ();
 b15zdnd11an1n04x5 FILLER_142_1789 ();
 b15zdnd11an1n64x5 FILLER_142_1796 ();
 b15zdnd11an1n08x5 FILLER_142_1860 ();
 b15zdnd11an1n32x5 FILLER_142_1872 ();
 b15zdnd11an1n16x5 FILLER_142_1904 ();
 b15zdnd11an1n04x5 FILLER_142_1920 ();
 b15zdnd00an1n02x5 FILLER_142_1924 ();
 b15zdnd00an1n01x5 FILLER_142_1926 ();
 b15zdnd11an1n64x5 FILLER_142_1943 ();
 b15zdnd11an1n64x5 FILLER_142_2007 ();
 b15zdnd11an1n64x5 FILLER_142_2071 ();
 b15zdnd11an1n16x5 FILLER_142_2135 ();
 b15zdnd00an1n02x5 FILLER_142_2151 ();
 b15zdnd00an1n01x5 FILLER_142_2153 ();
 b15zdnd00an1n02x5 FILLER_142_2162 ();
 b15zdnd11an1n32x5 FILLER_142_2206 ();
 b15zdnd11an1n16x5 FILLER_142_2238 ();
 b15zdnd11an1n08x5 FILLER_142_2254 ();
 b15zdnd11an1n04x5 FILLER_142_2262 ();
 b15zdnd11an1n04x5 FILLER_142_2270 ();
 b15zdnd00an1n02x5 FILLER_142_2274 ();
 b15zdnd11an1n64x5 FILLER_143_0 ();
 b15zdnd11an1n64x5 FILLER_143_64 ();
 b15zdnd11an1n64x5 FILLER_143_128 ();
 b15zdnd11an1n64x5 FILLER_143_192 ();
 b15zdnd11an1n64x5 FILLER_143_256 ();
 b15zdnd11an1n64x5 FILLER_143_320 ();
 b15zdnd11an1n64x5 FILLER_143_384 ();
 b15zdnd11an1n64x5 FILLER_143_448 ();
 b15zdnd11an1n64x5 FILLER_143_512 ();
 b15zdnd11an1n64x5 FILLER_143_576 ();
 b15zdnd11an1n64x5 FILLER_143_640 ();
 b15zdnd11an1n64x5 FILLER_143_704 ();
 b15zdnd11an1n32x5 FILLER_143_768 ();
 b15zdnd11an1n08x5 FILLER_143_800 ();
 b15zdnd11an1n04x5 FILLER_143_808 ();
 b15zdnd00an1n02x5 FILLER_143_812 ();
 b15zdnd11an1n04x5 FILLER_143_817 ();
 b15zdnd00an1n02x5 FILLER_143_821 ();
 b15zdnd00an1n01x5 FILLER_143_823 ();
 b15zdnd11an1n64x5 FILLER_143_827 ();
 b15zdnd11an1n64x5 FILLER_143_891 ();
 b15zdnd11an1n64x5 FILLER_143_955 ();
 b15zdnd11an1n64x5 FILLER_143_1019 ();
 b15zdnd11an1n16x5 FILLER_143_1083 ();
 b15zdnd11an1n08x5 FILLER_143_1099 ();
 b15zdnd11an1n04x5 FILLER_143_1107 ();
 b15zdnd00an1n02x5 FILLER_143_1111 ();
 b15zdnd11an1n64x5 FILLER_143_1165 ();
 b15zdnd11an1n08x5 FILLER_143_1229 ();
 b15zdnd11an1n04x5 FILLER_143_1237 ();
 b15zdnd00an1n02x5 FILLER_143_1241 ();
 b15zdnd00an1n01x5 FILLER_143_1243 ();
 b15zdnd11an1n64x5 FILLER_143_1247 ();
 b15zdnd11an1n32x5 FILLER_143_1311 ();
 b15zdnd11an1n16x5 FILLER_143_1343 ();
 b15zdnd00an1n02x5 FILLER_143_1359 ();
 b15zdnd11an1n64x5 FILLER_143_1369 ();
 b15zdnd11an1n64x5 FILLER_143_1433 ();
 b15zdnd11an1n64x5 FILLER_143_1497 ();
 b15zdnd11an1n64x5 FILLER_143_1561 ();
 b15zdnd11an1n64x5 FILLER_143_1625 ();
 b15zdnd11an1n64x5 FILLER_143_1689 ();
 b15zdnd11an1n32x5 FILLER_143_1753 ();
 b15zdnd11an1n04x5 FILLER_143_1785 ();
 b15zdnd00an1n01x5 FILLER_143_1789 ();
 b15zdnd11an1n64x5 FILLER_143_1793 ();
 b15zdnd11an1n08x5 FILLER_143_1857 ();
 b15zdnd11an1n04x5 FILLER_143_1865 ();
 b15zdnd00an1n02x5 FILLER_143_1869 ();
 b15zdnd00an1n01x5 FILLER_143_1871 ();
 b15zdnd11an1n64x5 FILLER_143_1876 ();
 b15zdnd11an1n64x5 FILLER_143_1940 ();
 b15zdnd11an1n64x5 FILLER_143_2004 ();
 b15zdnd11an1n64x5 FILLER_143_2068 ();
 b15zdnd11an1n08x5 FILLER_143_2132 ();
 b15zdnd11an1n04x5 FILLER_143_2140 ();
 b15zdnd00an1n02x5 FILLER_143_2144 ();
 b15zdnd11an1n64x5 FILLER_143_2164 ();
 b15zdnd11an1n08x5 FILLER_143_2228 ();
 b15zdnd00an1n02x5 FILLER_143_2236 ();
 b15zdnd11an1n04x5 FILLER_143_2280 ();
 b15zdnd11an1n64x5 FILLER_144_8 ();
 b15zdnd11an1n04x5 FILLER_144_72 ();
 b15zdnd11an1n64x5 FILLER_144_86 ();
 b15zdnd11an1n64x5 FILLER_144_150 ();
 b15zdnd11an1n64x5 FILLER_144_214 ();
 b15zdnd11an1n64x5 FILLER_144_278 ();
 b15zdnd11an1n64x5 FILLER_144_342 ();
 b15zdnd11an1n64x5 FILLER_144_406 ();
 b15zdnd11an1n64x5 FILLER_144_470 ();
 b15zdnd11an1n32x5 FILLER_144_534 ();
 b15zdnd11an1n16x5 FILLER_144_566 ();
 b15zdnd00an1n02x5 FILLER_144_582 ();
 b15zdnd00an1n01x5 FILLER_144_584 ();
 b15zdnd11an1n64x5 FILLER_144_600 ();
 b15zdnd11an1n32x5 FILLER_144_664 ();
 b15zdnd11an1n16x5 FILLER_144_696 ();
 b15zdnd11an1n04x5 FILLER_144_712 ();
 b15zdnd00an1n02x5 FILLER_144_716 ();
 b15zdnd11an1n04x5 FILLER_144_726 ();
 b15zdnd00an1n02x5 FILLER_144_730 ();
 b15zdnd11an1n32x5 FILLER_144_739 ();
 b15zdnd00an1n02x5 FILLER_144_771 ();
 b15zdnd00an1n01x5 FILLER_144_773 ();
 b15zdnd11an1n64x5 FILLER_144_819 ();
 b15zdnd11an1n64x5 FILLER_144_883 ();
 b15zdnd11an1n64x5 FILLER_144_947 ();
 b15zdnd11an1n64x5 FILLER_144_1011 ();
 b15zdnd11an1n16x5 FILLER_144_1075 ();
 b15zdnd11an1n08x5 FILLER_144_1091 ();
 b15zdnd11an1n04x5 FILLER_144_1099 ();
 b15zdnd00an1n02x5 FILLER_144_1103 ();
 b15zdnd00an1n01x5 FILLER_144_1105 ();
 b15zdnd11an1n04x5 FILLER_144_1148 ();
 b15zdnd00an1n02x5 FILLER_144_1152 ();
 b15zdnd11an1n32x5 FILLER_144_1157 ();
 b15zdnd11an1n16x5 FILLER_144_1189 ();
 b15zdnd11an1n08x5 FILLER_144_1205 ();
 b15zdnd11an1n04x5 FILLER_144_1213 ();
 b15zdnd00an1n02x5 FILLER_144_1217 ();
 b15zdnd11an1n64x5 FILLER_144_1271 ();
 b15zdnd11an1n64x5 FILLER_144_1335 ();
 b15zdnd11an1n64x5 FILLER_144_1399 ();
 b15zdnd11an1n64x5 FILLER_144_1463 ();
 b15zdnd11an1n32x5 FILLER_144_1527 ();
 b15zdnd11an1n16x5 FILLER_144_1559 ();
 b15zdnd11an1n08x5 FILLER_144_1575 ();
 b15zdnd11an1n04x5 FILLER_144_1583 ();
 b15zdnd11an1n32x5 FILLER_144_1602 ();
 b15zdnd11an1n16x5 FILLER_144_1634 ();
 b15zdnd11an1n04x5 FILLER_144_1650 ();
 b15zdnd00an1n01x5 FILLER_144_1654 ();
 b15zdnd11an1n64x5 FILLER_144_1663 ();
 b15zdnd11an1n64x5 FILLER_144_1727 ();
 b15zdnd11an1n64x5 FILLER_144_1791 ();
 b15zdnd11an1n64x5 FILLER_144_1855 ();
 b15zdnd11an1n64x5 FILLER_144_1919 ();
 b15zdnd11an1n64x5 FILLER_144_1983 ();
 b15zdnd11an1n64x5 FILLER_144_2047 ();
 b15zdnd11an1n32x5 FILLER_144_2111 ();
 b15zdnd11an1n08x5 FILLER_144_2143 ();
 b15zdnd00an1n02x5 FILLER_144_2151 ();
 b15zdnd00an1n01x5 FILLER_144_2153 ();
 b15zdnd11an1n32x5 FILLER_144_2162 ();
 b15zdnd11an1n16x5 FILLER_144_2194 ();
 b15zdnd11an1n04x5 FILLER_144_2210 ();
 b15zdnd00an1n01x5 FILLER_144_2214 ();
 b15zdnd11an1n04x5 FILLER_144_2257 ();
 b15zdnd11an1n04x5 FILLER_144_2265 ();
 b15zdnd00an1n02x5 FILLER_144_2273 ();
 b15zdnd00an1n01x5 FILLER_144_2275 ();
 b15zdnd11an1n64x5 FILLER_145_0 ();
 b15zdnd11an1n64x5 FILLER_145_64 ();
 b15zdnd11an1n64x5 FILLER_145_128 ();
 b15zdnd11an1n64x5 FILLER_145_192 ();
 b15zdnd11an1n64x5 FILLER_145_256 ();
 b15zdnd11an1n64x5 FILLER_145_320 ();
 b15zdnd11an1n64x5 FILLER_145_384 ();
 b15zdnd11an1n64x5 FILLER_145_448 ();
 b15zdnd11an1n64x5 FILLER_145_512 ();
 b15zdnd11an1n64x5 FILLER_145_576 ();
 b15zdnd11an1n64x5 FILLER_145_640 ();
 b15zdnd11an1n64x5 FILLER_145_704 ();
 b15zdnd11an1n64x5 FILLER_145_768 ();
 b15zdnd11an1n64x5 FILLER_145_832 ();
 b15zdnd11an1n64x5 FILLER_145_896 ();
 b15zdnd11an1n16x5 FILLER_145_960 ();
 b15zdnd00an1n02x5 FILLER_145_976 ();
 b15zdnd11an1n64x5 FILLER_145_986 ();
 b15zdnd11an1n64x5 FILLER_145_1050 ();
 b15zdnd11an1n08x5 FILLER_145_1114 ();
 b15zdnd00an1n01x5 FILLER_145_1122 ();
 b15zdnd11an1n04x5 FILLER_145_1126 ();
 b15zdnd11an1n04x5 FILLER_145_1133 ();
 b15zdnd11an1n04x5 FILLER_145_1140 ();
 b15zdnd00an1n02x5 FILLER_145_1144 ();
 b15zdnd00an1n01x5 FILLER_145_1146 ();
 b15zdnd11an1n64x5 FILLER_145_1150 ();
 b15zdnd00an1n01x5 FILLER_145_1214 ();
 b15zdnd11an1n64x5 FILLER_145_1267 ();
 b15zdnd11an1n16x5 FILLER_145_1331 ();
 b15zdnd11an1n04x5 FILLER_145_1347 ();
 b15zdnd11an1n64x5 FILLER_145_1363 ();
 b15zdnd11an1n64x5 FILLER_145_1427 ();
 b15zdnd11an1n64x5 FILLER_145_1491 ();
 b15zdnd11an1n32x5 FILLER_145_1555 ();
 b15zdnd11an1n16x5 FILLER_145_1587 ();
 b15zdnd11an1n04x5 FILLER_145_1603 ();
 b15zdnd11an1n64x5 FILLER_145_1615 ();
 b15zdnd11an1n32x5 FILLER_145_1679 ();
 b15zdnd11an1n16x5 FILLER_145_1711 ();
 b15zdnd11an1n08x5 FILLER_145_1727 ();
 b15zdnd00an1n02x5 FILLER_145_1735 ();
 b15zdnd00an1n01x5 FILLER_145_1737 ();
 b15zdnd11an1n64x5 FILLER_145_1747 ();
 b15zdnd11an1n64x5 FILLER_145_1811 ();
 b15zdnd11an1n64x5 FILLER_145_1875 ();
 b15zdnd11an1n64x5 FILLER_145_1939 ();
 b15zdnd11an1n32x5 FILLER_145_2003 ();
 b15zdnd11an1n04x5 FILLER_145_2041 ();
 b15zdnd11an1n64x5 FILLER_145_2097 ();
 b15zdnd11an1n64x5 FILLER_145_2161 ();
 b15zdnd11an1n08x5 FILLER_145_2225 ();
 b15zdnd11an1n04x5 FILLER_145_2233 ();
 b15zdnd00an1n02x5 FILLER_145_2237 ();
 b15zdnd00an1n01x5 FILLER_145_2239 ();
 b15zdnd00an1n02x5 FILLER_145_2282 ();
 b15zdnd11an1n16x5 FILLER_146_8 ();
 b15zdnd11an1n04x5 FILLER_146_24 ();
 b15zdnd00an1n02x5 FILLER_146_28 ();
 b15zdnd00an1n01x5 FILLER_146_30 ();
 b15zdnd11an1n64x5 FILLER_146_35 ();
 b15zdnd11an1n64x5 FILLER_146_99 ();
 b15zdnd11an1n64x5 FILLER_146_163 ();
 b15zdnd11an1n64x5 FILLER_146_227 ();
 b15zdnd11an1n64x5 FILLER_146_291 ();
 b15zdnd11an1n64x5 FILLER_146_355 ();
 b15zdnd11an1n64x5 FILLER_146_419 ();
 b15zdnd11an1n64x5 FILLER_146_483 ();
 b15zdnd11an1n64x5 FILLER_146_547 ();
 b15zdnd11an1n64x5 FILLER_146_611 ();
 b15zdnd11an1n32x5 FILLER_146_675 ();
 b15zdnd11an1n08x5 FILLER_146_707 ();
 b15zdnd00an1n02x5 FILLER_146_715 ();
 b15zdnd00an1n01x5 FILLER_146_717 ();
 b15zdnd11an1n64x5 FILLER_146_726 ();
 b15zdnd11an1n64x5 FILLER_146_790 ();
 b15zdnd11an1n64x5 FILLER_146_854 ();
 b15zdnd11an1n64x5 FILLER_146_918 ();
 b15zdnd11an1n64x5 FILLER_146_982 ();
 b15zdnd11an1n64x5 FILLER_146_1046 ();
 b15zdnd11an1n16x5 FILLER_146_1110 ();
 b15zdnd11an1n08x5 FILLER_146_1126 ();
 b15zdnd11an1n04x5 FILLER_146_1134 ();
 b15zdnd00an1n02x5 FILLER_146_1138 ();
 b15zdnd11an1n32x5 FILLER_146_1143 ();
 b15zdnd11an1n16x5 FILLER_146_1175 ();
 b15zdnd11an1n08x5 FILLER_146_1191 ();
 b15zdnd00an1n02x5 FILLER_146_1199 ();
 b15zdnd00an1n01x5 FILLER_146_1201 ();
 b15zdnd11an1n16x5 FILLER_146_1210 ();
 b15zdnd11an1n04x5 FILLER_146_1226 ();
 b15zdnd00an1n02x5 FILLER_146_1230 ();
 b15zdnd00an1n01x5 FILLER_146_1232 ();
 b15zdnd11an1n04x5 FILLER_146_1236 ();
 b15zdnd11an1n04x5 FILLER_146_1243 ();
 b15zdnd11an1n64x5 FILLER_146_1250 ();
 b15zdnd11an1n64x5 FILLER_146_1314 ();
 b15zdnd11an1n32x5 FILLER_146_1378 ();
 b15zdnd11an1n64x5 FILLER_146_1452 ();
 b15zdnd11an1n64x5 FILLER_146_1516 ();
 b15zdnd11an1n64x5 FILLER_146_1580 ();
 b15zdnd11an1n64x5 FILLER_146_1644 ();
 b15zdnd11an1n64x5 FILLER_146_1708 ();
 b15zdnd11an1n64x5 FILLER_146_1772 ();
 b15zdnd11an1n32x5 FILLER_146_1836 ();
 b15zdnd00an1n02x5 FILLER_146_1868 ();
 b15zdnd11an1n32x5 FILLER_146_1881 ();
 b15zdnd11an1n16x5 FILLER_146_1913 ();
 b15zdnd00an1n02x5 FILLER_146_1929 ();
 b15zdnd00an1n01x5 FILLER_146_1931 ();
 b15zdnd11an1n32x5 FILLER_146_1948 ();
 b15zdnd11an1n16x5 FILLER_146_1980 ();
 b15zdnd11an1n08x5 FILLER_146_1996 ();
 b15zdnd00an1n02x5 FILLER_146_2004 ();
 b15zdnd00an1n01x5 FILLER_146_2006 ();
 b15zdnd11an1n32x5 FILLER_146_2024 ();
 b15zdnd11an1n04x5 FILLER_146_2056 ();
 b15zdnd00an1n02x5 FILLER_146_2060 ();
 b15zdnd00an1n01x5 FILLER_146_2062 ();
 b15zdnd11an1n04x5 FILLER_146_2066 ();
 b15zdnd11an1n04x5 FILLER_146_2073 ();
 b15zdnd11an1n64x5 FILLER_146_2080 ();
 b15zdnd11an1n08x5 FILLER_146_2144 ();
 b15zdnd00an1n02x5 FILLER_146_2152 ();
 b15zdnd11an1n64x5 FILLER_146_2162 ();
 b15zdnd11an1n04x5 FILLER_146_2226 ();
 b15zdnd00an1n02x5 FILLER_146_2230 ();
 b15zdnd00an1n02x5 FILLER_146_2274 ();
 b15zdnd11an1n16x5 FILLER_147_0 ();
 b15zdnd00an1n02x5 FILLER_147_16 ();
 b15zdnd00an1n01x5 FILLER_147_18 ();
 b15zdnd11an1n32x5 FILLER_147_23 ();
 b15zdnd11an1n08x5 FILLER_147_55 ();
 b15zdnd11an1n04x5 FILLER_147_63 ();
 b15zdnd00an1n02x5 FILLER_147_67 ();
 b15zdnd11an1n64x5 FILLER_147_89 ();
 b15zdnd11an1n64x5 FILLER_147_153 ();
 b15zdnd11an1n64x5 FILLER_147_217 ();
 b15zdnd11an1n64x5 FILLER_147_281 ();
 b15zdnd11an1n64x5 FILLER_147_345 ();
 b15zdnd11an1n64x5 FILLER_147_409 ();
 b15zdnd11an1n64x5 FILLER_147_473 ();
 b15zdnd11an1n64x5 FILLER_147_537 ();
 b15zdnd11an1n64x5 FILLER_147_601 ();
 b15zdnd11an1n64x5 FILLER_147_665 ();
 b15zdnd11an1n32x5 FILLER_147_729 ();
 b15zdnd00an1n02x5 FILLER_147_761 ();
 b15zdnd00an1n01x5 FILLER_147_763 ();
 b15zdnd11an1n04x5 FILLER_147_767 ();
 b15zdnd11an1n64x5 FILLER_147_781 ();
 b15zdnd11an1n64x5 FILLER_147_845 ();
 b15zdnd11an1n64x5 FILLER_147_909 ();
 b15zdnd11an1n64x5 FILLER_147_973 ();
 b15zdnd11an1n64x5 FILLER_147_1037 ();
 b15zdnd11an1n64x5 FILLER_147_1101 ();
 b15zdnd11an1n64x5 FILLER_147_1165 ();
 b15zdnd11an1n08x5 FILLER_147_1229 ();
 b15zdnd11an1n04x5 FILLER_147_1237 ();
 b15zdnd11an1n04x5 FILLER_147_1244 ();
 b15zdnd11an1n64x5 FILLER_147_1251 ();
 b15zdnd11an1n64x5 FILLER_147_1315 ();
 b15zdnd11an1n16x5 FILLER_147_1379 ();
 b15zdnd00an1n02x5 FILLER_147_1395 ();
 b15zdnd11an1n64x5 FILLER_147_1413 ();
 b15zdnd11an1n32x5 FILLER_147_1477 ();
 b15zdnd11an1n16x5 FILLER_147_1509 ();
 b15zdnd11an1n08x5 FILLER_147_1525 ();
 b15zdnd00an1n02x5 FILLER_147_1533 ();
 b15zdnd00an1n01x5 FILLER_147_1535 ();
 b15zdnd11an1n04x5 FILLER_147_1539 ();
 b15zdnd11an1n04x5 FILLER_147_1546 ();
 b15zdnd11an1n64x5 FILLER_147_1553 ();
 b15zdnd11an1n64x5 FILLER_147_1617 ();
 b15zdnd11an1n64x5 FILLER_147_1681 ();
 b15zdnd11an1n64x5 FILLER_147_1745 ();
 b15zdnd11an1n64x5 FILLER_147_1809 ();
 b15zdnd11an1n64x5 FILLER_147_1873 ();
 b15zdnd11an1n64x5 FILLER_147_1937 ();
 b15zdnd00an1n02x5 FILLER_147_2001 ();
 b15zdnd11an1n64x5 FILLER_147_2048 ();
 b15zdnd11an1n16x5 FILLER_147_2112 ();
 b15zdnd11an1n08x5 FILLER_147_2128 ();
 b15zdnd11an1n04x5 FILLER_147_2136 ();
 b15zdnd00an1n02x5 FILLER_147_2140 ();
 b15zdnd11an1n64x5 FILLER_147_2184 ();
 b15zdnd11an1n32x5 FILLER_147_2248 ();
 b15zdnd11an1n04x5 FILLER_147_2280 ();
 b15zdnd11an1n64x5 FILLER_148_8 ();
 b15zdnd11an1n64x5 FILLER_148_72 ();
 b15zdnd11an1n64x5 FILLER_148_136 ();
 b15zdnd11an1n64x5 FILLER_148_200 ();
 b15zdnd11an1n64x5 FILLER_148_264 ();
 b15zdnd11an1n64x5 FILLER_148_328 ();
 b15zdnd11an1n64x5 FILLER_148_392 ();
 b15zdnd11an1n64x5 FILLER_148_456 ();
 b15zdnd11an1n64x5 FILLER_148_520 ();
 b15zdnd11an1n32x5 FILLER_148_584 ();
 b15zdnd11an1n16x5 FILLER_148_616 ();
 b15zdnd11an1n08x5 FILLER_148_632 ();
 b15zdnd11an1n04x5 FILLER_148_640 ();
 b15zdnd11an1n64x5 FILLER_148_651 ();
 b15zdnd00an1n02x5 FILLER_148_715 ();
 b15zdnd00an1n01x5 FILLER_148_717 ();
 b15zdnd11an1n16x5 FILLER_148_726 ();
 b15zdnd11an1n08x5 FILLER_148_742 ();
 b15zdnd11an1n04x5 FILLER_148_750 ();
 b15zdnd11an1n04x5 FILLER_148_757 ();
 b15zdnd00an1n02x5 FILLER_148_761 ();
 b15zdnd00an1n01x5 FILLER_148_763 ();
 b15zdnd11an1n64x5 FILLER_148_774 ();
 b15zdnd11an1n64x5 FILLER_148_838 ();
 b15zdnd11an1n16x5 FILLER_148_902 ();
 b15zdnd11an1n04x5 FILLER_148_918 ();
 b15zdnd00an1n02x5 FILLER_148_922 ();
 b15zdnd11an1n64x5 FILLER_148_938 ();
 b15zdnd11an1n64x5 FILLER_148_1002 ();
 b15zdnd11an1n64x5 FILLER_148_1066 ();
 b15zdnd11an1n64x5 FILLER_148_1130 ();
 b15zdnd11an1n64x5 FILLER_148_1194 ();
 b15zdnd11an1n64x5 FILLER_148_1258 ();
 b15zdnd11an1n16x5 FILLER_148_1322 ();
 b15zdnd11an1n08x5 FILLER_148_1338 ();
 b15zdnd11an1n04x5 FILLER_148_1346 ();
 b15zdnd00an1n01x5 FILLER_148_1350 ();
 b15zdnd11an1n64x5 FILLER_148_1362 ();
 b15zdnd11an1n64x5 FILLER_148_1426 ();
 b15zdnd11an1n16x5 FILLER_148_1490 ();
 b15zdnd00an1n02x5 FILLER_148_1506 ();
 b15zdnd00an1n01x5 FILLER_148_1508 ();
 b15zdnd11an1n04x5 FILLER_148_1561 ();
 b15zdnd11an1n08x5 FILLER_148_1571 ();
 b15zdnd11an1n04x5 FILLER_148_1579 ();
 b15zdnd11an1n08x5 FILLER_148_1590 ();
 b15zdnd11an1n64x5 FILLER_148_1650 ();
 b15zdnd11an1n64x5 FILLER_148_1714 ();
 b15zdnd11an1n64x5 FILLER_148_1778 ();
 b15zdnd11an1n64x5 FILLER_148_1842 ();
 b15zdnd11an1n64x5 FILLER_148_1906 ();
 b15zdnd11an1n64x5 FILLER_148_1970 ();
 b15zdnd11an1n64x5 FILLER_148_2034 ();
 b15zdnd11an1n32x5 FILLER_148_2098 ();
 b15zdnd11an1n04x5 FILLER_148_2130 ();
 b15zdnd00an1n02x5 FILLER_148_2134 ();
 b15zdnd11an1n04x5 FILLER_148_2150 ();
 b15zdnd11an1n64x5 FILLER_148_2162 ();
 b15zdnd11an1n32x5 FILLER_148_2226 ();
 b15zdnd11an1n16x5 FILLER_148_2258 ();
 b15zdnd00an1n02x5 FILLER_148_2274 ();
 b15zdnd11an1n64x5 FILLER_149_0 ();
 b15zdnd11an1n64x5 FILLER_149_64 ();
 b15zdnd11an1n32x5 FILLER_149_128 ();
 b15zdnd11an1n16x5 FILLER_149_160 ();
 b15zdnd11an1n08x5 FILLER_149_176 ();
 b15zdnd00an1n02x5 FILLER_149_184 ();
 b15zdnd00an1n01x5 FILLER_149_186 ();
 b15zdnd11an1n64x5 FILLER_149_207 ();
 b15zdnd11an1n32x5 FILLER_149_271 ();
 b15zdnd11an1n08x5 FILLER_149_303 ();
 b15zdnd11an1n04x5 FILLER_149_311 ();
 b15zdnd00an1n02x5 FILLER_149_315 ();
 b15zdnd11an1n32x5 FILLER_149_320 ();
 b15zdnd11an1n16x5 FILLER_149_352 ();
 b15zdnd11an1n04x5 FILLER_149_368 ();
 b15zdnd00an1n01x5 FILLER_149_372 ();
 b15zdnd11an1n64x5 FILLER_149_409 ();
 b15zdnd11an1n64x5 FILLER_149_473 ();
 b15zdnd11an1n64x5 FILLER_149_537 ();
 b15zdnd11an1n64x5 FILLER_149_601 ();
 b15zdnd11an1n64x5 FILLER_149_665 ();
 b15zdnd11an1n16x5 FILLER_149_729 ();
 b15zdnd11an1n08x5 FILLER_149_745 ();
 b15zdnd00an1n01x5 FILLER_149_753 ();
 b15zdnd11an1n08x5 FILLER_149_761 ();
 b15zdnd11an1n04x5 FILLER_149_769 ();
 b15zdnd11an1n64x5 FILLER_149_789 ();
 b15zdnd11an1n16x5 FILLER_149_853 ();
 b15zdnd11an1n04x5 FILLER_149_869 ();
 b15zdnd00an1n02x5 FILLER_149_873 ();
 b15zdnd11an1n32x5 FILLER_149_878 ();
 b15zdnd11an1n16x5 FILLER_149_910 ();
 b15zdnd11an1n04x5 FILLER_149_926 ();
 b15zdnd00an1n02x5 FILLER_149_930 ();
 b15zdnd11an1n64x5 FILLER_149_946 ();
 b15zdnd11an1n64x5 FILLER_149_1010 ();
 b15zdnd11an1n64x5 FILLER_149_1074 ();
 b15zdnd11an1n16x5 FILLER_149_1138 ();
 b15zdnd00an1n01x5 FILLER_149_1154 ();
 b15zdnd11an1n32x5 FILLER_149_1164 ();
 b15zdnd11an1n08x5 FILLER_149_1196 ();
 b15zdnd11an1n04x5 FILLER_149_1204 ();
 b15zdnd00an1n02x5 FILLER_149_1208 ();
 b15zdnd11an1n64x5 FILLER_149_1219 ();
 b15zdnd11an1n64x5 FILLER_149_1283 ();
 b15zdnd11an1n64x5 FILLER_149_1347 ();
 b15zdnd11an1n16x5 FILLER_149_1411 ();
 b15zdnd11an1n64x5 FILLER_149_1430 ();
 b15zdnd11an1n16x5 FILLER_149_1494 ();
 b15zdnd11an1n08x5 FILLER_149_1510 ();
 b15zdnd00an1n01x5 FILLER_149_1518 ();
 b15zdnd11an1n04x5 FILLER_149_1522 ();
 b15zdnd11an1n32x5 FILLER_149_1578 ();
 b15zdnd11an1n04x5 FILLER_149_1610 ();
 b15zdnd00an1n02x5 FILLER_149_1614 ();
 b15zdnd11an1n04x5 FILLER_149_1619 ();
 b15zdnd11an1n08x5 FILLER_149_1626 ();
 b15zdnd00an1n02x5 FILLER_149_1634 ();
 b15zdnd00an1n01x5 FILLER_149_1636 ();
 b15zdnd11an1n64x5 FILLER_149_1644 ();
 b15zdnd11an1n64x5 FILLER_149_1708 ();
 b15zdnd11an1n64x5 FILLER_149_1772 ();
 b15zdnd11an1n64x5 FILLER_149_1836 ();
 b15zdnd11an1n64x5 FILLER_149_1900 ();
 b15zdnd11an1n64x5 FILLER_149_1964 ();
 b15zdnd11an1n64x5 FILLER_149_2028 ();
 b15zdnd11an1n32x5 FILLER_149_2092 ();
 b15zdnd00an1n01x5 FILLER_149_2124 ();
 b15zdnd11an1n32x5 FILLER_149_2167 ();
 b15zdnd11an1n08x5 FILLER_149_2199 ();
 b15zdnd00an1n01x5 FILLER_149_2207 ();
 b15zdnd11an1n32x5 FILLER_149_2225 ();
 b15zdnd11an1n16x5 FILLER_149_2257 ();
 b15zdnd11an1n08x5 FILLER_149_2273 ();
 b15zdnd00an1n02x5 FILLER_149_2281 ();
 b15zdnd00an1n01x5 FILLER_149_2283 ();
 b15zdnd11an1n64x5 FILLER_150_8 ();
 b15zdnd11an1n64x5 FILLER_150_72 ();
 b15zdnd11an1n08x5 FILLER_150_136 ();
 b15zdnd11an1n04x5 FILLER_150_144 ();
 b15zdnd00an1n01x5 FILLER_150_148 ();
 b15zdnd11an1n04x5 FILLER_150_164 ();
 b15zdnd11an1n64x5 FILLER_150_208 ();
 b15zdnd11an1n16x5 FILLER_150_272 ();
 b15zdnd00an1n02x5 FILLER_150_288 ();
 b15zdnd11an1n64x5 FILLER_150_342 ();
 b15zdnd11an1n08x5 FILLER_150_406 ();
 b15zdnd11an1n04x5 FILLER_150_414 ();
 b15zdnd00an1n02x5 FILLER_150_418 ();
 b15zdnd00an1n01x5 FILLER_150_420 ();
 b15zdnd11an1n64x5 FILLER_150_463 ();
 b15zdnd11an1n64x5 FILLER_150_527 ();
 b15zdnd11an1n64x5 FILLER_150_591 ();
 b15zdnd11an1n32x5 FILLER_150_655 ();
 b15zdnd11an1n16x5 FILLER_150_687 ();
 b15zdnd11an1n08x5 FILLER_150_703 ();
 b15zdnd11an1n04x5 FILLER_150_711 ();
 b15zdnd00an1n02x5 FILLER_150_715 ();
 b15zdnd00an1n01x5 FILLER_150_717 ();
 b15zdnd11an1n16x5 FILLER_150_726 ();
 b15zdnd11an1n08x5 FILLER_150_742 ();
 b15zdnd00an1n01x5 FILLER_150_750 ();
 b15zdnd11an1n64x5 FILLER_150_775 ();
 b15zdnd11an1n64x5 FILLER_150_839 ();
 b15zdnd11an1n16x5 FILLER_150_903 ();
 b15zdnd00an1n02x5 FILLER_150_919 ();
 b15zdnd00an1n01x5 FILLER_150_921 ();
 b15zdnd11an1n04x5 FILLER_150_948 ();
 b15zdnd11an1n04x5 FILLER_150_963 ();
 b15zdnd00an1n02x5 FILLER_150_967 ();
 b15zdnd00an1n01x5 FILLER_150_969 ();
 b15zdnd11an1n32x5 FILLER_150_984 ();
 b15zdnd11an1n08x5 FILLER_150_1016 ();
 b15zdnd11an1n04x5 FILLER_150_1024 ();
 b15zdnd00an1n01x5 FILLER_150_1028 ();
 b15zdnd11an1n64x5 FILLER_150_1037 ();
 b15zdnd11an1n64x5 FILLER_150_1101 ();
 b15zdnd11an1n64x5 FILLER_150_1165 ();
 b15zdnd11an1n64x5 FILLER_150_1229 ();
 b15zdnd11an1n64x5 FILLER_150_1293 ();
 b15zdnd11an1n32x5 FILLER_150_1357 ();
 b15zdnd11an1n08x5 FILLER_150_1389 ();
 b15zdnd11an1n04x5 FILLER_150_1449 ();
 b15zdnd11an1n04x5 FILLER_150_1460 ();
 b15zdnd11an1n32x5 FILLER_150_1472 ();
 b15zdnd11an1n16x5 FILLER_150_1504 ();
 b15zdnd11an1n04x5 FILLER_150_1520 ();
 b15zdnd00an1n02x5 FILLER_150_1524 ();
 b15zdnd00an1n01x5 FILLER_150_1526 ();
 b15zdnd11an1n04x5 FILLER_150_1530 ();
 b15zdnd11an1n08x5 FILLER_150_1537 ();
 b15zdnd00an1n02x5 FILLER_150_1545 ();
 b15zdnd00an1n01x5 FILLER_150_1547 ();
 b15zdnd11an1n32x5 FILLER_150_1551 ();
 b15zdnd11an1n16x5 FILLER_150_1583 ();
 b15zdnd11an1n08x5 FILLER_150_1599 ();
 b15zdnd11an1n04x5 FILLER_150_1616 ();
 b15zdnd00an1n01x5 FILLER_150_1620 ();
 b15zdnd11an1n64x5 FILLER_150_1624 ();
 b15zdnd11an1n64x5 FILLER_150_1688 ();
 b15zdnd11an1n64x5 FILLER_150_1752 ();
 b15zdnd11an1n64x5 FILLER_150_1816 ();
 b15zdnd11an1n64x5 FILLER_150_1880 ();
 b15zdnd11an1n64x5 FILLER_150_1944 ();
 b15zdnd11an1n64x5 FILLER_150_2008 ();
 b15zdnd11an1n64x5 FILLER_150_2072 ();
 b15zdnd11an1n16x5 FILLER_150_2136 ();
 b15zdnd00an1n02x5 FILLER_150_2152 ();
 b15zdnd11an1n32x5 FILLER_150_2162 ();
 b15zdnd11an1n08x5 FILLER_150_2194 ();
 b15zdnd11an1n32x5 FILLER_150_2216 ();
 b15zdnd11an1n16x5 FILLER_150_2248 ();
 b15zdnd11an1n08x5 FILLER_150_2264 ();
 b15zdnd11an1n04x5 FILLER_150_2272 ();
 b15zdnd11an1n32x5 FILLER_151_0 ();
 b15zdnd00an1n02x5 FILLER_151_32 ();
 b15zdnd00an1n01x5 FILLER_151_34 ();
 b15zdnd11an1n32x5 FILLER_151_39 ();
 b15zdnd11an1n08x5 FILLER_151_71 ();
 b15zdnd11an1n04x5 FILLER_151_79 ();
 b15zdnd00an1n02x5 FILLER_151_83 ();
 b15zdnd11an1n04x5 FILLER_151_92 ();
 b15zdnd11an1n32x5 FILLER_151_104 ();
 b15zdnd11an1n04x5 FILLER_151_136 ();
 b15zdnd00an1n01x5 FILLER_151_140 ();
 b15zdnd11an1n16x5 FILLER_151_183 ();
 b15zdnd11an1n04x5 FILLER_151_202 ();
 b15zdnd11an1n64x5 FILLER_151_209 ();
 b15zdnd11an1n32x5 FILLER_151_273 ();
 b15zdnd00an1n02x5 FILLER_151_305 ();
 b15zdnd00an1n01x5 FILLER_151_307 ();
 b15zdnd11an1n04x5 FILLER_151_311 ();
 b15zdnd11an1n64x5 FILLER_151_318 ();
 b15zdnd11an1n64x5 FILLER_151_382 ();
 b15zdnd11an1n64x5 FILLER_151_446 ();
 b15zdnd11an1n64x5 FILLER_151_510 ();
 b15zdnd11an1n64x5 FILLER_151_574 ();
 b15zdnd11an1n64x5 FILLER_151_638 ();
 b15zdnd11an1n64x5 FILLER_151_702 ();
 b15zdnd11an1n32x5 FILLER_151_808 ();
 b15zdnd11an1n16x5 FILLER_151_840 ();
 b15zdnd11an1n08x5 FILLER_151_856 ();
 b15zdnd11an1n04x5 FILLER_151_864 ();
 b15zdnd00an1n01x5 FILLER_151_868 ();
 b15zdnd11an1n16x5 FILLER_151_883 ();
 b15zdnd11an1n08x5 FILLER_151_899 ();
 b15zdnd11an1n04x5 FILLER_151_907 ();
 b15zdnd00an1n02x5 FILLER_151_911 ();
 b15zdnd00an1n01x5 FILLER_151_913 ();
 b15zdnd11an1n08x5 FILLER_151_934 ();
 b15zdnd11an1n04x5 FILLER_151_942 ();
 b15zdnd00an1n02x5 FILLER_151_946 ();
 b15zdnd11an1n64x5 FILLER_151_962 ();
 b15zdnd11an1n16x5 FILLER_151_1026 ();
 b15zdnd11an1n04x5 FILLER_151_1042 ();
 b15zdnd00an1n02x5 FILLER_151_1046 ();
 b15zdnd00an1n01x5 FILLER_151_1048 ();
 b15zdnd11an1n64x5 FILLER_151_1070 ();
 b15zdnd11an1n64x5 FILLER_151_1134 ();
 b15zdnd11an1n64x5 FILLER_151_1207 ();
 b15zdnd11an1n64x5 FILLER_151_1271 ();
 b15zdnd11an1n64x5 FILLER_151_1335 ();
 b15zdnd00an1n02x5 FILLER_151_1399 ();
 b15zdnd11an1n32x5 FILLER_151_1453 ();
 b15zdnd11an1n08x5 FILLER_151_1485 ();
 b15zdnd11an1n04x5 FILLER_151_1493 ();
 b15zdnd00an1n01x5 FILLER_151_1497 ();
 b15zdnd11an1n04x5 FILLER_151_1509 ();
 b15zdnd11an1n16x5 FILLER_151_1565 ();
 b15zdnd11an1n08x5 FILLER_151_1581 ();
 b15zdnd00an1n02x5 FILLER_151_1589 ();
 b15zdnd11an1n64x5 FILLER_151_1602 ();
 b15zdnd11an1n64x5 FILLER_151_1666 ();
 b15zdnd11an1n64x5 FILLER_151_1730 ();
 b15zdnd11an1n64x5 FILLER_151_1794 ();
 b15zdnd11an1n64x5 FILLER_151_1858 ();
 b15zdnd11an1n64x5 FILLER_151_1922 ();
 b15zdnd11an1n16x5 FILLER_151_1986 ();
 b15zdnd11an1n08x5 FILLER_151_2002 ();
 b15zdnd00an1n02x5 FILLER_151_2010 ();
 b15zdnd00an1n01x5 FILLER_151_2012 ();
 b15zdnd11an1n64x5 FILLER_151_2016 ();
 b15zdnd11an1n16x5 FILLER_151_2080 ();
 b15zdnd11an1n08x5 FILLER_151_2096 ();
 b15zdnd11an1n04x5 FILLER_151_2104 ();
 b15zdnd00an1n02x5 FILLER_151_2108 ();
 b15zdnd11an1n04x5 FILLER_151_2122 ();
 b15zdnd11an1n64x5 FILLER_151_2140 ();
 b15zdnd11an1n64x5 FILLER_151_2204 ();
 b15zdnd11an1n16x5 FILLER_151_2268 ();
 b15zdnd00an1n02x5 FILLER_152_8 ();
 b15zdnd11an1n64x5 FILLER_152_52 ();
 b15zdnd11an1n64x5 FILLER_152_116 ();
 b15zdnd11an1n64x5 FILLER_152_222 ();
 b15zdnd00an1n02x5 FILLER_152_286 ();
 b15zdnd00an1n01x5 FILLER_152_288 ();
 b15zdnd11an1n64x5 FILLER_152_331 ();
 b15zdnd11an1n64x5 FILLER_152_395 ();
 b15zdnd11an1n64x5 FILLER_152_459 ();
 b15zdnd11an1n64x5 FILLER_152_523 ();
 b15zdnd11an1n64x5 FILLER_152_587 ();
 b15zdnd11an1n64x5 FILLER_152_651 ();
 b15zdnd00an1n02x5 FILLER_152_715 ();
 b15zdnd00an1n01x5 FILLER_152_717 ();
 b15zdnd11an1n16x5 FILLER_152_726 ();
 b15zdnd11an1n04x5 FILLER_152_742 ();
 b15zdnd00an1n02x5 FILLER_152_746 ();
 b15zdnd11an1n64x5 FILLER_152_751 ();
 b15zdnd11an1n32x5 FILLER_152_815 ();
 b15zdnd11an1n16x5 FILLER_152_847 ();
 b15zdnd11an1n08x5 FILLER_152_863 ();
 b15zdnd11an1n04x5 FILLER_152_885 ();
 b15zdnd00an1n02x5 FILLER_152_889 ();
 b15zdnd00an1n01x5 FILLER_152_891 ();
 b15zdnd11an1n04x5 FILLER_152_899 ();
 b15zdnd11an1n08x5 FILLER_152_908 ();
 b15zdnd11an1n04x5 FILLER_152_916 ();
 b15zdnd11an1n08x5 FILLER_152_934 ();
 b15zdnd11an1n04x5 FILLER_152_942 ();
 b15zdnd00an1n02x5 FILLER_152_946 ();
 b15zdnd11an1n64x5 FILLER_152_962 ();
 b15zdnd11an1n32x5 FILLER_152_1026 ();
 b15zdnd11an1n16x5 FILLER_152_1058 ();
 b15zdnd00an1n01x5 FILLER_152_1074 ();
 b15zdnd11an1n64x5 FILLER_152_1083 ();
 b15zdnd11an1n64x5 FILLER_152_1147 ();
 b15zdnd11an1n64x5 FILLER_152_1211 ();
 b15zdnd11an1n64x5 FILLER_152_1275 ();
 b15zdnd11an1n64x5 FILLER_152_1339 ();
 b15zdnd11an1n04x5 FILLER_152_1410 ();
 b15zdnd00an1n02x5 FILLER_152_1414 ();
 b15zdnd11an1n04x5 FILLER_152_1419 ();
 b15zdnd11an1n04x5 FILLER_152_1426 ();
 b15zdnd11an1n08x5 FILLER_152_1433 ();
 b15zdnd00an1n02x5 FILLER_152_1441 ();
 b15zdnd11an1n32x5 FILLER_152_1485 ();
 b15zdnd11an1n08x5 FILLER_152_1517 ();
 b15zdnd11an1n04x5 FILLER_152_1525 ();
 b15zdnd00an1n02x5 FILLER_152_1529 ();
 b15zdnd11an1n04x5 FILLER_152_1534 ();
 b15zdnd11an1n64x5 FILLER_152_1541 ();
 b15zdnd11an1n64x5 FILLER_152_1605 ();
 b15zdnd11an1n64x5 FILLER_152_1669 ();
 b15zdnd11an1n64x5 FILLER_152_1733 ();
 b15zdnd11an1n64x5 FILLER_152_1797 ();
 b15zdnd11an1n64x5 FILLER_152_1861 ();
 b15zdnd11an1n32x5 FILLER_152_1925 ();
 b15zdnd11an1n16x5 FILLER_152_1957 ();
 b15zdnd11an1n08x5 FILLER_152_1973 ();
 b15zdnd11an1n04x5 FILLER_152_1981 ();
 b15zdnd00an1n02x5 FILLER_152_1985 ();
 b15zdnd11an1n08x5 FILLER_152_2039 ();
 b15zdnd00an1n02x5 FILLER_152_2047 ();
 b15zdnd00an1n01x5 FILLER_152_2049 ();
 b15zdnd11an1n08x5 FILLER_152_2077 ();
 b15zdnd11an1n04x5 FILLER_152_2085 ();
 b15zdnd00an1n02x5 FILLER_152_2089 ();
 b15zdnd00an1n01x5 FILLER_152_2091 ();
 b15zdnd11an1n16x5 FILLER_152_2134 ();
 b15zdnd11an1n04x5 FILLER_152_2150 ();
 b15zdnd11an1n64x5 FILLER_152_2162 ();
 b15zdnd11an1n32x5 FILLER_152_2226 ();
 b15zdnd11an1n16x5 FILLER_152_2258 ();
 b15zdnd00an1n02x5 FILLER_152_2274 ();
 b15zdnd11an1n08x5 FILLER_153_0 ();
 b15zdnd11an1n04x5 FILLER_153_8 ();
 b15zdnd00an1n01x5 FILLER_153_12 ();
 b15zdnd11an1n64x5 FILLER_153_55 ();
 b15zdnd11an1n64x5 FILLER_153_119 ();
 b15zdnd11an1n64x5 FILLER_153_191 ();
 b15zdnd11an1n16x5 FILLER_153_255 ();
 b15zdnd00an1n02x5 FILLER_153_271 ();
 b15zdnd00an1n01x5 FILLER_153_273 ();
 b15zdnd11an1n64x5 FILLER_153_292 ();
 b15zdnd11an1n64x5 FILLER_153_356 ();
 b15zdnd11an1n64x5 FILLER_153_420 ();
 b15zdnd11an1n08x5 FILLER_153_484 ();
 b15zdnd11an1n64x5 FILLER_153_513 ();
 b15zdnd11an1n08x5 FILLER_153_577 ();
 b15zdnd11an1n04x5 FILLER_153_585 ();
 b15zdnd11an1n04x5 FILLER_153_617 ();
 b15zdnd11an1n64x5 FILLER_153_624 ();
 b15zdnd11an1n32x5 FILLER_153_688 ();
 b15zdnd11an1n04x5 FILLER_153_720 ();
 b15zdnd11an1n64x5 FILLER_153_768 ();
 b15zdnd11an1n32x5 FILLER_153_832 ();
 b15zdnd11an1n16x5 FILLER_153_864 ();
 b15zdnd00an1n01x5 FILLER_153_880 ();
 b15zdnd11an1n08x5 FILLER_153_926 ();
 b15zdnd11an1n04x5 FILLER_153_934 ();
 b15zdnd11an1n64x5 FILLER_153_944 ();
 b15zdnd11an1n32x5 FILLER_153_1008 ();
 b15zdnd11an1n04x5 FILLER_153_1040 ();
 b15zdnd00an1n02x5 FILLER_153_1044 ();
 b15zdnd00an1n01x5 FILLER_153_1046 ();
 b15zdnd11an1n64x5 FILLER_153_1056 ();
 b15zdnd11an1n64x5 FILLER_153_1120 ();
 b15zdnd11an1n64x5 FILLER_153_1184 ();
 b15zdnd11an1n64x5 FILLER_153_1248 ();
 b15zdnd11an1n64x5 FILLER_153_1312 ();
 b15zdnd11an1n32x5 FILLER_153_1376 ();
 b15zdnd11an1n08x5 FILLER_153_1408 ();
 b15zdnd00an1n01x5 FILLER_153_1416 ();
 b15zdnd11an1n04x5 FILLER_153_1420 ();
 b15zdnd11an1n08x5 FILLER_153_1427 ();
 b15zdnd00an1n02x5 FILLER_153_1435 ();
 b15zdnd11an1n64x5 FILLER_153_1444 ();
 b15zdnd11an1n64x5 FILLER_153_1508 ();
 b15zdnd11an1n64x5 FILLER_153_1572 ();
 b15zdnd11an1n64x5 FILLER_153_1636 ();
 b15zdnd11an1n32x5 FILLER_153_1700 ();
 b15zdnd11an1n04x5 FILLER_153_1732 ();
 b15zdnd00an1n02x5 FILLER_153_1736 ();
 b15zdnd11an1n16x5 FILLER_153_1747 ();
 b15zdnd00an1n01x5 FILLER_153_1763 ();
 b15zdnd11an1n64x5 FILLER_153_1773 ();
 b15zdnd11an1n64x5 FILLER_153_1837 ();
 b15zdnd11an1n32x5 FILLER_153_1901 ();
 b15zdnd11an1n16x5 FILLER_153_1933 ();
 b15zdnd11an1n08x5 FILLER_153_1949 ();
 b15zdnd11an1n04x5 FILLER_153_1957 ();
 b15zdnd00an1n02x5 FILLER_153_1961 ();
 b15zdnd00an1n01x5 FILLER_153_1963 ();
 b15zdnd11an1n16x5 FILLER_153_1988 ();
 b15zdnd00an1n01x5 FILLER_153_2004 ();
 b15zdnd11an1n04x5 FILLER_153_2008 ();
 b15zdnd11an1n32x5 FILLER_153_2015 ();
 b15zdnd00an1n02x5 FILLER_153_2047 ();
 b15zdnd11an1n64x5 FILLER_153_2052 ();
 b15zdnd11an1n64x5 FILLER_153_2116 ();
 b15zdnd11an1n64x5 FILLER_153_2180 ();
 b15zdnd11an1n32x5 FILLER_153_2244 ();
 b15zdnd11an1n08x5 FILLER_153_2276 ();
 b15zdnd00an1n02x5 FILLER_154_8 ();
 b15zdnd11an1n08x5 FILLER_154_15 ();
 b15zdnd11an1n04x5 FILLER_154_23 ();
 b15zdnd11an1n32x5 FILLER_154_31 ();
 b15zdnd11an1n08x5 FILLER_154_63 ();
 b15zdnd00an1n02x5 FILLER_154_71 ();
 b15zdnd11an1n64x5 FILLER_154_90 ();
 b15zdnd11an1n32x5 FILLER_154_154 ();
 b15zdnd11an1n08x5 FILLER_154_186 ();
 b15zdnd00an1n01x5 FILLER_154_194 ();
 b15zdnd11an1n32x5 FILLER_154_222 ();
 b15zdnd11an1n08x5 FILLER_154_254 ();
 b15zdnd11an1n04x5 FILLER_154_262 ();
 b15zdnd00an1n02x5 FILLER_154_266 ();
 b15zdnd00an1n01x5 FILLER_154_268 ();
 b15zdnd11an1n64x5 FILLER_154_283 ();
 b15zdnd11an1n64x5 FILLER_154_347 ();
 b15zdnd11an1n64x5 FILLER_154_411 ();
 b15zdnd11an1n32x5 FILLER_154_475 ();
 b15zdnd00an1n02x5 FILLER_154_507 ();
 b15zdnd00an1n01x5 FILLER_154_509 ();
 b15zdnd11an1n64x5 FILLER_154_517 ();
 b15zdnd11an1n16x5 FILLER_154_581 ();
 b15zdnd11an1n08x5 FILLER_154_597 ();
 b15zdnd00an1n02x5 FILLER_154_605 ();
 b15zdnd11an1n16x5 FILLER_154_610 ();
 b15zdnd11an1n08x5 FILLER_154_626 ();
 b15zdnd00an1n02x5 FILLER_154_634 ();
 b15zdnd00an1n01x5 FILLER_154_636 ();
 b15zdnd11an1n64x5 FILLER_154_648 ();
 b15zdnd11an1n04x5 FILLER_154_712 ();
 b15zdnd00an1n02x5 FILLER_154_716 ();
 b15zdnd11an1n08x5 FILLER_154_726 ();
 b15zdnd11an1n04x5 FILLER_154_734 ();
 b15zdnd00an1n02x5 FILLER_154_738 ();
 b15zdnd11an1n04x5 FILLER_154_743 ();
 b15zdnd11an1n64x5 FILLER_154_750 ();
 b15zdnd11an1n64x5 FILLER_154_814 ();
 b15zdnd11an1n32x5 FILLER_154_878 ();
 b15zdnd11an1n08x5 FILLER_154_910 ();
 b15zdnd11an1n04x5 FILLER_154_918 ();
 b15zdnd00an1n02x5 FILLER_154_922 ();
 b15zdnd11an1n64x5 FILLER_154_931 ();
 b15zdnd11an1n64x5 FILLER_154_995 ();
 b15zdnd11an1n04x5 FILLER_154_1059 ();
 b15zdnd11an1n64x5 FILLER_154_1073 ();
 b15zdnd11an1n64x5 FILLER_154_1137 ();
 b15zdnd11an1n64x5 FILLER_154_1201 ();
 b15zdnd11an1n64x5 FILLER_154_1265 ();
 b15zdnd11an1n64x5 FILLER_154_1329 ();
 b15zdnd11an1n64x5 FILLER_154_1393 ();
 b15zdnd00an1n02x5 FILLER_154_1457 ();
 b15zdnd00an1n01x5 FILLER_154_1459 ();
 b15zdnd11an1n32x5 FILLER_154_1469 ();
 b15zdnd11an1n08x5 FILLER_154_1501 ();
 b15zdnd11an1n04x5 FILLER_154_1509 ();
 b15zdnd00an1n02x5 FILLER_154_1513 ();
 b15zdnd00an1n01x5 FILLER_154_1515 ();
 b15zdnd11an1n64x5 FILLER_154_1525 ();
 b15zdnd11an1n64x5 FILLER_154_1589 ();
 b15zdnd11an1n64x5 FILLER_154_1653 ();
 b15zdnd11an1n16x5 FILLER_154_1717 ();
 b15zdnd11an1n08x5 FILLER_154_1733 ();
 b15zdnd00an1n02x5 FILLER_154_1741 ();
 b15zdnd11an1n64x5 FILLER_154_1770 ();
 b15zdnd11an1n32x5 FILLER_154_1834 ();
 b15zdnd11an1n08x5 FILLER_154_1866 ();
 b15zdnd00an1n02x5 FILLER_154_1874 ();
 b15zdnd00an1n01x5 FILLER_154_1876 ();
 b15zdnd11an1n64x5 FILLER_154_1919 ();
 b15zdnd11an1n64x5 FILLER_154_1983 ();
 b15zdnd11an1n64x5 FILLER_154_2047 ();
 b15zdnd11an1n32x5 FILLER_154_2111 ();
 b15zdnd11an1n08x5 FILLER_154_2143 ();
 b15zdnd00an1n02x5 FILLER_154_2151 ();
 b15zdnd00an1n01x5 FILLER_154_2153 ();
 b15zdnd11an1n64x5 FILLER_154_2162 ();
 b15zdnd11an1n32x5 FILLER_154_2226 ();
 b15zdnd11an1n16x5 FILLER_154_2258 ();
 b15zdnd00an1n02x5 FILLER_154_2274 ();
 b15zdnd11an1n64x5 FILLER_155_0 ();
 b15zdnd11an1n04x5 FILLER_155_64 ();
 b15zdnd11an1n64x5 FILLER_155_93 ();
 b15zdnd11an1n32x5 FILLER_155_157 ();
 b15zdnd11an1n08x5 FILLER_155_189 ();
 b15zdnd11an1n32x5 FILLER_155_201 ();
 b15zdnd11an1n16x5 FILLER_155_233 ();
 b15zdnd11an1n08x5 FILLER_155_249 ();
 b15zdnd11an1n04x5 FILLER_155_257 ();
 b15zdnd00an1n01x5 FILLER_155_261 ();
 b15zdnd11an1n64x5 FILLER_155_270 ();
 b15zdnd11an1n64x5 FILLER_155_334 ();
 b15zdnd11an1n64x5 FILLER_155_398 ();
 b15zdnd11an1n16x5 FILLER_155_462 ();
 b15zdnd11an1n08x5 FILLER_155_478 ();
 b15zdnd00an1n02x5 FILLER_155_486 ();
 b15zdnd00an1n01x5 FILLER_155_488 ();
 b15zdnd11an1n04x5 FILLER_155_496 ();
 b15zdnd11an1n64x5 FILLER_155_536 ();
 b15zdnd11an1n16x5 FILLER_155_600 ();
 b15zdnd11an1n08x5 FILLER_155_616 ();
 b15zdnd11an1n04x5 FILLER_155_624 ();
 b15zdnd00an1n02x5 FILLER_155_628 ();
 b15zdnd00an1n01x5 FILLER_155_630 ();
 b15zdnd11an1n04x5 FILLER_155_673 ();
 b15zdnd11an1n64x5 FILLER_155_691 ();
 b15zdnd11an1n64x5 FILLER_155_755 ();
 b15zdnd11an1n32x5 FILLER_155_819 ();
 b15zdnd11an1n04x5 FILLER_155_851 ();
 b15zdnd00an1n02x5 FILLER_155_855 ();
 b15zdnd00an1n01x5 FILLER_155_857 ();
 b15zdnd11an1n64x5 FILLER_155_872 ();
 b15zdnd11an1n32x5 FILLER_155_936 ();
 b15zdnd11an1n16x5 FILLER_155_968 ();
 b15zdnd11an1n08x5 FILLER_155_984 ();
 b15zdnd00an1n02x5 FILLER_155_992 ();
 b15zdnd00an1n01x5 FILLER_155_994 ();
 b15zdnd11an1n64x5 FILLER_155_1007 ();
 b15zdnd11an1n64x5 FILLER_155_1071 ();
 b15zdnd11an1n64x5 FILLER_155_1135 ();
 b15zdnd11an1n64x5 FILLER_155_1199 ();
 b15zdnd11an1n64x5 FILLER_155_1263 ();
 b15zdnd11an1n64x5 FILLER_155_1327 ();
 b15zdnd11an1n64x5 FILLER_155_1391 ();
 b15zdnd11an1n64x5 FILLER_155_1455 ();
 b15zdnd11an1n64x5 FILLER_155_1519 ();
 b15zdnd11an1n64x5 FILLER_155_1583 ();
 b15zdnd11an1n64x5 FILLER_155_1647 ();
 b15zdnd11an1n04x5 FILLER_155_1711 ();
 b15zdnd00an1n01x5 FILLER_155_1715 ();
 b15zdnd11an1n16x5 FILLER_155_1724 ();
 b15zdnd00an1n02x5 FILLER_155_1740 ();
 b15zdnd00an1n01x5 FILLER_155_1742 ();
 b15zdnd11an1n64x5 FILLER_155_1746 ();
 b15zdnd11an1n64x5 FILLER_155_1810 ();
 b15zdnd11an1n64x5 FILLER_155_1874 ();
 b15zdnd11an1n32x5 FILLER_155_1938 ();
 b15zdnd11an1n08x5 FILLER_155_1970 ();
 b15zdnd00an1n01x5 FILLER_155_1978 ();
 b15zdnd11an1n04x5 FILLER_155_1999 ();
 b15zdnd00an1n02x5 FILLER_155_2003 ();
 b15zdnd11an1n08x5 FILLER_155_2025 ();
 b15zdnd11an1n04x5 FILLER_155_2053 ();
 b15zdnd11an1n64x5 FILLER_155_2064 ();
 b15zdnd11an1n64x5 FILLER_155_2128 ();
 b15zdnd11an1n16x5 FILLER_155_2192 ();
 b15zdnd11an1n08x5 FILLER_155_2208 ();
 b15zdnd11an1n04x5 FILLER_155_2216 ();
 b15zdnd11an1n16x5 FILLER_155_2226 ();
 b15zdnd00an1n02x5 FILLER_155_2242 ();
 b15zdnd11an1n32x5 FILLER_155_2248 ();
 b15zdnd11an1n04x5 FILLER_155_2280 ();
 b15zdnd11an1n32x5 FILLER_156_8 ();
 b15zdnd11an1n16x5 FILLER_156_40 ();
 b15zdnd11an1n08x5 FILLER_156_56 ();
 b15zdnd11an1n04x5 FILLER_156_64 ();
 b15zdnd11an1n64x5 FILLER_156_99 ();
 b15zdnd11an1n64x5 FILLER_156_163 ();
 b15zdnd11an1n16x5 FILLER_156_227 ();
 b15zdnd11an1n08x5 FILLER_156_243 ();
 b15zdnd00an1n02x5 FILLER_156_251 ();
 b15zdnd00an1n01x5 FILLER_156_253 ();
 b15zdnd11an1n64x5 FILLER_156_296 ();
 b15zdnd11an1n64x5 FILLER_156_360 ();
 b15zdnd11an1n64x5 FILLER_156_424 ();
 b15zdnd11an1n64x5 FILLER_156_488 ();
 b15zdnd11an1n64x5 FILLER_156_552 ();
 b15zdnd11an1n16x5 FILLER_156_616 ();
 b15zdnd11an1n08x5 FILLER_156_632 ();
 b15zdnd11an1n64x5 FILLER_156_650 ();
 b15zdnd11an1n04x5 FILLER_156_714 ();
 b15zdnd11an1n32x5 FILLER_156_726 ();
 b15zdnd11an1n04x5 FILLER_156_758 ();
 b15zdnd11an1n08x5 FILLER_156_765 ();
 b15zdnd11an1n04x5 FILLER_156_773 ();
 b15zdnd00an1n01x5 FILLER_156_777 ();
 b15zdnd11an1n32x5 FILLER_156_791 ();
 b15zdnd11an1n04x5 FILLER_156_823 ();
 b15zdnd00an1n01x5 FILLER_156_827 ();
 b15zdnd11an1n64x5 FILLER_156_832 ();
 b15zdnd11an1n64x5 FILLER_156_896 ();
 b15zdnd11an1n64x5 FILLER_156_960 ();
 b15zdnd11an1n64x5 FILLER_156_1024 ();
 b15zdnd11an1n32x5 FILLER_156_1088 ();
 b15zdnd11an1n08x5 FILLER_156_1120 ();
 b15zdnd11an1n04x5 FILLER_156_1128 ();
 b15zdnd00an1n02x5 FILLER_156_1132 ();
 b15zdnd00an1n01x5 FILLER_156_1134 ();
 b15zdnd11an1n64x5 FILLER_156_1138 ();
 b15zdnd11an1n16x5 FILLER_156_1202 ();
 b15zdnd00an1n01x5 FILLER_156_1218 ();
 b15zdnd11an1n64x5 FILLER_156_1222 ();
 b15zdnd11an1n64x5 FILLER_156_1286 ();
 b15zdnd11an1n64x5 FILLER_156_1350 ();
 b15zdnd11an1n64x5 FILLER_156_1414 ();
 b15zdnd11an1n64x5 FILLER_156_1478 ();
 b15zdnd11an1n64x5 FILLER_156_1542 ();
 b15zdnd11an1n64x5 FILLER_156_1606 ();
 b15zdnd11an1n64x5 FILLER_156_1670 ();
 b15zdnd11an1n64x5 FILLER_156_1734 ();
 b15zdnd11an1n64x5 FILLER_156_1798 ();
 b15zdnd11an1n64x5 FILLER_156_1862 ();
 b15zdnd11an1n64x5 FILLER_156_1926 ();
 b15zdnd11an1n16x5 FILLER_156_1990 ();
 b15zdnd11an1n04x5 FILLER_156_2006 ();
 b15zdnd00an1n02x5 FILLER_156_2010 ();
 b15zdnd11an1n64x5 FILLER_156_2018 ();
 b15zdnd11an1n64x5 FILLER_156_2082 ();
 b15zdnd11an1n08x5 FILLER_156_2146 ();
 b15zdnd11an1n64x5 FILLER_156_2162 ();
 b15zdnd11an1n32x5 FILLER_156_2226 ();
 b15zdnd11an1n16x5 FILLER_156_2258 ();
 b15zdnd00an1n02x5 FILLER_156_2274 ();
 b15zdnd11an1n64x5 FILLER_157_0 ();
 b15zdnd11an1n64x5 FILLER_157_64 ();
 b15zdnd11an1n64x5 FILLER_157_128 ();
 b15zdnd11an1n64x5 FILLER_157_192 ();
 b15zdnd11an1n16x5 FILLER_157_256 ();
 b15zdnd11an1n08x5 FILLER_157_272 ();
 b15zdnd00an1n02x5 FILLER_157_280 ();
 b15zdnd11an1n64x5 FILLER_157_324 ();
 b15zdnd11an1n64x5 FILLER_157_388 ();
 b15zdnd11an1n64x5 FILLER_157_452 ();
 b15zdnd11an1n08x5 FILLER_157_516 ();
 b15zdnd00an1n01x5 FILLER_157_524 ();
 b15zdnd11an1n64x5 FILLER_157_567 ();
 b15zdnd11an1n64x5 FILLER_157_631 ();
 b15zdnd11an1n32x5 FILLER_157_695 ();
 b15zdnd11an1n16x5 FILLER_157_727 ();
 b15zdnd11an1n04x5 FILLER_157_743 ();
 b15zdnd11an1n32x5 FILLER_157_760 ();
 b15zdnd11an1n16x5 FILLER_157_792 ();
 b15zdnd11an1n04x5 FILLER_157_808 ();
 b15zdnd11an1n64x5 FILLER_157_828 ();
 b15zdnd11an1n64x5 FILLER_157_892 ();
 b15zdnd11an1n64x5 FILLER_157_956 ();
 b15zdnd11an1n64x5 FILLER_157_1020 ();
 b15zdnd11an1n32x5 FILLER_157_1084 ();
 b15zdnd11an1n08x5 FILLER_157_1116 ();
 b15zdnd11an1n04x5 FILLER_157_1124 ();
 b15zdnd00an1n02x5 FILLER_157_1128 ();
 b15zdnd11an1n04x5 FILLER_157_1133 ();
 b15zdnd11an1n64x5 FILLER_157_1140 ();
 b15zdnd11an1n16x5 FILLER_157_1204 ();
 b15zdnd11an1n04x5 FILLER_157_1223 ();
 b15zdnd11an1n64x5 FILLER_157_1230 ();
 b15zdnd11an1n64x5 FILLER_157_1294 ();
 b15zdnd11an1n64x5 FILLER_157_1358 ();
 b15zdnd11an1n64x5 FILLER_157_1422 ();
 b15zdnd11an1n64x5 FILLER_157_1486 ();
 b15zdnd11an1n64x5 FILLER_157_1550 ();
 b15zdnd11an1n64x5 FILLER_157_1614 ();
 b15zdnd11an1n64x5 FILLER_157_1678 ();
 b15zdnd11an1n64x5 FILLER_157_1742 ();
 b15zdnd11an1n32x5 FILLER_157_1806 ();
 b15zdnd11an1n16x5 FILLER_157_1838 ();
 b15zdnd11an1n04x5 FILLER_157_1854 ();
 b15zdnd00an1n01x5 FILLER_157_1858 ();
 b15zdnd11an1n64x5 FILLER_157_1876 ();
 b15zdnd11an1n64x5 FILLER_157_1940 ();
 b15zdnd11an1n64x5 FILLER_157_2004 ();
 b15zdnd11an1n64x5 FILLER_157_2068 ();
 b15zdnd11an1n64x5 FILLER_157_2132 ();
 b15zdnd11an1n64x5 FILLER_157_2196 ();
 b15zdnd11an1n16x5 FILLER_157_2260 ();
 b15zdnd11an1n08x5 FILLER_157_2276 ();
 b15zdnd11an1n08x5 FILLER_158_8 ();
 b15zdnd11an1n04x5 FILLER_158_16 ();
 b15zdnd00an1n02x5 FILLER_158_20 ();
 b15zdnd00an1n01x5 FILLER_158_22 ();
 b15zdnd11an1n64x5 FILLER_158_27 ();
 b15zdnd11an1n64x5 FILLER_158_91 ();
 b15zdnd11an1n64x5 FILLER_158_155 ();
 b15zdnd11an1n64x5 FILLER_158_219 ();
 b15zdnd11an1n64x5 FILLER_158_283 ();
 b15zdnd11an1n64x5 FILLER_158_347 ();
 b15zdnd11an1n64x5 FILLER_158_411 ();
 b15zdnd11an1n64x5 FILLER_158_475 ();
 b15zdnd11an1n64x5 FILLER_158_539 ();
 b15zdnd11an1n64x5 FILLER_158_603 ();
 b15zdnd11an1n32x5 FILLER_158_667 ();
 b15zdnd11an1n16x5 FILLER_158_699 ();
 b15zdnd00an1n02x5 FILLER_158_715 ();
 b15zdnd00an1n01x5 FILLER_158_717 ();
 b15zdnd11an1n16x5 FILLER_158_726 ();
 b15zdnd11an1n08x5 FILLER_158_742 ();
 b15zdnd00an1n02x5 FILLER_158_750 ();
 b15zdnd11an1n64x5 FILLER_158_755 ();
 b15zdnd11an1n64x5 FILLER_158_839 ();
 b15zdnd11an1n64x5 FILLER_158_903 ();
 b15zdnd11an1n64x5 FILLER_158_967 ();
 b15zdnd11an1n64x5 FILLER_158_1031 ();
 b15zdnd00an1n02x5 FILLER_158_1095 ();
 b15zdnd11an1n04x5 FILLER_158_1106 ();
 b15zdnd11an1n32x5 FILLER_158_1162 ();
 b15zdnd11an1n04x5 FILLER_158_1194 ();
 b15zdnd00an1n02x5 FILLER_158_1198 ();
 b15zdnd11an1n04x5 FILLER_158_1252 ();
 b15zdnd11an1n64x5 FILLER_158_1259 ();
 b15zdnd11an1n32x5 FILLER_158_1323 ();
 b15zdnd11an1n08x5 FILLER_158_1355 ();
 b15zdnd11an1n64x5 FILLER_158_1374 ();
 b15zdnd11an1n32x5 FILLER_158_1438 ();
 b15zdnd11an1n16x5 FILLER_158_1470 ();
 b15zdnd11an1n08x5 FILLER_158_1486 ();
 b15zdnd11an1n64x5 FILLER_158_1503 ();
 b15zdnd11an1n64x5 FILLER_158_1567 ();
 b15zdnd11an1n64x5 FILLER_158_1631 ();
 b15zdnd11an1n64x5 FILLER_158_1695 ();
 b15zdnd11an1n64x5 FILLER_158_1759 ();
 b15zdnd11an1n64x5 FILLER_158_1823 ();
 b15zdnd11an1n64x5 FILLER_158_1887 ();
 b15zdnd11an1n64x5 FILLER_158_1951 ();
 b15zdnd11an1n64x5 FILLER_158_2015 ();
 b15zdnd11an1n64x5 FILLER_158_2079 ();
 b15zdnd11an1n08x5 FILLER_158_2143 ();
 b15zdnd00an1n02x5 FILLER_158_2151 ();
 b15zdnd00an1n01x5 FILLER_158_2153 ();
 b15zdnd11an1n64x5 FILLER_158_2162 ();
 b15zdnd11an1n16x5 FILLER_158_2226 ();
 b15zdnd11an1n16x5 FILLER_158_2253 ();
 b15zdnd11an1n04x5 FILLER_158_2269 ();
 b15zdnd00an1n02x5 FILLER_158_2273 ();
 b15zdnd00an1n01x5 FILLER_158_2275 ();
 b15zdnd11an1n64x5 FILLER_159_0 ();
 b15zdnd11an1n64x5 FILLER_159_64 ();
 b15zdnd11an1n64x5 FILLER_159_128 ();
 b15zdnd11an1n64x5 FILLER_159_192 ();
 b15zdnd11an1n64x5 FILLER_159_256 ();
 b15zdnd11an1n64x5 FILLER_159_320 ();
 b15zdnd11an1n16x5 FILLER_159_384 ();
 b15zdnd11an1n04x5 FILLER_159_400 ();
 b15zdnd00an1n01x5 FILLER_159_404 ();
 b15zdnd11an1n64x5 FILLER_159_447 ();
 b15zdnd11an1n64x5 FILLER_159_511 ();
 b15zdnd11an1n32x5 FILLER_159_575 ();
 b15zdnd11an1n08x5 FILLER_159_607 ();
 b15zdnd11an1n04x5 FILLER_159_615 ();
 b15zdnd11an1n16x5 FILLER_159_627 ();
 b15zdnd11an1n04x5 FILLER_159_643 ();
 b15zdnd00an1n02x5 FILLER_159_647 ();
 b15zdnd00an1n01x5 FILLER_159_649 ();
 b15zdnd11an1n64x5 FILLER_159_653 ();
 b15zdnd11an1n64x5 FILLER_159_717 ();
 b15zdnd11an1n64x5 FILLER_159_781 ();
 b15zdnd11an1n64x5 FILLER_159_845 ();
 b15zdnd11an1n32x5 FILLER_159_909 ();
 b15zdnd11an1n08x5 FILLER_159_941 ();
 b15zdnd11an1n64x5 FILLER_159_952 ();
 b15zdnd11an1n32x5 FILLER_159_1016 ();
 b15zdnd00an1n02x5 FILLER_159_1048 ();
 b15zdnd11an1n32x5 FILLER_159_1059 ();
 b15zdnd11an1n16x5 FILLER_159_1091 ();
 b15zdnd00an1n02x5 FILLER_159_1107 ();
 b15zdnd00an1n01x5 FILLER_159_1109 ();
 b15zdnd11an1n64x5 FILLER_159_1162 ();
 b15zdnd11an1n16x5 FILLER_159_1226 ();
 b15zdnd00an1n01x5 FILLER_159_1242 ();
 b15zdnd11an1n64x5 FILLER_159_1270 ();
 b15zdnd11an1n64x5 FILLER_159_1334 ();
 b15zdnd11an1n64x5 FILLER_159_1398 ();
 b15zdnd11an1n64x5 FILLER_159_1462 ();
 b15zdnd11an1n64x5 FILLER_159_1526 ();
 b15zdnd11an1n64x5 FILLER_159_1590 ();
 b15zdnd11an1n64x5 FILLER_159_1654 ();
 b15zdnd11an1n64x5 FILLER_159_1718 ();
 b15zdnd11an1n64x5 FILLER_159_1782 ();
 b15zdnd11an1n64x5 FILLER_159_1846 ();
 b15zdnd11an1n64x5 FILLER_159_1910 ();
 b15zdnd11an1n64x5 FILLER_159_1974 ();
 b15zdnd11an1n64x5 FILLER_159_2038 ();
 b15zdnd11an1n32x5 FILLER_159_2102 ();
 b15zdnd11an1n04x5 FILLER_159_2134 ();
 b15zdnd00an1n01x5 FILLER_159_2138 ();
 b15zdnd11an1n64x5 FILLER_159_2147 ();
 b15zdnd11an1n64x5 FILLER_159_2211 ();
 b15zdnd11an1n08x5 FILLER_159_2275 ();
 b15zdnd00an1n01x5 FILLER_159_2283 ();
 b15zdnd11an1n64x5 FILLER_160_8 ();
 b15zdnd11an1n64x5 FILLER_160_72 ();
 b15zdnd11an1n64x5 FILLER_160_136 ();
 b15zdnd11an1n64x5 FILLER_160_200 ();
 b15zdnd11an1n16x5 FILLER_160_264 ();
 b15zdnd11an1n64x5 FILLER_160_286 ();
 b15zdnd11an1n32x5 FILLER_160_350 ();
 b15zdnd11an1n08x5 FILLER_160_382 ();
 b15zdnd11an1n04x5 FILLER_160_390 ();
 b15zdnd11an1n32x5 FILLER_160_446 ();
 b15zdnd11an1n16x5 FILLER_160_478 ();
 b15zdnd11an1n08x5 FILLER_160_494 ();
 b15zdnd00an1n01x5 FILLER_160_502 ();
 b15zdnd11an1n64x5 FILLER_160_506 ();
 b15zdnd11an1n32x5 FILLER_160_570 ();
 b15zdnd11an1n16x5 FILLER_160_602 ();
 b15zdnd11an1n04x5 FILLER_160_618 ();
 b15zdnd00an1n01x5 FILLER_160_622 ();
 b15zdnd11an1n32x5 FILLER_160_675 ();
 b15zdnd11an1n08x5 FILLER_160_707 ();
 b15zdnd00an1n02x5 FILLER_160_715 ();
 b15zdnd00an1n01x5 FILLER_160_717 ();
 b15zdnd11an1n64x5 FILLER_160_726 ();
 b15zdnd00an1n02x5 FILLER_160_790 ();
 b15zdnd11an1n64x5 FILLER_160_809 ();
 b15zdnd11an1n32x5 FILLER_160_873 ();
 b15zdnd00an1n02x5 FILLER_160_905 ();
 b15zdnd00an1n01x5 FILLER_160_907 ();
 b15zdnd11an1n04x5 FILLER_160_917 ();
 b15zdnd00an1n01x5 FILLER_160_921 ();
 b15zdnd11an1n32x5 FILLER_160_974 ();
 b15zdnd11an1n16x5 FILLER_160_1006 ();
 b15zdnd11an1n16x5 FILLER_160_1026 ();
 b15zdnd11an1n08x5 FILLER_160_1042 ();
 b15zdnd00an1n02x5 FILLER_160_1050 ();
 b15zdnd00an1n01x5 FILLER_160_1052 ();
 b15zdnd11an1n04x5 FILLER_160_1062 ();
 b15zdnd11an1n32x5 FILLER_160_1075 ();
 b15zdnd11an1n16x5 FILLER_160_1107 ();
 b15zdnd11an1n04x5 FILLER_160_1123 ();
 b15zdnd00an1n02x5 FILLER_160_1127 ();
 b15zdnd11an1n04x5 FILLER_160_1132 ();
 b15zdnd11an1n08x5 FILLER_160_1139 ();
 b15zdnd11an1n04x5 FILLER_160_1147 ();
 b15zdnd00an1n02x5 FILLER_160_1151 ();
 b15zdnd11an1n32x5 FILLER_160_1167 ();
 b15zdnd11an1n16x5 FILLER_160_1199 ();
 b15zdnd11an1n04x5 FILLER_160_1215 ();
 b15zdnd00an1n02x5 FILLER_160_1219 ();
 b15zdnd11an1n64x5 FILLER_160_1273 ();
 b15zdnd11an1n08x5 FILLER_160_1337 ();
 b15zdnd11an1n04x5 FILLER_160_1345 ();
 b15zdnd00an1n01x5 FILLER_160_1349 ();
 b15zdnd11an1n64x5 FILLER_160_1381 ();
 b15zdnd11an1n64x5 FILLER_160_1445 ();
 b15zdnd11an1n64x5 FILLER_160_1509 ();
 b15zdnd11an1n64x5 FILLER_160_1573 ();
 b15zdnd11an1n64x5 FILLER_160_1637 ();
 b15zdnd11an1n64x5 FILLER_160_1701 ();
 b15zdnd11an1n64x5 FILLER_160_1765 ();
 b15zdnd11an1n64x5 FILLER_160_1829 ();
 b15zdnd11an1n08x5 FILLER_160_1893 ();
 b15zdnd00an1n01x5 FILLER_160_1901 ();
 b15zdnd11an1n64x5 FILLER_160_1922 ();
 b15zdnd11an1n64x5 FILLER_160_1986 ();
 b15zdnd11an1n64x5 FILLER_160_2050 ();
 b15zdnd11an1n32x5 FILLER_160_2114 ();
 b15zdnd11an1n08x5 FILLER_160_2146 ();
 b15zdnd11an1n64x5 FILLER_160_2162 ();
 b15zdnd11an1n16x5 FILLER_160_2226 ();
 b15zdnd00an1n02x5 FILLER_160_2242 ();
 b15zdnd11an1n16x5 FILLER_160_2254 ();
 b15zdnd11an1n04x5 FILLER_160_2270 ();
 b15zdnd00an1n02x5 FILLER_160_2274 ();
 b15zdnd11an1n64x5 FILLER_161_0 ();
 b15zdnd11an1n32x5 FILLER_161_64 ();
 b15zdnd11an1n64x5 FILLER_161_138 ();
 b15zdnd11an1n64x5 FILLER_161_202 ();
 b15zdnd00an1n02x5 FILLER_161_266 ();
 b15zdnd11an1n64x5 FILLER_161_282 ();
 b15zdnd11an1n16x5 FILLER_161_346 ();
 b15zdnd11an1n04x5 FILLER_161_362 ();
 b15zdnd00an1n01x5 FILLER_161_366 ();
 b15zdnd11an1n04x5 FILLER_161_409 ();
 b15zdnd00an1n01x5 FILLER_161_413 ();
 b15zdnd11an1n04x5 FILLER_161_417 ();
 b15zdnd11an1n32x5 FILLER_161_424 ();
 b15zdnd11an1n16x5 FILLER_161_456 ();
 b15zdnd11an1n04x5 FILLER_161_472 ();
 b15zdnd11an1n64x5 FILLER_161_528 ();
 b15zdnd11an1n32x5 FILLER_161_592 ();
 b15zdnd11an1n16x5 FILLER_161_624 ();
 b15zdnd00an1n02x5 FILLER_161_640 ();
 b15zdnd11an1n04x5 FILLER_161_645 ();
 b15zdnd11an1n16x5 FILLER_161_652 ();
 b15zdnd11an1n08x5 FILLER_161_668 ();
 b15zdnd11an1n04x5 FILLER_161_676 ();
 b15zdnd11an1n64x5 FILLER_161_722 ();
 b15zdnd11an1n64x5 FILLER_161_786 ();
 b15zdnd11an1n64x5 FILLER_161_850 ();
 b15zdnd11an1n16x5 FILLER_161_914 ();
 b15zdnd11an1n08x5 FILLER_161_930 ();
 b15zdnd00an1n02x5 FILLER_161_938 ();
 b15zdnd00an1n01x5 FILLER_161_940 ();
 b15zdnd11an1n04x5 FILLER_161_944 ();
 b15zdnd11an1n64x5 FILLER_161_951 ();
 b15zdnd11an1n32x5 FILLER_161_1015 ();
 b15zdnd11an1n08x5 FILLER_161_1047 ();
 b15zdnd11an1n04x5 FILLER_161_1055 ();
 b15zdnd00an1n02x5 FILLER_161_1059 ();
 b15zdnd00an1n01x5 FILLER_161_1061 ();
 b15zdnd11an1n32x5 FILLER_161_1076 ();
 b15zdnd11an1n16x5 FILLER_161_1108 ();
 b15zdnd11an1n08x5 FILLER_161_1124 ();
 b15zdnd00an1n02x5 FILLER_161_1132 ();
 b15zdnd00an1n01x5 FILLER_161_1134 ();
 b15zdnd11an1n08x5 FILLER_161_1138 ();
 b15zdnd00an1n02x5 FILLER_161_1146 ();
 b15zdnd11an1n32x5 FILLER_161_1190 ();
 b15zdnd11an1n16x5 FILLER_161_1222 ();
 b15zdnd00an1n02x5 FILLER_161_1238 ();
 b15zdnd11an1n04x5 FILLER_161_1243 ();
 b15zdnd11an1n64x5 FILLER_161_1250 ();
 b15zdnd11an1n64x5 FILLER_161_1314 ();
 b15zdnd11an1n64x5 FILLER_161_1378 ();
 b15zdnd11an1n64x5 FILLER_161_1442 ();
 b15zdnd11an1n64x5 FILLER_161_1506 ();
 b15zdnd11an1n64x5 FILLER_161_1570 ();
 b15zdnd11an1n64x5 FILLER_161_1634 ();
 b15zdnd11an1n64x5 FILLER_161_1698 ();
 b15zdnd11an1n16x5 FILLER_161_1762 ();
 b15zdnd11an1n04x5 FILLER_161_1778 ();
 b15zdnd00an1n02x5 FILLER_161_1782 ();
 b15zdnd00an1n01x5 FILLER_161_1784 ();
 b15zdnd11an1n64x5 FILLER_161_1788 ();
 b15zdnd11an1n64x5 FILLER_161_1852 ();
 b15zdnd11an1n64x5 FILLER_161_1916 ();
 b15zdnd11an1n64x5 FILLER_161_1980 ();
 b15zdnd11an1n04x5 FILLER_161_2044 ();
 b15zdnd00an1n02x5 FILLER_161_2048 ();
 b15zdnd00an1n01x5 FILLER_161_2050 ();
 b15zdnd11an1n32x5 FILLER_161_2065 ();
 b15zdnd11an1n04x5 FILLER_161_2097 ();
 b15zdnd00an1n02x5 FILLER_161_2101 ();
 b15zdnd00an1n01x5 FILLER_161_2103 ();
 b15zdnd11an1n64x5 FILLER_161_2146 ();
 b15zdnd11an1n64x5 FILLER_161_2210 ();
 b15zdnd11an1n08x5 FILLER_161_2274 ();
 b15zdnd00an1n02x5 FILLER_161_2282 ();
 b15zdnd11an1n08x5 FILLER_162_8 ();
 b15zdnd00an1n02x5 FILLER_162_16 ();
 b15zdnd11an1n64x5 FILLER_162_22 ();
 b15zdnd11an1n04x5 FILLER_162_86 ();
 b15zdnd00an1n02x5 FILLER_162_90 ();
 b15zdnd11an1n04x5 FILLER_162_134 ();
 b15zdnd11an1n64x5 FILLER_162_141 ();
 b15zdnd11an1n64x5 FILLER_162_205 ();
 b15zdnd11an1n04x5 FILLER_162_284 ();
 b15zdnd11an1n64x5 FILLER_162_293 ();
 b15zdnd11an1n32x5 FILLER_162_357 ();
 b15zdnd11an1n16x5 FILLER_162_389 ();
 b15zdnd11an1n08x5 FILLER_162_405 ();
 b15zdnd11an1n04x5 FILLER_162_413 ();
 b15zdnd00an1n02x5 FILLER_162_417 ();
 b15zdnd11an1n64x5 FILLER_162_422 ();
 b15zdnd11an1n08x5 FILLER_162_486 ();
 b15zdnd00an1n01x5 FILLER_162_494 ();
 b15zdnd11an1n04x5 FILLER_162_498 ();
 b15zdnd11an1n64x5 FILLER_162_505 ();
 b15zdnd11an1n64x5 FILLER_162_569 ();
 b15zdnd11an1n64x5 FILLER_162_633 ();
 b15zdnd11an1n16x5 FILLER_162_697 ();
 b15zdnd11an1n04x5 FILLER_162_713 ();
 b15zdnd00an1n01x5 FILLER_162_717 ();
 b15zdnd11an1n64x5 FILLER_162_726 ();
 b15zdnd11an1n64x5 FILLER_162_790 ();
 b15zdnd11an1n16x5 FILLER_162_854 ();
 b15zdnd00an1n02x5 FILLER_162_870 ();
 b15zdnd11an1n64x5 FILLER_162_876 ();
 b15zdnd11an1n64x5 FILLER_162_940 ();
 b15zdnd11an1n64x5 FILLER_162_1004 ();
 b15zdnd11an1n64x5 FILLER_162_1068 ();
 b15zdnd11an1n64x5 FILLER_162_1132 ();
 b15zdnd11an1n32x5 FILLER_162_1196 ();
 b15zdnd11an1n16x5 FILLER_162_1228 ();
 b15zdnd00an1n02x5 FILLER_162_1244 ();
 b15zdnd11an1n64x5 FILLER_162_1249 ();
 b15zdnd11an1n64x5 FILLER_162_1313 ();
 b15zdnd11an1n16x5 FILLER_162_1377 ();
 b15zdnd11an1n08x5 FILLER_162_1393 ();
 b15zdnd11an1n04x5 FILLER_162_1401 ();
 b15zdnd11an1n64x5 FILLER_162_1432 ();
 b15zdnd11an1n64x5 FILLER_162_1496 ();
 b15zdnd11an1n64x5 FILLER_162_1560 ();
 b15zdnd11an1n64x5 FILLER_162_1624 ();
 b15zdnd11an1n64x5 FILLER_162_1688 ();
 b15zdnd11an1n04x5 FILLER_162_1752 ();
 b15zdnd00an1n02x5 FILLER_162_1756 ();
 b15zdnd11an1n64x5 FILLER_162_1810 ();
 b15zdnd11an1n64x5 FILLER_162_1874 ();
 b15zdnd11an1n64x5 FILLER_162_1938 ();
 b15zdnd11an1n32x5 FILLER_162_2002 ();
 b15zdnd11an1n16x5 FILLER_162_2034 ();
 b15zdnd00an1n01x5 FILLER_162_2050 ();
 b15zdnd11an1n64x5 FILLER_162_2058 ();
 b15zdnd11an1n32x5 FILLER_162_2122 ();
 b15zdnd11an1n64x5 FILLER_162_2162 ();
 b15zdnd11an1n32x5 FILLER_162_2226 ();
 b15zdnd11an1n16x5 FILLER_162_2258 ();
 b15zdnd00an1n02x5 FILLER_162_2274 ();
 b15zdnd11an1n16x5 FILLER_163_0 ();
 b15zdnd11an1n04x5 FILLER_163_16 ();
 b15zdnd00an1n02x5 FILLER_163_20 ();
 b15zdnd00an1n01x5 FILLER_163_22 ();
 b15zdnd11an1n04x5 FILLER_163_27 ();
 b15zdnd11an1n64x5 FILLER_163_35 ();
 b15zdnd11an1n08x5 FILLER_163_99 ();
 b15zdnd00an1n01x5 FILLER_163_107 ();
 b15zdnd11an1n64x5 FILLER_163_160 ();
 b15zdnd11an1n32x5 FILLER_163_224 ();
 b15zdnd00an1n01x5 FILLER_163_256 ();
 b15zdnd11an1n64x5 FILLER_163_299 ();
 b15zdnd11an1n64x5 FILLER_163_363 ();
 b15zdnd11an1n64x5 FILLER_163_427 ();
 b15zdnd11an1n64x5 FILLER_163_491 ();
 b15zdnd11an1n64x5 FILLER_163_555 ();
 b15zdnd11an1n64x5 FILLER_163_619 ();
 b15zdnd11an1n32x5 FILLER_163_683 ();
 b15zdnd11an1n16x5 FILLER_163_715 ();
 b15zdnd11an1n04x5 FILLER_163_731 ();
 b15zdnd00an1n01x5 FILLER_163_735 ();
 b15zdnd11an1n64x5 FILLER_163_741 ();
 b15zdnd11an1n64x5 FILLER_163_805 ();
 b15zdnd11an1n64x5 FILLER_163_869 ();
 b15zdnd11an1n64x5 FILLER_163_933 ();
 b15zdnd11an1n64x5 FILLER_163_997 ();
 b15zdnd11an1n64x5 FILLER_163_1061 ();
 b15zdnd11an1n64x5 FILLER_163_1125 ();
 b15zdnd11an1n64x5 FILLER_163_1189 ();
 b15zdnd11an1n64x5 FILLER_163_1253 ();
 b15zdnd11an1n64x5 FILLER_163_1317 ();
 b15zdnd11an1n16x5 FILLER_163_1381 ();
 b15zdnd11an1n08x5 FILLER_163_1397 ();
 b15zdnd00an1n02x5 FILLER_163_1405 ();
 b15zdnd00an1n01x5 FILLER_163_1407 ();
 b15zdnd11an1n16x5 FILLER_163_1411 ();
 b15zdnd11an1n04x5 FILLER_163_1427 ();
 b15zdnd00an1n02x5 FILLER_163_1431 ();
 b15zdnd11an1n64x5 FILLER_163_1441 ();
 b15zdnd11an1n64x5 FILLER_163_1505 ();
 b15zdnd11an1n64x5 FILLER_163_1569 ();
 b15zdnd11an1n64x5 FILLER_163_1633 ();
 b15zdnd11an1n32x5 FILLER_163_1697 ();
 b15zdnd11an1n08x5 FILLER_163_1729 ();
 b15zdnd11an1n04x5 FILLER_163_1740 ();
 b15zdnd00an1n02x5 FILLER_163_1744 ();
 b15zdnd11an1n16x5 FILLER_163_1798 ();
 b15zdnd11an1n04x5 FILLER_163_1814 ();
 b15zdnd00an1n02x5 FILLER_163_1818 ();
 b15zdnd11an1n16x5 FILLER_163_1834 ();
 b15zdnd11an1n08x5 FILLER_163_1850 ();
 b15zdnd00an1n01x5 FILLER_163_1858 ();
 b15zdnd11an1n64x5 FILLER_163_1863 ();
 b15zdnd11an1n64x5 FILLER_163_1927 ();
 b15zdnd11an1n16x5 FILLER_163_1991 ();
 b15zdnd00an1n02x5 FILLER_163_2007 ();
 b15zdnd00an1n01x5 FILLER_163_2009 ();
 b15zdnd11an1n64x5 FILLER_163_2016 ();
 b15zdnd11an1n64x5 FILLER_163_2080 ();
 b15zdnd11an1n64x5 FILLER_163_2144 ();
 b15zdnd11an1n64x5 FILLER_163_2208 ();
 b15zdnd11an1n08x5 FILLER_163_2272 ();
 b15zdnd11an1n04x5 FILLER_163_2280 ();
 b15zdnd11an1n32x5 FILLER_164_8 ();
 b15zdnd00an1n02x5 FILLER_164_40 ();
 b15zdnd00an1n01x5 FILLER_164_42 ();
 b15zdnd11an1n16x5 FILLER_164_85 ();
 b15zdnd00an1n02x5 FILLER_164_101 ();
 b15zdnd11an1n64x5 FILLER_164_145 ();
 b15zdnd11an1n64x5 FILLER_164_209 ();
 b15zdnd11an1n08x5 FILLER_164_273 ();
 b15zdnd11an1n04x5 FILLER_164_281 ();
 b15zdnd00an1n02x5 FILLER_164_285 ();
 b15zdnd00an1n01x5 FILLER_164_287 ();
 b15zdnd11an1n64x5 FILLER_164_291 ();
 b15zdnd11an1n64x5 FILLER_164_355 ();
 b15zdnd11an1n64x5 FILLER_164_419 ();
 b15zdnd11an1n64x5 FILLER_164_483 ();
 b15zdnd11an1n64x5 FILLER_164_547 ();
 b15zdnd11an1n64x5 FILLER_164_611 ();
 b15zdnd11an1n32x5 FILLER_164_675 ();
 b15zdnd11an1n08x5 FILLER_164_707 ();
 b15zdnd00an1n02x5 FILLER_164_715 ();
 b15zdnd00an1n01x5 FILLER_164_717 ();
 b15zdnd11an1n64x5 FILLER_164_726 ();
 b15zdnd11an1n64x5 FILLER_164_790 ();
 b15zdnd11an1n64x5 FILLER_164_854 ();
 b15zdnd11an1n64x5 FILLER_164_918 ();
 b15zdnd11an1n64x5 FILLER_164_982 ();
 b15zdnd11an1n64x5 FILLER_164_1046 ();
 b15zdnd11an1n64x5 FILLER_164_1110 ();
 b15zdnd11an1n64x5 FILLER_164_1174 ();
 b15zdnd11an1n64x5 FILLER_164_1238 ();
 b15zdnd11an1n16x5 FILLER_164_1302 ();
 b15zdnd11an1n64x5 FILLER_164_1349 ();
 b15zdnd11an1n64x5 FILLER_164_1413 ();
 b15zdnd11an1n64x5 FILLER_164_1477 ();
 b15zdnd11an1n64x5 FILLER_164_1541 ();
 b15zdnd11an1n64x5 FILLER_164_1605 ();
 b15zdnd11an1n32x5 FILLER_164_1669 ();
 b15zdnd11an1n08x5 FILLER_164_1701 ();
 b15zdnd11an1n08x5 FILLER_164_1761 ();
 b15zdnd11an1n04x5 FILLER_164_1772 ();
 b15zdnd11an1n04x5 FILLER_164_1779 ();
 b15zdnd11an1n32x5 FILLER_164_1786 ();
 b15zdnd11an1n16x5 FILLER_164_1818 ();
 b15zdnd00an1n02x5 FILLER_164_1834 ();
 b15zdnd00an1n01x5 FILLER_164_1836 ();
 b15zdnd11an1n04x5 FILLER_164_1845 ();
 b15zdnd11an1n04x5 FILLER_164_1853 ();
 b15zdnd11an1n64x5 FILLER_164_1861 ();
 b15zdnd11an1n64x5 FILLER_164_1925 ();
 b15zdnd11an1n64x5 FILLER_164_1989 ();
 b15zdnd11an1n64x5 FILLER_164_2053 ();
 b15zdnd11an1n04x5 FILLER_164_2117 ();
 b15zdnd00an1n02x5 FILLER_164_2121 ();
 b15zdnd00an1n01x5 FILLER_164_2123 ();
 b15zdnd00an1n02x5 FILLER_164_2152 ();
 b15zdnd00an1n02x5 FILLER_164_2162 ();
 b15zdnd11an1n64x5 FILLER_164_2182 ();
 b15zdnd11an1n16x5 FILLER_164_2246 ();
 b15zdnd11an1n08x5 FILLER_164_2262 ();
 b15zdnd11an1n04x5 FILLER_164_2270 ();
 b15zdnd00an1n02x5 FILLER_164_2274 ();
 b15zdnd11an1n64x5 FILLER_165_0 ();
 b15zdnd11an1n16x5 FILLER_165_64 ();
 b15zdnd11an1n08x5 FILLER_165_80 ();
 b15zdnd11an1n04x5 FILLER_165_88 ();
 b15zdnd00an1n01x5 FILLER_165_92 ();
 b15zdnd11an1n04x5 FILLER_165_135 ();
 b15zdnd11an1n64x5 FILLER_165_142 ();
 b15zdnd11an1n64x5 FILLER_165_206 ();
 b15zdnd11an1n08x5 FILLER_165_270 ();
 b15zdnd11an1n04x5 FILLER_165_278 ();
 b15zdnd00an1n01x5 FILLER_165_282 ();
 b15zdnd11an1n64x5 FILLER_165_289 ();
 b15zdnd11an1n64x5 FILLER_165_353 ();
 b15zdnd11an1n64x5 FILLER_165_417 ();
 b15zdnd11an1n64x5 FILLER_165_481 ();
 b15zdnd11an1n64x5 FILLER_165_545 ();
 b15zdnd11an1n64x5 FILLER_165_609 ();
 b15zdnd11an1n64x5 FILLER_165_673 ();
 b15zdnd11an1n64x5 FILLER_165_737 ();
 b15zdnd11an1n64x5 FILLER_165_801 ();
 b15zdnd11an1n64x5 FILLER_165_865 ();
 b15zdnd11an1n64x5 FILLER_165_929 ();
 b15zdnd11an1n64x5 FILLER_165_993 ();
 b15zdnd11an1n16x5 FILLER_165_1057 ();
 b15zdnd00an1n02x5 FILLER_165_1073 ();
 b15zdnd00an1n01x5 FILLER_165_1075 ();
 b15zdnd11an1n64x5 FILLER_165_1081 ();
 b15zdnd11an1n64x5 FILLER_165_1145 ();
 b15zdnd11an1n64x5 FILLER_165_1209 ();
 b15zdnd11an1n64x5 FILLER_165_1273 ();
 b15zdnd11an1n64x5 FILLER_165_1337 ();
 b15zdnd11an1n64x5 FILLER_165_1401 ();
 b15zdnd11an1n64x5 FILLER_165_1465 ();
 b15zdnd11an1n32x5 FILLER_165_1529 ();
 b15zdnd11an1n04x5 FILLER_165_1561 ();
 b15zdnd00an1n02x5 FILLER_165_1565 ();
 b15zdnd11an1n64x5 FILLER_165_1570 ();
 b15zdnd11an1n64x5 FILLER_165_1634 ();
 b15zdnd11an1n08x5 FILLER_165_1698 ();
 b15zdnd11an1n04x5 FILLER_165_1706 ();
 b15zdnd00an1n02x5 FILLER_165_1710 ();
 b15zdnd11an1n04x5 FILLER_165_1764 ();
 b15zdnd11an1n08x5 FILLER_165_1771 ();
 b15zdnd00an1n01x5 FILLER_165_1779 ();
 b15zdnd11an1n04x5 FILLER_165_1783 ();
 b15zdnd11an1n04x5 FILLER_165_1829 ();
 b15zdnd00an1n01x5 FILLER_165_1833 ();
 b15zdnd11an1n64x5 FILLER_165_1838 ();
 b15zdnd11an1n32x5 FILLER_165_1902 ();
 b15zdnd00an1n01x5 FILLER_165_1934 ();
 b15zdnd11an1n04x5 FILLER_165_1941 ();
 b15zdnd11an1n32x5 FILLER_165_1948 ();
 b15zdnd11an1n16x5 FILLER_165_1980 ();
 b15zdnd11an1n04x5 FILLER_165_1996 ();
 b15zdnd00an1n02x5 FILLER_165_2000 ();
 b15zdnd00an1n01x5 FILLER_165_2002 ();
 b15zdnd11an1n64x5 FILLER_165_2015 ();
 b15zdnd11an1n64x5 FILLER_165_2079 ();
 b15zdnd11an1n64x5 FILLER_165_2143 ();
 b15zdnd11an1n64x5 FILLER_165_2207 ();
 b15zdnd11an1n08x5 FILLER_165_2271 ();
 b15zdnd11an1n04x5 FILLER_165_2279 ();
 b15zdnd00an1n01x5 FILLER_165_2283 ();
 b15zdnd11an1n64x5 FILLER_166_8 ();
 b15zdnd00an1n01x5 FILLER_166_72 ();
 b15zdnd11an1n16x5 FILLER_166_104 ();
 b15zdnd11an1n04x5 FILLER_166_120 ();
 b15zdnd00an1n02x5 FILLER_166_124 ();
 b15zdnd11an1n64x5 FILLER_166_129 ();
 b15zdnd11an1n64x5 FILLER_166_193 ();
 b15zdnd11an1n16x5 FILLER_166_257 ();
 b15zdnd11an1n08x5 FILLER_166_273 ();
 b15zdnd11an1n04x5 FILLER_166_281 ();
 b15zdnd11an1n32x5 FILLER_166_295 ();
 b15zdnd11an1n04x5 FILLER_166_327 ();
 b15zdnd00an1n02x5 FILLER_166_331 ();
 b15zdnd00an1n01x5 FILLER_166_333 ();
 b15zdnd11an1n64x5 FILLER_166_340 ();
 b15zdnd11an1n64x5 FILLER_166_404 ();
 b15zdnd11an1n64x5 FILLER_166_468 ();
 b15zdnd11an1n64x5 FILLER_166_532 ();
 b15zdnd11an1n64x5 FILLER_166_596 ();
 b15zdnd11an1n08x5 FILLER_166_660 ();
 b15zdnd00an1n01x5 FILLER_166_668 ();
 b15zdnd11an1n16x5 FILLER_166_689 ();
 b15zdnd11an1n08x5 FILLER_166_705 ();
 b15zdnd11an1n04x5 FILLER_166_713 ();
 b15zdnd00an1n01x5 FILLER_166_717 ();
 b15zdnd11an1n64x5 FILLER_166_726 ();
 b15zdnd11an1n64x5 FILLER_166_790 ();
 b15zdnd11an1n64x5 FILLER_166_854 ();
 b15zdnd11an1n64x5 FILLER_166_918 ();
 b15zdnd11an1n16x5 FILLER_166_982 ();
 b15zdnd00an1n02x5 FILLER_166_998 ();
 b15zdnd00an1n01x5 FILLER_166_1000 ();
 b15zdnd11an1n64x5 FILLER_166_1021 ();
 b15zdnd11an1n64x5 FILLER_166_1085 ();
 b15zdnd11an1n64x5 FILLER_166_1149 ();
 b15zdnd11an1n32x5 FILLER_166_1213 ();
 b15zdnd11an1n16x5 FILLER_166_1245 ();
 b15zdnd11an1n08x5 FILLER_166_1261 ();
 b15zdnd00an1n02x5 FILLER_166_1269 ();
 b15zdnd11an1n64x5 FILLER_166_1313 ();
 b15zdnd11an1n32x5 FILLER_166_1377 ();
 b15zdnd11an1n08x5 FILLER_166_1409 ();
 b15zdnd00an1n01x5 FILLER_166_1417 ();
 b15zdnd11an1n04x5 FILLER_166_1421 ();
 b15zdnd11an1n64x5 FILLER_166_1428 ();
 b15zdnd11an1n32x5 FILLER_166_1492 ();
 b15zdnd11an1n16x5 FILLER_166_1524 ();
 b15zdnd00an1n01x5 FILLER_166_1540 ();
 b15zdnd11an1n64x5 FILLER_166_1593 ();
 b15zdnd11an1n64x5 FILLER_166_1657 ();
 b15zdnd11an1n04x5 FILLER_166_1721 ();
 b15zdnd00an1n02x5 FILLER_166_1725 ();
 b15zdnd11an1n04x5 FILLER_166_1730 ();
 b15zdnd11an1n04x5 FILLER_166_1737 ();
 b15zdnd11an1n04x5 FILLER_166_1744 ();
 b15zdnd11an1n16x5 FILLER_166_1751 ();
 b15zdnd11an1n08x5 FILLER_166_1767 ();
 b15zdnd00an1n01x5 FILLER_166_1775 ();
 b15zdnd11an1n64x5 FILLER_166_1783 ();
 b15zdnd11an1n64x5 FILLER_166_1847 ();
 b15zdnd11an1n08x5 FILLER_166_1911 ();
 b15zdnd11an1n04x5 FILLER_166_1919 ();
 b15zdnd00an1n02x5 FILLER_166_1923 ();
 b15zdnd00an1n01x5 FILLER_166_1925 ();
 b15zdnd11an1n64x5 FILLER_166_1968 ();
 b15zdnd11an1n16x5 FILLER_166_2032 ();
 b15zdnd11an1n08x5 FILLER_166_2048 ();
 b15zdnd11an1n04x5 FILLER_166_2056 ();
 b15zdnd00an1n02x5 FILLER_166_2060 ();
 b15zdnd00an1n01x5 FILLER_166_2062 ();
 b15zdnd11an1n08x5 FILLER_166_2068 ();
 b15zdnd00an1n01x5 FILLER_166_2076 ();
 b15zdnd11an1n64x5 FILLER_166_2089 ();
 b15zdnd00an1n01x5 FILLER_166_2153 ();
 b15zdnd11an1n04x5 FILLER_166_2162 ();
 b15zdnd00an1n02x5 FILLER_166_2166 ();
 b15zdnd00an1n01x5 FILLER_166_2168 ();
 b15zdnd11an1n16x5 FILLER_166_2181 ();
 b15zdnd00an1n01x5 FILLER_166_2197 ();
 b15zdnd11an1n64x5 FILLER_166_2206 ();
 b15zdnd11an1n04x5 FILLER_166_2270 ();
 b15zdnd00an1n02x5 FILLER_166_2274 ();
 b15zdnd11an1n64x5 FILLER_167_0 ();
 b15zdnd11an1n08x5 FILLER_167_64 ();
 b15zdnd11an1n16x5 FILLER_167_105 ();
 b15zdnd11an1n04x5 FILLER_167_121 ();
 b15zdnd00an1n02x5 FILLER_167_125 ();
 b15zdnd11an1n64x5 FILLER_167_138 ();
 b15zdnd11an1n64x5 FILLER_167_202 ();
 b15zdnd11an1n16x5 FILLER_167_266 ();
 b15zdnd11an1n08x5 FILLER_167_282 ();
 b15zdnd00an1n01x5 FILLER_167_290 ();
 b15zdnd11an1n32x5 FILLER_167_297 ();
 b15zdnd11an1n04x5 FILLER_167_329 ();
 b15zdnd00an1n02x5 FILLER_167_333 ();
 b15zdnd11an1n32x5 FILLER_167_344 ();
 b15zdnd11an1n16x5 FILLER_167_376 ();
 b15zdnd00an1n02x5 FILLER_167_392 ();
 b15zdnd00an1n01x5 FILLER_167_394 ();
 b15zdnd11an1n04x5 FILLER_167_398 ();
 b15zdnd11an1n04x5 FILLER_167_405 ();
 b15zdnd11an1n64x5 FILLER_167_412 ();
 b15zdnd11an1n64x5 FILLER_167_476 ();
 b15zdnd11an1n16x5 FILLER_167_540 ();
 b15zdnd00an1n02x5 FILLER_167_556 ();
 b15zdnd11an1n64x5 FILLER_167_597 ();
 b15zdnd11an1n04x5 FILLER_167_661 ();
 b15zdnd00an1n02x5 FILLER_167_665 ();
 b15zdnd00an1n01x5 FILLER_167_667 ();
 b15zdnd11an1n64x5 FILLER_167_682 ();
 b15zdnd11an1n64x5 FILLER_167_746 ();
 b15zdnd11an1n32x5 FILLER_167_810 ();
 b15zdnd11an1n04x5 FILLER_167_842 ();
 b15zdnd00an1n02x5 FILLER_167_846 ();
 b15zdnd11an1n32x5 FILLER_167_852 ();
 b15zdnd11an1n08x5 FILLER_167_884 ();
 b15zdnd11an1n04x5 FILLER_167_892 ();
 b15zdnd00an1n02x5 FILLER_167_896 ();
 b15zdnd11an1n08x5 FILLER_167_904 ();
 b15zdnd00an1n02x5 FILLER_167_912 ();
 b15zdnd11an1n64x5 FILLER_167_918 ();
 b15zdnd11an1n64x5 FILLER_167_982 ();
 b15zdnd11an1n64x5 FILLER_167_1046 ();
 b15zdnd11an1n64x5 FILLER_167_1110 ();
 b15zdnd11an1n64x5 FILLER_167_1174 ();
 b15zdnd11an1n64x5 FILLER_167_1238 ();
 b15zdnd11an1n64x5 FILLER_167_1302 ();
 b15zdnd11an1n32x5 FILLER_167_1366 ();
 b15zdnd11an1n16x5 FILLER_167_1398 ();
 b15zdnd00an1n02x5 FILLER_167_1414 ();
 b15zdnd11an1n04x5 FILLER_167_1419 ();
 b15zdnd11an1n64x5 FILLER_167_1430 ();
 b15zdnd11an1n32x5 FILLER_167_1494 ();
 b15zdnd11an1n04x5 FILLER_167_1526 ();
 b15zdnd00an1n02x5 FILLER_167_1530 ();
 b15zdnd00an1n01x5 FILLER_167_1532 ();
 b15zdnd11an1n16x5 FILLER_167_1536 ();
 b15zdnd11an1n08x5 FILLER_167_1552 ();
 b15zdnd00an1n02x5 FILLER_167_1560 ();
 b15zdnd11an1n16x5 FILLER_167_1565 ();
 b15zdnd00an1n01x5 FILLER_167_1581 ();
 b15zdnd11an1n64x5 FILLER_167_1591 ();
 b15zdnd11an1n64x5 FILLER_167_1655 ();
 b15zdnd11an1n16x5 FILLER_167_1719 ();
 b15zdnd00an1n02x5 FILLER_167_1735 ();
 b15zdnd11an1n64x5 FILLER_167_1740 ();
 b15zdnd11an1n64x5 FILLER_167_1804 ();
 b15zdnd11an1n32x5 FILLER_167_1868 ();
 b15zdnd11an1n08x5 FILLER_167_1900 ();
 b15zdnd11an1n04x5 FILLER_167_1908 ();
 b15zdnd11an1n64x5 FILLER_167_1964 ();
 b15zdnd11an1n04x5 FILLER_167_2028 ();
 b15zdnd11an1n16x5 FILLER_167_2043 ();
 b15zdnd00an1n01x5 FILLER_167_2059 ();
 b15zdnd11an1n64x5 FILLER_167_2063 ();
 b15zdnd11an1n64x5 FILLER_167_2127 ();
 b15zdnd11an1n64x5 FILLER_167_2191 ();
 b15zdnd11an1n16x5 FILLER_167_2255 ();
 b15zdnd11an1n08x5 FILLER_167_2271 ();
 b15zdnd11an1n04x5 FILLER_167_2279 ();
 b15zdnd00an1n01x5 FILLER_167_2283 ();
 b15zdnd11an1n32x5 FILLER_168_8 ();
 b15zdnd11an1n16x5 FILLER_168_40 ();
 b15zdnd11an1n08x5 FILLER_168_56 ();
 b15zdnd11an1n04x5 FILLER_168_64 ();
 b15zdnd00an1n02x5 FILLER_168_68 ();
 b15zdnd11an1n64x5 FILLER_168_74 ();
 b15zdnd11an1n64x5 FILLER_168_138 ();
 b15zdnd11an1n64x5 FILLER_168_202 ();
 b15zdnd11an1n64x5 FILLER_168_266 ();
 b15zdnd00an1n02x5 FILLER_168_330 ();
 b15zdnd11an1n32x5 FILLER_168_340 ();
 b15zdnd11an1n04x5 FILLER_168_372 ();
 b15zdnd00an1n02x5 FILLER_168_376 ();
 b15zdnd00an1n01x5 FILLER_168_378 ();
 b15zdnd11an1n64x5 FILLER_168_421 ();
 b15zdnd11an1n04x5 FILLER_168_485 ();
 b15zdnd00an1n02x5 FILLER_168_489 ();
 b15zdnd00an1n01x5 FILLER_168_491 ();
 b15zdnd11an1n08x5 FILLER_168_495 ();
 b15zdnd11an1n04x5 FILLER_168_503 ();
 b15zdnd00an1n01x5 FILLER_168_507 ();
 b15zdnd11an1n32x5 FILLER_168_529 ();
 b15zdnd11an1n16x5 FILLER_168_561 ();
 b15zdnd00an1n01x5 FILLER_168_577 ();
 b15zdnd11an1n64x5 FILLER_168_584 ();
 b15zdnd11an1n64x5 FILLER_168_648 ();
 b15zdnd11an1n04x5 FILLER_168_712 ();
 b15zdnd00an1n02x5 FILLER_168_716 ();
 b15zdnd11an1n64x5 FILLER_168_726 ();
 b15zdnd11an1n08x5 FILLER_168_790 ();
 b15zdnd11an1n04x5 FILLER_168_798 ();
 b15zdnd00an1n01x5 FILLER_168_802 ();
 b15zdnd11an1n32x5 FILLER_168_807 ();
 b15zdnd11an1n16x5 FILLER_168_839 ();
 b15zdnd11an1n04x5 FILLER_168_855 ();
 b15zdnd00an1n02x5 FILLER_168_859 ();
 b15zdnd11an1n32x5 FILLER_168_867 ();
 b15zdnd00an1n02x5 FILLER_168_899 ();
 b15zdnd11an1n64x5 FILLER_168_907 ();
 b15zdnd11an1n64x5 FILLER_168_971 ();
 b15zdnd11an1n16x5 FILLER_168_1035 ();
 b15zdnd00an1n01x5 FILLER_168_1051 ();
 b15zdnd11an1n08x5 FILLER_168_1064 ();
 b15zdnd11an1n64x5 FILLER_168_1079 ();
 b15zdnd11an1n64x5 FILLER_168_1143 ();
 b15zdnd11an1n64x5 FILLER_168_1207 ();
 b15zdnd11an1n64x5 FILLER_168_1271 ();
 b15zdnd11an1n32x5 FILLER_168_1335 ();
 b15zdnd11an1n16x5 FILLER_168_1367 ();
 b15zdnd11an1n08x5 FILLER_168_1383 ();
 b15zdnd11an1n04x5 FILLER_168_1391 ();
 b15zdnd11an1n32x5 FILLER_168_1447 ();
 b15zdnd11an1n16x5 FILLER_168_1479 ();
 b15zdnd11an1n08x5 FILLER_168_1495 ();
 b15zdnd00an1n02x5 FILLER_168_1503 ();
 b15zdnd00an1n01x5 FILLER_168_1505 ();
 b15zdnd11an1n08x5 FILLER_168_1558 ();
 b15zdnd11an1n04x5 FILLER_168_1566 ();
 b15zdnd00an1n02x5 FILLER_168_1570 ();
 b15zdnd11an1n64x5 FILLER_168_1614 ();
 b15zdnd11an1n64x5 FILLER_168_1678 ();
 b15zdnd11an1n64x5 FILLER_168_1742 ();
 b15zdnd11an1n64x5 FILLER_168_1806 ();
 b15zdnd11an1n32x5 FILLER_168_1870 ();
 b15zdnd11an1n16x5 FILLER_168_1902 ();
 b15zdnd11an1n08x5 FILLER_168_1918 ();
 b15zdnd11an1n04x5 FILLER_168_1926 ();
 b15zdnd11an1n04x5 FILLER_168_1933 ();
 b15zdnd11an1n64x5 FILLER_168_1940 ();
 b15zdnd11an1n32x5 FILLER_168_2004 ();
 b15zdnd11an1n16x5 FILLER_168_2036 ();
 b15zdnd11an1n08x5 FILLER_168_2052 ();
 b15zdnd11an1n64x5 FILLER_168_2063 ();
 b15zdnd11an1n16x5 FILLER_168_2127 ();
 b15zdnd11an1n08x5 FILLER_168_2143 ();
 b15zdnd00an1n02x5 FILLER_168_2151 ();
 b15zdnd00an1n01x5 FILLER_168_2153 ();
 b15zdnd11an1n32x5 FILLER_168_2162 ();
 b15zdnd11an1n16x5 FILLER_168_2194 ();
 b15zdnd00an1n01x5 FILLER_168_2210 ();
 b15zdnd11an1n16x5 FILLER_168_2223 ();
 b15zdnd11an1n04x5 FILLER_168_2239 ();
 b15zdnd00an1n02x5 FILLER_168_2243 ();
 b15zdnd11an1n16x5 FILLER_168_2257 ();
 b15zdnd00an1n02x5 FILLER_168_2273 ();
 b15zdnd00an1n01x5 FILLER_168_2275 ();
 b15zdnd11an1n64x5 FILLER_169_0 ();
 b15zdnd11an1n64x5 FILLER_169_64 ();
 b15zdnd11an1n64x5 FILLER_169_128 ();
 b15zdnd11an1n32x5 FILLER_169_192 ();
 b15zdnd11an1n08x5 FILLER_169_224 ();
 b15zdnd11an1n04x5 FILLER_169_232 ();
 b15zdnd11an1n64x5 FILLER_169_239 ();
 b15zdnd11an1n64x5 FILLER_169_303 ();
 b15zdnd11an1n04x5 FILLER_169_367 ();
 b15zdnd00an1n01x5 FILLER_169_371 ();
 b15zdnd11an1n16x5 FILLER_169_424 ();
 b15zdnd11an1n08x5 FILLER_169_440 ();
 b15zdnd11an1n04x5 FILLER_169_448 ();
 b15zdnd00an1n01x5 FILLER_169_452 ();
 b15zdnd11an1n64x5 FILLER_169_495 ();
 b15zdnd11an1n64x5 FILLER_169_559 ();
 b15zdnd11an1n64x5 FILLER_169_623 ();
 b15zdnd11an1n64x5 FILLER_169_687 ();
 b15zdnd11an1n16x5 FILLER_169_751 ();
 b15zdnd11an1n04x5 FILLER_169_767 ();
 b15zdnd00an1n01x5 FILLER_169_771 ();
 b15zdnd11an1n64x5 FILLER_169_776 ();
 b15zdnd11an1n64x5 FILLER_169_840 ();
 b15zdnd11an1n16x5 FILLER_169_904 ();
 b15zdnd11an1n04x5 FILLER_169_920 ();
 b15zdnd11an1n04x5 FILLER_169_936 ();
 b15zdnd11an1n08x5 FILLER_169_944 ();
 b15zdnd11an1n04x5 FILLER_169_952 ();
 b15zdnd11an1n32x5 FILLER_169_960 ();
 b15zdnd11an1n16x5 FILLER_169_992 ();
 b15zdnd11an1n04x5 FILLER_169_1008 ();
 b15zdnd11an1n04x5 FILLER_169_1043 ();
 b15zdnd11an1n04x5 FILLER_169_1059 ();
 b15zdnd11an1n64x5 FILLER_169_1070 ();
 b15zdnd11an1n64x5 FILLER_169_1134 ();
 b15zdnd11an1n64x5 FILLER_169_1198 ();
 b15zdnd11an1n64x5 FILLER_169_1262 ();
 b15zdnd11an1n08x5 FILLER_169_1326 ();
 b15zdnd11an1n04x5 FILLER_169_1334 ();
 b15zdnd00an1n01x5 FILLER_169_1338 ();
 b15zdnd11an1n64x5 FILLER_169_1343 ();
 b15zdnd11an1n08x5 FILLER_169_1407 ();
 b15zdnd00an1n02x5 FILLER_169_1415 ();
 b15zdnd00an1n01x5 FILLER_169_1417 ();
 b15zdnd11an1n64x5 FILLER_169_1434 ();
 b15zdnd11an1n16x5 FILLER_169_1498 ();
 b15zdnd11an1n08x5 FILLER_169_1514 ();
 b15zdnd00an1n02x5 FILLER_169_1522 ();
 b15zdnd00an1n01x5 FILLER_169_1524 ();
 b15zdnd11an1n04x5 FILLER_169_1528 ();
 b15zdnd11an1n16x5 FILLER_169_1535 ();
 b15zdnd11an1n08x5 FILLER_169_1551 ();
 b15zdnd11an1n04x5 FILLER_169_1559 ();
 b15zdnd11an1n16x5 FILLER_169_1566 ();
 b15zdnd11an1n08x5 FILLER_169_1582 ();
 b15zdnd00an1n02x5 FILLER_169_1590 ();
 b15zdnd00an1n01x5 FILLER_169_1592 ();
 b15zdnd11an1n64x5 FILLER_169_1602 ();
 b15zdnd11an1n64x5 FILLER_169_1666 ();
 b15zdnd11an1n64x5 FILLER_169_1730 ();
 b15zdnd11an1n64x5 FILLER_169_1794 ();
 b15zdnd11an1n32x5 FILLER_169_1858 ();
 b15zdnd11an1n08x5 FILLER_169_1890 ();
 b15zdnd00an1n02x5 FILLER_169_1898 ();
 b15zdnd00an1n01x5 FILLER_169_1900 ();
 b15zdnd11an1n64x5 FILLER_169_1912 ();
 b15zdnd11an1n32x5 FILLER_169_1976 ();
 b15zdnd11an1n08x5 FILLER_169_2008 ();
 b15zdnd11an1n04x5 FILLER_169_2016 ();
 b15zdnd11an1n08x5 FILLER_169_2026 ();
 b15zdnd00an1n02x5 FILLER_169_2034 ();
 b15zdnd11an1n64x5 FILLER_169_2088 ();
 b15zdnd00an1n01x5 FILLER_169_2152 ();
 b15zdnd11an1n16x5 FILLER_169_2179 ();
 b15zdnd11an1n08x5 FILLER_169_2195 ();
 b15zdnd11an1n04x5 FILLER_169_2203 ();
 b15zdnd00an1n01x5 FILLER_169_2207 ();
 b15zdnd11an1n32x5 FILLER_169_2245 ();
 b15zdnd11an1n04x5 FILLER_169_2277 ();
 b15zdnd00an1n02x5 FILLER_169_2281 ();
 b15zdnd00an1n01x5 FILLER_169_2283 ();
 b15zdnd11an1n64x5 FILLER_170_8 ();
 b15zdnd11an1n08x5 FILLER_170_72 ();
 b15zdnd00an1n02x5 FILLER_170_80 ();
 b15zdnd00an1n01x5 FILLER_170_82 ();
 b15zdnd11an1n64x5 FILLER_170_89 ();
 b15zdnd11an1n32x5 FILLER_170_153 ();
 b15zdnd11an1n16x5 FILLER_170_193 ();
 b15zdnd11an1n64x5 FILLER_170_261 ();
 b15zdnd11an1n08x5 FILLER_170_325 ();
 b15zdnd00an1n01x5 FILLER_170_333 ();
 b15zdnd11an1n64x5 FILLER_170_376 ();
 b15zdnd11an1n64x5 FILLER_170_440 ();
 b15zdnd11an1n64x5 FILLER_170_504 ();
 b15zdnd11an1n16x5 FILLER_170_568 ();
 b15zdnd11an1n04x5 FILLER_170_584 ();
 b15zdnd00an1n01x5 FILLER_170_588 ();
 b15zdnd11an1n64x5 FILLER_170_597 ();
 b15zdnd11an1n32x5 FILLER_170_661 ();
 b15zdnd11an1n16x5 FILLER_170_693 ();
 b15zdnd11an1n08x5 FILLER_170_709 ();
 b15zdnd00an1n01x5 FILLER_170_717 ();
 b15zdnd11an1n64x5 FILLER_170_726 ();
 b15zdnd11an1n64x5 FILLER_170_790 ();
 b15zdnd11an1n64x5 FILLER_170_854 ();
 b15zdnd11an1n64x5 FILLER_170_918 ();
 b15zdnd11an1n08x5 FILLER_170_982 ();
 b15zdnd11an1n04x5 FILLER_170_990 ();
 b15zdnd00an1n02x5 FILLER_170_994 ();
 b15zdnd11an1n64x5 FILLER_170_1018 ();
 b15zdnd11an1n64x5 FILLER_170_1082 ();
 b15zdnd11an1n64x5 FILLER_170_1146 ();
 b15zdnd11an1n64x5 FILLER_170_1210 ();
 b15zdnd11an1n64x5 FILLER_170_1274 ();
 b15zdnd11an1n32x5 FILLER_170_1338 ();
 b15zdnd11an1n08x5 FILLER_170_1370 ();
 b15zdnd11an1n04x5 FILLER_170_1378 ();
 b15zdnd00an1n02x5 FILLER_170_1382 ();
 b15zdnd00an1n01x5 FILLER_170_1384 ();
 b15zdnd11an1n16x5 FILLER_170_1394 ();
 b15zdnd00an1n02x5 FILLER_170_1410 ();
 b15zdnd11an1n64x5 FILLER_170_1432 ();
 b15zdnd11an1n64x5 FILLER_170_1496 ();
 b15zdnd11an1n32x5 FILLER_170_1560 ();
 b15zdnd11an1n16x5 FILLER_170_1592 ();
 b15zdnd00an1n02x5 FILLER_170_1608 ();
 b15zdnd00an1n01x5 FILLER_170_1610 ();
 b15zdnd11an1n64x5 FILLER_170_1617 ();
 b15zdnd11an1n64x5 FILLER_170_1681 ();
 b15zdnd11an1n64x5 FILLER_170_1745 ();
 b15zdnd11an1n16x5 FILLER_170_1809 ();
 b15zdnd11an1n04x5 FILLER_170_1825 ();
 b15zdnd11an1n64x5 FILLER_170_1833 ();
 b15zdnd11an1n64x5 FILLER_170_1897 ();
 b15zdnd11an1n32x5 FILLER_170_1961 ();
 b15zdnd11an1n04x5 FILLER_170_1993 ();
 b15zdnd00an1n02x5 FILLER_170_1997 ();
 b15zdnd11an1n32x5 FILLER_170_2023 ();
 b15zdnd11an1n04x5 FILLER_170_2055 ();
 b15zdnd00an1n02x5 FILLER_170_2059 ();
 b15zdnd11an1n64x5 FILLER_170_2064 ();
 b15zdnd11an1n04x5 FILLER_170_2128 ();
 b15zdnd00an1n02x5 FILLER_170_2132 ();
 b15zdnd11an1n08x5 FILLER_170_2143 ();
 b15zdnd00an1n02x5 FILLER_170_2151 ();
 b15zdnd00an1n01x5 FILLER_170_2153 ();
 b15zdnd00an1n02x5 FILLER_170_2162 ();
 b15zdnd11an1n64x5 FILLER_170_2178 ();
 b15zdnd11an1n04x5 FILLER_170_2256 ();
 b15zdnd00an1n02x5 FILLER_170_2274 ();
 b15zdnd11an1n64x5 FILLER_171_0 ();
 b15zdnd11an1n64x5 FILLER_171_64 ();
 b15zdnd11an1n32x5 FILLER_171_128 ();
 b15zdnd00an1n02x5 FILLER_171_160 ();
 b15zdnd11an1n16x5 FILLER_171_169 ();
 b15zdnd11an1n08x5 FILLER_171_185 ();
 b15zdnd11an1n04x5 FILLER_171_193 ();
 b15zdnd00an1n02x5 FILLER_171_197 ();
 b15zdnd11an1n64x5 FILLER_171_241 ();
 b15zdnd11an1n64x5 FILLER_171_305 ();
 b15zdnd11an1n64x5 FILLER_171_369 ();
 b15zdnd11an1n64x5 FILLER_171_433 ();
 b15zdnd11an1n64x5 FILLER_171_497 ();
 b15zdnd11an1n16x5 FILLER_171_561 ();
 b15zdnd11an1n08x5 FILLER_171_577 ();
 b15zdnd00an1n02x5 FILLER_171_585 ();
 b15zdnd11an1n04x5 FILLER_171_627 ();
 b15zdnd11an1n64x5 FILLER_171_634 ();
 b15zdnd11an1n64x5 FILLER_171_698 ();
 b15zdnd00an1n01x5 FILLER_171_762 ();
 b15zdnd11an1n04x5 FILLER_171_767 ();
 b15zdnd11an1n64x5 FILLER_171_775 ();
 b15zdnd11an1n64x5 FILLER_171_839 ();
 b15zdnd11an1n64x5 FILLER_171_903 ();
 b15zdnd11an1n64x5 FILLER_171_967 ();
 b15zdnd11an1n16x5 FILLER_171_1031 ();
 b15zdnd11an1n08x5 FILLER_171_1047 ();
 b15zdnd00an1n01x5 FILLER_171_1055 ();
 b15zdnd11an1n64x5 FILLER_171_1060 ();
 b15zdnd11an1n64x5 FILLER_171_1124 ();
 b15zdnd11an1n64x5 FILLER_171_1188 ();
 b15zdnd11an1n64x5 FILLER_171_1252 ();
 b15zdnd11an1n64x5 FILLER_171_1316 ();
 b15zdnd11an1n16x5 FILLER_171_1380 ();
 b15zdnd11an1n08x5 FILLER_171_1396 ();
 b15zdnd11an1n04x5 FILLER_171_1404 ();
 b15zdnd00an1n02x5 FILLER_171_1408 ();
 b15zdnd00an1n01x5 FILLER_171_1410 ();
 b15zdnd11an1n64x5 FILLER_171_1453 ();
 b15zdnd11an1n64x5 FILLER_171_1517 ();
 b15zdnd11an1n64x5 FILLER_171_1581 ();
 b15zdnd11an1n64x5 FILLER_171_1645 ();
 b15zdnd11an1n64x5 FILLER_171_1709 ();
 b15zdnd11an1n32x5 FILLER_171_1773 ();
 b15zdnd11an1n16x5 FILLER_171_1805 ();
 b15zdnd11an1n08x5 FILLER_171_1821 ();
 b15zdnd11an1n04x5 FILLER_171_1829 ();
 b15zdnd00an1n02x5 FILLER_171_1833 ();
 b15zdnd00an1n01x5 FILLER_171_1835 ();
 b15zdnd11an1n64x5 FILLER_171_1847 ();
 b15zdnd11an1n08x5 FILLER_171_1911 ();
 b15zdnd11an1n04x5 FILLER_171_1919 ();
 b15zdnd00an1n02x5 FILLER_171_1923 ();
 b15zdnd00an1n01x5 FILLER_171_1925 ();
 b15zdnd11an1n64x5 FILLER_171_1940 ();
 b15zdnd11an1n16x5 FILLER_171_2004 ();
 b15zdnd11an1n08x5 FILLER_171_2020 ();
 b15zdnd00an1n02x5 FILLER_171_2028 ();
 b15zdnd11an1n64x5 FILLER_171_2054 ();
 b15zdnd11an1n08x5 FILLER_171_2118 ();
 b15zdnd00an1n01x5 FILLER_171_2126 ();
 b15zdnd11an1n04x5 FILLER_171_2139 ();
 b15zdnd11an1n64x5 FILLER_171_2148 ();
 b15zdnd11an1n32x5 FILLER_171_2212 ();
 b15zdnd00an1n02x5 FILLER_171_2244 ();
 b15zdnd11an1n04x5 FILLER_171_2258 ();
 b15zdnd00an1n02x5 FILLER_171_2282 ();
 b15zdnd11an1n08x5 FILLER_172_8 ();
 b15zdnd11an1n04x5 FILLER_172_16 ();
 b15zdnd00an1n01x5 FILLER_172_20 ();
 b15zdnd11an1n04x5 FILLER_172_25 ();
 b15zdnd11an1n32x5 FILLER_172_33 ();
 b15zdnd11an1n04x5 FILLER_172_65 ();
 b15zdnd00an1n01x5 FILLER_172_69 ();
 b15zdnd11an1n64x5 FILLER_172_84 ();
 b15zdnd11an1n64x5 FILLER_172_148 ();
 b15zdnd11an1n16x5 FILLER_172_212 ();
 b15zdnd11an1n04x5 FILLER_172_228 ();
 b15zdnd11an1n04x5 FILLER_172_235 ();
 b15zdnd11an1n64x5 FILLER_172_242 ();
 b15zdnd11an1n64x5 FILLER_172_306 ();
 b15zdnd11an1n64x5 FILLER_172_370 ();
 b15zdnd11an1n64x5 FILLER_172_434 ();
 b15zdnd11an1n64x5 FILLER_172_498 ();
 b15zdnd11an1n16x5 FILLER_172_562 ();
 b15zdnd11an1n08x5 FILLER_172_578 ();
 b15zdnd11an1n04x5 FILLER_172_586 ();
 b15zdnd11an1n04x5 FILLER_172_632 ();
 b15zdnd11an1n16x5 FILLER_172_639 ();
 b15zdnd11an1n04x5 FILLER_172_655 ();
 b15zdnd00an1n02x5 FILLER_172_659 ();
 b15zdnd11an1n32x5 FILLER_172_667 ();
 b15zdnd11an1n16x5 FILLER_172_699 ();
 b15zdnd00an1n02x5 FILLER_172_715 ();
 b15zdnd00an1n01x5 FILLER_172_717 ();
 b15zdnd11an1n64x5 FILLER_172_726 ();
 b15zdnd11an1n64x5 FILLER_172_790 ();
 b15zdnd11an1n64x5 FILLER_172_854 ();
 b15zdnd11an1n64x5 FILLER_172_918 ();
 b15zdnd11an1n64x5 FILLER_172_982 ();
 b15zdnd11an1n64x5 FILLER_172_1046 ();
 b15zdnd11an1n64x5 FILLER_172_1110 ();
 b15zdnd11an1n64x5 FILLER_172_1174 ();
 b15zdnd11an1n16x5 FILLER_172_1238 ();
 b15zdnd11an1n08x5 FILLER_172_1254 ();
 b15zdnd11an1n04x5 FILLER_172_1262 ();
 b15zdnd00an1n02x5 FILLER_172_1266 ();
 b15zdnd00an1n01x5 FILLER_172_1268 ();
 b15zdnd11an1n64x5 FILLER_172_1275 ();
 b15zdnd11an1n16x5 FILLER_172_1339 ();
 b15zdnd11an1n04x5 FILLER_172_1355 ();
 b15zdnd00an1n02x5 FILLER_172_1359 ();
 b15zdnd00an1n01x5 FILLER_172_1361 ();
 b15zdnd11an1n08x5 FILLER_172_1373 ();
 b15zdnd00an1n02x5 FILLER_172_1381 ();
 b15zdnd00an1n01x5 FILLER_172_1383 ();
 b15zdnd11an1n64x5 FILLER_172_1423 ();
 b15zdnd11an1n64x5 FILLER_172_1487 ();
 b15zdnd11an1n64x5 FILLER_172_1551 ();
 b15zdnd11an1n64x5 FILLER_172_1615 ();
 b15zdnd11an1n64x5 FILLER_172_1679 ();
 b15zdnd11an1n64x5 FILLER_172_1743 ();
 b15zdnd11an1n64x5 FILLER_172_1807 ();
 b15zdnd11an1n32x5 FILLER_172_1871 ();
 b15zdnd11an1n16x5 FILLER_172_1903 ();
 b15zdnd11an1n08x5 FILLER_172_1919 ();
 b15zdnd00an1n02x5 FILLER_172_1927 ();
 b15zdnd11an1n64x5 FILLER_172_1932 ();
 b15zdnd11an1n64x5 FILLER_172_1996 ();
 b15zdnd11an1n64x5 FILLER_172_2060 ();
 b15zdnd11an1n16x5 FILLER_172_2124 ();
 b15zdnd11an1n08x5 FILLER_172_2140 ();
 b15zdnd11an1n04x5 FILLER_172_2148 ();
 b15zdnd00an1n02x5 FILLER_172_2152 ();
 b15zdnd11an1n64x5 FILLER_172_2162 ();
 b15zdnd11an1n16x5 FILLER_172_2226 ();
 b15zdnd11an1n08x5 FILLER_172_2242 ();
 b15zdnd11an1n04x5 FILLER_172_2250 ();
 b15zdnd11an1n08x5 FILLER_172_2268 ();
 b15zdnd11an1n64x5 FILLER_173_0 ();
 b15zdnd11an1n64x5 FILLER_173_64 ();
 b15zdnd11an1n64x5 FILLER_173_128 ();
 b15zdnd11an1n64x5 FILLER_173_192 ();
 b15zdnd11an1n64x5 FILLER_173_256 ();
 b15zdnd11an1n64x5 FILLER_173_320 ();
 b15zdnd11an1n64x5 FILLER_173_384 ();
 b15zdnd11an1n64x5 FILLER_173_448 ();
 b15zdnd11an1n32x5 FILLER_173_512 ();
 b15zdnd00an1n01x5 FILLER_173_544 ();
 b15zdnd11an1n64x5 FILLER_173_550 ();
 b15zdnd11an1n16x5 FILLER_173_614 ();
 b15zdnd00an1n02x5 FILLER_173_630 ();
 b15zdnd11an1n64x5 FILLER_173_636 ();
 b15zdnd11an1n64x5 FILLER_173_700 ();
 b15zdnd11an1n64x5 FILLER_173_764 ();
 b15zdnd11an1n64x5 FILLER_173_828 ();
 b15zdnd11an1n64x5 FILLER_173_892 ();
 b15zdnd11an1n64x5 FILLER_173_956 ();
 b15zdnd11an1n64x5 FILLER_173_1020 ();
 b15zdnd11an1n64x5 FILLER_173_1084 ();
 b15zdnd11an1n64x5 FILLER_173_1148 ();
 b15zdnd11an1n64x5 FILLER_173_1212 ();
 b15zdnd11an1n64x5 FILLER_173_1276 ();
 b15zdnd11an1n04x5 FILLER_173_1340 ();
 b15zdnd00an1n02x5 FILLER_173_1344 ();
 b15zdnd00an1n01x5 FILLER_173_1346 ();
 b15zdnd11an1n08x5 FILLER_173_1355 ();
 b15zdnd11an1n04x5 FILLER_173_1363 ();
 b15zdnd00an1n02x5 FILLER_173_1367 ();
 b15zdnd11an1n64x5 FILLER_173_1378 ();
 b15zdnd11an1n32x5 FILLER_173_1442 ();
 b15zdnd11an1n16x5 FILLER_173_1488 ();
 b15zdnd11an1n08x5 FILLER_173_1504 ();
 b15zdnd00an1n01x5 FILLER_173_1512 ();
 b15zdnd11an1n64x5 FILLER_173_1527 ();
 b15zdnd11an1n16x5 FILLER_173_1591 ();
 b15zdnd11an1n64x5 FILLER_173_1621 ();
 b15zdnd11an1n64x5 FILLER_173_1685 ();
 b15zdnd11an1n64x5 FILLER_173_1749 ();
 b15zdnd11an1n64x5 FILLER_173_1813 ();
 b15zdnd11an1n16x5 FILLER_173_1877 ();
 b15zdnd11an1n08x5 FILLER_173_1893 ();
 b15zdnd11an1n04x5 FILLER_173_1901 ();
 b15zdnd00an1n02x5 FILLER_173_1905 ();
 b15zdnd11an1n64x5 FILLER_173_1959 ();
 b15zdnd11an1n64x5 FILLER_173_2023 ();
 b15zdnd11an1n64x5 FILLER_173_2087 ();
 b15zdnd11an1n64x5 FILLER_173_2151 ();
 b15zdnd11an1n64x5 FILLER_173_2215 ();
 b15zdnd11an1n04x5 FILLER_173_2279 ();
 b15zdnd00an1n01x5 FILLER_173_2283 ();
 b15zdnd11an1n64x5 FILLER_174_8 ();
 b15zdnd11an1n64x5 FILLER_174_72 ();
 b15zdnd11an1n64x5 FILLER_174_136 ();
 b15zdnd11an1n64x5 FILLER_174_200 ();
 b15zdnd11an1n64x5 FILLER_174_264 ();
 b15zdnd11an1n64x5 FILLER_174_328 ();
 b15zdnd11an1n64x5 FILLER_174_392 ();
 b15zdnd11an1n64x5 FILLER_174_456 ();
 b15zdnd11an1n64x5 FILLER_174_520 ();
 b15zdnd11an1n32x5 FILLER_174_584 ();
 b15zdnd11an1n08x5 FILLER_174_616 ();
 b15zdnd00an1n02x5 FILLER_174_624 ();
 b15zdnd11an1n64x5 FILLER_174_630 ();
 b15zdnd11an1n16x5 FILLER_174_694 ();
 b15zdnd11an1n08x5 FILLER_174_710 ();
 b15zdnd11an1n64x5 FILLER_174_726 ();
 b15zdnd11an1n64x5 FILLER_174_790 ();
 b15zdnd11an1n64x5 FILLER_174_854 ();
 b15zdnd11an1n64x5 FILLER_174_918 ();
 b15zdnd11an1n64x5 FILLER_174_982 ();
 b15zdnd11an1n64x5 FILLER_174_1046 ();
 b15zdnd11an1n64x5 FILLER_174_1110 ();
 b15zdnd11an1n64x5 FILLER_174_1174 ();
 b15zdnd11an1n64x5 FILLER_174_1238 ();
 b15zdnd11an1n64x5 FILLER_174_1302 ();
 b15zdnd11an1n04x5 FILLER_174_1366 ();
 b15zdnd00an1n02x5 FILLER_174_1370 ();
 b15zdnd11an1n04x5 FILLER_174_1379 ();
 b15zdnd00an1n02x5 FILLER_174_1383 ();
 b15zdnd00an1n01x5 FILLER_174_1385 ();
 b15zdnd11an1n04x5 FILLER_174_1431 ();
 b15zdnd11an1n64x5 FILLER_174_1442 ();
 b15zdnd11an1n64x5 FILLER_174_1506 ();
 b15zdnd11an1n64x5 FILLER_174_1570 ();
 b15zdnd11an1n64x5 FILLER_174_1634 ();
 b15zdnd11an1n64x5 FILLER_174_1698 ();
 b15zdnd11an1n64x5 FILLER_174_1762 ();
 b15zdnd11an1n64x5 FILLER_174_1826 ();
 b15zdnd11an1n32x5 FILLER_174_1890 ();
 b15zdnd11an1n04x5 FILLER_174_1922 ();
 b15zdnd11an1n04x5 FILLER_174_1929 ();
 b15zdnd11an1n04x5 FILLER_174_1936 ();
 b15zdnd00an1n01x5 FILLER_174_1940 ();
 b15zdnd11an1n64x5 FILLER_174_1948 ();
 b15zdnd11an1n64x5 FILLER_174_2012 ();
 b15zdnd11an1n64x5 FILLER_174_2076 ();
 b15zdnd11an1n08x5 FILLER_174_2140 ();
 b15zdnd11an1n04x5 FILLER_174_2148 ();
 b15zdnd00an1n02x5 FILLER_174_2152 ();
 b15zdnd11an1n64x5 FILLER_174_2162 ();
 b15zdnd11an1n32x5 FILLER_174_2226 ();
 b15zdnd11an1n16x5 FILLER_174_2258 ();
 b15zdnd00an1n02x5 FILLER_174_2274 ();
 b15zdnd11an1n64x5 FILLER_175_0 ();
 b15zdnd11an1n64x5 FILLER_175_64 ();
 b15zdnd11an1n64x5 FILLER_175_128 ();
 b15zdnd11an1n64x5 FILLER_175_192 ();
 b15zdnd11an1n08x5 FILLER_175_256 ();
 b15zdnd11an1n04x5 FILLER_175_264 ();
 b15zdnd00an1n02x5 FILLER_175_268 ();
 b15zdnd11an1n64x5 FILLER_175_273 ();
 b15zdnd11an1n64x5 FILLER_175_337 ();
 b15zdnd11an1n64x5 FILLER_175_401 ();
 b15zdnd11an1n64x5 FILLER_175_465 ();
 b15zdnd11an1n64x5 FILLER_175_529 ();
 b15zdnd11an1n64x5 FILLER_175_593 ();
 b15zdnd11an1n64x5 FILLER_175_657 ();
 b15zdnd11an1n64x5 FILLER_175_721 ();
 b15zdnd11an1n64x5 FILLER_175_785 ();
 b15zdnd11an1n64x5 FILLER_175_849 ();
 b15zdnd11an1n64x5 FILLER_175_913 ();
 b15zdnd11an1n32x5 FILLER_175_977 ();
 b15zdnd11an1n16x5 FILLER_175_1009 ();
 b15zdnd11an1n08x5 FILLER_175_1025 ();
 b15zdnd11an1n04x5 FILLER_175_1033 ();
 b15zdnd00an1n02x5 FILLER_175_1037 ();
 b15zdnd00an1n01x5 FILLER_175_1039 ();
 b15zdnd11an1n64x5 FILLER_175_1044 ();
 b15zdnd11an1n64x5 FILLER_175_1108 ();
 b15zdnd11an1n64x5 FILLER_175_1172 ();
 b15zdnd11an1n64x5 FILLER_175_1236 ();
 b15zdnd11an1n64x5 FILLER_175_1300 ();
 b15zdnd11an1n64x5 FILLER_175_1364 ();
 b15zdnd11an1n64x5 FILLER_175_1428 ();
 b15zdnd11an1n32x5 FILLER_175_1492 ();
 b15zdnd00an1n01x5 FILLER_175_1524 ();
 b15zdnd11an1n04x5 FILLER_175_1534 ();
 b15zdnd11an1n16x5 FILLER_175_1549 ();
 b15zdnd11an1n08x5 FILLER_175_1565 ();
 b15zdnd00an1n02x5 FILLER_175_1573 ();
 b15zdnd11an1n32x5 FILLER_175_1584 ();
 b15zdnd11an1n16x5 FILLER_175_1616 ();
 b15zdnd11an1n08x5 FILLER_175_1632 ();
 b15zdnd00an1n01x5 FILLER_175_1640 ();
 b15zdnd11an1n32x5 FILLER_175_1661 ();
 b15zdnd11an1n16x5 FILLER_175_1693 ();
 b15zdnd11an1n08x5 FILLER_175_1709 ();
 b15zdnd11an1n04x5 FILLER_175_1717 ();
 b15zdnd00an1n02x5 FILLER_175_1721 ();
 b15zdnd11an1n64x5 FILLER_175_1731 ();
 b15zdnd11an1n64x5 FILLER_175_1795 ();
 b15zdnd11an1n64x5 FILLER_175_1859 ();
 b15zdnd11an1n64x5 FILLER_175_1923 ();
 b15zdnd11an1n64x5 FILLER_175_1987 ();
 b15zdnd11an1n64x5 FILLER_175_2057 ();
 b15zdnd11an1n64x5 FILLER_175_2121 ();
 b15zdnd11an1n16x5 FILLER_175_2185 ();
 b15zdnd00an1n02x5 FILLER_175_2201 ();
 b15zdnd00an1n01x5 FILLER_175_2203 ();
 b15zdnd11an1n64x5 FILLER_175_2218 ();
 b15zdnd00an1n02x5 FILLER_175_2282 ();
 b15zdnd11an1n32x5 FILLER_176_8 ();
 b15zdnd11an1n16x5 FILLER_176_40 ();
 b15zdnd11an1n08x5 FILLER_176_56 ();
 b15zdnd11an1n04x5 FILLER_176_64 ();
 b15zdnd00an1n02x5 FILLER_176_68 ();
 b15zdnd00an1n01x5 FILLER_176_70 ();
 b15zdnd11an1n64x5 FILLER_176_77 ();
 b15zdnd11an1n64x5 FILLER_176_141 ();
 b15zdnd11an1n32x5 FILLER_176_205 ();
 b15zdnd11an1n04x5 FILLER_176_237 ();
 b15zdnd00an1n02x5 FILLER_176_241 ();
 b15zdnd11an1n64x5 FILLER_176_295 ();
 b15zdnd11an1n64x5 FILLER_176_359 ();
 b15zdnd11an1n64x5 FILLER_176_423 ();
 b15zdnd11an1n32x5 FILLER_176_487 ();
 b15zdnd11an1n64x5 FILLER_176_525 ();
 b15zdnd11an1n64x5 FILLER_176_589 ();
 b15zdnd11an1n64x5 FILLER_176_653 ();
 b15zdnd00an1n01x5 FILLER_176_717 ();
 b15zdnd11an1n64x5 FILLER_176_726 ();
 b15zdnd11an1n64x5 FILLER_176_790 ();
 b15zdnd11an1n16x5 FILLER_176_854 ();
 b15zdnd11an1n08x5 FILLER_176_870 ();
 b15zdnd11an1n64x5 FILLER_176_881 ();
 b15zdnd11an1n64x5 FILLER_176_945 ();
 b15zdnd11an1n64x5 FILLER_176_1009 ();
 b15zdnd11an1n64x5 FILLER_176_1073 ();
 b15zdnd11an1n64x5 FILLER_176_1137 ();
 b15zdnd11an1n64x5 FILLER_176_1201 ();
 b15zdnd11an1n64x5 FILLER_176_1265 ();
 b15zdnd11an1n64x5 FILLER_176_1329 ();
 b15zdnd11an1n64x5 FILLER_176_1393 ();
 b15zdnd11an1n64x5 FILLER_176_1457 ();
 b15zdnd11an1n32x5 FILLER_176_1521 ();
 b15zdnd11an1n16x5 FILLER_176_1553 ();
 b15zdnd11an1n32x5 FILLER_176_1591 ();
 b15zdnd11an1n16x5 FILLER_176_1623 ();
 b15zdnd11an1n64x5 FILLER_176_1655 ();
 b15zdnd11an1n64x5 FILLER_176_1719 ();
 b15zdnd11an1n64x5 FILLER_176_1783 ();
 b15zdnd11an1n32x5 FILLER_176_1847 ();
 b15zdnd11an1n04x5 FILLER_176_1879 ();
 b15zdnd11an1n64x5 FILLER_176_1894 ();
 b15zdnd11an1n64x5 FILLER_176_1958 ();
 b15zdnd11an1n16x5 FILLER_176_2022 ();
 b15zdnd11an1n04x5 FILLER_176_2038 ();
 b15zdnd00an1n01x5 FILLER_176_2042 ();
 b15zdnd11an1n32x5 FILLER_176_2057 ();
 b15zdnd11an1n16x5 FILLER_176_2089 ();
 b15zdnd11an1n08x5 FILLER_176_2105 ();
 b15zdnd00an1n02x5 FILLER_176_2113 ();
 b15zdnd11an1n16x5 FILLER_176_2127 ();
 b15zdnd11an1n08x5 FILLER_176_2143 ();
 b15zdnd00an1n02x5 FILLER_176_2151 ();
 b15zdnd00an1n01x5 FILLER_176_2153 ();
 b15zdnd11an1n32x5 FILLER_176_2162 ();
 b15zdnd00an1n01x5 FILLER_176_2194 ();
 b15zdnd11an1n32x5 FILLER_176_2209 ();
 b15zdnd11an1n08x5 FILLER_176_2241 ();
 b15zdnd11an1n04x5 FILLER_176_2249 ();
 b15zdnd00an1n02x5 FILLER_176_2253 ();
 b15zdnd00an1n01x5 FILLER_176_2255 ();
 b15zdnd11an1n16x5 FILLER_176_2260 ();
 b15zdnd11an1n64x5 FILLER_177_0 ();
 b15zdnd11an1n64x5 FILLER_177_64 ();
 b15zdnd11an1n64x5 FILLER_177_128 ();
 b15zdnd11an1n32x5 FILLER_177_192 ();
 b15zdnd11an1n04x5 FILLER_177_257 ();
 b15zdnd11an1n04x5 FILLER_177_264 ();
 b15zdnd11an1n64x5 FILLER_177_271 ();
 b15zdnd11an1n64x5 FILLER_177_335 ();
 b15zdnd11an1n64x5 FILLER_177_399 ();
 b15zdnd11an1n64x5 FILLER_177_463 ();
 b15zdnd11an1n64x5 FILLER_177_527 ();
 b15zdnd11an1n64x5 FILLER_177_591 ();
 b15zdnd11an1n64x5 FILLER_177_655 ();
 b15zdnd11an1n64x5 FILLER_177_719 ();
 b15zdnd11an1n64x5 FILLER_177_783 ();
 b15zdnd11an1n04x5 FILLER_177_847 ();
 b15zdnd00an1n02x5 FILLER_177_851 ();
 b15zdnd11an1n64x5 FILLER_177_905 ();
 b15zdnd11an1n64x5 FILLER_177_969 ();
 b15zdnd11an1n64x5 FILLER_177_1033 ();
 b15zdnd11an1n64x5 FILLER_177_1097 ();
 b15zdnd11an1n64x5 FILLER_177_1161 ();
 b15zdnd11an1n64x5 FILLER_177_1225 ();
 b15zdnd11an1n64x5 FILLER_177_1289 ();
 b15zdnd11an1n64x5 FILLER_177_1353 ();
 b15zdnd11an1n64x5 FILLER_177_1417 ();
 b15zdnd11an1n64x5 FILLER_177_1481 ();
 b15zdnd11an1n64x5 FILLER_177_1545 ();
 b15zdnd11an1n32x5 FILLER_177_1609 ();
 b15zdnd11an1n08x5 FILLER_177_1641 ();
 b15zdnd11an1n04x5 FILLER_177_1659 ();
 b15zdnd11an1n64x5 FILLER_177_1666 ();
 b15zdnd11an1n32x5 FILLER_177_1730 ();
 b15zdnd11an1n16x5 FILLER_177_1762 ();
 b15zdnd11an1n08x5 FILLER_177_1778 ();
 b15zdnd00an1n02x5 FILLER_177_1786 ();
 b15zdnd00an1n01x5 FILLER_177_1788 ();
 b15zdnd11an1n64x5 FILLER_177_1793 ();
 b15zdnd11an1n64x5 FILLER_177_1857 ();
 b15zdnd11an1n64x5 FILLER_177_1921 ();
 b15zdnd11an1n32x5 FILLER_177_1985 ();
 b15zdnd11an1n16x5 FILLER_177_2017 ();
 b15zdnd11an1n08x5 FILLER_177_2033 ();
 b15zdnd11an1n04x5 FILLER_177_2041 ();
 b15zdnd00an1n02x5 FILLER_177_2045 ();
 b15zdnd11an1n08x5 FILLER_177_2059 ();
 b15zdnd11an1n04x5 FILLER_177_2067 ();
 b15zdnd00an1n02x5 FILLER_177_2071 ();
 b15zdnd11an1n08x5 FILLER_177_2095 ();
 b15zdnd00an1n02x5 FILLER_177_2103 ();
 b15zdnd00an1n01x5 FILLER_177_2105 ();
 b15zdnd11an1n64x5 FILLER_177_2148 ();
 b15zdnd11an1n64x5 FILLER_177_2212 ();
 b15zdnd11an1n08x5 FILLER_177_2276 ();
 b15zdnd11an1n64x5 FILLER_178_8 ();
 b15zdnd11an1n64x5 FILLER_178_72 ();
 b15zdnd11an1n64x5 FILLER_178_136 ();
 b15zdnd11an1n64x5 FILLER_178_200 ();
 b15zdnd11an1n32x5 FILLER_178_264 ();
 b15zdnd11an1n08x5 FILLER_178_296 ();
 b15zdnd11an1n04x5 FILLER_178_304 ();
 b15zdnd11an1n64x5 FILLER_178_350 ();
 b15zdnd11an1n64x5 FILLER_178_414 ();
 b15zdnd11an1n64x5 FILLER_178_478 ();
 b15zdnd11an1n64x5 FILLER_178_542 ();
 b15zdnd11an1n32x5 FILLER_178_606 ();
 b15zdnd11an1n16x5 FILLER_178_638 ();
 b15zdnd11an1n08x5 FILLER_178_654 ();
 b15zdnd11an1n32x5 FILLER_178_666 ();
 b15zdnd11an1n16x5 FILLER_178_698 ();
 b15zdnd11an1n04x5 FILLER_178_714 ();
 b15zdnd11an1n64x5 FILLER_178_726 ();
 b15zdnd11an1n64x5 FILLER_178_790 ();
 b15zdnd11an1n16x5 FILLER_178_854 ();
 b15zdnd00an1n01x5 FILLER_178_870 ();
 b15zdnd11an1n64x5 FILLER_178_923 ();
 b15zdnd11an1n64x5 FILLER_178_987 ();
 b15zdnd11an1n64x5 FILLER_178_1051 ();
 b15zdnd11an1n64x5 FILLER_178_1115 ();
 b15zdnd11an1n64x5 FILLER_178_1179 ();
 b15zdnd11an1n64x5 FILLER_178_1243 ();
 b15zdnd11an1n64x5 FILLER_178_1307 ();
 b15zdnd11an1n64x5 FILLER_178_1371 ();
 b15zdnd11an1n64x5 FILLER_178_1435 ();
 b15zdnd11an1n64x5 FILLER_178_1499 ();
 b15zdnd11an1n64x5 FILLER_178_1563 ();
 b15zdnd11an1n16x5 FILLER_178_1627 ();
 b15zdnd11an1n08x5 FILLER_178_1643 ();
 b15zdnd00an1n02x5 FILLER_178_1651 ();
 b15zdnd11an1n04x5 FILLER_178_1656 ();
 b15zdnd11an1n64x5 FILLER_178_1670 ();
 b15zdnd11an1n64x5 FILLER_178_1734 ();
 b15zdnd11an1n64x5 FILLER_178_1798 ();
 b15zdnd11an1n64x5 FILLER_178_1862 ();
 b15zdnd11an1n64x5 FILLER_178_1926 ();
 b15zdnd11an1n64x5 FILLER_178_1990 ();
 b15zdnd11an1n64x5 FILLER_178_2054 ();
 b15zdnd11an1n32x5 FILLER_178_2118 ();
 b15zdnd11an1n04x5 FILLER_178_2150 ();
 b15zdnd11an1n32x5 FILLER_178_2162 ();
 b15zdnd11an1n16x5 FILLER_178_2194 ();
 b15zdnd00an1n01x5 FILLER_178_2210 ();
 b15zdnd11an1n32x5 FILLER_178_2217 ();
 b15zdnd11an1n16x5 FILLER_178_2249 ();
 b15zdnd11an1n08x5 FILLER_178_2265 ();
 b15zdnd00an1n02x5 FILLER_178_2273 ();
 b15zdnd00an1n01x5 FILLER_178_2275 ();
 b15zdnd11an1n64x5 FILLER_179_0 ();
 b15zdnd11an1n64x5 FILLER_179_64 ();
 b15zdnd11an1n64x5 FILLER_179_128 ();
 b15zdnd11an1n64x5 FILLER_179_192 ();
 b15zdnd11an1n64x5 FILLER_179_256 ();
 b15zdnd11an1n64x5 FILLER_179_320 ();
 b15zdnd11an1n64x5 FILLER_179_384 ();
 b15zdnd11an1n64x5 FILLER_179_448 ();
 b15zdnd11an1n64x5 FILLER_179_512 ();
 b15zdnd11an1n32x5 FILLER_179_576 ();
 b15zdnd11an1n08x5 FILLER_179_608 ();
 b15zdnd00an1n02x5 FILLER_179_616 ();
 b15zdnd11an1n16x5 FILLER_179_622 ();
 b15zdnd11an1n08x5 FILLER_179_638 ();
 b15zdnd00an1n02x5 FILLER_179_646 ();
 b15zdnd11an1n64x5 FILLER_179_652 ();
 b15zdnd11an1n32x5 FILLER_179_716 ();
 b15zdnd11an1n16x5 FILLER_179_748 ();
 b15zdnd11an1n08x5 FILLER_179_764 ();
 b15zdnd00an1n02x5 FILLER_179_772 ();
 b15zdnd11an1n64x5 FILLER_179_777 ();
 b15zdnd11an1n16x5 FILLER_179_841 ();
 b15zdnd11an1n08x5 FILLER_179_857 ();
 b15zdnd11an1n04x5 FILLER_179_865 ();
 b15zdnd00an1n02x5 FILLER_179_869 ();
 b15zdnd11an1n04x5 FILLER_179_874 ();
 b15zdnd11an1n08x5 FILLER_179_881 ();
 b15zdnd00an1n01x5 FILLER_179_889 ();
 b15zdnd11an1n04x5 FILLER_179_893 ();
 b15zdnd11an1n04x5 FILLER_179_900 ();
 b15zdnd00an1n02x5 FILLER_179_904 ();
 b15zdnd00an1n01x5 FILLER_179_906 ();
 b15zdnd11an1n64x5 FILLER_179_915 ();
 b15zdnd11an1n64x5 FILLER_179_979 ();
 b15zdnd11an1n64x5 FILLER_179_1043 ();
 b15zdnd11an1n64x5 FILLER_179_1146 ();
 b15zdnd11an1n64x5 FILLER_179_1210 ();
 b15zdnd11an1n08x5 FILLER_179_1274 ();
 b15zdnd11an1n04x5 FILLER_179_1282 ();
 b15zdnd00an1n01x5 FILLER_179_1286 ();
 b15zdnd11an1n64x5 FILLER_179_1291 ();
 b15zdnd11an1n64x5 FILLER_179_1355 ();
 b15zdnd11an1n64x5 FILLER_179_1419 ();
 b15zdnd11an1n64x5 FILLER_179_1483 ();
 b15zdnd11an1n64x5 FILLER_179_1547 ();
 b15zdnd11an1n64x5 FILLER_179_1611 ();
 b15zdnd11an1n64x5 FILLER_179_1675 ();
 b15zdnd11an1n64x5 FILLER_179_1739 ();
 b15zdnd11an1n64x5 FILLER_179_1803 ();
 b15zdnd11an1n64x5 FILLER_179_1867 ();
 b15zdnd11an1n64x5 FILLER_179_1931 ();
 b15zdnd11an1n16x5 FILLER_179_1995 ();
 b15zdnd11an1n08x5 FILLER_179_2011 ();
 b15zdnd00an1n01x5 FILLER_179_2019 ();
 b15zdnd11an1n64x5 FILLER_179_2031 ();
 b15zdnd11an1n64x5 FILLER_179_2095 ();
 b15zdnd11an1n16x5 FILLER_179_2159 ();
 b15zdnd11an1n04x5 FILLER_179_2175 ();
 b15zdnd00an1n01x5 FILLER_179_2179 ();
 b15zdnd11an1n16x5 FILLER_179_2206 ();
 b15zdnd00an1n01x5 FILLER_179_2222 ();
 b15zdnd11an1n16x5 FILLER_179_2249 ();
 b15zdnd11an1n08x5 FILLER_179_2269 ();
 b15zdnd11an1n04x5 FILLER_179_2277 ();
 b15zdnd00an1n02x5 FILLER_179_2281 ();
 b15zdnd00an1n01x5 FILLER_179_2283 ();
 b15zdnd11an1n64x5 FILLER_180_8 ();
 b15zdnd11an1n64x5 FILLER_180_72 ();
 b15zdnd11an1n64x5 FILLER_180_136 ();
 b15zdnd11an1n64x5 FILLER_180_200 ();
 b15zdnd11an1n64x5 FILLER_180_264 ();
 b15zdnd11an1n64x5 FILLER_180_328 ();
 b15zdnd11an1n32x5 FILLER_180_392 ();
 b15zdnd11an1n04x5 FILLER_180_424 ();
 b15zdnd00an1n01x5 FILLER_180_428 ();
 b15zdnd11an1n64x5 FILLER_180_436 ();
 b15zdnd11an1n64x5 FILLER_180_500 ();
 b15zdnd11an1n64x5 FILLER_180_564 ();
 b15zdnd11an1n64x5 FILLER_180_628 ();
 b15zdnd11an1n16x5 FILLER_180_692 ();
 b15zdnd11an1n08x5 FILLER_180_708 ();
 b15zdnd00an1n02x5 FILLER_180_716 ();
 b15zdnd11an1n16x5 FILLER_180_726 ();
 b15zdnd11an1n04x5 FILLER_180_742 ();
 b15zdnd00an1n01x5 FILLER_180_746 ();
 b15zdnd11an1n64x5 FILLER_180_799 ();
 b15zdnd11an1n32x5 FILLER_180_863 ();
 b15zdnd00an1n02x5 FILLER_180_895 ();
 b15zdnd00an1n01x5 FILLER_180_897 ();
 b15zdnd11an1n64x5 FILLER_180_901 ();
 b15zdnd11an1n64x5 FILLER_180_965 ();
 b15zdnd11an1n64x5 FILLER_180_1029 ();
 b15zdnd11an1n64x5 FILLER_180_1093 ();
 b15zdnd11an1n64x5 FILLER_180_1157 ();
 b15zdnd11an1n32x5 FILLER_180_1221 ();
 b15zdnd11an1n04x5 FILLER_180_1253 ();
 b15zdnd11an1n64x5 FILLER_180_1273 ();
 b15zdnd11an1n64x5 FILLER_180_1337 ();
 b15zdnd11an1n64x5 FILLER_180_1401 ();
 b15zdnd11an1n64x5 FILLER_180_1465 ();
 b15zdnd11an1n64x5 FILLER_180_1529 ();
 b15zdnd11an1n08x5 FILLER_180_1593 ();
 b15zdnd11an1n04x5 FILLER_180_1601 ();
 b15zdnd00an1n02x5 FILLER_180_1605 ();
 b15zdnd00an1n01x5 FILLER_180_1607 ();
 b15zdnd11an1n64x5 FILLER_180_1650 ();
 b15zdnd11an1n64x5 FILLER_180_1714 ();
 b15zdnd11an1n64x5 FILLER_180_1778 ();
 b15zdnd11an1n64x5 FILLER_180_1842 ();
 b15zdnd11an1n64x5 FILLER_180_1906 ();
 b15zdnd11an1n08x5 FILLER_180_1970 ();
 b15zdnd11an1n04x5 FILLER_180_1978 ();
 b15zdnd00an1n02x5 FILLER_180_1982 ();
 b15zdnd11an1n64x5 FILLER_180_2004 ();
 b15zdnd11an1n64x5 FILLER_180_2068 ();
 b15zdnd11an1n16x5 FILLER_180_2132 ();
 b15zdnd11an1n04x5 FILLER_180_2148 ();
 b15zdnd00an1n02x5 FILLER_180_2152 ();
 b15zdnd11an1n16x5 FILLER_180_2162 ();
 b15zdnd11an1n04x5 FILLER_180_2178 ();
 b15zdnd11an1n04x5 FILLER_180_2202 ();
 b15zdnd11an1n16x5 FILLER_180_2220 ();
 b15zdnd11an1n08x5 FILLER_180_2236 ();
 b15zdnd11an1n04x5 FILLER_180_2248 ();
 b15zdnd11an1n04x5 FILLER_180_2256 ();
 b15zdnd00an1n02x5 FILLER_180_2260 ();
 b15zdnd11an1n08x5 FILLER_180_2266 ();
 b15zdnd00an1n02x5 FILLER_180_2274 ();
 b15zdnd11an1n64x5 FILLER_181_0 ();
 b15zdnd11an1n32x5 FILLER_181_64 ();
 b15zdnd11an1n16x5 FILLER_181_96 ();
 b15zdnd11an1n08x5 FILLER_181_112 ();
 b15zdnd11an1n04x5 FILLER_181_120 ();
 b15zdnd00an1n02x5 FILLER_181_124 ();
 b15zdnd11an1n04x5 FILLER_181_129 ();
 b15zdnd11an1n04x5 FILLER_181_140 ();
 b15zdnd11an1n64x5 FILLER_181_151 ();
 b15zdnd11an1n64x5 FILLER_181_215 ();
 b15zdnd11an1n64x5 FILLER_181_279 ();
 b15zdnd11an1n64x5 FILLER_181_343 ();
 b15zdnd11an1n64x5 FILLER_181_407 ();
 b15zdnd11an1n64x5 FILLER_181_471 ();
 b15zdnd11an1n64x5 FILLER_181_535 ();
 b15zdnd11an1n64x5 FILLER_181_599 ();
 b15zdnd11an1n64x5 FILLER_181_663 ();
 b15zdnd00an1n02x5 FILLER_181_727 ();
 b15zdnd11an1n08x5 FILLER_181_737 ();
 b15zdnd11an1n64x5 FILLER_181_797 ();
 b15zdnd11an1n64x5 FILLER_181_861 ();
 b15zdnd11an1n64x5 FILLER_181_925 ();
 b15zdnd11an1n64x5 FILLER_181_989 ();
 b15zdnd11an1n64x5 FILLER_181_1053 ();
 b15zdnd11an1n64x5 FILLER_181_1117 ();
 b15zdnd11an1n32x5 FILLER_181_1181 ();
 b15zdnd11an1n16x5 FILLER_181_1213 ();
 b15zdnd11an1n04x5 FILLER_181_1229 ();
 b15zdnd00an1n02x5 FILLER_181_1233 ();
 b15zdnd00an1n01x5 FILLER_181_1235 ();
 b15zdnd11an1n64x5 FILLER_181_1240 ();
 b15zdnd11an1n64x5 FILLER_181_1304 ();
 b15zdnd11an1n32x5 FILLER_181_1368 ();
 b15zdnd11an1n04x5 FILLER_181_1400 ();
 b15zdnd00an1n01x5 FILLER_181_1404 ();
 b15zdnd11an1n16x5 FILLER_181_1429 ();
 b15zdnd11an1n08x5 FILLER_181_1445 ();
 b15zdnd11an1n04x5 FILLER_181_1453 ();
 b15zdnd00an1n01x5 FILLER_181_1457 ();
 b15zdnd11an1n64x5 FILLER_181_1478 ();
 b15zdnd11an1n64x5 FILLER_181_1542 ();
 b15zdnd11an1n64x5 FILLER_181_1606 ();
 b15zdnd11an1n32x5 FILLER_181_1670 ();
 b15zdnd11an1n16x5 FILLER_181_1702 ();
 b15zdnd11an1n08x5 FILLER_181_1718 ();
 b15zdnd00an1n02x5 FILLER_181_1726 ();
 b15zdnd00an1n01x5 FILLER_181_1728 ();
 b15zdnd11an1n32x5 FILLER_181_1733 ();
 b15zdnd11an1n08x5 FILLER_181_1765 ();
 b15zdnd00an1n02x5 FILLER_181_1773 ();
 b15zdnd11an1n64x5 FILLER_181_1817 ();
 b15zdnd11an1n64x5 FILLER_181_1881 ();
 b15zdnd11an1n64x5 FILLER_181_1945 ();
 b15zdnd11an1n64x5 FILLER_181_2009 ();
 b15zdnd11an1n64x5 FILLER_181_2073 ();
 b15zdnd11an1n64x5 FILLER_181_2137 ();
 b15zdnd11an1n32x5 FILLER_181_2201 ();
 b15zdnd11an1n04x5 FILLER_181_2233 ();
 b15zdnd00an1n02x5 FILLER_181_2237 ();
 b15zdnd00an1n01x5 FILLER_181_2239 ();
 b15zdnd00an1n02x5 FILLER_181_2282 ();
 b15zdnd11an1n32x5 FILLER_182_8 ();
 b15zdnd00an1n02x5 FILLER_182_40 ();
 b15zdnd11an1n16x5 FILLER_182_57 ();
 b15zdnd00an1n01x5 FILLER_182_73 ();
 b15zdnd11an1n04x5 FILLER_182_119 ();
 b15zdnd11an1n04x5 FILLER_182_126 ();
 b15zdnd11an1n16x5 FILLER_182_133 ();
 b15zdnd11an1n64x5 FILLER_182_191 ();
 b15zdnd11an1n64x5 FILLER_182_255 ();
 b15zdnd11an1n64x5 FILLER_182_319 ();
 b15zdnd11an1n64x5 FILLER_182_383 ();
 b15zdnd11an1n32x5 FILLER_182_447 ();
 b15zdnd11an1n08x5 FILLER_182_479 ();
 b15zdnd00an1n02x5 FILLER_182_487 ();
 b15zdnd11an1n64x5 FILLER_182_492 ();
 b15zdnd11an1n64x5 FILLER_182_556 ();
 b15zdnd11an1n64x5 FILLER_182_620 ();
 b15zdnd11an1n32x5 FILLER_182_684 ();
 b15zdnd00an1n02x5 FILLER_182_716 ();
 b15zdnd11an1n32x5 FILLER_182_726 ();
 b15zdnd11an1n04x5 FILLER_182_758 ();
 b15zdnd00an1n02x5 FILLER_182_762 ();
 b15zdnd00an1n01x5 FILLER_182_764 ();
 b15zdnd11an1n04x5 FILLER_182_768 ();
 b15zdnd11an1n04x5 FILLER_182_775 ();
 b15zdnd11an1n64x5 FILLER_182_782 ();
 b15zdnd11an1n64x5 FILLER_182_846 ();
 b15zdnd11an1n64x5 FILLER_182_910 ();
 b15zdnd11an1n64x5 FILLER_182_974 ();
 b15zdnd11an1n64x5 FILLER_182_1038 ();
 b15zdnd11an1n64x5 FILLER_182_1102 ();
 b15zdnd11an1n64x5 FILLER_182_1166 ();
 b15zdnd11an1n08x5 FILLER_182_1230 ();
 b15zdnd00an1n02x5 FILLER_182_1238 ();
 b15zdnd00an1n01x5 FILLER_182_1240 ();
 b15zdnd11an1n64x5 FILLER_182_1245 ();
 b15zdnd11an1n32x5 FILLER_182_1309 ();
 b15zdnd11an1n04x5 FILLER_182_1341 ();
 b15zdnd00an1n02x5 FILLER_182_1345 ();
 b15zdnd00an1n01x5 FILLER_182_1347 ();
 b15zdnd11an1n64x5 FILLER_182_1364 ();
 b15zdnd11an1n64x5 FILLER_182_1428 ();
 b15zdnd11an1n64x5 FILLER_182_1492 ();
 b15zdnd11an1n64x5 FILLER_182_1556 ();
 b15zdnd11an1n64x5 FILLER_182_1620 ();
 b15zdnd11an1n64x5 FILLER_182_1684 ();
 b15zdnd11an1n64x5 FILLER_182_1748 ();
 b15zdnd11an1n64x5 FILLER_182_1812 ();
 b15zdnd11an1n64x5 FILLER_182_1876 ();
 b15zdnd11an1n64x5 FILLER_182_1940 ();
 b15zdnd11an1n64x5 FILLER_182_2004 ();
 b15zdnd11an1n32x5 FILLER_182_2068 ();
 b15zdnd11an1n16x5 FILLER_182_2100 ();
 b15zdnd11an1n08x5 FILLER_182_2116 ();
 b15zdnd11an1n04x5 FILLER_182_2124 ();
 b15zdnd00an1n01x5 FILLER_182_2128 ();
 b15zdnd11an1n08x5 FILLER_182_2146 ();
 b15zdnd11an1n64x5 FILLER_182_2162 ();
 b15zdnd11an1n32x5 FILLER_182_2226 ();
 b15zdnd11an1n16x5 FILLER_182_2258 ();
 b15zdnd00an1n02x5 FILLER_182_2274 ();
 b15zdnd11an1n64x5 FILLER_183_0 ();
 b15zdnd11an1n16x5 FILLER_183_64 ();
 b15zdnd11an1n04x5 FILLER_183_80 ();
 b15zdnd00an1n01x5 FILLER_183_84 ();
 b15zdnd11an1n08x5 FILLER_183_92 ();
 b15zdnd00an1n02x5 FILLER_183_100 ();
 b15zdnd00an1n01x5 FILLER_183_102 ();
 b15zdnd11an1n64x5 FILLER_183_155 ();
 b15zdnd11an1n64x5 FILLER_183_219 ();
 b15zdnd11an1n64x5 FILLER_183_283 ();
 b15zdnd11an1n64x5 FILLER_183_347 ();
 b15zdnd11an1n32x5 FILLER_183_411 ();
 b15zdnd11an1n16x5 FILLER_183_443 ();
 b15zdnd11an1n04x5 FILLER_183_459 ();
 b15zdnd00an1n02x5 FILLER_183_463 ();
 b15zdnd00an1n01x5 FILLER_183_465 ();
 b15zdnd11an1n64x5 FILLER_183_508 ();
 b15zdnd11an1n64x5 FILLER_183_572 ();
 b15zdnd11an1n64x5 FILLER_183_636 ();
 b15zdnd11an1n64x5 FILLER_183_700 ();
 b15zdnd00an1n02x5 FILLER_183_764 ();
 b15zdnd11an1n04x5 FILLER_183_769 ();
 b15zdnd11an1n16x5 FILLER_183_776 ();
 b15zdnd00an1n02x5 FILLER_183_792 ();
 b15zdnd11an1n32x5 FILLER_183_803 ();
 b15zdnd11an1n08x5 FILLER_183_835 ();
 b15zdnd11an1n04x5 FILLER_183_843 ();
 b15zdnd00an1n02x5 FILLER_183_847 ();
 b15zdnd11an1n64x5 FILLER_183_858 ();
 b15zdnd11an1n64x5 FILLER_183_922 ();
 b15zdnd11an1n64x5 FILLER_183_986 ();
 b15zdnd11an1n64x5 FILLER_183_1050 ();
 b15zdnd11an1n64x5 FILLER_183_1114 ();
 b15zdnd11an1n32x5 FILLER_183_1178 ();
 b15zdnd11an1n04x5 FILLER_183_1210 ();
 b15zdnd00an1n02x5 FILLER_183_1214 ();
 b15zdnd00an1n01x5 FILLER_183_1216 ();
 b15zdnd11an1n16x5 FILLER_183_1228 ();
 b15zdnd11an1n08x5 FILLER_183_1244 ();
 b15zdnd00an1n02x5 FILLER_183_1252 ();
 b15zdnd00an1n01x5 FILLER_183_1254 ();
 b15zdnd11an1n32x5 FILLER_183_1261 ();
 b15zdnd11an1n16x5 FILLER_183_1293 ();
 b15zdnd11an1n04x5 FILLER_183_1309 ();
 b15zdnd00an1n01x5 FILLER_183_1313 ();
 b15zdnd11an1n64x5 FILLER_183_1322 ();
 b15zdnd11an1n32x5 FILLER_183_1386 ();
 b15zdnd11an1n16x5 FILLER_183_1418 ();
 b15zdnd00an1n01x5 FILLER_183_1434 ();
 b15zdnd11an1n04x5 FILLER_183_1446 ();
 b15zdnd00an1n02x5 FILLER_183_1450 ();
 b15zdnd00an1n01x5 FILLER_183_1452 ();
 b15zdnd11an1n64x5 FILLER_183_1480 ();
 b15zdnd11an1n64x5 FILLER_183_1544 ();
 b15zdnd11an1n64x5 FILLER_183_1608 ();
 b15zdnd11an1n64x5 FILLER_183_1672 ();
 b15zdnd11an1n64x5 FILLER_183_1736 ();
 b15zdnd11an1n32x5 FILLER_183_1800 ();
 b15zdnd00an1n02x5 FILLER_183_1832 ();
 b15zdnd00an1n01x5 FILLER_183_1834 ();
 b15zdnd11an1n16x5 FILLER_183_1855 ();
 b15zdnd00an1n01x5 FILLER_183_1871 ();
 b15zdnd11an1n04x5 FILLER_183_1875 ();
 b15zdnd11an1n64x5 FILLER_183_1882 ();
 b15zdnd11an1n64x5 FILLER_183_1946 ();
 b15zdnd11an1n64x5 FILLER_183_2010 ();
 b15zdnd11an1n16x5 FILLER_183_2074 ();
 b15zdnd11an1n04x5 FILLER_183_2090 ();
 b15zdnd00an1n02x5 FILLER_183_2094 ();
 b15zdnd11an1n64x5 FILLER_183_2121 ();
 b15zdnd11an1n08x5 FILLER_183_2185 ();
 b15zdnd00an1n02x5 FILLER_183_2193 ();
 b15zdnd00an1n01x5 FILLER_183_2195 ();
 b15zdnd11an1n32x5 FILLER_183_2202 ();
 b15zdnd11an1n16x5 FILLER_183_2234 ();
 b15zdnd11an1n04x5 FILLER_183_2250 ();
 b15zdnd00an1n02x5 FILLER_183_2254 ();
 b15zdnd11an1n16x5 FILLER_183_2267 ();
 b15zdnd00an1n01x5 FILLER_183_2283 ();
 b15zdnd11an1n32x5 FILLER_184_8 ();
 b15zdnd11an1n16x5 FILLER_184_40 ();
 b15zdnd11an1n08x5 FILLER_184_56 ();
 b15zdnd11an1n04x5 FILLER_184_64 ();
 b15zdnd00an1n01x5 FILLER_184_68 ();
 b15zdnd11an1n04x5 FILLER_184_100 ();
 b15zdnd11an1n64x5 FILLER_184_156 ();
 b15zdnd11an1n16x5 FILLER_184_220 ();
 b15zdnd11an1n08x5 FILLER_184_236 ();
 b15zdnd11an1n04x5 FILLER_184_244 ();
 b15zdnd11an1n64x5 FILLER_184_290 ();
 b15zdnd11an1n16x5 FILLER_184_385 ();
 b15zdnd00an1n02x5 FILLER_184_401 ();
 b15zdnd11an1n04x5 FILLER_184_414 ();
 b15zdnd11an1n16x5 FILLER_184_432 ();
 b15zdnd11an1n08x5 FILLER_184_448 ();
 b15zdnd00an1n02x5 FILLER_184_456 ();
 b15zdnd00an1n01x5 FILLER_184_458 ();
 b15zdnd11an1n04x5 FILLER_184_466 ();
 b15zdnd00an1n02x5 FILLER_184_470 ();
 b15zdnd11an1n04x5 FILLER_184_476 ();
 b15zdnd00an1n02x5 FILLER_184_480 ();
 b15zdnd11an1n64x5 FILLER_184_524 ();
 b15zdnd11an1n64x5 FILLER_184_588 ();
 b15zdnd11an1n64x5 FILLER_184_652 ();
 b15zdnd00an1n02x5 FILLER_184_716 ();
 b15zdnd11an1n64x5 FILLER_184_726 ();
 b15zdnd11an1n64x5 FILLER_184_790 ();
 b15zdnd11an1n64x5 FILLER_184_854 ();
 b15zdnd11an1n64x5 FILLER_184_918 ();
 b15zdnd11an1n64x5 FILLER_184_982 ();
 b15zdnd11an1n04x5 FILLER_184_1046 ();
 b15zdnd00an1n01x5 FILLER_184_1050 ();
 b15zdnd11an1n04x5 FILLER_184_1054 ();
 b15zdnd11an1n64x5 FILLER_184_1061 ();
 b15zdnd11an1n32x5 FILLER_184_1125 ();
 b15zdnd11an1n16x5 FILLER_184_1157 ();
 b15zdnd11an1n08x5 FILLER_184_1173 ();
 b15zdnd11an1n04x5 FILLER_184_1184 ();
 b15zdnd11an1n64x5 FILLER_184_1191 ();
 b15zdnd00an1n02x5 FILLER_184_1255 ();
 b15zdnd11an1n32x5 FILLER_184_1271 ();
 b15zdnd00an1n01x5 FILLER_184_1303 ();
 b15zdnd11an1n64x5 FILLER_184_1331 ();
 b15zdnd11an1n64x5 FILLER_184_1395 ();
 b15zdnd11an1n64x5 FILLER_184_1459 ();
 b15zdnd11an1n08x5 FILLER_184_1523 ();
 b15zdnd00an1n01x5 FILLER_184_1531 ();
 b15zdnd11an1n08x5 FILLER_184_1539 ();
 b15zdnd11an1n04x5 FILLER_184_1547 ();
 b15zdnd00an1n01x5 FILLER_184_1551 ();
 b15zdnd11an1n64x5 FILLER_184_1564 ();
 b15zdnd11an1n16x5 FILLER_184_1628 ();
 b15zdnd11an1n08x5 FILLER_184_1644 ();
 b15zdnd11an1n64x5 FILLER_184_1669 ();
 b15zdnd11an1n64x5 FILLER_184_1733 ();
 b15zdnd11an1n16x5 FILLER_184_1797 ();
 b15zdnd11an1n08x5 FILLER_184_1813 ();
 b15zdnd00an1n02x5 FILLER_184_1821 ();
 b15zdnd00an1n01x5 FILLER_184_1823 ();
 b15zdnd11an1n08x5 FILLER_184_1848 ();
 b15zdnd00an1n01x5 FILLER_184_1856 ();
 b15zdnd11an1n64x5 FILLER_184_1901 ();
 b15zdnd11an1n64x5 FILLER_184_1965 ();
 b15zdnd11an1n64x5 FILLER_184_2029 ();
 b15zdnd11an1n32x5 FILLER_184_2093 ();
 b15zdnd11an1n16x5 FILLER_184_2125 ();
 b15zdnd11an1n08x5 FILLER_184_2141 ();
 b15zdnd11an1n04x5 FILLER_184_2149 ();
 b15zdnd00an1n01x5 FILLER_184_2153 ();
 b15zdnd11an1n64x5 FILLER_184_2162 ();
 b15zdnd11an1n32x5 FILLER_184_2226 ();
 b15zdnd11an1n16x5 FILLER_184_2258 ();
 b15zdnd00an1n02x5 FILLER_184_2274 ();
 b15zdnd11an1n32x5 FILLER_185_0 ();
 b15zdnd11an1n16x5 FILLER_185_32 ();
 b15zdnd11an1n08x5 FILLER_185_48 ();
 b15zdnd00an1n02x5 FILLER_185_56 ();
 b15zdnd00an1n01x5 FILLER_185_58 ();
 b15zdnd11an1n04x5 FILLER_185_79 ();
 b15zdnd11an1n08x5 FILLER_185_89 ();
 b15zdnd00an1n02x5 FILLER_185_97 ();
 b15zdnd11an1n04x5 FILLER_185_141 ();
 b15zdnd11an1n64x5 FILLER_185_148 ();
 b15zdnd11an1n64x5 FILLER_185_212 ();
 b15zdnd11an1n64x5 FILLER_185_276 ();
 b15zdnd11an1n64x5 FILLER_185_340 ();
 b15zdnd11an1n08x5 FILLER_185_404 ();
 b15zdnd00an1n02x5 FILLER_185_412 ();
 b15zdnd11an1n16x5 FILLER_185_421 ();
 b15zdnd11an1n04x5 FILLER_185_437 ();
 b15zdnd00an1n01x5 FILLER_185_441 ();
 b15zdnd11an1n04x5 FILLER_185_456 ();
 b15zdnd11an1n08x5 FILLER_185_465 ();
 b15zdnd00an1n02x5 FILLER_185_473 ();
 b15zdnd11an1n04x5 FILLER_185_481 ();
 b15zdnd11an1n64x5 FILLER_185_527 ();
 b15zdnd11an1n64x5 FILLER_185_591 ();
 b15zdnd11an1n64x5 FILLER_185_655 ();
 b15zdnd11an1n64x5 FILLER_185_719 ();
 b15zdnd11an1n64x5 FILLER_185_783 ();
 b15zdnd11an1n64x5 FILLER_185_847 ();
 b15zdnd11an1n64x5 FILLER_185_911 ();
 b15zdnd11an1n32x5 FILLER_185_975 ();
 b15zdnd11an1n16x5 FILLER_185_1007 ();
 b15zdnd11an1n08x5 FILLER_185_1023 ();
 b15zdnd11an1n32x5 FILLER_185_1083 ();
 b15zdnd11an1n16x5 FILLER_185_1115 ();
 b15zdnd00an1n01x5 FILLER_185_1131 ();
 b15zdnd11an1n16x5 FILLER_185_1139 ();
 b15zdnd00an1n01x5 FILLER_185_1155 ();
 b15zdnd11an1n32x5 FILLER_185_1208 ();
 b15zdnd11an1n08x5 FILLER_185_1240 ();
 b15zdnd00an1n01x5 FILLER_185_1248 ();
 b15zdnd11an1n04x5 FILLER_185_1253 ();
 b15zdnd11an1n04x5 FILLER_185_1299 ();
 b15zdnd11an1n16x5 FILLER_185_1314 ();
 b15zdnd11an1n08x5 FILLER_185_1330 ();
 b15zdnd11an1n04x5 FILLER_185_1338 ();
 b15zdnd00an1n02x5 FILLER_185_1342 ();
 b15zdnd00an1n01x5 FILLER_185_1344 ();
 b15zdnd11an1n64x5 FILLER_185_1358 ();
 b15zdnd11an1n64x5 FILLER_185_1422 ();
 b15zdnd11an1n32x5 FILLER_185_1486 ();
 b15zdnd11an1n08x5 FILLER_185_1518 ();
 b15zdnd11an1n04x5 FILLER_185_1526 ();
 b15zdnd11an1n64x5 FILLER_185_1575 ();
 b15zdnd11an1n64x5 FILLER_185_1639 ();
 b15zdnd11an1n64x5 FILLER_185_1703 ();
 b15zdnd11an1n64x5 FILLER_185_1767 ();
 b15zdnd11an1n32x5 FILLER_185_1831 ();
 b15zdnd11an1n16x5 FILLER_185_1863 ();
 b15zdnd00an1n01x5 FILLER_185_1879 ();
 b15zdnd11an1n64x5 FILLER_185_1883 ();
 b15zdnd11an1n64x5 FILLER_185_1947 ();
 b15zdnd11an1n64x5 FILLER_185_2011 ();
 b15zdnd11an1n16x5 FILLER_185_2075 ();
 b15zdnd11an1n64x5 FILLER_185_2133 ();
 b15zdnd11an1n64x5 FILLER_185_2197 ();
 b15zdnd11an1n16x5 FILLER_185_2261 ();
 b15zdnd11an1n04x5 FILLER_185_2277 ();
 b15zdnd00an1n02x5 FILLER_185_2281 ();
 b15zdnd00an1n01x5 FILLER_185_2283 ();
 b15zdnd11an1n64x5 FILLER_186_8 ();
 b15zdnd00an1n02x5 FILLER_186_72 ();
 b15zdnd00an1n01x5 FILLER_186_74 ();
 b15zdnd11an1n16x5 FILLER_186_95 ();
 b15zdnd11an1n08x5 FILLER_186_111 ();
 b15zdnd11an1n04x5 FILLER_186_119 ();
 b15zdnd00an1n01x5 FILLER_186_123 ();
 b15zdnd11an1n04x5 FILLER_186_127 ();
 b15zdnd11an1n64x5 FILLER_186_134 ();
 b15zdnd11an1n64x5 FILLER_186_198 ();
 b15zdnd11an1n64x5 FILLER_186_262 ();
 b15zdnd11an1n64x5 FILLER_186_326 ();
 b15zdnd11an1n64x5 FILLER_186_390 ();
 b15zdnd11an1n16x5 FILLER_186_454 ();
 b15zdnd11an1n04x5 FILLER_186_470 ();
 b15zdnd00an1n01x5 FILLER_186_474 ();
 b15zdnd11an1n04x5 FILLER_186_478 ();
 b15zdnd11an1n04x5 FILLER_186_487 ();
 b15zdnd11an1n04x5 FILLER_186_533 ();
 b15zdnd11an1n64x5 FILLER_186_545 ();
 b15zdnd11an1n64x5 FILLER_186_609 ();
 b15zdnd11an1n32x5 FILLER_186_673 ();
 b15zdnd11an1n08x5 FILLER_186_705 ();
 b15zdnd11an1n04x5 FILLER_186_713 ();
 b15zdnd00an1n01x5 FILLER_186_717 ();
 b15zdnd11an1n64x5 FILLER_186_726 ();
 b15zdnd11an1n64x5 FILLER_186_790 ();
 b15zdnd11an1n16x5 FILLER_186_854 ();
 b15zdnd11an1n08x5 FILLER_186_870 ();
 b15zdnd11an1n04x5 FILLER_186_878 ();
 b15zdnd00an1n02x5 FILLER_186_882 ();
 b15zdnd00an1n01x5 FILLER_186_884 ();
 b15zdnd11an1n64x5 FILLER_186_893 ();
 b15zdnd11an1n64x5 FILLER_186_957 ();
 b15zdnd11an1n08x5 FILLER_186_1021 ();
 b15zdnd00an1n02x5 FILLER_186_1029 ();
 b15zdnd00an1n01x5 FILLER_186_1031 ();
 b15zdnd11an1n64x5 FILLER_186_1084 ();
 b15zdnd11an1n16x5 FILLER_186_1148 ();
 b15zdnd11an1n08x5 FILLER_186_1164 ();
 b15zdnd11an1n04x5 FILLER_186_1172 ();
 b15zdnd11an1n04x5 FILLER_186_1179 ();
 b15zdnd11an1n04x5 FILLER_186_1186 ();
 b15zdnd11an1n04x5 FILLER_186_1193 ();
 b15zdnd11an1n64x5 FILLER_186_1204 ();
 b15zdnd11an1n32x5 FILLER_186_1268 ();
 b15zdnd11an1n16x5 FILLER_186_1300 ();
 b15zdnd11an1n04x5 FILLER_186_1316 ();
 b15zdnd00an1n01x5 FILLER_186_1320 ();
 b15zdnd11an1n16x5 FILLER_186_1327 ();
 b15zdnd11an1n04x5 FILLER_186_1343 ();
 b15zdnd00an1n02x5 FILLER_186_1347 ();
 b15zdnd00an1n01x5 FILLER_186_1349 ();
 b15zdnd11an1n64x5 FILLER_186_1363 ();
 b15zdnd11an1n64x5 FILLER_186_1427 ();
 b15zdnd11an1n64x5 FILLER_186_1491 ();
 b15zdnd11an1n64x5 FILLER_186_1555 ();
 b15zdnd11an1n64x5 FILLER_186_1619 ();
 b15zdnd11an1n64x5 FILLER_186_1683 ();
 b15zdnd11an1n16x5 FILLER_186_1747 ();
 b15zdnd11an1n64x5 FILLER_186_1767 ();
 b15zdnd11an1n64x5 FILLER_186_1831 ();
 b15zdnd11an1n64x5 FILLER_186_1895 ();
 b15zdnd11an1n64x5 FILLER_186_1959 ();
 b15zdnd11an1n32x5 FILLER_186_2023 ();
 b15zdnd11an1n04x5 FILLER_186_2055 ();
 b15zdnd00an1n02x5 FILLER_186_2059 ();
 b15zdnd11an1n64x5 FILLER_186_2085 ();
 b15zdnd11an1n04x5 FILLER_186_2149 ();
 b15zdnd00an1n01x5 FILLER_186_2153 ();
 b15zdnd11an1n64x5 FILLER_186_2162 ();
 b15zdnd11an1n16x5 FILLER_186_2226 ();
 b15zdnd11an1n08x5 FILLER_186_2242 ();
 b15zdnd11an1n04x5 FILLER_186_2250 ();
 b15zdnd00an1n01x5 FILLER_186_2254 ();
 b15zdnd11an1n08x5 FILLER_186_2261 ();
 b15zdnd11an1n04x5 FILLER_186_2269 ();
 b15zdnd00an1n02x5 FILLER_186_2273 ();
 b15zdnd00an1n01x5 FILLER_186_2275 ();
 b15zdnd11an1n64x5 FILLER_187_0 ();
 b15zdnd11an1n08x5 FILLER_187_64 ();
 b15zdnd00an1n02x5 FILLER_187_72 ();
 b15zdnd11an1n08x5 FILLER_187_119 ();
 b15zdnd00an1n01x5 FILLER_187_127 ();
 b15zdnd11an1n64x5 FILLER_187_161 ();
 b15zdnd11an1n64x5 FILLER_187_225 ();
 b15zdnd11an1n64x5 FILLER_187_289 ();
 b15zdnd11an1n64x5 FILLER_187_353 ();
 b15zdnd11an1n32x5 FILLER_187_417 ();
 b15zdnd11an1n16x5 FILLER_187_449 ();
 b15zdnd00an1n01x5 FILLER_187_465 ();
 b15zdnd11an1n64x5 FILLER_187_518 ();
 b15zdnd11an1n64x5 FILLER_187_582 ();
 b15zdnd11an1n64x5 FILLER_187_646 ();
 b15zdnd11an1n64x5 FILLER_187_710 ();
 b15zdnd11an1n64x5 FILLER_187_774 ();
 b15zdnd11an1n32x5 FILLER_187_847 ();
 b15zdnd11an1n08x5 FILLER_187_879 ();
 b15zdnd11an1n04x5 FILLER_187_887 ();
 b15zdnd00an1n02x5 FILLER_187_891 ();
 b15zdnd11an1n64x5 FILLER_187_896 ();
 b15zdnd11an1n64x5 FILLER_187_960 ();
 b15zdnd11an1n16x5 FILLER_187_1024 ();
 b15zdnd11an1n08x5 FILLER_187_1040 ();
 b15zdnd11an1n04x5 FILLER_187_1048 ();
 b15zdnd11an1n04x5 FILLER_187_1055 ();
 b15zdnd11an1n04x5 FILLER_187_1062 ();
 b15zdnd11an1n32x5 FILLER_187_1069 ();
 b15zdnd11an1n16x5 FILLER_187_1101 ();
 b15zdnd11an1n08x5 FILLER_187_1117 ();
 b15zdnd00an1n02x5 FILLER_187_1125 ();
 b15zdnd11an1n16x5 FILLER_187_1136 ();
 b15zdnd11an1n04x5 FILLER_187_1152 ();
 b15zdnd00an1n02x5 FILLER_187_1156 ();
 b15zdnd11an1n64x5 FILLER_187_1210 ();
 b15zdnd11an1n32x5 FILLER_187_1274 ();
 b15zdnd11an1n08x5 FILLER_187_1306 ();
 b15zdnd11an1n04x5 FILLER_187_1314 ();
 b15zdnd00an1n01x5 FILLER_187_1318 ();
 b15zdnd11an1n08x5 FILLER_187_1342 ();
 b15zdnd00an1n02x5 FILLER_187_1350 ();
 b15zdnd00an1n01x5 FILLER_187_1352 ();
 b15zdnd11an1n64x5 FILLER_187_1356 ();
 b15zdnd11an1n64x5 FILLER_187_1420 ();
 b15zdnd11an1n64x5 FILLER_187_1484 ();
 b15zdnd11an1n64x5 FILLER_187_1548 ();
 b15zdnd11an1n32x5 FILLER_187_1612 ();
 b15zdnd11an1n16x5 FILLER_187_1644 ();
 b15zdnd11an1n08x5 FILLER_187_1660 ();
 b15zdnd11an1n04x5 FILLER_187_1668 ();
 b15zdnd00an1n01x5 FILLER_187_1672 ();
 b15zdnd11an1n32x5 FILLER_187_1677 ();
 b15zdnd11an1n16x5 FILLER_187_1709 ();
 b15zdnd11an1n08x5 FILLER_187_1725 ();
 b15zdnd00an1n01x5 FILLER_187_1733 ();
 b15zdnd11an1n16x5 FILLER_187_1748 ();
 b15zdnd11an1n08x5 FILLER_187_1764 ();
 b15zdnd00an1n02x5 FILLER_187_1772 ();
 b15zdnd00an1n01x5 FILLER_187_1774 ();
 b15zdnd11an1n32x5 FILLER_187_1778 ();
 b15zdnd11an1n16x5 FILLER_187_1810 ();
 b15zdnd11an1n08x5 FILLER_187_1826 ();
 b15zdnd00an1n02x5 FILLER_187_1834 ();
 b15zdnd00an1n01x5 FILLER_187_1836 ();
 b15zdnd11an1n64x5 FILLER_187_1879 ();
 b15zdnd11an1n64x5 FILLER_187_1943 ();
 b15zdnd11an1n32x5 FILLER_187_2007 ();
 b15zdnd00an1n01x5 FILLER_187_2039 ();
 b15zdnd11an1n32x5 FILLER_187_2054 ();
 b15zdnd11an1n08x5 FILLER_187_2086 ();
 b15zdnd11an1n04x5 FILLER_187_2094 ();
 b15zdnd00an1n02x5 FILLER_187_2098 ();
 b15zdnd00an1n01x5 FILLER_187_2100 ();
 b15zdnd11an1n32x5 FILLER_187_2121 ();
 b15zdnd11an1n16x5 FILLER_187_2153 ();
 b15zdnd00an1n02x5 FILLER_187_2169 ();
 b15zdnd00an1n01x5 FILLER_187_2171 ();
 b15zdnd11an1n32x5 FILLER_187_2190 ();
 b15zdnd11an1n16x5 FILLER_187_2222 ();
 b15zdnd11an1n08x5 FILLER_187_2238 ();
 b15zdnd11an1n04x5 FILLER_187_2246 ();
 b15zdnd11an1n16x5 FILLER_187_2264 ();
 b15zdnd11an1n04x5 FILLER_187_2280 ();
 b15zdnd11an1n32x5 FILLER_188_8 ();
 b15zdnd11an1n16x5 FILLER_188_40 ();
 b15zdnd11an1n08x5 FILLER_188_56 ();
 b15zdnd00an1n02x5 FILLER_188_64 ();
 b15zdnd00an1n01x5 FILLER_188_66 ();
 b15zdnd11an1n04x5 FILLER_188_109 ();
 b15zdnd11an1n64x5 FILLER_188_120 ();
 b15zdnd11an1n64x5 FILLER_188_184 ();
 b15zdnd00an1n02x5 FILLER_188_248 ();
 b15zdnd11an1n64x5 FILLER_188_253 ();
 b15zdnd11an1n64x5 FILLER_188_317 ();
 b15zdnd11an1n32x5 FILLER_188_381 ();
 b15zdnd11an1n16x5 FILLER_188_413 ();
 b15zdnd11an1n04x5 FILLER_188_429 ();
 b15zdnd11an1n16x5 FILLER_188_437 ();
 b15zdnd11an1n08x5 FILLER_188_453 ();
 b15zdnd11an1n04x5 FILLER_188_461 ();
 b15zdnd00an1n01x5 FILLER_188_465 ();
 b15zdnd11an1n64x5 FILLER_188_508 ();
 b15zdnd11an1n64x5 FILLER_188_572 ();
 b15zdnd11an1n64x5 FILLER_188_636 ();
 b15zdnd11an1n16x5 FILLER_188_700 ();
 b15zdnd00an1n02x5 FILLER_188_716 ();
 b15zdnd11an1n64x5 FILLER_188_726 ();
 b15zdnd11an1n64x5 FILLER_188_790 ();
 b15zdnd11an1n08x5 FILLER_188_854 ();
 b15zdnd11an1n04x5 FILLER_188_862 ();
 b15zdnd11an1n64x5 FILLER_188_918 ();
 b15zdnd11an1n64x5 FILLER_188_982 ();
 b15zdnd11an1n08x5 FILLER_188_1046 ();
 b15zdnd00an1n02x5 FILLER_188_1054 ();
 b15zdnd00an1n01x5 FILLER_188_1056 ();
 b15zdnd11an1n64x5 FILLER_188_1060 ();
 b15zdnd11an1n32x5 FILLER_188_1124 ();
 b15zdnd11an1n16x5 FILLER_188_1156 ();
 b15zdnd11an1n08x5 FILLER_188_1172 ();
 b15zdnd00an1n02x5 FILLER_188_1180 ();
 b15zdnd00an1n01x5 FILLER_188_1182 ();
 b15zdnd11an1n64x5 FILLER_188_1186 ();
 b15zdnd11an1n32x5 FILLER_188_1250 ();
 b15zdnd11an1n16x5 FILLER_188_1282 ();
 b15zdnd11an1n08x5 FILLER_188_1298 ();
 b15zdnd00an1n02x5 FILLER_188_1306 ();
 b15zdnd00an1n01x5 FILLER_188_1308 ();
 b15zdnd11an1n08x5 FILLER_188_1325 ();
 b15zdnd11an1n04x5 FILLER_188_1333 ();
 b15zdnd00an1n01x5 FILLER_188_1337 ();
 b15zdnd11an1n64x5 FILLER_188_1345 ();
 b15zdnd11an1n32x5 FILLER_188_1409 ();
 b15zdnd11an1n04x5 FILLER_188_1441 ();
 b15zdnd00an1n02x5 FILLER_188_1445 ();
 b15zdnd00an1n01x5 FILLER_188_1447 ();
 b15zdnd11an1n64x5 FILLER_188_1465 ();
 b15zdnd11an1n32x5 FILLER_188_1529 ();
 b15zdnd11an1n16x5 FILLER_188_1561 ();
 b15zdnd00an1n01x5 FILLER_188_1577 ();
 b15zdnd11an1n64x5 FILLER_188_1594 ();
 b15zdnd11an1n04x5 FILLER_188_1658 ();
 b15zdnd00an1n01x5 FILLER_188_1662 ();
 b15zdnd11an1n16x5 FILLER_188_1671 ();
 b15zdnd11an1n04x5 FILLER_188_1687 ();
 b15zdnd00an1n02x5 FILLER_188_1691 ();
 b15zdnd11an1n08x5 FILLER_188_1700 ();
 b15zdnd00an1n02x5 FILLER_188_1708 ();
 b15zdnd00an1n01x5 FILLER_188_1710 ();
 b15zdnd11an1n64x5 FILLER_188_1725 ();
 b15zdnd11an1n16x5 FILLER_188_1789 ();
 b15zdnd11an1n08x5 FILLER_188_1805 ();
 b15zdnd00an1n01x5 FILLER_188_1813 ();
 b15zdnd11an1n64x5 FILLER_188_1828 ();
 b15zdnd11an1n64x5 FILLER_188_1892 ();
 b15zdnd11an1n64x5 FILLER_188_1956 ();
 b15zdnd11an1n64x5 FILLER_188_2020 ();
 b15zdnd11an1n64x5 FILLER_188_2084 ();
 b15zdnd11an1n04x5 FILLER_188_2148 ();
 b15zdnd00an1n02x5 FILLER_188_2152 ();
 b15zdnd11an1n64x5 FILLER_188_2162 ();
 b15zdnd11an1n32x5 FILLER_188_2226 ();
 b15zdnd11an1n16x5 FILLER_188_2258 ();
 b15zdnd00an1n02x5 FILLER_188_2274 ();
 b15zdnd00an1n02x5 FILLER_189_0 ();
 b15zdnd11an1n16x5 FILLER_189_6 ();
 b15zdnd11an1n08x5 FILLER_189_22 ();
 b15zdnd00an1n01x5 FILLER_189_30 ();
 b15zdnd11an1n16x5 FILLER_189_35 ();
 b15zdnd11an1n08x5 FILLER_189_51 ();
 b15zdnd11an1n04x5 FILLER_189_59 ();
 b15zdnd00an1n02x5 FILLER_189_63 ();
 b15zdnd00an1n01x5 FILLER_189_65 ();
 b15zdnd11an1n64x5 FILLER_189_108 ();
 b15zdnd11an1n32x5 FILLER_189_172 ();
 b15zdnd11an1n08x5 FILLER_189_204 ();
 b15zdnd00an1n02x5 FILLER_189_212 ();
 b15zdnd11an1n04x5 FILLER_189_254 ();
 b15zdnd11an1n64x5 FILLER_189_261 ();
 b15zdnd11an1n64x5 FILLER_189_325 ();
 b15zdnd11an1n64x5 FILLER_189_389 ();
 b15zdnd11an1n32x5 FILLER_189_453 ();
 b15zdnd00an1n01x5 FILLER_189_485 ();
 b15zdnd11an1n04x5 FILLER_189_489 ();
 b15zdnd11an1n64x5 FILLER_189_496 ();
 b15zdnd11an1n64x5 FILLER_189_560 ();
 b15zdnd11an1n64x5 FILLER_189_624 ();
 b15zdnd11an1n64x5 FILLER_189_688 ();
 b15zdnd11an1n64x5 FILLER_189_752 ();
 b15zdnd11an1n64x5 FILLER_189_816 ();
 b15zdnd11an1n04x5 FILLER_189_880 ();
 b15zdnd00an1n01x5 FILLER_189_884 ();
 b15zdnd11an1n04x5 FILLER_189_888 ();
 b15zdnd11an1n64x5 FILLER_189_895 ();
 b15zdnd11an1n64x5 FILLER_189_959 ();
 b15zdnd11an1n32x5 FILLER_189_1023 ();
 b15zdnd11an1n16x5 FILLER_189_1055 ();
 b15zdnd11an1n08x5 FILLER_189_1071 ();
 b15zdnd11an1n04x5 FILLER_189_1082 ();
 b15zdnd11an1n64x5 FILLER_189_1113 ();
 b15zdnd11an1n08x5 FILLER_189_1177 ();
 b15zdnd00an1n01x5 FILLER_189_1185 ();
 b15zdnd11an1n64x5 FILLER_189_1189 ();
 b15zdnd11an1n64x5 FILLER_189_1253 ();
 b15zdnd11an1n64x5 FILLER_189_1317 ();
 b15zdnd11an1n64x5 FILLER_189_1381 ();
 b15zdnd11an1n64x5 FILLER_189_1487 ();
 b15zdnd11an1n64x5 FILLER_189_1551 ();
 b15zdnd11an1n64x5 FILLER_189_1615 ();
 b15zdnd11an1n64x5 FILLER_189_1679 ();
 b15zdnd11an1n64x5 FILLER_189_1743 ();
 b15zdnd11an1n16x5 FILLER_189_1807 ();
 b15zdnd11an1n08x5 FILLER_189_1823 ();
 b15zdnd00an1n02x5 FILLER_189_1831 ();
 b15zdnd00an1n01x5 FILLER_189_1833 ();
 b15zdnd11an1n64x5 FILLER_189_1837 ();
 b15zdnd11an1n64x5 FILLER_189_1901 ();
 b15zdnd11an1n32x5 FILLER_189_1965 ();
 b15zdnd00an1n02x5 FILLER_189_1997 ();
 b15zdnd11an1n64x5 FILLER_189_2023 ();
 b15zdnd11an1n64x5 FILLER_189_2087 ();
 b15zdnd11an1n32x5 FILLER_189_2151 ();
 b15zdnd11an1n16x5 FILLER_189_2183 ();
 b15zdnd11an1n04x5 FILLER_189_2199 ();
 b15zdnd11an1n32x5 FILLER_189_2221 ();
 b15zdnd11an1n16x5 FILLER_189_2253 ();
 b15zdnd11an1n08x5 FILLER_189_2269 ();
 b15zdnd11an1n04x5 FILLER_189_2277 ();
 b15zdnd00an1n02x5 FILLER_189_2281 ();
 b15zdnd00an1n01x5 FILLER_189_2283 ();
 b15zdnd11an1n04x5 FILLER_190_8 ();
 b15zdnd00an1n02x5 FILLER_190_12 ();
 b15zdnd11an1n04x5 FILLER_190_18 ();
 b15zdnd11an1n04x5 FILLER_190_26 ();
 b15zdnd11an1n64x5 FILLER_190_34 ();
 b15zdnd11an1n08x5 FILLER_190_98 ();
 b15zdnd11an1n64x5 FILLER_190_148 ();
 b15zdnd11an1n16x5 FILLER_190_212 ();
 b15zdnd11an1n04x5 FILLER_190_228 ();
 b15zdnd11an1n04x5 FILLER_190_235 ();
 b15zdnd11an1n64x5 FILLER_190_257 ();
 b15zdnd11an1n64x5 FILLER_190_321 ();
 b15zdnd11an1n64x5 FILLER_190_385 ();
 b15zdnd11an1n64x5 FILLER_190_449 ();
 b15zdnd11an1n64x5 FILLER_190_513 ();
 b15zdnd11an1n16x5 FILLER_190_577 ();
 b15zdnd11an1n08x5 FILLER_190_593 ();
 b15zdnd00an1n02x5 FILLER_190_601 ();
 b15zdnd11an1n64x5 FILLER_190_611 ();
 b15zdnd11an1n32x5 FILLER_190_675 ();
 b15zdnd11an1n08x5 FILLER_190_707 ();
 b15zdnd00an1n02x5 FILLER_190_715 ();
 b15zdnd00an1n01x5 FILLER_190_717 ();
 b15zdnd11an1n64x5 FILLER_190_726 ();
 b15zdnd11an1n64x5 FILLER_190_790 ();
 b15zdnd11an1n64x5 FILLER_190_854 ();
 b15zdnd11an1n64x5 FILLER_190_918 ();
 b15zdnd11an1n64x5 FILLER_190_982 ();
 b15zdnd11an1n64x5 FILLER_190_1046 ();
 b15zdnd11an1n64x5 FILLER_190_1110 ();
 b15zdnd11an1n08x5 FILLER_190_1174 ();
 b15zdnd11an1n04x5 FILLER_190_1182 ();
 b15zdnd11an1n64x5 FILLER_190_1189 ();
 b15zdnd11an1n64x5 FILLER_190_1253 ();
 b15zdnd11an1n16x5 FILLER_190_1317 ();
 b15zdnd11an1n08x5 FILLER_190_1333 ();
 b15zdnd11an1n04x5 FILLER_190_1341 ();
 b15zdnd00an1n02x5 FILLER_190_1345 ();
 b15zdnd00an1n01x5 FILLER_190_1347 ();
 b15zdnd11an1n64x5 FILLER_190_1351 ();
 b15zdnd11an1n32x5 FILLER_190_1415 ();
 b15zdnd11an1n16x5 FILLER_190_1447 ();
 b15zdnd11an1n04x5 FILLER_190_1463 ();
 b15zdnd00an1n02x5 FILLER_190_1467 ();
 b15zdnd11an1n32x5 FILLER_190_1489 ();
 b15zdnd11an1n08x5 FILLER_190_1521 ();
 b15zdnd11an1n04x5 FILLER_190_1529 ();
 b15zdnd00an1n02x5 FILLER_190_1533 ();
 b15zdnd11an1n32x5 FILLER_190_1549 ();
 b15zdnd00an1n01x5 FILLER_190_1581 ();
 b15zdnd11an1n32x5 FILLER_190_1594 ();
 b15zdnd11an1n16x5 FILLER_190_1626 ();
 b15zdnd11an1n04x5 FILLER_190_1642 ();
 b15zdnd00an1n01x5 FILLER_190_1646 ();
 b15zdnd11an1n64x5 FILLER_190_1651 ();
 b15zdnd11an1n04x5 FILLER_190_1715 ();
 b15zdnd00an1n02x5 FILLER_190_1719 ();
 b15zdnd11an1n64x5 FILLER_190_1738 ();
 b15zdnd11an1n64x5 FILLER_190_1802 ();
 b15zdnd11an1n64x5 FILLER_190_1866 ();
 b15zdnd11an1n64x5 FILLER_190_1930 ();
 b15zdnd11an1n64x5 FILLER_190_1994 ();
 b15zdnd11an1n08x5 FILLER_190_2058 ();
 b15zdnd11an1n04x5 FILLER_190_2066 ();
 b15zdnd00an1n02x5 FILLER_190_2070 ();
 b15zdnd11an1n64x5 FILLER_190_2089 ();
 b15zdnd00an1n01x5 FILLER_190_2153 ();
 b15zdnd11an1n32x5 FILLER_190_2162 ();
 b15zdnd11an1n16x5 FILLER_190_2194 ();
 b15zdnd00an1n02x5 FILLER_190_2210 ();
 b15zdnd00an1n01x5 FILLER_190_2212 ();
 b15zdnd11an1n04x5 FILLER_190_2228 ();
 b15zdnd11an1n16x5 FILLER_190_2254 ();
 b15zdnd11an1n04x5 FILLER_190_2270 ();
 b15zdnd00an1n02x5 FILLER_190_2274 ();
 b15zdnd11an1n04x5 FILLER_191_0 ();
 b15zdnd00an1n02x5 FILLER_191_4 ();
 b15zdnd00an1n01x5 FILLER_191_6 ();
 b15zdnd11an1n16x5 FILLER_191_49 ();
 b15zdnd11an1n04x5 FILLER_191_65 ();
 b15zdnd00an1n02x5 FILLER_191_69 ();
 b15zdnd11an1n16x5 FILLER_191_113 ();
 b15zdnd11an1n08x5 FILLER_191_129 ();
 b15zdnd00an1n02x5 FILLER_191_137 ();
 b15zdnd00an1n01x5 FILLER_191_139 ();
 b15zdnd11an1n16x5 FILLER_191_182 ();
 b15zdnd11an1n04x5 FILLER_191_198 ();
 b15zdnd00an1n02x5 FILLER_191_202 ();
 b15zdnd00an1n01x5 FILLER_191_204 ();
 b15zdnd11an1n64x5 FILLER_191_257 ();
 b15zdnd11an1n64x5 FILLER_191_321 ();
 b15zdnd11an1n64x5 FILLER_191_385 ();
 b15zdnd11an1n64x5 FILLER_191_449 ();
 b15zdnd11an1n64x5 FILLER_191_513 ();
 b15zdnd11an1n32x5 FILLER_191_577 ();
 b15zdnd11an1n08x5 FILLER_191_609 ();
 b15zdnd00an1n02x5 FILLER_191_617 ();
 b15zdnd11an1n64x5 FILLER_191_622 ();
 b15zdnd11an1n64x5 FILLER_191_686 ();
 b15zdnd11an1n16x5 FILLER_191_750 ();
 b15zdnd11an1n08x5 FILLER_191_766 ();
 b15zdnd11an1n04x5 FILLER_191_774 ();
 b15zdnd00an1n02x5 FILLER_191_778 ();
 b15zdnd00an1n01x5 FILLER_191_780 ();
 b15zdnd11an1n08x5 FILLER_191_784 ();
 b15zdnd11an1n64x5 FILLER_191_819 ();
 b15zdnd11an1n64x5 FILLER_191_883 ();
 b15zdnd11an1n64x5 FILLER_191_947 ();
 b15zdnd11an1n64x5 FILLER_191_1011 ();
 b15zdnd11an1n64x5 FILLER_191_1075 ();
 b15zdnd11an1n16x5 FILLER_191_1139 ();
 b15zdnd11an1n04x5 FILLER_191_1155 ();
 b15zdnd00an1n02x5 FILLER_191_1159 ();
 b15zdnd11an1n64x5 FILLER_191_1213 ();
 b15zdnd11an1n64x5 FILLER_191_1277 ();
 b15zdnd11an1n64x5 FILLER_191_1341 ();
 b15zdnd11an1n16x5 FILLER_191_1405 ();
 b15zdnd11an1n08x5 FILLER_191_1421 ();
 b15zdnd11an1n04x5 FILLER_191_1429 ();
 b15zdnd11an1n64x5 FILLER_191_1447 ();
 b15zdnd11an1n64x5 FILLER_191_1511 ();
 b15zdnd11an1n64x5 FILLER_191_1575 ();
 b15zdnd11an1n16x5 FILLER_191_1639 ();
 b15zdnd00an1n02x5 FILLER_191_1655 ();
 b15zdnd11an1n16x5 FILLER_191_1665 ();
 b15zdnd11an1n04x5 FILLER_191_1681 ();
 b15zdnd00an1n02x5 FILLER_191_1685 ();
 b15zdnd00an1n01x5 FILLER_191_1687 ();
 b15zdnd11an1n16x5 FILLER_191_1713 ();
 b15zdnd00an1n02x5 FILLER_191_1729 ();
 b15zdnd11an1n32x5 FILLER_191_1751 ();
 b15zdnd11an1n16x5 FILLER_191_1783 ();
 b15zdnd11an1n04x5 FILLER_191_1799 ();
 b15zdnd00an1n01x5 FILLER_191_1803 ();
 b15zdnd11an1n32x5 FILLER_191_1829 ();
 b15zdnd11an1n16x5 FILLER_191_1861 ();
 b15zdnd11an1n04x5 FILLER_191_1877 ();
 b15zdnd00an1n01x5 FILLER_191_1881 ();
 b15zdnd11an1n32x5 FILLER_191_1885 ();
 b15zdnd11an1n08x5 FILLER_191_1917 ();
 b15zdnd11an1n04x5 FILLER_191_1925 ();
 b15zdnd00an1n02x5 FILLER_191_1929 ();
 b15zdnd11an1n08x5 FILLER_191_1934 ();
 b15zdnd00an1n02x5 FILLER_191_1942 ();
 b15zdnd00an1n01x5 FILLER_191_1944 ();
 b15zdnd11an1n64x5 FILLER_191_1948 ();
 b15zdnd11an1n16x5 FILLER_191_2012 ();
 b15zdnd11an1n08x5 FILLER_191_2028 ();
 b15zdnd11an1n04x5 FILLER_191_2036 ();
 b15zdnd00an1n02x5 FILLER_191_2040 ();
 b15zdnd00an1n01x5 FILLER_191_2042 ();
 b15zdnd11an1n04x5 FILLER_191_2050 ();
 b15zdnd11an1n64x5 FILLER_191_2068 ();
 b15zdnd11an1n32x5 FILLER_191_2132 ();
 b15zdnd00an1n02x5 FILLER_191_2164 ();
 b15zdnd00an1n01x5 FILLER_191_2166 ();
 b15zdnd11an1n64x5 FILLER_191_2182 ();
 b15zdnd11an1n08x5 FILLER_191_2246 ();
 b15zdnd11an1n04x5 FILLER_191_2254 ();
 b15zdnd00an1n02x5 FILLER_191_2258 ();
 b15zdnd00an1n01x5 FILLER_191_2260 ();
 b15zdnd11an1n16x5 FILLER_191_2267 ();
 b15zdnd00an1n01x5 FILLER_191_2283 ();
 b15zdnd00an1n02x5 FILLER_192_8 ();
 b15zdnd11an1n32x5 FILLER_192_52 ();
 b15zdnd11an1n08x5 FILLER_192_84 ();
 b15zdnd11an1n04x5 FILLER_192_92 ();
 b15zdnd00an1n02x5 FILLER_192_96 ();
 b15zdnd11an1n08x5 FILLER_192_140 ();
 b15zdnd11an1n04x5 FILLER_192_148 ();
 b15zdnd11an1n04x5 FILLER_192_194 ();
 b15zdnd11an1n64x5 FILLER_192_240 ();
 b15zdnd11an1n64x5 FILLER_192_304 ();
 b15zdnd11an1n64x5 FILLER_192_368 ();
 b15zdnd11an1n64x5 FILLER_192_432 ();
 b15zdnd11an1n64x5 FILLER_192_496 ();
 b15zdnd11an1n32x5 FILLER_192_560 ();
 b15zdnd11an1n16x5 FILLER_192_592 ();
 b15zdnd00an1n02x5 FILLER_192_608 ();
 b15zdnd00an1n01x5 FILLER_192_610 ();
 b15zdnd11an1n04x5 FILLER_192_620 ();
 b15zdnd00an1n02x5 FILLER_192_624 ();
 b15zdnd11an1n08x5 FILLER_192_629 ();
 b15zdnd11an1n04x5 FILLER_192_640 ();
 b15zdnd11an1n64x5 FILLER_192_647 ();
 b15zdnd11an1n04x5 FILLER_192_711 ();
 b15zdnd00an1n02x5 FILLER_192_715 ();
 b15zdnd00an1n01x5 FILLER_192_717 ();
 b15zdnd11an1n64x5 FILLER_192_726 ();
 b15zdnd11an1n64x5 FILLER_192_790 ();
 b15zdnd11an1n64x5 FILLER_192_854 ();
 b15zdnd11an1n64x5 FILLER_192_918 ();
 b15zdnd11an1n64x5 FILLER_192_982 ();
 b15zdnd11an1n16x5 FILLER_192_1046 ();
 b15zdnd11an1n08x5 FILLER_192_1062 ();
 b15zdnd00an1n01x5 FILLER_192_1070 ();
 b15zdnd11an1n32x5 FILLER_192_1080 ();
 b15zdnd11an1n08x5 FILLER_192_1112 ();
 b15zdnd11an1n04x5 FILLER_192_1120 ();
 b15zdnd11an1n32x5 FILLER_192_1133 ();
 b15zdnd11an1n16x5 FILLER_192_1165 ();
 b15zdnd11an1n04x5 FILLER_192_1181 ();
 b15zdnd00an1n01x5 FILLER_192_1185 ();
 b15zdnd11an1n64x5 FILLER_192_1189 ();
 b15zdnd11an1n08x5 FILLER_192_1253 ();
 b15zdnd11an1n04x5 FILLER_192_1261 ();
 b15zdnd00an1n02x5 FILLER_192_1265 ();
 b15zdnd11an1n32x5 FILLER_192_1273 ();
 b15zdnd00an1n02x5 FILLER_192_1305 ();
 b15zdnd00an1n01x5 FILLER_192_1307 ();
 b15zdnd11an1n64x5 FILLER_192_1322 ();
 b15zdnd11an1n32x5 FILLER_192_1386 ();
 b15zdnd11an1n04x5 FILLER_192_1460 ();
 b15zdnd11an1n08x5 FILLER_192_1476 ();
 b15zdnd11an1n32x5 FILLER_192_1491 ();
 b15zdnd11an1n16x5 FILLER_192_1523 ();
 b15zdnd11an1n04x5 FILLER_192_1539 ();
 b15zdnd00an1n02x5 FILLER_192_1543 ();
 b15zdnd00an1n01x5 FILLER_192_1545 ();
 b15zdnd11an1n64x5 FILLER_192_1564 ();
 b15zdnd11an1n32x5 FILLER_192_1628 ();
 b15zdnd00an1n02x5 FILLER_192_1660 ();
 b15zdnd11an1n08x5 FILLER_192_1679 ();
 b15zdnd11an1n04x5 FILLER_192_1687 ();
 b15zdnd11an1n16x5 FILLER_192_1711 ();
 b15zdnd11an1n08x5 FILLER_192_1727 ();
 b15zdnd11an1n04x5 FILLER_192_1735 ();
 b15zdnd11an1n64x5 FILLER_192_1753 ();
 b15zdnd00an1n01x5 FILLER_192_1817 ();
 b15zdnd11an1n04x5 FILLER_192_1836 ();
 b15zdnd11an1n16x5 FILLER_192_1857 ();
 b15zdnd11an1n08x5 FILLER_192_1873 ();
 b15zdnd00an1n01x5 FILLER_192_1881 ();
 b15zdnd11an1n16x5 FILLER_192_1909 ();
 b15zdnd11an1n08x5 FILLER_192_1925 ();
 b15zdnd11an1n04x5 FILLER_192_1933 ();
 b15zdnd11an1n64x5 FILLER_192_1940 ();
 b15zdnd11an1n04x5 FILLER_192_2004 ();
 b15zdnd11an1n32x5 FILLER_192_2053 ();
 b15zdnd11an1n08x5 FILLER_192_2085 ();
 b15zdnd00an1n01x5 FILLER_192_2093 ();
 b15zdnd11an1n08x5 FILLER_192_2112 ();
 b15zdnd11an1n16x5 FILLER_192_2135 ();
 b15zdnd00an1n02x5 FILLER_192_2151 ();
 b15zdnd00an1n01x5 FILLER_192_2153 ();
 b15zdnd00an1n02x5 FILLER_192_2162 ();
 b15zdnd11an1n32x5 FILLER_192_2184 ();
 b15zdnd00an1n01x5 FILLER_192_2216 ();
 b15zdnd11an1n32x5 FILLER_192_2228 ();
 b15zdnd11an1n16x5 FILLER_192_2260 ();
 b15zdnd11an1n08x5 FILLER_193_0 ();
 b15zdnd11an1n04x5 FILLER_193_8 ();
 b15zdnd00an1n01x5 FILLER_193_12 ();
 b15zdnd11an1n04x5 FILLER_193_19 ();
 b15zdnd00an1n02x5 FILLER_193_23 ();
 b15zdnd00an1n01x5 FILLER_193_25 ();
 b15zdnd11an1n64x5 FILLER_193_30 ();
 b15zdnd11an1n64x5 FILLER_193_94 ();
 b15zdnd11an1n64x5 FILLER_193_158 ();
 b15zdnd00an1n01x5 FILLER_193_222 ();
 b15zdnd11an1n04x5 FILLER_193_226 ();
 b15zdnd11an1n64x5 FILLER_193_233 ();
 b15zdnd11an1n08x5 FILLER_193_297 ();
 b15zdnd00an1n02x5 FILLER_193_305 ();
 b15zdnd11an1n64x5 FILLER_193_359 ();
 b15zdnd11an1n64x5 FILLER_193_423 ();
 b15zdnd11an1n64x5 FILLER_193_487 ();
 b15zdnd11an1n32x5 FILLER_193_551 ();
 b15zdnd11an1n08x5 FILLER_193_583 ();
 b15zdnd11an1n04x5 FILLER_193_591 ();
 b15zdnd00an1n02x5 FILLER_193_595 ();
 b15zdnd00an1n01x5 FILLER_193_597 ();
 b15zdnd11an1n64x5 FILLER_193_650 ();
 b15zdnd11an1n64x5 FILLER_193_714 ();
 b15zdnd11an1n64x5 FILLER_193_778 ();
 b15zdnd11an1n32x5 FILLER_193_842 ();
 b15zdnd11an1n16x5 FILLER_193_874 ();
 b15zdnd00an1n01x5 FILLER_193_890 ();
 b15zdnd11an1n04x5 FILLER_193_894 ();
 b15zdnd11an1n04x5 FILLER_193_901 ();
 b15zdnd11an1n64x5 FILLER_193_908 ();
 b15zdnd11an1n64x5 FILLER_193_972 ();
 b15zdnd11an1n64x5 FILLER_193_1036 ();
 b15zdnd11an1n16x5 FILLER_193_1100 ();
 b15zdnd11an1n04x5 FILLER_193_1116 ();
 b15zdnd00an1n02x5 FILLER_193_1120 ();
 b15zdnd00an1n01x5 FILLER_193_1122 ();
 b15zdnd11an1n64x5 FILLER_193_1132 ();
 b15zdnd11an1n64x5 FILLER_193_1196 ();
 b15zdnd11an1n64x5 FILLER_193_1260 ();
 b15zdnd11an1n64x5 FILLER_193_1324 ();
 b15zdnd11an1n16x5 FILLER_193_1388 ();
 b15zdnd11an1n04x5 FILLER_193_1404 ();
 b15zdnd00an1n02x5 FILLER_193_1408 ();
 b15zdnd11an1n64x5 FILLER_193_1455 ();
 b15zdnd11an1n16x5 FILLER_193_1519 ();
 b15zdnd11an1n08x5 FILLER_193_1535 ();
 b15zdnd00an1n02x5 FILLER_193_1543 ();
 b15zdnd11an1n64x5 FILLER_193_1557 ();
 b15zdnd00an1n02x5 FILLER_193_1621 ();
 b15zdnd00an1n01x5 FILLER_193_1623 ();
 b15zdnd11an1n16x5 FILLER_193_1630 ();
 b15zdnd11an1n08x5 FILLER_193_1646 ();
 b15zdnd00an1n01x5 FILLER_193_1654 ();
 b15zdnd11an1n32x5 FILLER_193_1672 ();
 b15zdnd11an1n08x5 FILLER_193_1704 ();
 b15zdnd00an1n02x5 FILLER_193_1712 ();
 b15zdnd11an1n64x5 FILLER_193_1745 ();
 b15zdnd11an1n08x5 FILLER_193_1809 ();
 b15zdnd11an1n04x5 FILLER_193_1817 ();
 b15zdnd11an1n64x5 FILLER_193_1838 ();
 b15zdnd11an1n08x5 FILLER_193_1902 ();
 b15zdnd11an1n04x5 FILLER_193_1910 ();
 b15zdnd00an1n02x5 FILLER_193_1914 ();
 b15zdnd00an1n01x5 FILLER_193_1916 ();
 b15zdnd11an1n16x5 FILLER_193_1969 ();
 b15zdnd11an1n08x5 FILLER_193_1985 ();
 b15zdnd11an1n64x5 FILLER_193_1999 ();
 b15zdnd11an1n32x5 FILLER_193_2063 ();
 b15zdnd11an1n16x5 FILLER_193_2095 ();
 b15zdnd00an1n02x5 FILLER_193_2111 ();
 b15zdnd11an1n64x5 FILLER_193_2153 ();
 b15zdnd11an1n64x5 FILLER_193_2217 ();
 b15zdnd00an1n02x5 FILLER_193_2281 ();
 b15zdnd00an1n01x5 FILLER_193_2283 ();
 b15zdnd00an1n02x5 FILLER_194_8 ();
 b15zdnd11an1n08x5 FILLER_194_52 ();
 b15zdnd11an1n64x5 FILLER_194_65 ();
 b15zdnd11an1n64x5 FILLER_194_129 ();
 b15zdnd11an1n64x5 FILLER_194_193 ();
 b15zdnd11an1n64x5 FILLER_194_257 ();
 b15zdnd11an1n08x5 FILLER_194_321 ();
 b15zdnd00an1n02x5 FILLER_194_329 ();
 b15zdnd11an1n64x5 FILLER_194_334 ();
 b15zdnd11an1n64x5 FILLER_194_398 ();
 b15zdnd11an1n64x5 FILLER_194_462 ();
 b15zdnd11an1n64x5 FILLER_194_526 ();
 b15zdnd11an1n08x5 FILLER_194_590 ();
 b15zdnd00an1n01x5 FILLER_194_598 ();
 b15zdnd11an1n04x5 FILLER_194_651 ();
 b15zdnd11an1n04x5 FILLER_194_658 ();
 b15zdnd11an1n32x5 FILLER_194_669 ();
 b15zdnd11an1n16x5 FILLER_194_701 ();
 b15zdnd00an1n01x5 FILLER_194_717 ();
 b15zdnd11an1n32x5 FILLER_194_726 ();
 b15zdnd11an1n16x5 FILLER_194_758 ();
 b15zdnd11an1n04x5 FILLER_194_774 ();
 b15zdnd00an1n02x5 FILLER_194_778 ();
 b15zdnd11an1n64x5 FILLER_194_783 ();
 b15zdnd11an1n16x5 FILLER_194_847 ();
 b15zdnd11an1n08x5 FILLER_194_863 ();
 b15zdnd11an1n64x5 FILLER_194_923 ();
 b15zdnd11an1n64x5 FILLER_194_987 ();
 b15zdnd11an1n64x5 FILLER_194_1051 ();
 b15zdnd11an1n64x5 FILLER_194_1115 ();
 b15zdnd11an1n64x5 FILLER_194_1179 ();
 b15zdnd11an1n32x5 FILLER_194_1243 ();
 b15zdnd11an1n08x5 FILLER_194_1275 ();
 b15zdnd11an1n04x5 FILLER_194_1283 ();
 b15zdnd00an1n02x5 FILLER_194_1287 ();
 b15zdnd00an1n01x5 FILLER_194_1289 ();
 b15zdnd11an1n32x5 FILLER_194_1304 ();
 b15zdnd11an1n16x5 FILLER_194_1336 ();
 b15zdnd11an1n08x5 FILLER_194_1352 ();
 b15zdnd11an1n04x5 FILLER_194_1360 ();
 b15zdnd00an1n02x5 FILLER_194_1364 ();
 b15zdnd11an1n32x5 FILLER_194_1374 ();
 b15zdnd11an1n04x5 FILLER_194_1406 ();
 b15zdnd11an1n64x5 FILLER_194_1413 ();
 b15zdnd11an1n16x5 FILLER_194_1477 ();
 b15zdnd11an1n08x5 FILLER_194_1493 ();
 b15zdnd00an1n01x5 FILLER_194_1501 ();
 b15zdnd11an1n04x5 FILLER_194_1522 ();
 b15zdnd11an1n16x5 FILLER_194_1540 ();
 b15zdnd00an1n02x5 FILLER_194_1556 ();
 b15zdnd11an1n64x5 FILLER_194_1563 ();
 b15zdnd11an1n64x5 FILLER_194_1627 ();
 b15zdnd11an1n64x5 FILLER_194_1691 ();
 b15zdnd11an1n64x5 FILLER_194_1755 ();
 b15zdnd11an1n64x5 FILLER_194_1819 ();
 b15zdnd11an1n64x5 FILLER_194_1883 ();
 b15zdnd11an1n64x5 FILLER_194_1947 ();
 b15zdnd11an1n64x5 FILLER_194_2011 ();
 b15zdnd11an1n64x5 FILLER_194_2075 ();
 b15zdnd11an1n08x5 FILLER_194_2139 ();
 b15zdnd11an1n04x5 FILLER_194_2147 ();
 b15zdnd00an1n02x5 FILLER_194_2151 ();
 b15zdnd00an1n01x5 FILLER_194_2153 ();
 b15zdnd11an1n64x5 FILLER_194_2162 ();
 b15zdnd11an1n32x5 FILLER_194_2226 ();
 b15zdnd11an1n16x5 FILLER_194_2258 ();
 b15zdnd00an1n02x5 FILLER_194_2274 ();
 b15zdnd11an1n08x5 FILLER_195_0 ();
 b15zdnd11an1n04x5 FILLER_195_8 ();
 b15zdnd00an1n01x5 FILLER_195_12 ();
 b15zdnd11an1n04x5 FILLER_195_17 ();
 b15zdnd11an1n04x5 FILLER_195_25 ();
 b15zdnd11an1n64x5 FILLER_195_33 ();
 b15zdnd11an1n64x5 FILLER_195_97 ();
 b15zdnd11an1n64x5 FILLER_195_161 ();
 b15zdnd11an1n64x5 FILLER_195_225 ();
 b15zdnd11an1n32x5 FILLER_195_289 ();
 b15zdnd11an1n08x5 FILLER_195_321 ();
 b15zdnd11an1n04x5 FILLER_195_329 ();
 b15zdnd11an1n08x5 FILLER_195_336 ();
 b15zdnd00an1n02x5 FILLER_195_344 ();
 b15zdnd00an1n01x5 FILLER_195_346 ();
 b15zdnd11an1n64x5 FILLER_195_350 ();
 b15zdnd11an1n64x5 FILLER_195_414 ();
 b15zdnd11an1n64x5 FILLER_195_478 ();
 b15zdnd11an1n32x5 FILLER_195_542 ();
 b15zdnd11an1n16x5 FILLER_195_574 ();
 b15zdnd11an1n08x5 FILLER_195_590 ();
 b15zdnd00an1n01x5 FILLER_195_598 ();
 b15zdnd11an1n08x5 FILLER_195_605 ();
 b15zdnd11an1n04x5 FILLER_195_613 ();
 b15zdnd11an1n64x5 FILLER_195_669 ();
 b15zdnd11an1n16x5 FILLER_195_733 ();
 b15zdnd11an1n04x5 FILLER_195_749 ();
 b15zdnd11an1n32x5 FILLER_195_805 ();
 b15zdnd11an1n16x5 FILLER_195_837 ();
 b15zdnd11an1n08x5 FILLER_195_853 ();
 b15zdnd11an1n04x5 FILLER_195_861 ();
 b15zdnd11an1n16x5 FILLER_195_917 ();
 b15zdnd11an1n08x5 FILLER_195_933 ();
 b15zdnd00an1n02x5 FILLER_195_941 ();
 b15zdnd11an1n64x5 FILLER_195_949 ();
 b15zdnd11an1n64x5 FILLER_195_1013 ();
 b15zdnd11an1n64x5 FILLER_195_1077 ();
 b15zdnd11an1n64x5 FILLER_195_1141 ();
 b15zdnd11an1n64x5 FILLER_195_1205 ();
 b15zdnd11an1n16x5 FILLER_195_1269 ();
 b15zdnd11an1n08x5 FILLER_195_1285 ();
 b15zdnd00an1n02x5 FILLER_195_1293 ();
 b15zdnd11an1n04x5 FILLER_195_1306 ();
 b15zdnd11an1n04x5 FILLER_195_1326 ();
 b15zdnd00an1n02x5 FILLER_195_1330 ();
 b15zdnd11an1n32x5 FILLER_195_1346 ();
 b15zdnd11an1n04x5 FILLER_195_1378 ();
 b15zdnd00an1n02x5 FILLER_195_1382 ();
 b15zdnd11an1n64x5 FILLER_195_1436 ();
 b15zdnd11an1n16x5 FILLER_195_1500 ();
 b15zdnd11an1n08x5 FILLER_195_1536 ();
 b15zdnd11an1n64x5 FILLER_195_1563 ();
 b15zdnd11an1n32x5 FILLER_195_1627 ();
 b15zdnd11an1n08x5 FILLER_195_1659 ();
 b15zdnd00an1n02x5 FILLER_195_1667 ();
 b15zdnd00an1n01x5 FILLER_195_1669 ();
 b15zdnd11an1n04x5 FILLER_195_1674 ();
 b15zdnd11an1n64x5 FILLER_195_1709 ();
 b15zdnd11an1n64x5 FILLER_195_1773 ();
 b15zdnd11an1n64x5 FILLER_195_1851 ();
 b15zdnd11an1n64x5 FILLER_195_1915 ();
 b15zdnd11an1n64x5 FILLER_195_1979 ();
 b15zdnd11an1n64x5 FILLER_195_2043 ();
 b15zdnd11an1n16x5 FILLER_195_2138 ();
 b15zdnd00an1n02x5 FILLER_195_2154 ();
 b15zdnd11an1n32x5 FILLER_195_2201 ();
 b15zdnd11an1n16x5 FILLER_195_2233 ();
 b15zdnd00an1n01x5 FILLER_195_2249 ();
 b15zdnd11an1n16x5 FILLER_195_2264 ();
 b15zdnd11an1n04x5 FILLER_195_2280 ();
 b15zdnd00an1n02x5 FILLER_196_8 ();
 b15zdnd11an1n64x5 FILLER_196_52 ();
 b15zdnd11an1n64x5 FILLER_196_116 ();
 b15zdnd11an1n64x5 FILLER_196_180 ();
 b15zdnd11an1n16x5 FILLER_196_244 ();
 b15zdnd11an1n04x5 FILLER_196_260 ();
 b15zdnd00an1n02x5 FILLER_196_264 ();
 b15zdnd11an1n64x5 FILLER_196_308 ();
 b15zdnd11an1n64x5 FILLER_196_372 ();
 b15zdnd11an1n64x5 FILLER_196_436 ();
 b15zdnd11an1n64x5 FILLER_196_500 ();
 b15zdnd11an1n32x5 FILLER_196_564 ();
 b15zdnd11an1n08x5 FILLER_196_596 ();
 b15zdnd11an1n32x5 FILLER_196_656 ();
 b15zdnd11an1n16x5 FILLER_196_688 ();
 b15zdnd11an1n08x5 FILLER_196_704 ();
 b15zdnd11an1n04x5 FILLER_196_712 ();
 b15zdnd00an1n02x5 FILLER_196_716 ();
 b15zdnd11an1n32x5 FILLER_196_726 ();
 b15zdnd11an1n08x5 FILLER_196_758 ();
 b15zdnd11an1n04x5 FILLER_196_766 ();
 b15zdnd00an1n01x5 FILLER_196_770 ();
 b15zdnd11an1n04x5 FILLER_196_774 ();
 b15zdnd11an1n64x5 FILLER_196_781 ();
 b15zdnd11an1n32x5 FILLER_196_845 ();
 b15zdnd11an1n08x5 FILLER_196_877 ();
 b15zdnd11an1n04x5 FILLER_196_888 ();
 b15zdnd11an1n04x5 FILLER_196_895 ();
 b15zdnd11an1n64x5 FILLER_196_902 ();
 b15zdnd11an1n64x5 FILLER_196_966 ();
 b15zdnd11an1n16x5 FILLER_196_1030 ();
 b15zdnd11an1n04x5 FILLER_196_1046 ();
 b15zdnd11an1n64x5 FILLER_196_1053 ();
 b15zdnd11an1n64x5 FILLER_196_1117 ();
 b15zdnd11an1n64x5 FILLER_196_1181 ();
 b15zdnd11an1n32x5 FILLER_196_1245 ();
 b15zdnd11an1n16x5 FILLER_196_1277 ();
 b15zdnd11an1n08x5 FILLER_196_1293 ();
 b15zdnd11an1n04x5 FILLER_196_1301 ();
 b15zdnd00an1n02x5 FILLER_196_1305 ();
 b15zdnd11an1n04x5 FILLER_196_1318 ();
 b15zdnd00an1n02x5 FILLER_196_1322 ();
 b15zdnd11an1n64x5 FILLER_196_1332 ();
 b15zdnd11an1n08x5 FILLER_196_1396 ();
 b15zdnd11an1n04x5 FILLER_196_1404 ();
 b15zdnd00an1n01x5 FILLER_196_1408 ();
 b15zdnd11an1n64x5 FILLER_196_1412 ();
 b15zdnd11an1n32x5 FILLER_196_1476 ();
 b15zdnd11an1n08x5 FILLER_196_1508 ();
 b15zdnd00an1n01x5 FILLER_196_1516 ();
 b15zdnd11an1n04x5 FILLER_196_1542 ();
 b15zdnd11an1n08x5 FILLER_196_1561 ();
 b15zdnd11an1n64x5 FILLER_196_1578 ();
 b15zdnd11an1n64x5 FILLER_196_1642 ();
 b15zdnd11an1n16x5 FILLER_196_1706 ();
 b15zdnd11an1n08x5 FILLER_196_1730 ();
 b15zdnd11an1n04x5 FILLER_196_1738 ();
 b15zdnd00an1n02x5 FILLER_196_1742 ();
 b15zdnd11an1n32x5 FILLER_196_1762 ();
 b15zdnd11an1n16x5 FILLER_196_1794 ();
 b15zdnd00an1n02x5 FILLER_196_1810 ();
 b15zdnd11an1n64x5 FILLER_196_1823 ();
 b15zdnd11an1n64x5 FILLER_196_1887 ();
 b15zdnd11an1n64x5 FILLER_196_1951 ();
 b15zdnd11an1n64x5 FILLER_196_2015 ();
 b15zdnd11an1n16x5 FILLER_196_2079 ();
 b15zdnd11an1n04x5 FILLER_196_2095 ();
 b15zdnd11an1n16x5 FILLER_196_2130 ();
 b15zdnd11an1n08x5 FILLER_196_2146 ();
 b15zdnd11an1n64x5 FILLER_196_2162 ();
 b15zdnd11an1n16x5 FILLER_196_2226 ();
 b15zdnd11an1n08x5 FILLER_196_2242 ();
 b15zdnd11an1n04x5 FILLER_196_2250 ();
 b15zdnd11an1n08x5 FILLER_196_2268 ();
 b15zdnd11an1n16x5 FILLER_197_0 ();
 b15zdnd11an1n04x5 FILLER_197_16 ();
 b15zdnd00an1n02x5 FILLER_197_20 ();
 b15zdnd11an1n64x5 FILLER_197_26 ();
 b15zdnd11an1n64x5 FILLER_197_90 ();
 b15zdnd11an1n64x5 FILLER_197_154 ();
 b15zdnd11an1n64x5 FILLER_197_218 ();
 b15zdnd11an1n64x5 FILLER_197_282 ();
 b15zdnd11an1n64x5 FILLER_197_346 ();
 b15zdnd11an1n64x5 FILLER_197_410 ();
 b15zdnd11an1n64x5 FILLER_197_474 ();
 b15zdnd11an1n64x5 FILLER_197_538 ();
 b15zdnd11an1n04x5 FILLER_197_602 ();
 b15zdnd11an1n08x5 FILLER_197_613 ();
 b15zdnd00an1n01x5 FILLER_197_621 ();
 b15zdnd11an1n04x5 FILLER_197_625 ();
 b15zdnd11an1n04x5 FILLER_197_632 ();
 b15zdnd11an1n08x5 FILLER_197_639 ();
 b15zdnd11an1n64x5 FILLER_197_650 ();
 b15zdnd11an1n64x5 FILLER_197_714 ();
 b15zdnd11an1n64x5 FILLER_197_778 ();
 b15zdnd11an1n64x5 FILLER_197_842 ();
 b15zdnd11an1n04x5 FILLER_197_906 ();
 b15zdnd00an1n02x5 FILLER_197_910 ();
 b15zdnd11an1n64x5 FILLER_197_916 ();
 b15zdnd11an1n32x5 FILLER_197_980 ();
 b15zdnd11an1n16x5 FILLER_197_1012 ();
 b15zdnd11an1n04x5 FILLER_197_1028 ();
 b15zdnd11an1n64x5 FILLER_197_1084 ();
 b15zdnd11an1n16x5 FILLER_197_1148 ();
 b15zdnd11an1n08x5 FILLER_197_1164 ();
 b15zdnd11an1n04x5 FILLER_197_1172 ();
 b15zdnd00an1n02x5 FILLER_197_1176 ();
 b15zdnd11an1n64x5 FILLER_197_1181 ();
 b15zdnd11an1n64x5 FILLER_197_1245 ();
 b15zdnd11an1n08x5 FILLER_197_1309 ();
 b15zdnd11an1n04x5 FILLER_197_1317 ();
 b15zdnd11an1n64x5 FILLER_197_1324 ();
 b15zdnd11an1n16x5 FILLER_197_1388 ();
 b15zdnd11an1n04x5 FILLER_197_1404 ();
 b15zdnd11an1n32x5 FILLER_197_1411 ();
 b15zdnd11an1n08x5 FILLER_197_1443 ();
 b15zdnd00an1n02x5 FILLER_197_1451 ();
 b15zdnd11an1n64x5 FILLER_197_1460 ();
 b15zdnd11an1n64x5 FILLER_197_1524 ();
 b15zdnd11an1n16x5 FILLER_197_1588 ();
 b15zdnd11an1n08x5 FILLER_197_1604 ();
 b15zdnd11an1n64x5 FILLER_197_1616 ();
 b15zdnd11an1n04x5 FILLER_197_1680 ();
 b15zdnd00an1n02x5 FILLER_197_1684 ();
 b15zdnd00an1n01x5 FILLER_197_1686 ();
 b15zdnd11an1n32x5 FILLER_197_1705 ();
 b15zdnd11an1n16x5 FILLER_197_1737 ();
 b15zdnd00an1n02x5 FILLER_197_1753 ();
 b15zdnd00an1n01x5 FILLER_197_1755 ();
 b15zdnd11an1n64x5 FILLER_197_1770 ();
 b15zdnd00an1n02x5 FILLER_197_1834 ();
 b15zdnd00an1n01x5 FILLER_197_1836 ();
 b15zdnd11an1n64x5 FILLER_197_1882 ();
 b15zdnd11an1n64x5 FILLER_197_1946 ();
 b15zdnd11an1n64x5 FILLER_197_2010 ();
 b15zdnd11an1n64x5 FILLER_197_2074 ();
 b15zdnd11an1n64x5 FILLER_197_2138 ();
 b15zdnd11an1n64x5 FILLER_197_2202 ();
 b15zdnd11an1n04x5 FILLER_197_2266 ();
 b15zdnd00an1n01x5 FILLER_197_2270 ();
 b15zdnd11an1n08x5 FILLER_197_2275 ();
 b15zdnd00an1n01x5 FILLER_197_2283 ();
 b15zdnd11an1n64x5 FILLER_198_8 ();
 b15zdnd11an1n64x5 FILLER_198_72 ();
 b15zdnd11an1n64x5 FILLER_198_136 ();
 b15zdnd11an1n16x5 FILLER_198_200 ();
 b15zdnd11an1n08x5 FILLER_198_216 ();
 b15zdnd11an1n04x5 FILLER_198_224 ();
 b15zdnd00an1n01x5 FILLER_198_228 ();
 b15zdnd11an1n04x5 FILLER_198_232 ();
 b15zdnd11an1n64x5 FILLER_198_256 ();
 b15zdnd11an1n64x5 FILLER_198_320 ();
 b15zdnd11an1n64x5 FILLER_198_384 ();
 b15zdnd11an1n32x5 FILLER_198_448 ();
 b15zdnd11an1n16x5 FILLER_198_480 ();
 b15zdnd11an1n04x5 FILLER_198_496 ();
 b15zdnd00an1n02x5 FILLER_198_500 ();
 b15zdnd11an1n64x5 FILLER_198_533 ();
 b15zdnd11an1n16x5 FILLER_198_597 ();
 b15zdnd11an1n04x5 FILLER_198_613 ();
 b15zdnd11an1n04x5 FILLER_198_620 ();
 b15zdnd11an1n04x5 FILLER_198_627 ();
 b15zdnd11an1n04x5 FILLER_198_634 ();
 b15zdnd11an1n32x5 FILLER_198_664 ();
 b15zdnd11an1n16x5 FILLER_198_696 ();
 b15zdnd11an1n04x5 FILLER_198_712 ();
 b15zdnd00an1n02x5 FILLER_198_716 ();
 b15zdnd11an1n64x5 FILLER_198_726 ();
 b15zdnd11an1n64x5 FILLER_198_790 ();
 b15zdnd11an1n64x5 FILLER_198_854 ();
 b15zdnd11an1n64x5 FILLER_198_918 ();
 b15zdnd11an1n32x5 FILLER_198_982 ();
 b15zdnd11an1n08x5 FILLER_198_1014 ();
 b15zdnd00an1n02x5 FILLER_198_1022 ();
 b15zdnd11an1n64x5 FILLER_198_1076 ();
 b15zdnd11an1n16x5 FILLER_198_1140 ();
 b15zdnd11an1n08x5 FILLER_198_1156 ();
 b15zdnd11an1n04x5 FILLER_198_1164 ();
 b15zdnd00an1n02x5 FILLER_198_1168 ();
 b15zdnd11an1n04x5 FILLER_198_1173 ();
 b15zdnd11an1n64x5 FILLER_198_1180 ();
 b15zdnd11an1n32x5 FILLER_198_1244 ();
 b15zdnd11an1n08x5 FILLER_198_1276 ();
 b15zdnd11an1n04x5 FILLER_198_1284 ();
 b15zdnd00an1n01x5 FILLER_198_1288 ();
 b15zdnd11an1n04x5 FILLER_198_1305 ();
 b15zdnd11an1n64x5 FILLER_198_1323 ();
 b15zdnd11an1n32x5 FILLER_198_1387 ();
 b15zdnd00an1n02x5 FILLER_198_1419 ();
 b15zdnd11an1n64x5 FILLER_198_1430 ();
 b15zdnd11an1n64x5 FILLER_198_1494 ();
 b15zdnd11an1n32x5 FILLER_198_1558 ();
 b15zdnd11an1n16x5 FILLER_198_1590 ();
 b15zdnd00an1n02x5 FILLER_198_1606 ();
 b15zdnd00an1n01x5 FILLER_198_1608 ();
 b15zdnd11an1n64x5 FILLER_198_1613 ();
 b15zdnd11an1n64x5 FILLER_198_1677 ();
 b15zdnd11an1n32x5 FILLER_198_1741 ();
 b15zdnd11an1n16x5 FILLER_198_1773 ();
 b15zdnd11an1n08x5 FILLER_198_1789 ();
 b15zdnd11an1n04x5 FILLER_198_1797 ();
 b15zdnd00an1n01x5 FILLER_198_1801 ();
 b15zdnd11an1n16x5 FILLER_198_1822 ();
 b15zdnd00an1n01x5 FILLER_198_1838 ();
 b15zdnd11an1n64x5 FILLER_198_1847 ();
 b15zdnd11an1n64x5 FILLER_198_1911 ();
 b15zdnd11an1n64x5 FILLER_198_1975 ();
 b15zdnd11an1n64x5 FILLER_198_2039 ();
 b15zdnd11an1n32x5 FILLER_198_2103 ();
 b15zdnd11an1n16x5 FILLER_198_2135 ();
 b15zdnd00an1n02x5 FILLER_198_2151 ();
 b15zdnd00an1n01x5 FILLER_198_2153 ();
 b15zdnd11an1n64x5 FILLER_198_2162 ();
 b15zdnd11an1n32x5 FILLER_198_2226 ();
 b15zdnd00an1n02x5 FILLER_198_2258 ();
 b15zdnd11an1n04x5 FILLER_198_2271 ();
 b15zdnd00an1n01x5 FILLER_198_2275 ();
 b15zdnd11an1n64x5 FILLER_199_0 ();
 b15zdnd11an1n64x5 FILLER_199_64 ();
 b15zdnd11an1n64x5 FILLER_199_128 ();
 b15zdnd11an1n08x5 FILLER_199_192 ();
 b15zdnd00an1n02x5 FILLER_199_200 ();
 b15zdnd00an1n01x5 FILLER_199_202 ();
 b15zdnd11an1n64x5 FILLER_199_255 ();
 b15zdnd11an1n64x5 FILLER_199_319 ();
 b15zdnd11an1n64x5 FILLER_199_383 ();
 b15zdnd11an1n64x5 FILLER_199_447 ();
 b15zdnd11an1n64x5 FILLER_199_511 ();
 b15zdnd11an1n64x5 FILLER_199_575 ();
 b15zdnd11an1n64x5 FILLER_199_639 ();
 b15zdnd11an1n64x5 FILLER_199_703 ();
 b15zdnd11an1n64x5 FILLER_199_767 ();
 b15zdnd11an1n64x5 FILLER_199_831 ();
 b15zdnd11an1n64x5 FILLER_199_895 ();
 b15zdnd11an1n64x5 FILLER_199_959 ();
 b15zdnd11an1n16x5 FILLER_199_1023 ();
 b15zdnd11an1n04x5 FILLER_199_1039 ();
 b15zdnd11an1n04x5 FILLER_199_1046 ();
 b15zdnd11an1n04x5 FILLER_199_1053 ();
 b15zdnd11an1n04x5 FILLER_199_1060 ();
 b15zdnd11an1n64x5 FILLER_199_1067 ();
 b15zdnd11an1n16x5 FILLER_199_1131 ();
 b15zdnd11an1n04x5 FILLER_199_1147 ();
 b15zdnd00an1n01x5 FILLER_199_1151 ();
 b15zdnd11an1n64x5 FILLER_199_1204 ();
 b15zdnd11an1n32x5 FILLER_199_1268 ();
 b15zdnd11an1n08x5 FILLER_199_1300 ();
 b15zdnd00an1n02x5 FILLER_199_1308 ();
 b15zdnd11an1n64x5 FILLER_199_1317 ();
 b15zdnd11an1n64x5 FILLER_199_1381 ();
 b15zdnd11an1n32x5 FILLER_199_1445 ();
 b15zdnd11an1n16x5 FILLER_199_1477 ();
 b15zdnd11an1n08x5 FILLER_199_1493 ();
 b15zdnd00an1n02x5 FILLER_199_1501 ();
 b15zdnd11an1n64x5 FILLER_199_1519 ();
 b15zdnd11an1n64x5 FILLER_199_1583 ();
 b15zdnd11an1n64x5 FILLER_199_1647 ();
 b15zdnd11an1n64x5 FILLER_199_1711 ();
 b15zdnd11an1n32x5 FILLER_199_1775 ();
 b15zdnd11an1n16x5 FILLER_199_1807 ();
 b15zdnd11an1n04x5 FILLER_199_1823 ();
 b15zdnd00an1n01x5 FILLER_199_1827 ();
 b15zdnd11an1n64x5 FILLER_199_1840 ();
 b15zdnd11an1n64x5 FILLER_199_1904 ();
 b15zdnd11an1n64x5 FILLER_199_1968 ();
 b15zdnd11an1n64x5 FILLER_199_2032 ();
 b15zdnd11an1n64x5 FILLER_199_2096 ();
 b15zdnd11an1n64x5 FILLER_199_2160 ();
 b15zdnd11an1n08x5 FILLER_199_2224 ();
 b15zdnd11an1n04x5 FILLER_199_2232 ();
 b15zdnd00an1n01x5 FILLER_199_2236 ();
 b15zdnd11an1n16x5 FILLER_199_2245 ();
 b15zdnd11an1n08x5 FILLER_199_2261 ();
 b15zdnd11an1n04x5 FILLER_199_2269 ();
 b15zdnd00an1n02x5 FILLER_199_2273 ();
 b15zdnd00an1n01x5 FILLER_199_2275 ();
 b15zdnd00an1n02x5 FILLER_199_2282 ();
 b15zdnd11an1n64x5 FILLER_200_8 ();
 b15zdnd11an1n64x5 FILLER_200_72 ();
 b15zdnd11an1n64x5 FILLER_200_136 ();
 b15zdnd11an1n16x5 FILLER_200_200 ();
 b15zdnd11an1n08x5 FILLER_200_216 ();
 b15zdnd00an1n01x5 FILLER_200_224 ();
 b15zdnd11an1n04x5 FILLER_200_228 ();
 b15zdnd11an1n16x5 FILLER_200_235 ();
 b15zdnd11an1n08x5 FILLER_200_251 ();
 b15zdnd00an1n02x5 FILLER_200_259 ();
 b15zdnd11an1n64x5 FILLER_200_281 ();
 b15zdnd11an1n64x5 FILLER_200_345 ();
 b15zdnd11an1n64x5 FILLER_200_409 ();
 b15zdnd11an1n64x5 FILLER_200_473 ();
 b15zdnd11an1n64x5 FILLER_200_537 ();
 b15zdnd11an1n64x5 FILLER_200_601 ();
 b15zdnd11an1n32x5 FILLER_200_665 ();
 b15zdnd11an1n16x5 FILLER_200_697 ();
 b15zdnd11an1n04x5 FILLER_200_713 ();
 b15zdnd00an1n01x5 FILLER_200_717 ();
 b15zdnd11an1n64x5 FILLER_200_726 ();
 b15zdnd11an1n64x5 FILLER_200_790 ();
 b15zdnd11an1n64x5 FILLER_200_854 ();
 b15zdnd11an1n64x5 FILLER_200_918 ();
 b15zdnd11an1n64x5 FILLER_200_982 ();
 b15zdnd11an1n08x5 FILLER_200_1046 ();
 b15zdnd00an1n02x5 FILLER_200_1054 ();
 b15zdnd00an1n01x5 FILLER_200_1056 ();
 b15zdnd11an1n64x5 FILLER_200_1060 ();
 b15zdnd11an1n32x5 FILLER_200_1124 ();
 b15zdnd11an1n64x5 FILLER_200_1182 ();
 b15zdnd11an1n64x5 FILLER_200_1246 ();
 b15zdnd11an1n64x5 FILLER_200_1310 ();
 b15zdnd11an1n64x5 FILLER_200_1374 ();
 b15zdnd11an1n64x5 FILLER_200_1438 ();
 b15zdnd11an1n64x5 FILLER_200_1502 ();
 b15zdnd11an1n64x5 FILLER_200_1566 ();
 b15zdnd11an1n64x5 FILLER_200_1630 ();
 b15zdnd11an1n64x5 FILLER_200_1694 ();
 b15zdnd11an1n64x5 FILLER_200_1758 ();
 b15zdnd11an1n08x5 FILLER_200_1822 ();
 b15zdnd11an1n04x5 FILLER_200_1830 ();
 b15zdnd11an1n64x5 FILLER_200_1876 ();
 b15zdnd11an1n64x5 FILLER_200_1940 ();
 b15zdnd11an1n64x5 FILLER_200_2004 ();
 b15zdnd11an1n64x5 FILLER_200_2068 ();
 b15zdnd11an1n16x5 FILLER_200_2132 ();
 b15zdnd11an1n04x5 FILLER_200_2148 ();
 b15zdnd00an1n02x5 FILLER_200_2152 ();
 b15zdnd00an1n02x5 FILLER_200_2162 ();
 b15zdnd00an1n01x5 FILLER_200_2164 ();
 b15zdnd11an1n64x5 FILLER_200_2179 ();
 b15zdnd11an1n08x5 FILLER_200_2243 ();
 b15zdnd00an1n02x5 FILLER_200_2251 ();
 b15zdnd00an1n01x5 FILLER_200_2253 ();
 b15zdnd11an1n08x5 FILLER_200_2262 ();
 b15zdnd11an1n04x5 FILLER_200_2270 ();
 b15zdnd00an1n02x5 FILLER_200_2274 ();
 b15zdnd11an1n16x5 FILLER_201_0 ();
 b15zdnd00an1n02x5 FILLER_201_16 ();
 b15zdnd00an1n01x5 FILLER_201_18 ();
 b15zdnd11an1n64x5 FILLER_201_23 ();
 b15zdnd11an1n64x5 FILLER_201_87 ();
 b15zdnd11an1n64x5 FILLER_201_151 ();
 b15zdnd11an1n64x5 FILLER_201_215 ();
 b15zdnd11an1n64x5 FILLER_201_279 ();
 b15zdnd11an1n08x5 FILLER_201_343 ();
 b15zdnd11an1n04x5 FILLER_201_351 ();
 b15zdnd00an1n01x5 FILLER_201_355 ();
 b15zdnd11an1n04x5 FILLER_201_361 ();
 b15zdnd11an1n64x5 FILLER_201_369 ();
 b15zdnd11an1n32x5 FILLER_201_433 ();
 b15zdnd11an1n08x5 FILLER_201_465 ();
 b15zdnd00an1n01x5 FILLER_201_473 ();
 b15zdnd11an1n64x5 FILLER_201_516 ();
 b15zdnd11an1n64x5 FILLER_201_580 ();
 b15zdnd11an1n64x5 FILLER_201_644 ();
 b15zdnd11an1n64x5 FILLER_201_708 ();
 b15zdnd11an1n64x5 FILLER_201_772 ();
 b15zdnd11an1n64x5 FILLER_201_836 ();
 b15zdnd11an1n64x5 FILLER_201_900 ();
 b15zdnd11an1n64x5 FILLER_201_964 ();
 b15zdnd11an1n64x5 FILLER_201_1028 ();
 b15zdnd11an1n64x5 FILLER_201_1092 ();
 b15zdnd11an1n16x5 FILLER_201_1156 ();
 b15zdnd11an1n08x5 FILLER_201_1172 ();
 b15zdnd00an1n02x5 FILLER_201_1180 ();
 b15zdnd11an1n64x5 FILLER_201_1208 ();
 b15zdnd11an1n64x5 FILLER_201_1272 ();
 b15zdnd11an1n64x5 FILLER_201_1336 ();
 b15zdnd11an1n64x5 FILLER_201_1400 ();
 b15zdnd11an1n64x5 FILLER_201_1464 ();
 b15zdnd11an1n64x5 FILLER_201_1528 ();
 b15zdnd11an1n64x5 FILLER_201_1592 ();
 b15zdnd11an1n64x5 FILLER_201_1656 ();
 b15zdnd11an1n64x5 FILLER_201_1720 ();
 b15zdnd11an1n16x5 FILLER_201_1784 ();
 b15zdnd11an1n08x5 FILLER_201_1800 ();
 b15zdnd11an1n04x5 FILLER_201_1808 ();
 b15zdnd00an1n02x5 FILLER_201_1812 ();
 b15zdnd11an1n64x5 FILLER_201_1822 ();
 b15zdnd11an1n64x5 FILLER_201_1886 ();
 b15zdnd11an1n64x5 FILLER_201_1950 ();
 b15zdnd11an1n64x5 FILLER_201_2014 ();
 b15zdnd11an1n64x5 FILLER_201_2078 ();
 b15zdnd11an1n64x5 FILLER_201_2156 ();
 b15zdnd11an1n64x5 FILLER_201_2220 ();
 b15zdnd11an1n08x5 FILLER_202_8 ();
 b15zdnd11an1n04x5 FILLER_202_16 ();
 b15zdnd00an1n01x5 FILLER_202_20 ();
 b15zdnd11an1n64x5 FILLER_202_25 ();
 b15zdnd11an1n64x5 FILLER_202_89 ();
 b15zdnd11an1n64x5 FILLER_202_153 ();
 b15zdnd11an1n64x5 FILLER_202_217 ();
 b15zdnd11an1n16x5 FILLER_202_281 ();
 b15zdnd11an1n04x5 FILLER_202_297 ();
 b15zdnd11an1n16x5 FILLER_202_343 ();
 b15zdnd11an1n04x5 FILLER_202_359 ();
 b15zdnd11an1n32x5 FILLER_202_368 ();
 b15zdnd00an1n02x5 FILLER_202_400 ();
 b15zdnd11an1n04x5 FILLER_202_444 ();
 b15zdnd00an1n02x5 FILLER_202_448 ();
 b15zdnd11an1n04x5 FILLER_202_453 ();
 b15zdnd11an1n64x5 FILLER_202_460 ();
 b15zdnd11an1n64x5 FILLER_202_524 ();
 b15zdnd11an1n32x5 FILLER_202_588 ();
 b15zdnd11an1n04x5 FILLER_202_620 ();
 b15zdnd00an1n02x5 FILLER_202_624 ();
 b15zdnd00an1n01x5 FILLER_202_626 ();
 b15zdnd11an1n64x5 FILLER_202_636 ();
 b15zdnd11an1n16x5 FILLER_202_700 ();
 b15zdnd00an1n02x5 FILLER_202_716 ();
 b15zdnd11an1n64x5 FILLER_202_726 ();
 b15zdnd11an1n64x5 FILLER_202_790 ();
 b15zdnd11an1n64x5 FILLER_202_854 ();
 b15zdnd11an1n64x5 FILLER_202_918 ();
 b15zdnd11an1n16x5 FILLER_202_982 ();
 b15zdnd11an1n08x5 FILLER_202_998 ();
 b15zdnd00an1n02x5 FILLER_202_1006 ();
 b15zdnd00an1n01x5 FILLER_202_1008 ();
 b15zdnd11an1n64x5 FILLER_202_1013 ();
 b15zdnd11an1n64x5 FILLER_202_1077 ();
 b15zdnd11an1n64x5 FILLER_202_1141 ();
 b15zdnd11an1n64x5 FILLER_202_1205 ();
 b15zdnd11an1n32x5 FILLER_202_1269 ();
 b15zdnd11an1n08x5 FILLER_202_1301 ();
 b15zdnd11an1n64x5 FILLER_202_1312 ();
 b15zdnd11an1n64x5 FILLER_202_1376 ();
 b15zdnd11an1n64x5 FILLER_202_1440 ();
 b15zdnd11an1n64x5 FILLER_202_1504 ();
 b15zdnd00an1n02x5 FILLER_202_1568 ();
 b15zdnd00an1n01x5 FILLER_202_1570 ();
 b15zdnd11an1n64x5 FILLER_202_1580 ();
 b15zdnd11an1n16x5 FILLER_202_1644 ();
 b15zdnd11an1n04x5 FILLER_202_1660 ();
 b15zdnd11an1n64x5 FILLER_202_1706 ();
 b15zdnd11an1n32x5 FILLER_202_1770 ();
 b15zdnd11an1n16x5 FILLER_202_1802 ();
 b15zdnd11an1n04x5 FILLER_202_1818 ();
 b15zdnd00an1n01x5 FILLER_202_1822 ();
 b15zdnd11an1n64x5 FILLER_202_1841 ();
 b15zdnd11an1n16x5 FILLER_202_1905 ();
 b15zdnd11an1n08x5 FILLER_202_1921 ();
 b15zdnd11an1n04x5 FILLER_202_1929 ();
 b15zdnd00an1n01x5 FILLER_202_1933 ();
 b15zdnd11an1n64x5 FILLER_202_1939 ();
 b15zdnd11an1n64x5 FILLER_202_2003 ();
 b15zdnd11an1n16x5 FILLER_202_2067 ();
 b15zdnd11an1n08x5 FILLER_202_2083 ();
 b15zdnd11an1n04x5 FILLER_202_2091 ();
 b15zdnd11an1n32x5 FILLER_202_2107 ();
 b15zdnd11an1n08x5 FILLER_202_2139 ();
 b15zdnd11an1n04x5 FILLER_202_2147 ();
 b15zdnd00an1n02x5 FILLER_202_2151 ();
 b15zdnd00an1n01x5 FILLER_202_2153 ();
 b15zdnd11an1n16x5 FILLER_202_2162 ();
 b15zdnd11an1n08x5 FILLER_202_2178 ();
 b15zdnd11an1n04x5 FILLER_202_2186 ();
 b15zdnd00an1n02x5 FILLER_202_2190 ();
 b15zdnd11an1n04x5 FILLER_202_2206 ();
 b15zdnd00an1n01x5 FILLER_202_2210 ();
 b15zdnd11an1n32x5 FILLER_202_2237 ();
 b15zdnd11an1n04x5 FILLER_202_2269 ();
 b15zdnd00an1n02x5 FILLER_202_2273 ();
 b15zdnd00an1n01x5 FILLER_202_2275 ();
 b15zdnd11an1n64x5 FILLER_203_0 ();
 b15zdnd11an1n64x5 FILLER_203_64 ();
 b15zdnd11an1n64x5 FILLER_203_128 ();
 b15zdnd11an1n64x5 FILLER_203_192 ();
 b15zdnd11an1n64x5 FILLER_203_256 ();
 b15zdnd11an1n32x5 FILLER_203_320 ();
 b15zdnd11an1n04x5 FILLER_203_352 ();
 b15zdnd00an1n02x5 FILLER_203_356 ();
 b15zdnd00an1n01x5 FILLER_203_358 ();
 b15zdnd11an1n32x5 FILLER_203_369 ();
 b15zdnd11an1n16x5 FILLER_203_401 ();
 b15zdnd11an1n04x5 FILLER_203_417 ();
 b15zdnd00an1n01x5 FILLER_203_421 ();
 b15zdnd11an1n64x5 FILLER_203_464 ();
 b15zdnd11an1n64x5 FILLER_203_528 ();
 b15zdnd11an1n64x5 FILLER_203_592 ();
 b15zdnd11an1n64x5 FILLER_203_656 ();
 b15zdnd11an1n64x5 FILLER_203_720 ();
 b15zdnd11an1n64x5 FILLER_203_784 ();
 b15zdnd11an1n64x5 FILLER_203_848 ();
 b15zdnd11an1n64x5 FILLER_203_912 ();
 b15zdnd11an1n64x5 FILLER_203_976 ();
 b15zdnd11an1n64x5 FILLER_203_1040 ();
 b15zdnd11an1n64x5 FILLER_203_1104 ();
 b15zdnd11an1n64x5 FILLER_203_1168 ();
 b15zdnd11an1n64x5 FILLER_203_1232 ();
 b15zdnd11an1n64x5 FILLER_203_1296 ();
 b15zdnd11an1n64x5 FILLER_203_1360 ();
 b15zdnd11an1n64x5 FILLER_203_1424 ();
 b15zdnd11an1n64x5 FILLER_203_1488 ();
 b15zdnd11an1n64x5 FILLER_203_1552 ();
 b15zdnd11an1n08x5 FILLER_203_1616 ();
 b15zdnd00an1n02x5 FILLER_203_1624 ();
 b15zdnd11an1n64x5 FILLER_203_1634 ();
 b15zdnd11an1n64x5 FILLER_203_1698 ();
 b15zdnd11an1n64x5 FILLER_203_1762 ();
 b15zdnd11an1n64x5 FILLER_203_1826 ();
 b15zdnd11an1n64x5 FILLER_203_1890 ();
 b15zdnd11an1n64x5 FILLER_203_1954 ();
 b15zdnd11an1n64x5 FILLER_203_2018 ();
 b15zdnd11an1n64x5 FILLER_203_2082 ();
 b15zdnd11an1n64x5 FILLER_203_2146 ();
 b15zdnd11an1n64x5 FILLER_203_2210 ();
 b15zdnd11an1n08x5 FILLER_203_2274 ();
 b15zdnd00an1n02x5 FILLER_203_2282 ();
 b15zdnd11an1n64x5 FILLER_204_8 ();
 b15zdnd11an1n64x5 FILLER_204_72 ();
 b15zdnd11an1n64x5 FILLER_204_136 ();
 b15zdnd11an1n64x5 FILLER_204_200 ();
 b15zdnd11an1n64x5 FILLER_204_264 ();
 b15zdnd11an1n16x5 FILLER_204_328 ();
 b15zdnd11an1n08x5 FILLER_204_344 ();
 b15zdnd00an1n02x5 FILLER_204_352 ();
 b15zdnd11an1n04x5 FILLER_204_367 ();
 b15zdnd11an1n32x5 FILLER_204_386 ();
 b15zdnd11an1n08x5 FILLER_204_418 ();
 b15zdnd00an1n01x5 FILLER_204_426 ();
 b15zdnd11an1n64x5 FILLER_204_479 ();
 b15zdnd11an1n64x5 FILLER_204_543 ();
 b15zdnd11an1n64x5 FILLER_204_607 ();
 b15zdnd11an1n32x5 FILLER_204_671 ();
 b15zdnd11an1n08x5 FILLER_204_703 ();
 b15zdnd11an1n04x5 FILLER_204_711 ();
 b15zdnd00an1n02x5 FILLER_204_715 ();
 b15zdnd00an1n01x5 FILLER_204_717 ();
 b15zdnd11an1n64x5 FILLER_204_726 ();
 b15zdnd11an1n64x5 FILLER_204_790 ();
 b15zdnd11an1n64x5 FILLER_204_854 ();
 b15zdnd11an1n64x5 FILLER_204_918 ();
 b15zdnd11an1n32x5 FILLER_204_982 ();
 b15zdnd00an1n01x5 FILLER_204_1014 ();
 b15zdnd11an1n64x5 FILLER_204_1029 ();
 b15zdnd11an1n64x5 FILLER_204_1093 ();
 b15zdnd11an1n64x5 FILLER_204_1157 ();
 b15zdnd11an1n64x5 FILLER_204_1221 ();
 b15zdnd11an1n64x5 FILLER_204_1285 ();
 b15zdnd11an1n64x5 FILLER_204_1349 ();
 b15zdnd11an1n32x5 FILLER_204_1413 ();
 b15zdnd11an1n08x5 FILLER_204_1445 ();
 b15zdnd11an1n32x5 FILLER_204_1466 ();
 b15zdnd11an1n16x5 FILLER_204_1498 ();
 b15zdnd11an1n64x5 FILLER_204_1522 ();
 b15zdnd11an1n64x5 FILLER_204_1586 ();
 b15zdnd11an1n64x5 FILLER_204_1650 ();
 b15zdnd11an1n64x5 FILLER_204_1714 ();
 b15zdnd11an1n64x5 FILLER_204_1778 ();
 b15zdnd11an1n64x5 FILLER_204_1842 ();
 b15zdnd11an1n64x5 FILLER_204_1906 ();
 b15zdnd11an1n32x5 FILLER_204_1970 ();
 b15zdnd00an1n02x5 FILLER_204_2002 ();
 b15zdnd00an1n01x5 FILLER_204_2004 ();
 b15zdnd11an1n64x5 FILLER_204_2011 ();
 b15zdnd11an1n32x5 FILLER_204_2075 ();
 b15zdnd11an1n16x5 FILLER_204_2138 ();
 b15zdnd11an1n64x5 FILLER_204_2162 ();
 b15zdnd11an1n32x5 FILLER_204_2226 ();
 b15zdnd11an1n16x5 FILLER_204_2258 ();
 b15zdnd00an1n02x5 FILLER_204_2274 ();
 b15zdnd11an1n64x5 FILLER_205_0 ();
 b15zdnd11an1n64x5 FILLER_205_64 ();
 b15zdnd11an1n64x5 FILLER_205_128 ();
 b15zdnd11an1n64x5 FILLER_205_192 ();
 b15zdnd11an1n64x5 FILLER_205_256 ();
 b15zdnd11an1n16x5 FILLER_205_320 ();
 b15zdnd11an1n08x5 FILLER_205_336 ();
 b15zdnd11an1n04x5 FILLER_205_357 ();
 b15zdnd00an1n02x5 FILLER_205_361 ();
 b15zdnd00an1n01x5 FILLER_205_363 ();
 b15zdnd11an1n32x5 FILLER_205_369 ();
 b15zdnd11an1n08x5 FILLER_205_401 ();
 b15zdnd11an1n04x5 FILLER_205_409 ();
 b15zdnd00an1n02x5 FILLER_205_413 ();
 b15zdnd00an1n01x5 FILLER_205_415 ();
 b15zdnd11an1n04x5 FILLER_205_458 ();
 b15zdnd11an1n16x5 FILLER_205_465 ();
 b15zdnd11an1n32x5 FILLER_205_523 ();
 b15zdnd11an1n16x5 FILLER_205_555 ();
 b15zdnd11an1n08x5 FILLER_205_571 ();
 b15zdnd11an1n04x5 FILLER_205_579 ();
 b15zdnd00an1n02x5 FILLER_205_583 ();
 b15zdnd00an1n01x5 FILLER_205_585 ();
 b15zdnd11an1n64x5 FILLER_205_628 ();
 b15zdnd11an1n64x5 FILLER_205_692 ();
 b15zdnd11an1n64x5 FILLER_205_756 ();
 b15zdnd11an1n64x5 FILLER_205_820 ();
 b15zdnd11an1n16x5 FILLER_205_884 ();
 b15zdnd11an1n08x5 FILLER_205_900 ();
 b15zdnd11an1n04x5 FILLER_205_908 ();
 b15zdnd00an1n02x5 FILLER_205_912 ();
 b15zdnd00an1n01x5 FILLER_205_914 ();
 b15zdnd11an1n64x5 FILLER_205_924 ();
 b15zdnd11an1n64x5 FILLER_205_988 ();
 b15zdnd11an1n64x5 FILLER_205_1052 ();
 b15zdnd11an1n64x5 FILLER_205_1116 ();
 b15zdnd11an1n64x5 FILLER_205_1180 ();
 b15zdnd11an1n64x5 FILLER_205_1244 ();
 b15zdnd11an1n64x5 FILLER_205_1308 ();
 b15zdnd11an1n64x5 FILLER_205_1372 ();
 b15zdnd11an1n64x5 FILLER_205_1436 ();
 b15zdnd11an1n64x5 FILLER_205_1500 ();
 b15zdnd11an1n32x5 FILLER_205_1564 ();
 b15zdnd11an1n16x5 FILLER_205_1596 ();
 b15zdnd11an1n64x5 FILLER_205_1621 ();
 b15zdnd11an1n64x5 FILLER_205_1685 ();
 b15zdnd11an1n64x5 FILLER_205_1749 ();
 b15zdnd11an1n64x5 FILLER_205_1813 ();
 b15zdnd11an1n64x5 FILLER_205_1877 ();
 b15zdnd11an1n64x5 FILLER_205_1941 ();
 b15zdnd11an1n04x5 FILLER_205_2005 ();
 b15zdnd00an1n01x5 FILLER_205_2009 ();
 b15zdnd11an1n04x5 FILLER_205_2013 ();
 b15zdnd11an1n64x5 FILLER_205_2020 ();
 b15zdnd11an1n64x5 FILLER_205_2084 ();
 b15zdnd11an1n16x5 FILLER_205_2148 ();
 b15zdnd00an1n01x5 FILLER_205_2164 ();
 b15zdnd11an1n64x5 FILLER_205_2210 ();
 b15zdnd11an1n08x5 FILLER_205_2274 ();
 b15zdnd00an1n02x5 FILLER_205_2282 ();
 b15zdnd11an1n64x5 FILLER_206_8 ();
 b15zdnd11an1n64x5 FILLER_206_72 ();
 b15zdnd11an1n64x5 FILLER_206_136 ();
 b15zdnd11an1n64x5 FILLER_206_200 ();
 b15zdnd11an1n64x5 FILLER_206_264 ();
 b15zdnd11an1n32x5 FILLER_206_328 ();
 b15zdnd11an1n64x5 FILLER_206_363 ();
 b15zdnd11an1n64x5 FILLER_206_427 ();
 b15zdnd11an1n64x5 FILLER_206_491 ();
 b15zdnd11an1n64x5 FILLER_206_555 ();
 b15zdnd11an1n64x5 FILLER_206_619 ();
 b15zdnd11an1n32x5 FILLER_206_683 ();
 b15zdnd00an1n02x5 FILLER_206_715 ();
 b15zdnd00an1n01x5 FILLER_206_717 ();
 b15zdnd11an1n64x5 FILLER_206_726 ();
 b15zdnd11an1n64x5 FILLER_206_790 ();
 b15zdnd11an1n64x5 FILLER_206_854 ();
 b15zdnd11an1n16x5 FILLER_206_918 ();
 b15zdnd11an1n64x5 FILLER_206_957 ();
 b15zdnd11an1n64x5 FILLER_206_1021 ();
 b15zdnd11an1n64x5 FILLER_206_1085 ();
 b15zdnd11an1n64x5 FILLER_206_1149 ();
 b15zdnd11an1n64x5 FILLER_206_1213 ();
 b15zdnd11an1n64x5 FILLER_206_1277 ();
 b15zdnd11an1n16x5 FILLER_206_1341 ();
 b15zdnd00an1n02x5 FILLER_206_1357 ();
 b15zdnd00an1n01x5 FILLER_206_1359 ();
 b15zdnd11an1n64x5 FILLER_206_1371 ();
 b15zdnd11an1n64x5 FILLER_206_1435 ();
 b15zdnd11an1n08x5 FILLER_206_1499 ();
 b15zdnd11an1n04x5 FILLER_206_1507 ();
 b15zdnd00an1n01x5 FILLER_206_1511 ();
 b15zdnd11an1n32x5 FILLER_206_1519 ();
 b15zdnd11an1n04x5 FILLER_206_1551 ();
 b15zdnd00an1n02x5 FILLER_206_1555 ();
 b15zdnd00an1n01x5 FILLER_206_1557 ();
 b15zdnd11an1n64x5 FILLER_206_1575 ();
 b15zdnd11an1n64x5 FILLER_206_1639 ();
 b15zdnd11an1n64x5 FILLER_206_1703 ();
 b15zdnd11an1n64x5 FILLER_206_1767 ();
 b15zdnd11an1n64x5 FILLER_206_1831 ();
 b15zdnd11an1n64x5 FILLER_206_1895 ();
 b15zdnd11an1n32x5 FILLER_206_1959 ();
 b15zdnd11an1n08x5 FILLER_206_1991 ();
 b15zdnd11an1n04x5 FILLER_206_1999 ();
 b15zdnd00an1n02x5 FILLER_206_2003 ();
 b15zdnd00an1n01x5 FILLER_206_2005 ();
 b15zdnd11an1n64x5 FILLER_206_2048 ();
 b15zdnd00an1n02x5 FILLER_206_2112 ();
 b15zdnd11an1n32x5 FILLER_206_2119 ();
 b15zdnd00an1n02x5 FILLER_206_2151 ();
 b15zdnd00an1n01x5 FILLER_206_2153 ();
 b15zdnd11an1n64x5 FILLER_206_2162 ();
 b15zdnd11an1n32x5 FILLER_206_2226 ();
 b15zdnd11an1n16x5 FILLER_206_2258 ();
 b15zdnd00an1n02x5 FILLER_206_2274 ();
 b15zdnd11an1n64x5 FILLER_207_0 ();
 b15zdnd11an1n64x5 FILLER_207_64 ();
 b15zdnd11an1n64x5 FILLER_207_128 ();
 b15zdnd11an1n64x5 FILLER_207_192 ();
 b15zdnd11an1n64x5 FILLER_207_256 ();
 b15zdnd11an1n32x5 FILLER_207_320 ();
 b15zdnd11an1n04x5 FILLER_207_352 ();
 b15zdnd00an1n02x5 FILLER_207_356 ();
 b15zdnd00an1n01x5 FILLER_207_358 ();
 b15zdnd11an1n64x5 FILLER_207_401 ();
 b15zdnd11an1n64x5 FILLER_207_465 ();
 b15zdnd11an1n64x5 FILLER_207_529 ();
 b15zdnd11an1n64x5 FILLER_207_593 ();
 b15zdnd11an1n64x5 FILLER_207_657 ();
 b15zdnd11an1n64x5 FILLER_207_721 ();
 b15zdnd11an1n64x5 FILLER_207_785 ();
 b15zdnd11an1n64x5 FILLER_207_849 ();
 b15zdnd11an1n32x5 FILLER_207_913 ();
 b15zdnd11an1n16x5 FILLER_207_945 ();
 b15zdnd00an1n02x5 FILLER_207_961 ();
 b15zdnd00an1n01x5 FILLER_207_963 ();
 b15zdnd11an1n32x5 FILLER_207_972 ();
 b15zdnd11an1n04x5 FILLER_207_1004 ();
 b15zdnd00an1n01x5 FILLER_207_1008 ();
 b15zdnd11an1n64x5 FILLER_207_1013 ();
 b15zdnd11an1n64x5 FILLER_207_1077 ();
 b15zdnd11an1n64x5 FILLER_207_1141 ();
 b15zdnd11an1n64x5 FILLER_207_1205 ();
 b15zdnd11an1n16x5 FILLER_207_1277 ();
 b15zdnd11an1n08x5 FILLER_207_1293 ();
 b15zdnd00an1n02x5 FILLER_207_1301 ();
 b15zdnd00an1n01x5 FILLER_207_1303 ();
 b15zdnd11an1n16x5 FILLER_207_1321 ();
 b15zdnd11an1n08x5 FILLER_207_1337 ();
 b15zdnd00an1n01x5 FILLER_207_1345 ();
 b15zdnd11an1n08x5 FILLER_207_1370 ();
 b15zdnd00an1n02x5 FILLER_207_1378 ();
 b15zdnd11an1n64x5 FILLER_207_1402 ();
 b15zdnd11an1n64x5 FILLER_207_1466 ();
 b15zdnd11an1n64x5 FILLER_207_1530 ();
 b15zdnd11an1n64x5 FILLER_207_1594 ();
 b15zdnd11an1n64x5 FILLER_207_1658 ();
 b15zdnd11an1n64x5 FILLER_207_1722 ();
 b15zdnd11an1n64x5 FILLER_207_1786 ();
 b15zdnd11an1n64x5 FILLER_207_1850 ();
 b15zdnd11an1n64x5 FILLER_207_1914 ();
 b15zdnd11an1n04x5 FILLER_207_1978 ();
 b15zdnd00an1n02x5 FILLER_207_1982 ();
 b15zdnd00an1n01x5 FILLER_207_1984 ();
 b15zdnd11an1n64x5 FILLER_207_2037 ();
 b15zdnd11an1n16x5 FILLER_207_2101 ();
 b15zdnd11an1n08x5 FILLER_207_2159 ();
 b15zdnd00an1n01x5 FILLER_207_2167 ();
 b15zdnd11an1n64x5 FILLER_207_2186 ();
 b15zdnd11an1n08x5 FILLER_207_2250 ();
 b15zdnd11an1n04x5 FILLER_207_2264 ();
 b15zdnd11an1n08x5 FILLER_207_2272 ();
 b15zdnd11an1n04x5 FILLER_207_2280 ();
 b15zdnd11an1n64x5 FILLER_208_8 ();
 b15zdnd11an1n64x5 FILLER_208_72 ();
 b15zdnd11an1n64x5 FILLER_208_136 ();
 b15zdnd11an1n64x5 FILLER_208_200 ();
 b15zdnd11an1n64x5 FILLER_208_264 ();
 b15zdnd11an1n32x5 FILLER_208_328 ();
 b15zdnd11an1n04x5 FILLER_208_360 ();
 b15zdnd00an1n02x5 FILLER_208_364 ();
 b15zdnd11an1n64x5 FILLER_208_372 ();
 b15zdnd11an1n64x5 FILLER_208_436 ();
 b15zdnd11an1n64x5 FILLER_208_500 ();
 b15zdnd11an1n64x5 FILLER_208_564 ();
 b15zdnd11an1n08x5 FILLER_208_628 ();
 b15zdnd00an1n02x5 FILLER_208_636 ();
 b15zdnd00an1n01x5 FILLER_208_638 ();
 b15zdnd11an1n64x5 FILLER_208_648 ();
 b15zdnd11an1n04x5 FILLER_208_712 ();
 b15zdnd00an1n02x5 FILLER_208_716 ();
 b15zdnd11an1n64x5 FILLER_208_726 ();
 b15zdnd11an1n64x5 FILLER_208_790 ();
 b15zdnd11an1n64x5 FILLER_208_854 ();
 b15zdnd11an1n64x5 FILLER_208_918 ();
 b15zdnd11an1n04x5 FILLER_208_982 ();
 b15zdnd00an1n02x5 FILLER_208_986 ();
 b15zdnd11an1n64x5 FILLER_208_996 ();
 b15zdnd11an1n64x5 FILLER_208_1060 ();
 b15zdnd11an1n64x5 FILLER_208_1124 ();
 b15zdnd11an1n64x5 FILLER_208_1188 ();
 b15zdnd11an1n32x5 FILLER_208_1252 ();
 b15zdnd11an1n16x5 FILLER_208_1284 ();
 b15zdnd11an1n64x5 FILLER_208_1310 ();
 b15zdnd11an1n64x5 FILLER_208_1374 ();
 b15zdnd11an1n08x5 FILLER_208_1438 ();
 b15zdnd11an1n04x5 FILLER_208_1446 ();
 b15zdnd11an1n64x5 FILLER_208_1459 ();
 b15zdnd11an1n64x5 FILLER_208_1523 ();
 b15zdnd11an1n64x5 FILLER_208_1587 ();
 b15zdnd11an1n64x5 FILLER_208_1651 ();
 b15zdnd11an1n32x5 FILLER_208_1715 ();
 b15zdnd11an1n16x5 FILLER_208_1747 ();
 b15zdnd11an1n04x5 FILLER_208_1763 ();
 b15zdnd00an1n01x5 FILLER_208_1767 ();
 b15zdnd11an1n64x5 FILLER_208_1783 ();
 b15zdnd11an1n64x5 FILLER_208_1847 ();
 b15zdnd11an1n64x5 FILLER_208_1911 ();
 b15zdnd11an1n32x5 FILLER_208_1975 ();
 b15zdnd00an1n02x5 FILLER_208_2007 ();
 b15zdnd00an1n01x5 FILLER_208_2009 ();
 b15zdnd11an1n32x5 FILLER_208_2013 ();
 b15zdnd11an1n08x5 FILLER_208_2045 ();
 b15zdnd11an1n04x5 FILLER_208_2095 ();
 b15zdnd11an1n08x5 FILLER_208_2141 ();
 b15zdnd11an1n04x5 FILLER_208_2149 ();
 b15zdnd00an1n01x5 FILLER_208_2153 ();
 b15zdnd11an1n64x5 FILLER_208_2162 ();
 b15zdnd11an1n04x5 FILLER_208_2226 ();
 b15zdnd00an1n02x5 FILLER_208_2230 ();
 b15zdnd00an1n02x5 FILLER_208_2274 ();
 b15zdnd11an1n16x5 FILLER_209_0 ();
 b15zdnd11an1n08x5 FILLER_209_16 ();
 b15zdnd00an1n02x5 FILLER_209_24 ();
 b15zdnd00an1n01x5 FILLER_209_26 ();
 b15zdnd11an1n04x5 FILLER_209_35 ();
 b15zdnd00an1n02x5 FILLER_209_39 ();
 b15zdnd00an1n01x5 FILLER_209_41 ();
 b15zdnd11an1n64x5 FILLER_209_62 ();
 b15zdnd11an1n64x5 FILLER_209_126 ();
 b15zdnd11an1n64x5 FILLER_209_190 ();
 b15zdnd11an1n64x5 FILLER_209_254 ();
 b15zdnd11an1n64x5 FILLER_209_318 ();
 b15zdnd11an1n64x5 FILLER_209_382 ();
 b15zdnd11an1n64x5 FILLER_209_446 ();
 b15zdnd11an1n64x5 FILLER_209_510 ();
 b15zdnd11an1n64x5 FILLER_209_574 ();
 b15zdnd11an1n64x5 FILLER_209_638 ();
 b15zdnd11an1n64x5 FILLER_209_702 ();
 b15zdnd11an1n16x5 FILLER_209_766 ();
 b15zdnd00an1n02x5 FILLER_209_782 ();
 b15zdnd00an1n01x5 FILLER_209_784 ();
 b15zdnd11an1n64x5 FILLER_209_789 ();
 b15zdnd11an1n64x5 FILLER_209_853 ();
 b15zdnd11an1n64x5 FILLER_209_917 ();
 b15zdnd11an1n32x5 FILLER_209_981 ();
 b15zdnd11an1n08x5 FILLER_209_1013 ();
 b15zdnd00an1n01x5 FILLER_209_1021 ();
 b15zdnd11an1n32x5 FILLER_209_1028 ();
 b15zdnd11an1n16x5 FILLER_209_1060 ();
 b15zdnd11an1n08x5 FILLER_209_1076 ();
 b15zdnd00an1n02x5 FILLER_209_1084 ();
 b15zdnd11an1n64x5 FILLER_209_1099 ();
 b15zdnd11an1n32x5 FILLER_209_1163 ();
 b15zdnd11an1n04x5 FILLER_209_1195 ();
 b15zdnd00an1n01x5 FILLER_209_1199 ();
 b15zdnd11an1n04x5 FILLER_209_1211 ();
 b15zdnd11an1n16x5 FILLER_209_1235 ();
 b15zdnd00an1n02x5 FILLER_209_1251 ();
 b15zdnd11an1n64x5 FILLER_209_1270 ();
 b15zdnd11an1n64x5 FILLER_209_1334 ();
 b15zdnd11an1n64x5 FILLER_209_1398 ();
 b15zdnd11an1n08x5 FILLER_209_1462 ();
 b15zdnd00an1n01x5 FILLER_209_1470 ();
 b15zdnd11an1n64x5 FILLER_209_1477 ();
 b15zdnd11an1n64x5 FILLER_209_1541 ();
 b15zdnd11an1n16x5 FILLER_209_1605 ();
 b15zdnd11an1n08x5 FILLER_209_1621 ();
 b15zdnd00an1n02x5 FILLER_209_1629 ();
 b15zdnd11an1n64x5 FILLER_209_1673 ();
 b15zdnd11an1n32x5 FILLER_209_1737 ();
 b15zdnd11an1n08x5 FILLER_209_1769 ();
 b15zdnd11an1n32x5 FILLER_209_1794 ();
 b15zdnd11an1n64x5 FILLER_209_1857 ();
 b15zdnd11an1n64x5 FILLER_209_1921 ();
 b15zdnd11an1n64x5 FILLER_209_1985 ();
 b15zdnd11an1n32x5 FILLER_209_2049 ();
 b15zdnd11an1n16x5 FILLER_209_2081 ();
 b15zdnd11an1n04x5 FILLER_209_2097 ();
 b15zdnd00an1n01x5 FILLER_209_2101 ();
 b15zdnd11an1n32x5 FILLER_209_2121 ();
 b15zdnd11an1n32x5 FILLER_209_2195 ();
 b15zdnd11an1n08x5 FILLER_209_2227 ();
 b15zdnd11an1n04x5 FILLER_209_2235 ();
 b15zdnd00an1n01x5 FILLER_209_2239 ();
 b15zdnd00an1n02x5 FILLER_209_2282 ();
 b15zdnd11an1n64x5 FILLER_210_8 ();
 b15zdnd11an1n64x5 FILLER_210_72 ();
 b15zdnd11an1n64x5 FILLER_210_136 ();
 b15zdnd11an1n64x5 FILLER_210_200 ();
 b15zdnd11an1n64x5 FILLER_210_264 ();
 b15zdnd11an1n64x5 FILLER_210_328 ();
 b15zdnd11an1n64x5 FILLER_210_392 ();
 b15zdnd11an1n16x5 FILLER_210_456 ();
 b15zdnd11an1n64x5 FILLER_210_514 ();
 b15zdnd11an1n64x5 FILLER_210_578 ();
 b15zdnd11an1n64x5 FILLER_210_642 ();
 b15zdnd11an1n08x5 FILLER_210_706 ();
 b15zdnd11an1n04x5 FILLER_210_714 ();
 b15zdnd11an1n64x5 FILLER_210_726 ();
 b15zdnd11an1n64x5 FILLER_210_790 ();
 b15zdnd11an1n32x5 FILLER_210_854 ();
 b15zdnd11an1n16x5 FILLER_210_886 ();
 b15zdnd00an1n01x5 FILLER_210_902 ();
 b15zdnd11an1n64x5 FILLER_210_907 ();
 b15zdnd11an1n32x5 FILLER_210_971 ();
 b15zdnd11an1n16x5 FILLER_210_1003 ();
 b15zdnd11an1n08x5 FILLER_210_1019 ();
 b15zdnd11an1n04x5 FILLER_210_1027 ();
 b15zdnd00an1n02x5 FILLER_210_1031 ();
 b15zdnd00an1n01x5 FILLER_210_1033 ();
 b15zdnd11an1n32x5 FILLER_210_1038 ();
 b15zdnd11an1n16x5 FILLER_210_1070 ();
 b15zdnd00an1n01x5 FILLER_210_1086 ();
 b15zdnd11an1n64x5 FILLER_210_1094 ();
 b15zdnd11an1n32x5 FILLER_210_1158 ();
 b15zdnd11an1n16x5 FILLER_210_1190 ();
 b15zdnd11an1n08x5 FILLER_210_1206 ();
 b15zdnd11an1n64x5 FILLER_210_1225 ();
 b15zdnd11an1n04x5 FILLER_210_1289 ();
 b15zdnd11an1n32x5 FILLER_210_1304 ();
 b15zdnd11an1n16x5 FILLER_210_1336 ();
 b15zdnd11an1n08x5 FILLER_210_1352 ();
 b15zdnd11an1n04x5 FILLER_210_1360 ();
 b15zdnd00an1n01x5 FILLER_210_1364 ();
 b15zdnd11an1n16x5 FILLER_210_1373 ();
 b15zdnd11an1n08x5 FILLER_210_1389 ();
 b15zdnd00an1n02x5 FILLER_210_1397 ();
 b15zdnd00an1n01x5 FILLER_210_1399 ();
 b15zdnd11an1n64x5 FILLER_210_1425 ();
 b15zdnd00an1n02x5 FILLER_210_1489 ();
 b15zdnd00an1n01x5 FILLER_210_1491 ();
 b15zdnd11an1n64x5 FILLER_210_1509 ();
 b15zdnd11an1n64x5 FILLER_210_1573 ();
 b15zdnd11an1n64x5 FILLER_210_1637 ();
 b15zdnd11an1n08x5 FILLER_210_1701 ();
 b15zdnd11an1n04x5 FILLER_210_1709 ();
 b15zdnd00an1n01x5 FILLER_210_1713 ();
 b15zdnd11an1n64x5 FILLER_210_1718 ();
 b15zdnd11an1n08x5 FILLER_210_1782 ();
 b15zdnd11an1n04x5 FILLER_210_1810 ();
 b15zdnd11an1n64x5 FILLER_210_1829 ();
 b15zdnd11an1n16x5 FILLER_210_1893 ();
 b15zdnd00an1n02x5 FILLER_210_1909 ();
 b15zdnd00an1n01x5 FILLER_210_1911 ();
 b15zdnd11an1n64x5 FILLER_210_1924 ();
 b15zdnd11an1n64x5 FILLER_210_1988 ();
 b15zdnd11an1n16x5 FILLER_210_2052 ();
 b15zdnd11an1n08x5 FILLER_210_2068 ();
 b15zdnd11an1n04x5 FILLER_210_2076 ();
 b15zdnd00an1n02x5 FILLER_210_2080 ();
 b15zdnd00an1n01x5 FILLER_210_2082 ();
 b15zdnd11an1n08x5 FILLER_210_2125 ();
 b15zdnd00an1n01x5 FILLER_210_2133 ();
 b15zdnd11an1n08x5 FILLER_210_2141 ();
 b15zdnd11an1n04x5 FILLER_210_2149 ();
 b15zdnd00an1n01x5 FILLER_210_2153 ();
 b15zdnd11an1n64x5 FILLER_210_2162 ();
 b15zdnd11an1n16x5 FILLER_210_2226 ();
 b15zdnd00an1n02x5 FILLER_210_2242 ();
 b15zdnd11an1n04x5 FILLER_210_2248 ();
 b15zdnd11an1n16x5 FILLER_210_2256 ();
 b15zdnd11an1n04x5 FILLER_210_2272 ();
 b15zdnd11an1n64x5 FILLER_211_0 ();
 b15zdnd11an1n64x5 FILLER_211_64 ();
 b15zdnd11an1n64x5 FILLER_211_128 ();
 b15zdnd11an1n16x5 FILLER_211_192 ();
 b15zdnd11an1n08x5 FILLER_211_208 ();
 b15zdnd11an1n64x5 FILLER_211_219 ();
 b15zdnd11an1n64x5 FILLER_211_283 ();
 b15zdnd11an1n04x5 FILLER_211_347 ();
 b15zdnd00an1n02x5 FILLER_211_351 ();
 b15zdnd00an1n01x5 FILLER_211_353 ();
 b15zdnd11an1n64x5 FILLER_211_359 ();
 b15zdnd11an1n32x5 FILLER_211_423 ();
 b15zdnd11an1n08x5 FILLER_211_455 ();
 b15zdnd11an1n04x5 FILLER_211_463 ();
 b15zdnd00an1n02x5 FILLER_211_467 ();
 b15zdnd00an1n01x5 FILLER_211_469 ();
 b15zdnd11an1n64x5 FILLER_211_473 ();
 b15zdnd11an1n64x5 FILLER_211_537 ();
 b15zdnd11an1n16x5 FILLER_211_601 ();
 b15zdnd11an1n08x5 FILLER_211_617 ();
 b15zdnd00an1n02x5 FILLER_211_625 ();
 b15zdnd11an1n64x5 FILLER_211_636 ();
 b15zdnd11an1n64x5 FILLER_211_700 ();
 b15zdnd11an1n16x5 FILLER_211_764 ();
 b15zdnd11an1n64x5 FILLER_211_784 ();
 b15zdnd11an1n64x5 FILLER_211_848 ();
 b15zdnd11an1n64x5 FILLER_211_912 ();
 b15zdnd11an1n64x5 FILLER_211_976 ();
 b15zdnd11an1n16x5 FILLER_211_1040 ();
 b15zdnd00an1n02x5 FILLER_211_1056 ();
 b15zdnd00an1n01x5 FILLER_211_1058 ();
 b15zdnd11an1n64x5 FILLER_211_1063 ();
 b15zdnd11an1n32x5 FILLER_211_1127 ();
 b15zdnd11an1n16x5 FILLER_211_1159 ();
 b15zdnd11an1n08x5 FILLER_211_1175 ();
 b15zdnd00an1n01x5 FILLER_211_1183 ();
 b15zdnd11an1n64x5 FILLER_211_1195 ();
 b15zdnd11an1n64x5 FILLER_211_1259 ();
 b15zdnd11an1n64x5 FILLER_211_1323 ();
 b15zdnd11an1n64x5 FILLER_211_1387 ();
 b15zdnd11an1n64x5 FILLER_211_1451 ();
 b15zdnd11an1n64x5 FILLER_211_1515 ();
 b15zdnd11an1n64x5 FILLER_211_1579 ();
 b15zdnd11an1n64x5 FILLER_211_1643 ();
 b15zdnd11an1n64x5 FILLER_211_1707 ();
 b15zdnd11an1n64x5 FILLER_211_1771 ();
 b15zdnd11an1n64x5 FILLER_211_1835 ();
 b15zdnd11an1n16x5 FILLER_211_1899 ();
 b15zdnd11an1n04x5 FILLER_211_1915 ();
 b15zdnd00an1n02x5 FILLER_211_1919 ();
 b15zdnd00an1n01x5 FILLER_211_1921 ();
 b15zdnd11an1n16x5 FILLER_211_1974 ();
 b15zdnd11an1n08x5 FILLER_211_1990 ();
 b15zdnd11an1n64x5 FILLER_211_2012 ();
 b15zdnd11an1n32x5 FILLER_211_2076 ();
 b15zdnd11an1n08x5 FILLER_211_2108 ();
 b15zdnd11an1n04x5 FILLER_211_2116 ();
 b15zdnd11an1n08x5 FILLER_211_2162 ();
 b15zdnd11an1n04x5 FILLER_211_2170 ();
 b15zdnd00an1n02x5 FILLER_211_2174 ();
 b15zdnd11an1n64x5 FILLER_211_2194 ();
 b15zdnd11an1n16x5 FILLER_211_2258 ();
 b15zdnd11an1n08x5 FILLER_211_2274 ();
 b15zdnd00an1n02x5 FILLER_211_2282 ();
 b15zdnd11an1n64x5 FILLER_212_8 ();
 b15zdnd11an1n64x5 FILLER_212_72 ();
 b15zdnd11an1n64x5 FILLER_212_136 ();
 b15zdnd11an1n64x5 FILLER_212_200 ();
 b15zdnd11an1n64x5 FILLER_212_264 ();
 b15zdnd11an1n64x5 FILLER_212_328 ();
 b15zdnd11an1n32x5 FILLER_212_392 ();
 b15zdnd11an1n08x5 FILLER_212_424 ();
 b15zdnd00an1n01x5 FILLER_212_432 ();
 b15zdnd11an1n64x5 FILLER_212_473 ();
 b15zdnd11an1n64x5 FILLER_212_537 ();
 b15zdnd11an1n64x5 FILLER_212_601 ();
 b15zdnd11an1n32x5 FILLER_212_665 ();
 b15zdnd11an1n16x5 FILLER_212_697 ();
 b15zdnd11an1n04x5 FILLER_212_713 ();
 b15zdnd00an1n01x5 FILLER_212_717 ();
 b15zdnd00an1n02x5 FILLER_212_726 ();
 b15zdnd11an1n16x5 FILLER_212_734 ();
 b15zdnd11an1n04x5 FILLER_212_750 ();
 b15zdnd11an1n16x5 FILLER_212_761 ();
 b15zdnd11an1n08x5 FILLER_212_777 ();
 b15zdnd00an1n02x5 FILLER_212_785 ();
 b15zdnd11an1n16x5 FILLER_212_797 ();
 b15zdnd00an1n02x5 FILLER_212_813 ();
 b15zdnd00an1n01x5 FILLER_212_815 ();
 b15zdnd11an1n64x5 FILLER_212_825 ();
 b15zdnd11an1n64x5 FILLER_212_889 ();
 b15zdnd11an1n64x5 FILLER_212_953 ();
 b15zdnd11an1n32x5 FILLER_212_1017 ();
 b15zdnd11an1n08x5 FILLER_212_1049 ();
 b15zdnd11an1n04x5 FILLER_212_1057 ();
 b15zdnd00an1n02x5 FILLER_212_1061 ();
 b15zdnd11an1n64x5 FILLER_212_1067 ();
 b15zdnd11an1n64x5 FILLER_212_1131 ();
 b15zdnd11an1n64x5 FILLER_212_1195 ();
 b15zdnd11an1n64x5 FILLER_212_1259 ();
 b15zdnd11an1n32x5 FILLER_212_1323 ();
 b15zdnd00an1n01x5 FILLER_212_1355 ();
 b15zdnd11an1n32x5 FILLER_212_1370 ();
 b15zdnd11an1n16x5 FILLER_212_1402 ();
 b15zdnd11an1n08x5 FILLER_212_1418 ();
 b15zdnd11an1n04x5 FILLER_212_1426 ();
 b15zdnd00an1n01x5 FILLER_212_1430 ();
 b15zdnd11an1n64x5 FILLER_212_1440 ();
 b15zdnd11an1n64x5 FILLER_212_1504 ();
 b15zdnd11an1n64x5 FILLER_212_1568 ();
 b15zdnd11an1n16x5 FILLER_212_1632 ();
 b15zdnd11an1n04x5 FILLER_212_1648 ();
 b15zdnd00an1n01x5 FILLER_212_1652 ();
 b15zdnd11an1n64x5 FILLER_212_1705 ();
 b15zdnd11an1n64x5 FILLER_212_1769 ();
 b15zdnd11an1n64x5 FILLER_212_1833 ();
 b15zdnd11an1n32x5 FILLER_212_1897 ();
 b15zdnd11an1n08x5 FILLER_212_1929 ();
 b15zdnd00an1n02x5 FILLER_212_1937 ();
 b15zdnd00an1n01x5 FILLER_212_1939 ();
 b15zdnd11an1n04x5 FILLER_212_1943 ();
 b15zdnd11an1n16x5 FILLER_212_1950 ();
 b15zdnd11an1n08x5 FILLER_212_1966 ();
 b15zdnd00an1n02x5 FILLER_212_1974 ();
 b15zdnd11an1n32x5 FILLER_212_2018 ();
 b15zdnd00an1n02x5 FILLER_212_2050 ();
 b15zdnd00an1n01x5 FILLER_212_2052 ();
 b15zdnd11an1n64x5 FILLER_212_2067 ();
 b15zdnd11an1n16x5 FILLER_212_2131 ();
 b15zdnd11an1n04x5 FILLER_212_2147 ();
 b15zdnd00an1n02x5 FILLER_212_2151 ();
 b15zdnd00an1n01x5 FILLER_212_2153 ();
 b15zdnd11an1n64x5 FILLER_212_2162 ();
 b15zdnd11an1n16x5 FILLER_212_2226 ();
 b15zdnd11an1n08x5 FILLER_212_2242 ();
 b15zdnd11an1n04x5 FILLER_212_2250 ();
 b15zdnd11an1n16x5 FILLER_212_2259 ();
 b15zdnd00an1n01x5 FILLER_212_2275 ();
 b15zdnd11an1n64x5 FILLER_213_0 ();
 b15zdnd11an1n64x5 FILLER_213_64 ();
 b15zdnd11an1n64x5 FILLER_213_128 ();
 b15zdnd11an1n64x5 FILLER_213_192 ();
 b15zdnd11an1n64x5 FILLER_213_256 ();
 b15zdnd11an1n64x5 FILLER_213_320 ();
 b15zdnd11an1n64x5 FILLER_213_384 ();
 b15zdnd11an1n16x5 FILLER_213_448 ();
 b15zdnd00an1n01x5 FILLER_213_464 ();
 b15zdnd11an1n64x5 FILLER_213_468 ();
 b15zdnd11an1n64x5 FILLER_213_532 ();
 b15zdnd11an1n64x5 FILLER_213_596 ();
 b15zdnd11an1n64x5 FILLER_213_660 ();
 b15zdnd11an1n64x5 FILLER_213_724 ();
 b15zdnd11an1n16x5 FILLER_213_788 ();
 b15zdnd11an1n08x5 FILLER_213_804 ();
 b15zdnd11an1n04x5 FILLER_213_812 ();
 b15zdnd00an1n01x5 FILLER_213_816 ();
 b15zdnd11an1n04x5 FILLER_213_829 ();
 b15zdnd00an1n02x5 FILLER_213_833 ();
 b15zdnd00an1n01x5 FILLER_213_835 ();
 b15zdnd11an1n64x5 FILLER_213_850 ();
 b15zdnd11an1n64x5 FILLER_213_914 ();
 b15zdnd11an1n64x5 FILLER_213_978 ();
 b15zdnd11an1n64x5 FILLER_213_1042 ();
 b15zdnd11an1n64x5 FILLER_213_1106 ();
 b15zdnd11an1n64x5 FILLER_213_1170 ();
 b15zdnd11an1n64x5 FILLER_213_1234 ();
 b15zdnd11an1n64x5 FILLER_213_1298 ();
 b15zdnd11an1n64x5 FILLER_213_1362 ();
 b15zdnd11an1n16x5 FILLER_213_1426 ();
 b15zdnd11an1n04x5 FILLER_213_1442 ();
 b15zdnd00an1n01x5 FILLER_213_1446 ();
 b15zdnd11an1n64x5 FILLER_213_1462 ();
 b15zdnd11an1n64x5 FILLER_213_1526 ();
 b15zdnd11an1n64x5 FILLER_213_1590 ();
 b15zdnd11an1n64x5 FILLER_213_1654 ();
 b15zdnd11an1n64x5 FILLER_213_1718 ();
 b15zdnd11an1n64x5 FILLER_213_1782 ();
 b15zdnd11an1n64x5 FILLER_213_1846 ();
 b15zdnd11an1n32x5 FILLER_213_1910 ();
 b15zdnd11an1n04x5 FILLER_213_1942 ();
 b15zdnd00an1n02x5 FILLER_213_1946 ();
 b15zdnd11an1n64x5 FILLER_213_1951 ();
 b15zdnd11an1n32x5 FILLER_213_2015 ();
 b15zdnd00an1n02x5 FILLER_213_2047 ();
 b15zdnd11an1n04x5 FILLER_213_2060 ();
 b15zdnd00an1n02x5 FILLER_213_2064 ();
 b15zdnd11an1n64x5 FILLER_213_2073 ();
 b15zdnd11an1n64x5 FILLER_213_2137 ();
 b15zdnd11an1n32x5 FILLER_213_2201 ();
 b15zdnd11an1n04x5 FILLER_213_2233 ();
 b15zdnd00an1n01x5 FILLER_213_2237 ();
 b15zdnd11an1n16x5 FILLER_213_2258 ();
 b15zdnd11an1n08x5 FILLER_213_2274 ();
 b15zdnd00an1n02x5 FILLER_213_2282 ();
 b15zdnd11an1n64x5 FILLER_214_8 ();
 b15zdnd11an1n64x5 FILLER_214_72 ();
 b15zdnd11an1n64x5 FILLER_214_136 ();
 b15zdnd11an1n16x5 FILLER_214_200 ();
 b15zdnd00an1n02x5 FILLER_214_216 ();
 b15zdnd00an1n01x5 FILLER_214_218 ();
 b15zdnd11an1n64x5 FILLER_214_226 ();
 b15zdnd11an1n64x5 FILLER_214_290 ();
 b15zdnd11an1n64x5 FILLER_214_354 ();
 b15zdnd11an1n64x5 FILLER_214_418 ();
 b15zdnd11an1n64x5 FILLER_214_482 ();
 b15zdnd11an1n32x5 FILLER_214_546 ();
 b15zdnd11an1n16x5 FILLER_214_578 ();
 b15zdnd11an1n08x5 FILLER_214_594 ();
 b15zdnd11an1n08x5 FILLER_214_609 ();
 b15zdnd11an1n04x5 FILLER_214_617 ();
 b15zdnd00an1n02x5 FILLER_214_621 ();
 b15zdnd11an1n64x5 FILLER_214_626 ();
 b15zdnd11an1n16x5 FILLER_214_690 ();
 b15zdnd11an1n08x5 FILLER_214_706 ();
 b15zdnd11an1n04x5 FILLER_214_714 ();
 b15zdnd11an1n32x5 FILLER_214_726 ();
 b15zdnd11an1n16x5 FILLER_214_758 ();
 b15zdnd11an1n04x5 FILLER_214_774 ();
 b15zdnd11an1n64x5 FILLER_214_784 ();
 b15zdnd11an1n64x5 FILLER_214_848 ();
 b15zdnd11an1n32x5 FILLER_214_912 ();
 b15zdnd11an1n08x5 FILLER_214_944 ();
 b15zdnd11an1n04x5 FILLER_214_952 ();
 b15zdnd00an1n02x5 FILLER_214_956 ();
 b15zdnd00an1n01x5 FILLER_214_958 ();
 b15zdnd11an1n64x5 FILLER_214_990 ();
 b15zdnd11an1n32x5 FILLER_214_1054 ();
 b15zdnd11an1n16x5 FILLER_214_1086 ();
 b15zdnd11an1n04x5 FILLER_214_1102 ();
 b15zdnd00an1n01x5 FILLER_214_1106 ();
 b15zdnd11an1n32x5 FILLER_214_1121 ();
 b15zdnd11an1n16x5 FILLER_214_1153 ();
 b15zdnd11an1n04x5 FILLER_214_1169 ();
 b15zdnd11an1n16x5 FILLER_214_1180 ();
 b15zdnd11an1n08x5 FILLER_214_1196 ();
 b15zdnd11an1n04x5 FILLER_214_1204 ();
 b15zdnd00an1n02x5 FILLER_214_1208 ();
 b15zdnd11an1n64x5 FILLER_214_1241 ();
 b15zdnd11an1n64x5 FILLER_214_1305 ();
 b15zdnd11an1n32x5 FILLER_214_1369 ();
 b15zdnd11an1n16x5 FILLER_214_1401 ();
 b15zdnd11an1n04x5 FILLER_214_1417 ();
 b15zdnd11an1n08x5 FILLER_214_1433 ();
 b15zdnd11an1n04x5 FILLER_214_1441 ();
 b15zdnd00an1n01x5 FILLER_214_1445 ();
 b15zdnd11an1n64x5 FILLER_214_1458 ();
 b15zdnd11an1n08x5 FILLER_214_1522 ();
 b15zdnd00an1n02x5 FILLER_214_1530 ();
 b15zdnd00an1n01x5 FILLER_214_1532 ();
 b15zdnd11an1n64x5 FILLER_214_1541 ();
 b15zdnd11an1n16x5 FILLER_214_1605 ();
 b15zdnd11an1n08x5 FILLER_214_1621 ();
 b15zdnd11an1n04x5 FILLER_214_1629 ();
 b15zdnd11an1n04x5 FILLER_214_1685 ();
 b15zdnd11an1n64x5 FILLER_214_1692 ();
 b15zdnd11an1n64x5 FILLER_214_1756 ();
 b15zdnd11an1n64x5 FILLER_214_1820 ();
 b15zdnd11an1n64x5 FILLER_214_1884 ();
 b15zdnd11an1n64x5 FILLER_214_1948 ();
 b15zdnd11an1n64x5 FILLER_214_2012 ();
 b15zdnd11an1n64x5 FILLER_214_2076 ();
 b15zdnd11an1n08x5 FILLER_214_2140 ();
 b15zdnd11an1n04x5 FILLER_214_2148 ();
 b15zdnd00an1n02x5 FILLER_214_2152 ();
 b15zdnd11an1n32x5 FILLER_214_2162 ();
 b15zdnd11an1n08x5 FILLER_214_2194 ();
 b15zdnd00an1n01x5 FILLER_214_2202 ();
 b15zdnd11an1n08x5 FILLER_214_2227 ();
 b15zdnd11an1n04x5 FILLER_214_2235 ();
 b15zdnd00an1n02x5 FILLER_214_2239 ();
 b15zdnd11an1n16x5 FILLER_214_2255 ();
 b15zdnd11an1n04x5 FILLER_214_2271 ();
 b15zdnd00an1n01x5 FILLER_214_2275 ();
 b15zdnd11an1n64x5 FILLER_215_0 ();
 b15zdnd11an1n64x5 FILLER_215_64 ();
 b15zdnd11an1n64x5 FILLER_215_128 ();
 b15zdnd11an1n16x5 FILLER_215_192 ();
 b15zdnd11an1n04x5 FILLER_215_208 ();
 b15zdnd00an1n01x5 FILLER_215_212 ();
 b15zdnd11an1n04x5 FILLER_215_223 ();
 b15zdnd11an1n64x5 FILLER_215_231 ();
 b15zdnd11an1n64x5 FILLER_215_295 ();
 b15zdnd11an1n64x5 FILLER_215_359 ();
 b15zdnd11an1n16x5 FILLER_215_423 ();
 b15zdnd11an1n04x5 FILLER_215_439 ();
 b15zdnd00an1n01x5 FILLER_215_443 ();
 b15zdnd11an1n64x5 FILLER_215_496 ();
 b15zdnd11an1n32x5 FILLER_215_560 ();
 b15zdnd11an1n04x5 FILLER_215_592 ();
 b15zdnd11an1n64x5 FILLER_215_648 ();
 b15zdnd11an1n64x5 FILLER_215_712 ();
 b15zdnd11an1n32x5 FILLER_215_776 ();
 b15zdnd11an1n08x5 FILLER_215_808 ();
 b15zdnd11an1n04x5 FILLER_215_816 ();
 b15zdnd00an1n02x5 FILLER_215_820 ();
 b15zdnd11an1n04x5 FILLER_215_842 ();
 b15zdnd11an1n16x5 FILLER_215_860 ();
 b15zdnd11an1n08x5 FILLER_215_876 ();
 b15zdnd00an1n01x5 FILLER_215_884 ();
 b15zdnd11an1n08x5 FILLER_215_894 ();
 b15zdnd11an1n64x5 FILLER_215_909 ();
 b15zdnd11an1n08x5 FILLER_215_973 ();
 b15zdnd11an1n04x5 FILLER_215_981 ();
 b15zdnd00an1n02x5 FILLER_215_985 ();
 b15zdnd11an1n04x5 FILLER_215_990 ();
 b15zdnd11an1n32x5 FILLER_215_997 ();
 b15zdnd11an1n08x5 FILLER_215_1029 ();
 b15zdnd11an1n04x5 FILLER_215_1037 ();
 b15zdnd00an1n02x5 FILLER_215_1041 ();
 b15zdnd11an1n64x5 FILLER_215_1052 ();
 b15zdnd00an1n02x5 FILLER_215_1116 ();
 b15zdnd00an1n01x5 FILLER_215_1118 ();
 b15zdnd11an1n04x5 FILLER_215_1129 ();
 b15zdnd11an1n16x5 FILLER_215_1139 ();
 b15zdnd11an1n08x5 FILLER_215_1155 ();
 b15zdnd11an1n04x5 FILLER_215_1163 ();
 b15zdnd00an1n01x5 FILLER_215_1167 ();
 b15zdnd11an1n04x5 FILLER_215_1188 ();
 b15zdnd11an1n32x5 FILLER_215_1206 ();
 b15zdnd11an1n16x5 FILLER_215_1238 ();
 b15zdnd11an1n04x5 FILLER_215_1254 ();
 b15zdnd00an1n02x5 FILLER_215_1258 ();
 b15zdnd11an1n64x5 FILLER_215_1280 ();
 b15zdnd11an1n08x5 FILLER_215_1344 ();
 b15zdnd11an1n04x5 FILLER_215_1352 ();
 b15zdnd11an1n64x5 FILLER_215_1398 ();
 b15zdnd11an1n08x5 FILLER_215_1478 ();
 b15zdnd00an1n01x5 FILLER_215_1486 ();
 b15zdnd11an1n04x5 FILLER_215_1491 ();
 b15zdnd00an1n02x5 FILLER_215_1495 ();
 b15zdnd11an1n64x5 FILLER_215_1514 ();
 b15zdnd11an1n32x5 FILLER_215_1578 ();
 b15zdnd11an1n04x5 FILLER_215_1610 ();
 b15zdnd11an1n04x5 FILLER_215_1666 ();
 b15zdnd11an1n04x5 FILLER_215_1673 ();
 b15zdnd00an1n01x5 FILLER_215_1677 ();
 b15zdnd11an1n04x5 FILLER_215_1681 ();
 b15zdnd00an1n01x5 FILLER_215_1685 ();
 b15zdnd11an1n64x5 FILLER_215_1689 ();
 b15zdnd11an1n32x5 FILLER_215_1753 ();
 b15zdnd11an1n16x5 FILLER_215_1785 ();
 b15zdnd00an1n01x5 FILLER_215_1801 ();
 b15zdnd11an1n64x5 FILLER_215_1810 ();
 b15zdnd11an1n64x5 FILLER_215_1874 ();
 b15zdnd11an1n64x5 FILLER_215_1938 ();
 b15zdnd11an1n64x5 FILLER_215_2002 ();
 b15zdnd11an1n64x5 FILLER_215_2066 ();
 b15zdnd11an1n64x5 FILLER_215_2130 ();
 b15zdnd11an1n32x5 FILLER_215_2194 ();
 b15zdnd11an1n16x5 FILLER_215_2226 ();
 b15zdnd11an1n04x5 FILLER_215_2242 ();
 b15zdnd00an1n02x5 FILLER_215_2246 ();
 b15zdnd11an1n16x5 FILLER_215_2254 ();
 b15zdnd11an1n08x5 FILLER_215_2270 ();
 b15zdnd11an1n04x5 FILLER_215_2278 ();
 b15zdnd00an1n02x5 FILLER_215_2282 ();
 b15zdnd11an1n64x5 FILLER_216_8 ();
 b15zdnd11an1n64x5 FILLER_216_72 ();
 b15zdnd11an1n64x5 FILLER_216_136 ();
 b15zdnd11an1n08x5 FILLER_216_200 ();
 b15zdnd11an1n04x5 FILLER_216_221 ();
 b15zdnd11an1n04x5 FILLER_216_230 ();
 b15zdnd00an1n02x5 FILLER_216_234 ();
 b15zdnd00an1n01x5 FILLER_216_236 ();
 b15zdnd11an1n32x5 FILLER_216_279 ();
 b15zdnd11an1n08x5 FILLER_216_311 ();
 b15zdnd11an1n04x5 FILLER_216_319 ();
 b15zdnd00an1n02x5 FILLER_216_323 ();
 b15zdnd11an1n08x5 FILLER_216_329 ();
 b15zdnd11an1n04x5 FILLER_216_337 ();
 b15zdnd00an1n01x5 FILLER_216_341 ();
 b15zdnd11an1n64x5 FILLER_216_384 ();
 b15zdnd11an1n16x5 FILLER_216_448 ();
 b15zdnd11an1n04x5 FILLER_216_467 ();
 b15zdnd11an1n64x5 FILLER_216_474 ();
 b15zdnd11an1n64x5 FILLER_216_538 ();
 b15zdnd11an1n08x5 FILLER_216_602 ();
 b15zdnd11an1n04x5 FILLER_216_610 ();
 b15zdnd11an1n04x5 FILLER_216_617 ();
 b15zdnd11an1n64x5 FILLER_216_624 ();
 b15zdnd11an1n16x5 FILLER_216_688 ();
 b15zdnd11an1n08x5 FILLER_216_704 ();
 b15zdnd11an1n04x5 FILLER_216_712 ();
 b15zdnd00an1n02x5 FILLER_216_716 ();
 b15zdnd11an1n64x5 FILLER_216_726 ();
 b15zdnd11an1n16x5 FILLER_216_790 ();
 b15zdnd00an1n01x5 FILLER_216_806 ();
 b15zdnd11an1n04x5 FILLER_216_827 ();
 b15zdnd11an1n16x5 FILLER_216_849 ();
 b15zdnd11an1n08x5 FILLER_216_865 ();
 b15zdnd11an1n16x5 FILLER_216_880 ();
 b15zdnd11an1n32x5 FILLER_216_910 ();
 b15zdnd11an1n16x5 FILLER_216_942 ();
 b15zdnd11an1n08x5 FILLER_216_958 ();
 b15zdnd11an1n04x5 FILLER_216_966 ();
 b15zdnd11an1n16x5 FILLER_216_1014 ();
 b15zdnd11an1n64x5 FILLER_216_1046 ();
 b15zdnd11an1n64x5 FILLER_216_1110 ();
 b15zdnd11an1n08x5 FILLER_216_1174 ();
 b15zdnd11an1n04x5 FILLER_216_1182 ();
 b15zdnd00an1n02x5 FILLER_216_1186 ();
 b15zdnd11an1n32x5 FILLER_216_1208 ();
 b15zdnd11an1n16x5 FILLER_216_1240 ();
 b15zdnd11an1n08x5 FILLER_216_1256 ();
 b15zdnd00an1n01x5 FILLER_216_1264 ();
 b15zdnd11an1n04x5 FILLER_216_1281 ();
 b15zdnd11an1n64x5 FILLER_216_1307 ();
 b15zdnd11an1n64x5 FILLER_216_1371 ();
 b15zdnd11an1n32x5 FILLER_216_1435 ();
 b15zdnd11an1n04x5 FILLER_216_1467 ();
 b15zdnd00an1n02x5 FILLER_216_1471 ();
 b15zdnd00an1n01x5 FILLER_216_1473 ();
 b15zdnd11an1n04x5 FILLER_216_1478 ();
 b15zdnd11an1n64x5 FILLER_216_1486 ();
 b15zdnd11an1n32x5 FILLER_216_1550 ();
 b15zdnd11an1n16x5 FILLER_216_1582 ();
 b15zdnd11an1n08x5 FILLER_216_1598 ();
 b15zdnd11an1n04x5 FILLER_216_1606 ();
 b15zdnd00an1n01x5 FILLER_216_1610 ();
 b15zdnd11an1n04x5 FILLER_216_1663 ();
 b15zdnd11an1n04x5 FILLER_216_1670 ();
 b15zdnd11an1n64x5 FILLER_216_1679 ();
 b15zdnd11an1n08x5 FILLER_216_1743 ();
 b15zdnd00an1n01x5 FILLER_216_1751 ();
 b15zdnd11an1n64x5 FILLER_216_1772 ();
 b15zdnd11an1n64x5 FILLER_216_1836 ();
 b15zdnd11an1n64x5 FILLER_216_1900 ();
 b15zdnd11an1n64x5 FILLER_216_1964 ();
 b15zdnd11an1n64x5 FILLER_216_2028 ();
 b15zdnd11an1n32x5 FILLER_216_2092 ();
 b15zdnd11an1n16x5 FILLER_216_2124 ();
 b15zdnd11an1n08x5 FILLER_216_2140 ();
 b15zdnd11an1n04x5 FILLER_216_2148 ();
 b15zdnd00an1n02x5 FILLER_216_2152 ();
 b15zdnd11an1n64x5 FILLER_216_2162 ();
 b15zdnd11an1n16x5 FILLER_216_2226 ();
 b15zdnd11an1n04x5 FILLER_216_2242 ();
 b15zdnd11an1n16x5 FILLER_216_2250 ();
 b15zdnd11an1n08x5 FILLER_216_2266 ();
 b15zdnd00an1n02x5 FILLER_216_2274 ();
 b15zdnd11an1n64x5 FILLER_217_0 ();
 b15zdnd11an1n64x5 FILLER_217_64 ();
 b15zdnd11an1n64x5 FILLER_217_128 ();
 b15zdnd11an1n08x5 FILLER_217_192 ();
 b15zdnd11an1n04x5 FILLER_217_200 ();
 b15zdnd00an1n01x5 FILLER_217_204 ();
 b15zdnd11an1n16x5 FILLER_217_247 ();
 b15zdnd11an1n04x5 FILLER_217_263 ();
 b15zdnd11an1n64x5 FILLER_217_309 ();
 b15zdnd11an1n08x5 FILLER_217_373 ();
 b15zdnd00an1n01x5 FILLER_217_381 ();
 b15zdnd11an1n32x5 FILLER_217_424 ();
 b15zdnd11an1n08x5 FILLER_217_456 ();
 b15zdnd11an1n64x5 FILLER_217_467 ();
 b15zdnd11an1n64x5 FILLER_217_531 ();
 b15zdnd11an1n16x5 FILLER_217_595 ();
 b15zdnd11an1n08x5 FILLER_217_611 ();
 b15zdnd00an1n01x5 FILLER_217_619 ();
 b15zdnd11an1n64x5 FILLER_217_623 ();
 b15zdnd11an1n64x5 FILLER_217_687 ();
 b15zdnd11an1n32x5 FILLER_217_751 ();
 b15zdnd00an1n01x5 FILLER_217_783 ();
 b15zdnd11an1n16x5 FILLER_217_804 ();
 b15zdnd11an1n04x5 FILLER_217_820 ();
 b15zdnd00an1n02x5 FILLER_217_824 ();
 b15zdnd11an1n64x5 FILLER_217_868 ();
 b15zdnd11an1n32x5 FILLER_217_932 ();
 b15zdnd11an1n04x5 FILLER_217_964 ();
 b15zdnd00an1n01x5 FILLER_217_968 ();
 b15zdnd11an1n04x5 FILLER_217_995 ();
 b15zdnd11an1n08x5 FILLER_217_1013 ();
 b15zdnd00an1n02x5 FILLER_217_1021 ();
 b15zdnd11an1n64x5 FILLER_217_1043 ();
 b15zdnd11an1n32x5 FILLER_217_1107 ();
 b15zdnd11an1n16x5 FILLER_217_1139 ();
 b15zdnd00an1n01x5 FILLER_217_1155 ();
 b15zdnd11an1n64x5 FILLER_217_1198 ();
 b15zdnd11an1n64x5 FILLER_217_1262 ();
 b15zdnd00an1n01x5 FILLER_217_1326 ();
 b15zdnd11an1n64x5 FILLER_217_1335 ();
 b15zdnd11an1n64x5 FILLER_217_1399 ();
 b15zdnd11an1n16x5 FILLER_217_1463 ();
 b15zdnd11an1n04x5 FILLER_217_1479 ();
 b15zdnd00an1n01x5 FILLER_217_1483 ();
 b15zdnd11an1n64x5 FILLER_217_1488 ();
 b15zdnd11an1n64x5 FILLER_217_1552 ();
 b15zdnd11an1n08x5 FILLER_217_1616 ();
 b15zdnd11an1n04x5 FILLER_217_1624 ();
 b15zdnd00an1n02x5 FILLER_217_1628 ();
 b15zdnd11an1n04x5 FILLER_217_1633 ();
 b15zdnd11an1n04x5 FILLER_217_1640 ();
 b15zdnd11an1n08x5 FILLER_217_1647 ();
 b15zdnd11an1n16x5 FILLER_217_1664 ();
 b15zdnd11an1n08x5 FILLER_217_1680 ();
 b15zdnd00an1n02x5 FILLER_217_1688 ();
 b15zdnd11an1n64x5 FILLER_217_1732 ();
 b15zdnd11an1n16x5 FILLER_217_1796 ();
 b15zdnd11an1n04x5 FILLER_217_1812 ();
 b15zdnd00an1n01x5 FILLER_217_1816 ();
 b15zdnd11an1n64x5 FILLER_217_1821 ();
 b15zdnd11an1n64x5 FILLER_217_1885 ();
 b15zdnd11an1n64x5 FILLER_217_1949 ();
 b15zdnd11an1n64x5 FILLER_217_2013 ();
 b15zdnd11an1n64x5 FILLER_217_2077 ();
 b15zdnd11an1n64x5 FILLER_217_2141 ();
 b15zdnd11an1n32x5 FILLER_217_2205 ();
 b15zdnd00an1n02x5 FILLER_217_2237 ();
 b15zdnd00an1n01x5 FILLER_217_2239 ();
 b15zdnd00an1n02x5 FILLER_217_2282 ();
 b15zdnd11an1n16x5 FILLER_218_8 ();
 b15zdnd00an1n01x5 FILLER_218_24 ();
 b15zdnd11an1n08x5 FILLER_218_29 ();
 b15zdnd00an1n01x5 FILLER_218_37 ();
 b15zdnd11an1n64x5 FILLER_218_42 ();
 b15zdnd11an1n64x5 FILLER_218_106 ();
 b15zdnd11an1n32x5 FILLER_218_170 ();
 b15zdnd00an1n02x5 FILLER_218_202 ();
 b15zdnd11an1n04x5 FILLER_218_213 ();
 b15zdnd11an1n64x5 FILLER_218_259 ();
 b15zdnd11an1n16x5 FILLER_218_323 ();
 b15zdnd11an1n08x5 FILLER_218_339 ();
 b15zdnd00an1n02x5 FILLER_218_347 ();
 b15zdnd11an1n64x5 FILLER_218_352 ();
 b15zdnd11an1n64x5 FILLER_218_416 ();
 b15zdnd11an1n64x5 FILLER_218_480 ();
 b15zdnd11an1n32x5 FILLER_218_544 ();
 b15zdnd11an1n16x5 FILLER_218_576 ();
 b15zdnd11an1n08x5 FILLER_218_592 ();
 b15zdnd11an1n04x5 FILLER_218_600 ();
 b15zdnd00an1n01x5 FILLER_218_604 ();
 b15zdnd11an1n04x5 FILLER_218_632 ();
 b15zdnd11an1n04x5 FILLER_218_639 ();
 b15zdnd11an1n64x5 FILLER_218_646 ();
 b15zdnd11an1n08x5 FILLER_218_710 ();
 b15zdnd11an1n64x5 FILLER_218_726 ();
 b15zdnd11an1n32x5 FILLER_218_790 ();
 b15zdnd11an1n08x5 FILLER_218_822 ();
 b15zdnd00an1n02x5 FILLER_218_830 ();
 b15zdnd11an1n04x5 FILLER_218_849 ();
 b15zdnd11an1n32x5 FILLER_218_867 ();
 b15zdnd11an1n04x5 FILLER_218_899 ();
 b15zdnd00an1n02x5 FILLER_218_903 ();
 b15zdnd00an1n01x5 FILLER_218_905 ();
 b15zdnd11an1n04x5 FILLER_218_920 ();
 b15zdnd11an1n32x5 FILLER_218_938 ();
 b15zdnd11an1n16x5 FILLER_218_970 ();
 b15zdnd11an1n04x5 FILLER_218_986 ();
 b15zdnd00an1n01x5 FILLER_218_990 ();
 b15zdnd11an1n16x5 FILLER_218_994 ();
 b15zdnd00an1n01x5 FILLER_218_1010 ();
 b15zdnd11an1n04x5 FILLER_218_1016 ();
 b15zdnd11an1n64x5 FILLER_218_1032 ();
 b15zdnd11an1n64x5 FILLER_218_1096 ();
 b15zdnd11an1n64x5 FILLER_218_1160 ();
 b15zdnd11an1n64x5 FILLER_218_1224 ();
 b15zdnd11an1n64x5 FILLER_218_1288 ();
 b15zdnd11an1n64x5 FILLER_218_1352 ();
 b15zdnd11an1n32x5 FILLER_218_1416 ();
 b15zdnd11an1n16x5 FILLER_218_1448 ();
 b15zdnd00an1n02x5 FILLER_218_1464 ();
 b15zdnd00an1n01x5 FILLER_218_1466 ();
 b15zdnd11an1n64x5 FILLER_218_1475 ();
 b15zdnd11an1n16x5 FILLER_218_1539 ();
 b15zdnd11an1n08x5 FILLER_218_1555 ();
 b15zdnd11an1n04x5 FILLER_218_1563 ();
 b15zdnd11an1n32x5 FILLER_218_1578 ();
 b15zdnd00an1n02x5 FILLER_218_1610 ();
 b15zdnd00an1n01x5 FILLER_218_1612 ();
 b15zdnd11an1n04x5 FILLER_218_1639 ();
 b15zdnd11an1n04x5 FILLER_218_1646 ();
 b15zdnd00an1n01x5 FILLER_218_1650 ();
 b15zdnd11an1n04x5 FILLER_218_1654 ();
 b15zdnd11an1n64x5 FILLER_218_1661 ();
 b15zdnd11an1n64x5 FILLER_218_1725 ();
 b15zdnd11an1n16x5 FILLER_218_1789 ();
 b15zdnd11an1n08x5 FILLER_218_1805 ();
 b15zdnd00an1n01x5 FILLER_218_1813 ();
 b15zdnd11an1n32x5 FILLER_218_1819 ();
 b15zdnd00an1n01x5 FILLER_218_1851 ();
 b15zdnd11an1n32x5 FILLER_218_1866 ();
 b15zdnd11an1n16x5 FILLER_218_1898 ();
 b15zdnd11an1n08x5 FILLER_218_1914 ();
 b15zdnd00an1n02x5 FILLER_218_1922 ();
 b15zdnd11an1n64x5 FILLER_218_1931 ();
 b15zdnd11an1n64x5 FILLER_218_1995 ();
 b15zdnd11an1n64x5 FILLER_218_2059 ();
 b15zdnd11an1n16x5 FILLER_218_2123 ();
 b15zdnd11an1n08x5 FILLER_218_2139 ();
 b15zdnd11an1n04x5 FILLER_218_2147 ();
 b15zdnd00an1n02x5 FILLER_218_2151 ();
 b15zdnd00an1n01x5 FILLER_218_2153 ();
 b15zdnd11an1n64x5 FILLER_218_2162 ();
 b15zdnd11an1n16x5 FILLER_218_2226 ();
 b15zdnd11an1n04x5 FILLER_218_2242 ();
 b15zdnd11an1n08x5 FILLER_218_2266 ();
 b15zdnd00an1n02x5 FILLER_218_2274 ();
 b15zdnd11an1n08x5 FILLER_219_0 ();
 b15zdnd11an1n64x5 FILLER_219_50 ();
 b15zdnd11an1n64x5 FILLER_219_114 ();
 b15zdnd11an1n16x5 FILLER_219_178 ();
 b15zdnd11an1n08x5 FILLER_219_194 ();
 b15zdnd11an1n04x5 FILLER_219_202 ();
 b15zdnd11an1n04x5 FILLER_219_216 ();
 b15zdnd11an1n32x5 FILLER_219_262 ();
 b15zdnd11an1n16x5 FILLER_219_294 ();
 b15zdnd11an1n08x5 FILLER_219_310 ();
 b15zdnd11an1n04x5 FILLER_219_318 ();
 b15zdnd00an1n02x5 FILLER_219_322 ();
 b15zdnd00an1n01x5 FILLER_219_324 ();
 b15zdnd11an1n04x5 FILLER_219_367 ();
 b15zdnd11an1n64x5 FILLER_219_389 ();
 b15zdnd11an1n64x5 FILLER_219_453 ();
 b15zdnd11an1n64x5 FILLER_219_517 ();
 b15zdnd11an1n16x5 FILLER_219_581 ();
 b15zdnd11an1n04x5 FILLER_219_597 ();
 b15zdnd00an1n02x5 FILLER_219_601 ();
 b15zdnd00an1n01x5 FILLER_219_603 ();
 b15zdnd11an1n04x5 FILLER_219_607 ();
 b15zdnd11an1n64x5 FILLER_219_663 ();
 b15zdnd11an1n32x5 FILLER_219_727 ();
 b15zdnd11an1n16x5 FILLER_219_759 ();
 b15zdnd00an1n01x5 FILLER_219_775 ();
 b15zdnd11an1n16x5 FILLER_219_780 ();
 b15zdnd11an1n08x5 FILLER_219_796 ();
 b15zdnd00an1n01x5 FILLER_219_804 ();
 b15zdnd11an1n08x5 FILLER_219_817 ();
 b15zdnd00an1n02x5 FILLER_219_825 ();
 b15zdnd00an1n01x5 FILLER_219_827 ();
 b15zdnd11an1n64x5 FILLER_219_845 ();
 b15zdnd11an1n32x5 FILLER_219_909 ();
 b15zdnd11an1n16x5 FILLER_219_941 ();
 b15zdnd11an1n08x5 FILLER_219_957 ();
 b15zdnd11an1n04x5 FILLER_219_965 ();
 b15zdnd00an1n02x5 FILLER_219_969 ();
 b15zdnd00an1n01x5 FILLER_219_971 ();
 b15zdnd11an1n64x5 FILLER_219_979 ();
 b15zdnd11an1n64x5 FILLER_219_1043 ();
 b15zdnd11an1n16x5 FILLER_219_1107 ();
 b15zdnd11an1n08x5 FILLER_219_1123 ();
 b15zdnd11an1n04x5 FILLER_219_1131 ();
 b15zdnd00an1n01x5 FILLER_219_1135 ();
 b15zdnd11an1n64x5 FILLER_219_1188 ();
 b15zdnd11an1n32x5 FILLER_219_1252 ();
 b15zdnd11an1n16x5 FILLER_219_1284 ();
 b15zdnd11an1n04x5 FILLER_219_1300 ();
 b15zdnd00an1n01x5 FILLER_219_1304 ();
 b15zdnd11an1n64x5 FILLER_219_1311 ();
 b15zdnd11an1n64x5 FILLER_219_1375 ();
 b15zdnd11an1n64x5 FILLER_219_1439 ();
 b15zdnd11an1n16x5 FILLER_219_1503 ();
 b15zdnd11an1n32x5 FILLER_219_1533 ();
 b15zdnd11an1n64x5 FILLER_219_1571 ();
 b15zdnd00an1n01x5 FILLER_219_1635 ();
 b15zdnd11an1n64x5 FILLER_219_1639 ();
 b15zdnd11an1n64x5 FILLER_219_1703 ();
 b15zdnd11an1n64x5 FILLER_219_1767 ();
 b15zdnd11an1n64x5 FILLER_219_1831 ();
 b15zdnd11an1n04x5 FILLER_219_1895 ();
 b15zdnd11an1n04x5 FILLER_219_1905 ();
 b15zdnd00an1n01x5 FILLER_219_1909 ();
 b15zdnd11an1n64x5 FILLER_219_1927 ();
 b15zdnd11an1n64x5 FILLER_219_1991 ();
 b15zdnd11an1n64x5 FILLER_219_2055 ();
 b15zdnd11an1n64x5 FILLER_219_2119 ();
 b15zdnd11an1n64x5 FILLER_219_2183 ();
 b15zdnd11an1n04x5 FILLER_219_2247 ();
 b15zdnd00an1n02x5 FILLER_219_2251 ();
 b15zdnd11an1n16x5 FILLER_219_2259 ();
 b15zdnd11an1n08x5 FILLER_219_2275 ();
 b15zdnd00an1n01x5 FILLER_219_2283 ();
 b15zdnd11an1n04x5 FILLER_220_8 ();
 b15zdnd00an1n02x5 FILLER_220_12 ();
 b15zdnd00an1n01x5 FILLER_220_14 ();
 b15zdnd11an1n64x5 FILLER_220_57 ();
 b15zdnd11an1n64x5 FILLER_220_121 ();
 b15zdnd11an1n16x5 FILLER_220_185 ();
 b15zdnd11an1n04x5 FILLER_220_201 ();
 b15zdnd00an1n02x5 FILLER_220_205 ();
 b15zdnd00an1n01x5 FILLER_220_207 ();
 b15zdnd11an1n04x5 FILLER_220_218 ();
 b15zdnd00an1n02x5 FILLER_220_222 ();
 b15zdnd00an1n01x5 FILLER_220_224 ();
 b15zdnd11an1n04x5 FILLER_220_230 ();
 b15zdnd11an1n64x5 FILLER_220_237 ();
 b15zdnd11an1n16x5 FILLER_220_301 ();
 b15zdnd11an1n04x5 FILLER_220_317 ();
 b15zdnd00an1n01x5 FILLER_220_321 ();
 b15zdnd11an1n04x5 FILLER_220_374 ();
 b15zdnd11an1n64x5 FILLER_220_420 ();
 b15zdnd11an1n64x5 FILLER_220_484 ();
 b15zdnd11an1n32x5 FILLER_220_548 ();
 b15zdnd11an1n16x5 FILLER_220_580 ();
 b15zdnd11an1n08x5 FILLER_220_596 ();
 b15zdnd11an1n04x5 FILLER_220_607 ();
 b15zdnd11an1n04x5 FILLER_220_614 ();
 b15zdnd11an1n08x5 FILLER_220_670 ();
 b15zdnd11an1n32x5 FILLER_220_685 ();
 b15zdnd00an1n01x5 FILLER_220_717 ();
 b15zdnd11an1n08x5 FILLER_220_726 ();
 b15zdnd00an1n02x5 FILLER_220_734 ();
 b15zdnd11an1n32x5 FILLER_220_740 ();
 b15zdnd00an1n02x5 FILLER_220_772 ();
 b15zdnd00an1n01x5 FILLER_220_774 ();
 b15zdnd11an1n32x5 FILLER_220_779 ();
 b15zdnd11an1n16x5 FILLER_220_811 ();
 b15zdnd11an1n08x5 FILLER_220_827 ();
 b15zdnd00an1n02x5 FILLER_220_835 ();
 b15zdnd11an1n64x5 FILLER_220_843 ();
 b15zdnd11an1n32x5 FILLER_220_907 ();
 b15zdnd11an1n08x5 FILLER_220_939 ();
 b15zdnd00an1n02x5 FILLER_220_947 ();
 b15zdnd00an1n01x5 FILLER_220_949 ();
 b15zdnd11an1n64x5 FILLER_220_958 ();
 b15zdnd11an1n32x5 FILLER_220_1022 ();
 b15zdnd11an1n08x5 FILLER_220_1054 ();
 b15zdnd11an1n04x5 FILLER_220_1062 ();
 b15zdnd00an1n02x5 FILLER_220_1066 ();
 b15zdnd00an1n01x5 FILLER_220_1068 ();
 b15zdnd11an1n32x5 FILLER_220_1111 ();
 b15zdnd11an1n08x5 FILLER_220_1143 ();
 b15zdnd00an1n02x5 FILLER_220_1151 ();
 b15zdnd00an1n01x5 FILLER_220_1153 ();
 b15zdnd11an1n04x5 FILLER_220_1157 ();
 b15zdnd11an1n04x5 FILLER_220_1164 ();
 b15zdnd11an1n64x5 FILLER_220_1171 ();
 b15zdnd11an1n16x5 FILLER_220_1235 ();
 b15zdnd11an1n08x5 FILLER_220_1251 ();
 b15zdnd00an1n01x5 FILLER_220_1259 ();
 b15zdnd11an1n16x5 FILLER_220_1263 ();
 b15zdnd11an1n08x5 FILLER_220_1279 ();
 b15zdnd11an1n04x5 FILLER_220_1287 ();
 b15zdnd00an1n02x5 FILLER_220_1291 ();
 b15zdnd11an1n64x5 FILLER_220_1345 ();
 b15zdnd11an1n32x5 FILLER_220_1409 ();
 b15zdnd11an1n08x5 FILLER_220_1441 ();
 b15zdnd11an1n04x5 FILLER_220_1449 ();
 b15zdnd00an1n02x5 FILLER_220_1453 ();
 b15zdnd11an1n32x5 FILLER_220_1461 ();
 b15zdnd11an1n16x5 FILLER_220_1493 ();
 b15zdnd11an1n08x5 FILLER_220_1509 ();
 b15zdnd11an1n64x5 FILLER_220_1541 ();
 b15zdnd11an1n64x5 FILLER_220_1605 ();
 b15zdnd11an1n64x5 FILLER_220_1669 ();
 b15zdnd11an1n64x5 FILLER_220_1733 ();
 b15zdnd11an1n64x5 FILLER_220_1797 ();
 b15zdnd11an1n32x5 FILLER_220_1861 ();
 b15zdnd11an1n16x5 FILLER_220_1893 ();
 b15zdnd00an1n01x5 FILLER_220_1909 ();
 b15zdnd11an1n64x5 FILLER_220_1930 ();
 b15zdnd11an1n64x5 FILLER_220_1994 ();
 b15zdnd11an1n32x5 FILLER_220_2058 ();
 b15zdnd11an1n16x5 FILLER_220_2090 ();
 b15zdnd00an1n01x5 FILLER_220_2106 ();
 b15zdnd11an1n04x5 FILLER_220_2149 ();
 b15zdnd00an1n01x5 FILLER_220_2153 ();
 b15zdnd11an1n64x5 FILLER_220_2162 ();
 b15zdnd11an1n32x5 FILLER_220_2226 ();
 b15zdnd11an1n16x5 FILLER_220_2258 ();
 b15zdnd00an1n02x5 FILLER_220_2274 ();
 b15zdnd11an1n16x5 FILLER_221_0 ();
 b15zdnd11an1n04x5 FILLER_221_16 ();
 b15zdnd00an1n02x5 FILLER_221_20 ();
 b15zdnd11an1n04x5 FILLER_221_26 ();
 b15zdnd11an1n64x5 FILLER_221_37 ();
 b15zdnd11an1n64x5 FILLER_221_101 ();
 b15zdnd11an1n16x5 FILLER_221_165 ();
 b15zdnd11an1n08x5 FILLER_221_181 ();
 b15zdnd00an1n02x5 FILLER_221_189 ();
 b15zdnd00an1n01x5 FILLER_221_191 ();
 b15zdnd11an1n64x5 FILLER_221_244 ();
 b15zdnd11an1n32x5 FILLER_221_308 ();
 b15zdnd11an1n04x5 FILLER_221_343 ();
 b15zdnd11an1n64x5 FILLER_221_350 ();
 b15zdnd11an1n64x5 FILLER_221_414 ();
 b15zdnd11an1n04x5 FILLER_221_486 ();
 b15zdnd11an1n32x5 FILLER_221_532 ();
 b15zdnd11an1n16x5 FILLER_221_564 ();
 b15zdnd11an1n08x5 FILLER_221_580 ();
 b15zdnd11an1n04x5 FILLER_221_588 ();
 b15zdnd00an1n02x5 FILLER_221_592 ();
 b15zdnd00an1n01x5 FILLER_221_594 ();
 b15zdnd11an1n04x5 FILLER_221_647 ();
 b15zdnd11an1n64x5 FILLER_221_654 ();
 b15zdnd11an1n64x5 FILLER_221_718 ();
 b15zdnd11an1n64x5 FILLER_221_782 ();
 b15zdnd11an1n64x5 FILLER_221_846 ();
 b15zdnd11an1n64x5 FILLER_221_910 ();
 b15zdnd11an1n64x5 FILLER_221_974 ();
 b15zdnd11an1n64x5 FILLER_221_1038 ();
 b15zdnd11an1n32x5 FILLER_221_1102 ();
 b15zdnd11an1n16x5 FILLER_221_1134 ();
 b15zdnd11an1n04x5 FILLER_221_1150 ();
 b15zdnd00an1n02x5 FILLER_221_1154 ();
 b15zdnd00an1n01x5 FILLER_221_1156 ();
 b15zdnd11an1n08x5 FILLER_221_1164 ();
 b15zdnd11an1n04x5 FILLER_221_1172 ();
 b15zdnd00an1n02x5 FILLER_221_1176 ();
 b15zdnd00an1n01x5 FILLER_221_1178 ();
 b15zdnd11an1n64x5 FILLER_221_1183 ();
 b15zdnd11an1n08x5 FILLER_221_1247 ();
 b15zdnd11an1n04x5 FILLER_221_1255 ();
 b15zdnd00an1n01x5 FILLER_221_1259 ();
 b15zdnd11an1n32x5 FILLER_221_1263 ();
 b15zdnd11an1n16x5 FILLER_221_1295 ();
 b15zdnd11an1n04x5 FILLER_221_1314 ();
 b15zdnd11an1n64x5 FILLER_221_1321 ();
 b15zdnd11an1n64x5 FILLER_221_1385 ();
 b15zdnd11an1n32x5 FILLER_221_1449 ();
 b15zdnd11an1n16x5 FILLER_221_1481 ();
 b15zdnd11an1n64x5 FILLER_221_1517 ();
 b15zdnd11an1n32x5 FILLER_221_1581 ();
 b15zdnd11an1n08x5 FILLER_221_1613 ();
 b15zdnd11an1n04x5 FILLER_221_1648 ();
 b15zdnd00an1n02x5 FILLER_221_1652 ();
 b15zdnd00an1n01x5 FILLER_221_1654 ();
 b15zdnd11an1n64x5 FILLER_221_1664 ();
 b15zdnd11an1n32x5 FILLER_221_1728 ();
 b15zdnd11an1n16x5 FILLER_221_1760 ();
 b15zdnd11an1n64x5 FILLER_221_1791 ();
 b15zdnd11an1n64x5 FILLER_221_1855 ();
 b15zdnd11an1n64x5 FILLER_221_1919 ();
 b15zdnd11an1n64x5 FILLER_221_1983 ();
 b15zdnd11an1n08x5 FILLER_221_2047 ();
 b15zdnd11an1n04x5 FILLER_221_2055 ();
 b15zdnd00an1n02x5 FILLER_221_2059 ();
 b15zdnd11an1n64x5 FILLER_221_2103 ();
 b15zdnd11an1n64x5 FILLER_221_2167 ();
 b15zdnd11an1n16x5 FILLER_221_2231 ();
 b15zdnd11an1n08x5 FILLER_221_2247 ();
 b15zdnd00an1n02x5 FILLER_221_2255 ();
 b15zdnd00an1n01x5 FILLER_221_2257 ();
 b15zdnd11an1n16x5 FILLER_221_2263 ();
 b15zdnd11an1n04x5 FILLER_221_2279 ();
 b15zdnd00an1n01x5 FILLER_221_2283 ();
 b15zdnd11an1n64x5 FILLER_222_8 ();
 b15zdnd11an1n64x5 FILLER_222_72 ();
 b15zdnd11an1n64x5 FILLER_222_136 ();
 b15zdnd11an1n08x5 FILLER_222_200 ();
 b15zdnd11an1n04x5 FILLER_222_208 ();
 b15zdnd11an1n04x5 FILLER_222_215 ();
 b15zdnd11an1n64x5 FILLER_222_222 ();
 b15zdnd11an1n64x5 FILLER_222_286 ();
 b15zdnd11an1n64x5 FILLER_222_350 ();
 b15zdnd11an1n64x5 FILLER_222_414 ();
 b15zdnd11an1n64x5 FILLER_222_478 ();
 b15zdnd11an1n64x5 FILLER_222_542 ();
 b15zdnd11an1n08x5 FILLER_222_606 ();
 b15zdnd11an1n04x5 FILLER_222_614 ();
 b15zdnd00an1n02x5 FILLER_222_618 ();
 b15zdnd11an1n04x5 FILLER_222_627 ();
 b15zdnd00an1n02x5 FILLER_222_631 ();
 b15zdnd00an1n01x5 FILLER_222_633 ();
 b15zdnd11an1n04x5 FILLER_222_637 ();
 b15zdnd00an1n02x5 FILLER_222_641 ();
 b15zdnd11an1n64x5 FILLER_222_646 ();
 b15zdnd11an1n08x5 FILLER_222_710 ();
 b15zdnd11an1n64x5 FILLER_222_726 ();
 b15zdnd11an1n64x5 FILLER_222_790 ();
 b15zdnd11an1n08x5 FILLER_222_854 ();
 b15zdnd11an1n04x5 FILLER_222_862 ();
 b15zdnd00an1n02x5 FILLER_222_866 ();
 b15zdnd00an1n01x5 FILLER_222_868 ();
 b15zdnd11an1n32x5 FILLER_222_875 ();
 b15zdnd11an1n16x5 FILLER_222_907 ();
 b15zdnd11an1n08x5 FILLER_222_923 ();
 b15zdnd11an1n04x5 FILLER_222_931 ();
 b15zdnd11an1n64x5 FILLER_222_942 ();
 b15zdnd11an1n32x5 FILLER_222_1006 ();
 b15zdnd11an1n04x5 FILLER_222_1038 ();
 b15zdnd11an1n64x5 FILLER_222_1065 ();
 b15zdnd11an1n64x5 FILLER_222_1129 ();
 b15zdnd11an1n04x5 FILLER_222_1193 ();
 b15zdnd00an1n01x5 FILLER_222_1197 ();
 b15zdnd11an1n16x5 FILLER_222_1209 ();
 b15zdnd11an1n08x5 FILLER_222_1225 ();
 b15zdnd11an1n04x5 FILLER_222_1233 ();
 b15zdnd00an1n01x5 FILLER_222_1237 ();
 b15zdnd11an1n32x5 FILLER_222_1282 ();
 b15zdnd00an1n02x5 FILLER_222_1314 ();
 b15zdnd00an1n01x5 FILLER_222_1316 ();
 b15zdnd11an1n64x5 FILLER_222_1320 ();
 b15zdnd11an1n64x5 FILLER_222_1384 ();
 b15zdnd11an1n32x5 FILLER_222_1448 ();
 b15zdnd11an1n16x5 FILLER_222_1480 ();
 b15zdnd11an1n04x5 FILLER_222_1496 ();
 b15zdnd00an1n01x5 FILLER_222_1500 ();
 b15zdnd11an1n64x5 FILLER_222_1521 ();
 b15zdnd11an1n32x5 FILLER_222_1585 ();
 b15zdnd11an1n04x5 FILLER_222_1617 ();
 b15zdnd00an1n02x5 FILLER_222_1621 ();
 b15zdnd00an1n01x5 FILLER_222_1623 ();
 b15zdnd11an1n64x5 FILLER_222_1627 ();
 b15zdnd11an1n64x5 FILLER_222_1691 ();
 b15zdnd11an1n16x5 FILLER_222_1755 ();
 b15zdnd11an1n04x5 FILLER_222_1771 ();
 b15zdnd00an1n02x5 FILLER_222_1775 ();
 b15zdnd00an1n01x5 FILLER_222_1777 ();
 b15zdnd11an1n64x5 FILLER_222_1796 ();
 b15zdnd11an1n64x5 FILLER_222_1860 ();
 b15zdnd11an1n64x5 FILLER_222_1924 ();
 b15zdnd11an1n32x5 FILLER_222_1988 ();
 b15zdnd11an1n04x5 FILLER_222_2020 ();
 b15zdnd00an1n02x5 FILLER_222_2024 ();
 b15zdnd11an1n64x5 FILLER_222_2050 ();
 b15zdnd11an1n32x5 FILLER_222_2114 ();
 b15zdnd11an1n08x5 FILLER_222_2146 ();
 b15zdnd11an1n16x5 FILLER_222_2162 ();
 b15zdnd00an1n02x5 FILLER_222_2178 ();
 b15zdnd00an1n01x5 FILLER_222_2180 ();
 b15zdnd11an1n64x5 FILLER_222_2207 ();
 b15zdnd11an1n04x5 FILLER_222_2271 ();
 b15zdnd00an1n01x5 FILLER_222_2275 ();
 b15zdnd11an1n64x5 FILLER_223_0 ();
 b15zdnd11an1n64x5 FILLER_223_64 ();
 b15zdnd11an1n64x5 FILLER_223_128 ();
 b15zdnd11an1n16x5 FILLER_223_192 ();
 b15zdnd11an1n08x5 FILLER_223_208 ();
 b15zdnd00an1n02x5 FILLER_223_216 ();
 b15zdnd11an1n64x5 FILLER_223_221 ();
 b15zdnd11an1n64x5 FILLER_223_285 ();
 b15zdnd11an1n64x5 FILLER_223_349 ();
 b15zdnd11an1n64x5 FILLER_223_413 ();
 b15zdnd11an1n64x5 FILLER_223_477 ();
 b15zdnd11an1n64x5 FILLER_223_541 ();
 b15zdnd11an1n32x5 FILLER_223_605 ();
 b15zdnd11an1n64x5 FILLER_223_640 ();
 b15zdnd11an1n64x5 FILLER_223_704 ();
 b15zdnd11an1n64x5 FILLER_223_768 ();
 b15zdnd11an1n64x5 FILLER_223_832 ();
 b15zdnd11an1n16x5 FILLER_223_896 ();
 b15zdnd11an1n08x5 FILLER_223_912 ();
 b15zdnd00an1n02x5 FILLER_223_920 ();
 b15zdnd11an1n64x5 FILLER_223_942 ();
 b15zdnd11an1n32x5 FILLER_223_1006 ();
 b15zdnd11an1n04x5 FILLER_223_1038 ();
 b15zdnd11an1n04x5 FILLER_223_1062 ();
 b15zdnd11an1n64x5 FILLER_223_1097 ();
 b15zdnd11an1n16x5 FILLER_223_1161 ();
 b15zdnd11an1n08x5 FILLER_223_1177 ();
 b15zdnd11an1n64x5 FILLER_223_1193 ();
 b15zdnd11an1n04x5 FILLER_223_1257 ();
 b15zdnd11an1n64x5 FILLER_223_1264 ();
 b15zdnd11an1n64x5 FILLER_223_1328 ();
 b15zdnd11an1n64x5 FILLER_223_1392 ();
 b15zdnd11an1n64x5 FILLER_223_1456 ();
 b15zdnd11an1n64x5 FILLER_223_1520 ();
 b15zdnd11an1n64x5 FILLER_223_1584 ();
 b15zdnd11an1n64x5 FILLER_223_1648 ();
 b15zdnd11an1n64x5 FILLER_223_1712 ();
 b15zdnd11an1n64x5 FILLER_223_1776 ();
 b15zdnd11an1n64x5 FILLER_223_1840 ();
 b15zdnd11an1n64x5 FILLER_223_1904 ();
 b15zdnd11an1n64x5 FILLER_223_1968 ();
 b15zdnd11an1n32x5 FILLER_223_2032 ();
 b15zdnd11an1n16x5 FILLER_223_2064 ();
 b15zdnd11an1n08x5 FILLER_223_2080 ();
 b15zdnd00an1n02x5 FILLER_223_2088 ();
 b15zdnd00an1n01x5 FILLER_223_2090 ();
 b15zdnd11an1n32x5 FILLER_223_2105 ();
 b15zdnd11an1n08x5 FILLER_223_2137 ();
 b15zdnd00an1n02x5 FILLER_223_2145 ();
 b15zdnd00an1n01x5 FILLER_223_2147 ();
 b15zdnd11an1n08x5 FILLER_223_2184 ();
 b15zdnd00an1n02x5 FILLER_223_2192 ();
 b15zdnd11an1n64x5 FILLER_223_2216 ();
 b15zdnd11an1n04x5 FILLER_223_2280 ();
 b15zdnd11an1n64x5 FILLER_224_8 ();
 b15zdnd11an1n64x5 FILLER_224_72 ();
 b15zdnd11an1n64x5 FILLER_224_136 ();
 b15zdnd11an1n08x5 FILLER_224_200 ();
 b15zdnd00an1n02x5 FILLER_224_208 ();
 b15zdnd11an1n64x5 FILLER_224_216 ();
 b15zdnd11an1n64x5 FILLER_224_280 ();
 b15zdnd11an1n64x5 FILLER_224_344 ();
 b15zdnd11an1n32x5 FILLER_224_408 ();
 b15zdnd11an1n16x5 FILLER_224_440 ();
 b15zdnd11an1n08x5 FILLER_224_456 ();
 b15zdnd11an1n64x5 FILLER_224_485 ();
 b15zdnd11an1n64x5 FILLER_224_549 ();
 b15zdnd11an1n64x5 FILLER_224_613 ();
 b15zdnd11an1n32x5 FILLER_224_677 ();
 b15zdnd11an1n08x5 FILLER_224_709 ();
 b15zdnd00an1n01x5 FILLER_224_717 ();
 b15zdnd11an1n64x5 FILLER_224_726 ();
 b15zdnd11an1n32x5 FILLER_224_790 ();
 b15zdnd11an1n08x5 FILLER_224_822 ();
 b15zdnd00an1n01x5 FILLER_224_830 ();
 b15zdnd11an1n64x5 FILLER_224_851 ();
 b15zdnd11an1n16x5 FILLER_224_915 ();
 b15zdnd11an1n64x5 FILLER_224_949 ();
 b15zdnd11an1n64x5 FILLER_224_1013 ();
 b15zdnd11an1n32x5 FILLER_224_1077 ();
 b15zdnd00an1n01x5 FILLER_224_1109 ();
 b15zdnd11an1n64x5 FILLER_224_1133 ();
 b15zdnd11an1n64x5 FILLER_224_1197 ();
 b15zdnd11an1n64x5 FILLER_224_1261 ();
 b15zdnd11an1n64x5 FILLER_224_1325 ();
 b15zdnd11an1n32x5 FILLER_224_1389 ();
 b15zdnd11an1n08x5 FILLER_224_1421 ();
 b15zdnd00an1n02x5 FILLER_224_1429 ();
 b15zdnd00an1n01x5 FILLER_224_1431 ();
 b15zdnd11an1n64x5 FILLER_224_1445 ();
 b15zdnd11an1n64x5 FILLER_224_1509 ();
 b15zdnd11an1n64x5 FILLER_224_1573 ();
 b15zdnd11an1n64x5 FILLER_224_1637 ();
 b15zdnd11an1n64x5 FILLER_224_1701 ();
 b15zdnd11an1n32x5 FILLER_224_1765 ();
 b15zdnd11an1n16x5 FILLER_224_1797 ();
 b15zdnd11an1n04x5 FILLER_224_1813 ();
 b15zdnd11an1n64x5 FILLER_224_1829 ();
 b15zdnd11an1n64x5 FILLER_224_1893 ();
 b15zdnd11an1n64x5 FILLER_224_1957 ();
 b15zdnd11an1n64x5 FILLER_224_2021 ();
 b15zdnd11an1n64x5 FILLER_224_2085 ();
 b15zdnd11an1n04x5 FILLER_224_2149 ();
 b15zdnd00an1n01x5 FILLER_224_2153 ();
 b15zdnd11an1n64x5 FILLER_224_2162 ();
 b15zdnd11an1n32x5 FILLER_224_2226 ();
 b15zdnd11an1n16x5 FILLER_224_2258 ();
 b15zdnd00an1n02x5 FILLER_224_2274 ();
 b15zdnd11an1n16x5 FILLER_225_0 ();
 b15zdnd11an1n08x5 FILLER_225_16 ();
 b15zdnd11an1n04x5 FILLER_225_24 ();
 b15zdnd00an1n02x5 FILLER_225_28 ();
 b15zdnd00an1n01x5 FILLER_225_30 ();
 b15zdnd11an1n64x5 FILLER_225_35 ();
 b15zdnd11an1n64x5 FILLER_225_99 ();
 b15zdnd11an1n64x5 FILLER_225_163 ();
 b15zdnd11an1n64x5 FILLER_225_227 ();
 b15zdnd11an1n64x5 FILLER_225_291 ();
 b15zdnd11an1n64x5 FILLER_225_355 ();
 b15zdnd11an1n32x5 FILLER_225_419 ();
 b15zdnd11an1n08x5 FILLER_225_451 ();
 b15zdnd11an1n04x5 FILLER_225_459 ();
 b15zdnd00an1n02x5 FILLER_225_463 ();
 b15zdnd00an1n01x5 FILLER_225_465 ();
 b15zdnd11an1n64x5 FILLER_225_469 ();
 b15zdnd11an1n64x5 FILLER_225_533 ();
 b15zdnd11an1n64x5 FILLER_225_597 ();
 b15zdnd11an1n64x5 FILLER_225_661 ();
 b15zdnd11an1n64x5 FILLER_225_725 ();
 b15zdnd11an1n32x5 FILLER_225_789 ();
 b15zdnd00an1n01x5 FILLER_225_821 ();
 b15zdnd11an1n64x5 FILLER_225_839 ();
 b15zdnd11an1n16x5 FILLER_225_903 ();
 b15zdnd11an1n08x5 FILLER_225_919 ();
 b15zdnd11an1n04x5 FILLER_225_927 ();
 b15zdnd00an1n02x5 FILLER_225_931 ();
 b15zdnd11an1n32x5 FILLER_225_945 ();
 b15zdnd11an1n08x5 FILLER_225_977 ();
 b15zdnd11an1n64x5 FILLER_225_996 ();
 b15zdnd11an1n16x5 FILLER_225_1060 ();
 b15zdnd00an1n01x5 FILLER_225_1076 ();
 b15zdnd11an1n32x5 FILLER_225_1095 ();
 b15zdnd11an1n04x5 FILLER_225_1127 ();
 b15zdnd00an1n02x5 FILLER_225_1131 ();
 b15zdnd00an1n01x5 FILLER_225_1133 ();
 b15zdnd11an1n32x5 FILLER_225_1148 ();
 b15zdnd11an1n08x5 FILLER_225_1180 ();
 b15zdnd11an1n64x5 FILLER_225_1211 ();
 b15zdnd11an1n64x5 FILLER_225_1275 ();
 b15zdnd00an1n02x5 FILLER_225_1339 ();
 b15zdnd11an1n32x5 FILLER_225_1347 ();
 b15zdnd11an1n04x5 FILLER_225_1379 ();
 b15zdnd00an1n01x5 FILLER_225_1383 ();
 b15zdnd11an1n64x5 FILLER_225_1391 ();
 b15zdnd11an1n64x5 FILLER_225_1455 ();
 b15zdnd11an1n64x5 FILLER_225_1519 ();
 b15zdnd11an1n64x5 FILLER_225_1583 ();
 b15zdnd11an1n64x5 FILLER_225_1647 ();
 b15zdnd11an1n64x5 FILLER_225_1711 ();
 b15zdnd11an1n64x5 FILLER_225_1775 ();
 b15zdnd11an1n32x5 FILLER_225_1839 ();
 b15zdnd11an1n32x5 FILLER_225_1923 ();
 b15zdnd11an1n16x5 FILLER_225_1955 ();
 b15zdnd11an1n08x5 FILLER_225_1971 ();
 b15zdnd11an1n64x5 FILLER_225_1990 ();
 b15zdnd11an1n64x5 FILLER_225_2054 ();
 b15zdnd11an1n64x5 FILLER_225_2118 ();
 b15zdnd11an1n32x5 FILLER_225_2182 ();
 b15zdnd11an1n16x5 FILLER_225_2214 ();
 b15zdnd11an1n08x5 FILLER_225_2230 ();
 b15zdnd11an1n04x5 FILLER_225_2238 ();
 b15zdnd00an1n02x5 FILLER_225_2242 ();
 b15zdnd11an1n32x5 FILLER_225_2248 ();
 b15zdnd11an1n04x5 FILLER_225_2280 ();
 b15zdnd11an1n64x5 FILLER_226_8 ();
 b15zdnd11an1n64x5 FILLER_226_72 ();
 b15zdnd11an1n64x5 FILLER_226_136 ();
 b15zdnd11an1n64x5 FILLER_226_200 ();
 b15zdnd11an1n64x5 FILLER_226_264 ();
 b15zdnd11an1n64x5 FILLER_226_328 ();
 b15zdnd11an1n64x5 FILLER_226_392 ();
 b15zdnd11an1n64x5 FILLER_226_456 ();
 b15zdnd11an1n64x5 FILLER_226_520 ();
 b15zdnd11an1n64x5 FILLER_226_584 ();
 b15zdnd11an1n64x5 FILLER_226_648 ();
 b15zdnd11an1n04x5 FILLER_226_712 ();
 b15zdnd00an1n02x5 FILLER_226_716 ();
 b15zdnd11an1n64x5 FILLER_226_726 ();
 b15zdnd11an1n32x5 FILLER_226_790 ();
 b15zdnd11an1n08x5 FILLER_226_822 ();
 b15zdnd11an1n04x5 FILLER_226_830 ();
 b15zdnd00an1n01x5 FILLER_226_834 ();
 b15zdnd11an1n04x5 FILLER_226_861 ();
 b15zdnd11an1n64x5 FILLER_226_879 ();
 b15zdnd11an1n64x5 FILLER_226_943 ();
 b15zdnd11an1n04x5 FILLER_226_1007 ();
 b15zdnd00an1n02x5 FILLER_226_1011 ();
 b15zdnd00an1n01x5 FILLER_226_1013 ();
 b15zdnd11an1n08x5 FILLER_226_1031 ();
 b15zdnd00an1n02x5 FILLER_226_1039 ();
 b15zdnd00an1n01x5 FILLER_226_1041 ();
 b15zdnd11an1n16x5 FILLER_226_1062 ();
 b15zdnd11an1n08x5 FILLER_226_1078 ();
 b15zdnd11an1n04x5 FILLER_226_1086 ();
 b15zdnd00an1n02x5 FILLER_226_1090 ();
 b15zdnd00an1n01x5 FILLER_226_1092 ();
 b15zdnd11an1n16x5 FILLER_226_1107 ();
 b15zdnd11an1n08x5 FILLER_226_1123 ();
 b15zdnd11an1n04x5 FILLER_226_1131 ();
 b15zdnd00an1n02x5 FILLER_226_1135 ();
 b15zdnd00an1n01x5 FILLER_226_1137 ();
 b15zdnd11an1n16x5 FILLER_226_1150 ();
 b15zdnd11an1n64x5 FILLER_226_1182 ();
 b15zdnd11an1n04x5 FILLER_226_1246 ();
 b15zdnd00an1n02x5 FILLER_226_1250 ();
 b15zdnd11an1n08x5 FILLER_226_1294 ();
 b15zdnd11an1n04x5 FILLER_226_1302 ();
 b15zdnd00an1n02x5 FILLER_226_1306 ();
 b15zdnd11an1n64x5 FILLER_226_1328 ();
 b15zdnd11an1n64x5 FILLER_226_1392 ();
 b15zdnd11an1n64x5 FILLER_226_1456 ();
 b15zdnd11an1n64x5 FILLER_226_1520 ();
 b15zdnd11an1n64x5 FILLER_226_1584 ();
 b15zdnd11an1n16x5 FILLER_226_1648 ();
 b15zdnd11an1n64x5 FILLER_226_1673 ();
 b15zdnd11an1n64x5 FILLER_226_1737 ();
 b15zdnd11an1n64x5 FILLER_226_1801 ();
 b15zdnd11an1n16x5 FILLER_226_1865 ();
 b15zdnd11an1n08x5 FILLER_226_1881 ();
 b15zdnd11an1n04x5 FILLER_226_1892 ();
 b15zdnd11an1n04x5 FILLER_226_1899 ();
 b15zdnd11an1n64x5 FILLER_226_1906 ();
 b15zdnd11an1n64x5 FILLER_226_1970 ();
 b15zdnd11an1n64x5 FILLER_226_2034 ();
 b15zdnd11an1n32x5 FILLER_226_2098 ();
 b15zdnd11an1n16x5 FILLER_226_2130 ();
 b15zdnd11an1n08x5 FILLER_226_2146 ();
 b15zdnd11an1n64x5 FILLER_226_2162 ();
 b15zdnd11an1n04x5 FILLER_226_2226 ();
 b15zdnd00an1n02x5 FILLER_226_2230 ();
 b15zdnd00an1n02x5 FILLER_226_2274 ();
 b15zdnd11an1n64x5 FILLER_227_0 ();
 b15zdnd11an1n64x5 FILLER_227_64 ();
 b15zdnd11an1n64x5 FILLER_227_128 ();
 b15zdnd11an1n64x5 FILLER_227_192 ();
 b15zdnd11an1n64x5 FILLER_227_256 ();
 b15zdnd11an1n32x5 FILLER_227_320 ();
 b15zdnd11an1n16x5 FILLER_227_352 ();
 b15zdnd11an1n04x5 FILLER_227_368 ();
 b15zdnd00an1n01x5 FILLER_227_372 ();
 b15zdnd11an1n64x5 FILLER_227_415 ();
 b15zdnd11an1n64x5 FILLER_227_479 ();
 b15zdnd11an1n64x5 FILLER_227_543 ();
 b15zdnd11an1n64x5 FILLER_227_607 ();
 b15zdnd11an1n64x5 FILLER_227_671 ();
 b15zdnd11an1n64x5 FILLER_227_735 ();
 b15zdnd11an1n64x5 FILLER_227_799 ();
 b15zdnd11an1n64x5 FILLER_227_863 ();
 b15zdnd11an1n64x5 FILLER_227_927 ();
 b15zdnd11an1n16x5 FILLER_227_991 ();
 b15zdnd00an1n02x5 FILLER_227_1007 ();
 b15zdnd11an1n04x5 FILLER_227_1023 ();
 b15zdnd11an1n32x5 FILLER_227_1069 ();
 b15zdnd11an1n16x5 FILLER_227_1101 ();
 b15zdnd11an1n04x5 FILLER_227_1117 ();
 b15zdnd00an1n02x5 FILLER_227_1121 ();
 b15zdnd00an1n01x5 FILLER_227_1123 ();
 b15zdnd11an1n64x5 FILLER_227_1144 ();
 b15zdnd11an1n64x5 FILLER_227_1208 ();
 b15zdnd11an1n16x5 FILLER_227_1272 ();
 b15zdnd11an1n64x5 FILLER_227_1333 ();
 b15zdnd11an1n64x5 FILLER_227_1397 ();
 b15zdnd11an1n16x5 FILLER_227_1461 ();
 b15zdnd00an1n02x5 FILLER_227_1477 ();
 b15zdnd11an1n64x5 FILLER_227_1483 ();
 b15zdnd11an1n64x5 FILLER_227_1547 ();
 b15zdnd11an1n64x5 FILLER_227_1611 ();
 b15zdnd11an1n64x5 FILLER_227_1675 ();
 b15zdnd11an1n64x5 FILLER_227_1739 ();
 b15zdnd11an1n64x5 FILLER_227_1803 ();
 b15zdnd11an1n64x5 FILLER_227_1867 ();
 b15zdnd11an1n64x5 FILLER_227_1931 ();
 b15zdnd11an1n16x5 FILLER_227_1995 ();
 b15zdnd11an1n04x5 FILLER_227_2011 ();
 b15zdnd11an1n64x5 FILLER_227_2067 ();
 b15zdnd11an1n64x5 FILLER_227_2131 ();
 b15zdnd11an1n04x5 FILLER_227_2195 ();
 b15zdnd00an1n02x5 FILLER_227_2199 ();
 b15zdnd00an1n01x5 FILLER_227_2201 ();
 b15zdnd11an1n04x5 FILLER_227_2247 ();
 b15zdnd11an1n04x5 FILLER_227_2255 ();
 b15zdnd11an1n04x5 FILLER_227_2263 ();
 b15zdnd00an1n02x5 FILLER_227_2267 ();
 b15zdnd00an1n01x5 FILLER_227_2269 ();
 b15zdnd11an1n08x5 FILLER_227_2274 ();
 b15zdnd00an1n02x5 FILLER_227_2282 ();
 b15zdnd11an1n64x5 FILLER_228_8 ();
 b15zdnd11an1n64x5 FILLER_228_72 ();
 b15zdnd11an1n64x5 FILLER_228_136 ();
 b15zdnd11an1n16x5 FILLER_228_200 ();
 b15zdnd11an1n08x5 FILLER_228_216 ();
 b15zdnd00an1n02x5 FILLER_228_224 ();
 b15zdnd00an1n01x5 FILLER_228_226 ();
 b15zdnd11an1n64x5 FILLER_228_269 ();
 b15zdnd11an1n64x5 FILLER_228_333 ();
 b15zdnd11an1n64x5 FILLER_228_397 ();
 b15zdnd11an1n64x5 FILLER_228_461 ();
 b15zdnd11an1n64x5 FILLER_228_525 ();
 b15zdnd11an1n64x5 FILLER_228_589 ();
 b15zdnd11an1n64x5 FILLER_228_653 ();
 b15zdnd00an1n01x5 FILLER_228_717 ();
 b15zdnd11an1n64x5 FILLER_228_726 ();
 b15zdnd11an1n64x5 FILLER_228_790 ();
 b15zdnd11an1n64x5 FILLER_228_854 ();
 b15zdnd11an1n64x5 FILLER_228_918 ();
 b15zdnd11an1n16x5 FILLER_228_982 ();
 b15zdnd11an1n08x5 FILLER_228_998 ();
 b15zdnd00an1n02x5 FILLER_228_1006 ();
 b15zdnd00an1n01x5 FILLER_228_1008 ();
 b15zdnd11an1n04x5 FILLER_228_1012 ();
 b15zdnd00an1n02x5 FILLER_228_1016 ();
 b15zdnd11an1n64x5 FILLER_228_1044 ();
 b15zdnd11an1n08x5 FILLER_228_1108 ();
 b15zdnd11an1n04x5 FILLER_228_1116 ();
 b15zdnd11an1n04x5 FILLER_228_1140 ();
 b15zdnd11an1n64x5 FILLER_228_1155 ();
 b15zdnd11an1n16x5 FILLER_228_1219 ();
 b15zdnd11an1n04x5 FILLER_228_1235 ();
 b15zdnd00an1n02x5 FILLER_228_1239 ();
 b15zdnd11an1n64x5 FILLER_228_1255 ();
 b15zdnd11an1n64x5 FILLER_228_1319 ();
 b15zdnd11an1n64x5 FILLER_228_1383 ();
 b15zdnd11an1n32x5 FILLER_228_1447 ();
 b15zdnd11an1n16x5 FILLER_228_1479 ();
 b15zdnd11an1n04x5 FILLER_228_1495 ();
 b15zdnd11an1n64x5 FILLER_228_1503 ();
 b15zdnd11an1n64x5 FILLER_228_1567 ();
 b15zdnd11an1n64x5 FILLER_228_1631 ();
 b15zdnd11an1n64x5 FILLER_228_1695 ();
 b15zdnd11an1n32x5 FILLER_228_1759 ();
 b15zdnd11an1n16x5 FILLER_228_1791 ();
 b15zdnd11an1n08x5 FILLER_228_1807 ();
 b15zdnd11an1n04x5 FILLER_228_1815 ();
 b15zdnd11an1n64x5 FILLER_228_1834 ();
 b15zdnd11an1n64x5 FILLER_228_1898 ();
 b15zdnd11an1n08x5 FILLER_228_1962 ();
 b15zdnd11an1n32x5 FILLER_228_1982 ();
 b15zdnd11an1n16x5 FILLER_228_2014 ();
 b15zdnd00an1n02x5 FILLER_228_2030 ();
 b15zdnd00an1n01x5 FILLER_228_2032 ();
 b15zdnd11an1n04x5 FILLER_228_2036 ();
 b15zdnd11an1n04x5 FILLER_228_2043 ();
 b15zdnd11an1n04x5 FILLER_228_2050 ();
 b15zdnd11an1n64x5 FILLER_228_2057 ();
 b15zdnd11an1n32x5 FILLER_228_2121 ();
 b15zdnd00an1n01x5 FILLER_228_2153 ();
 b15zdnd11an1n64x5 FILLER_228_2162 ();
 b15zdnd11an1n04x5 FILLER_228_2226 ();
 b15zdnd00an1n02x5 FILLER_228_2230 ();
 b15zdnd00an1n02x5 FILLER_228_2274 ();
 b15zdnd11an1n64x5 FILLER_229_0 ();
 b15zdnd11an1n64x5 FILLER_229_64 ();
 b15zdnd11an1n64x5 FILLER_229_128 ();
 b15zdnd11an1n32x5 FILLER_229_192 ();
 b15zdnd11an1n64x5 FILLER_229_266 ();
 b15zdnd11an1n64x5 FILLER_229_330 ();
 b15zdnd11an1n64x5 FILLER_229_394 ();
 b15zdnd11an1n64x5 FILLER_229_458 ();
 b15zdnd11an1n64x5 FILLER_229_522 ();
 b15zdnd11an1n64x5 FILLER_229_586 ();
 b15zdnd11an1n64x5 FILLER_229_650 ();
 b15zdnd11an1n64x5 FILLER_229_714 ();
 b15zdnd11an1n64x5 FILLER_229_778 ();
 b15zdnd11an1n16x5 FILLER_229_842 ();
 b15zdnd11an1n08x5 FILLER_229_858 ();
 b15zdnd11an1n04x5 FILLER_229_866 ();
 b15zdnd00an1n02x5 FILLER_229_870 ();
 b15zdnd00an1n01x5 FILLER_229_872 ();
 b15zdnd11an1n64x5 FILLER_229_889 ();
 b15zdnd11an1n32x5 FILLER_229_953 ();
 b15zdnd11an1n16x5 FILLER_229_985 ();
 b15zdnd11an1n08x5 FILLER_229_1001 ();
 b15zdnd00an1n02x5 FILLER_229_1009 ();
 b15zdnd11an1n04x5 FILLER_229_1021 ();
 b15zdnd00an1n01x5 FILLER_229_1025 ();
 b15zdnd11an1n04x5 FILLER_229_1042 ();
 b15zdnd00an1n02x5 FILLER_229_1046 ();
 b15zdnd11an1n64x5 FILLER_229_1068 ();
 b15zdnd11an1n64x5 FILLER_229_1132 ();
 b15zdnd11an1n32x5 FILLER_229_1196 ();
 b15zdnd11an1n16x5 FILLER_229_1228 ();
 b15zdnd00an1n01x5 FILLER_229_1244 ();
 b15zdnd11an1n32x5 FILLER_229_1259 ();
 b15zdnd11an1n04x5 FILLER_229_1291 ();
 b15zdnd11an1n64x5 FILLER_229_1299 ();
 b15zdnd11an1n64x5 FILLER_229_1363 ();
 b15zdnd11an1n64x5 FILLER_229_1427 ();
 b15zdnd11an1n64x5 FILLER_229_1491 ();
 b15zdnd11an1n64x5 FILLER_229_1555 ();
 b15zdnd11an1n64x5 FILLER_229_1619 ();
 b15zdnd11an1n64x5 FILLER_229_1683 ();
 b15zdnd11an1n64x5 FILLER_229_1747 ();
 b15zdnd11an1n64x5 FILLER_229_1811 ();
 b15zdnd11an1n64x5 FILLER_229_1875 ();
 b15zdnd11an1n16x5 FILLER_229_1939 ();
 b15zdnd11an1n08x5 FILLER_229_1955 ();
 b15zdnd11an1n04x5 FILLER_229_1963 ();
 b15zdnd00an1n02x5 FILLER_229_1967 ();
 b15zdnd00an1n01x5 FILLER_229_1969 ();
 b15zdnd11an1n32x5 FILLER_229_1990 ();
 b15zdnd11an1n04x5 FILLER_229_2022 ();
 b15zdnd11an1n04x5 FILLER_229_2078 ();
 b15zdnd11an1n64x5 FILLER_229_2089 ();
 b15zdnd11an1n08x5 FILLER_229_2153 ();
 b15zdnd00an1n01x5 FILLER_229_2161 ();
 b15zdnd11an1n32x5 FILLER_229_2204 ();
 b15zdnd11an1n04x5 FILLER_229_2236 ();
 b15zdnd00an1n02x5 FILLER_229_2282 ();
 b15zdnd11an1n64x5 FILLER_230_8 ();
 b15zdnd11an1n64x5 FILLER_230_72 ();
 b15zdnd11an1n64x5 FILLER_230_136 ();
 b15zdnd11an1n64x5 FILLER_230_200 ();
 b15zdnd11an1n64x5 FILLER_230_264 ();
 b15zdnd11an1n64x5 FILLER_230_328 ();
 b15zdnd11an1n64x5 FILLER_230_392 ();
 b15zdnd11an1n64x5 FILLER_230_456 ();
 b15zdnd11an1n64x5 FILLER_230_520 ();
 b15zdnd11an1n64x5 FILLER_230_584 ();
 b15zdnd11an1n64x5 FILLER_230_648 ();
 b15zdnd11an1n04x5 FILLER_230_712 ();
 b15zdnd00an1n02x5 FILLER_230_716 ();
 b15zdnd11an1n64x5 FILLER_230_726 ();
 b15zdnd11an1n08x5 FILLER_230_790 ();
 b15zdnd11an1n16x5 FILLER_230_809 ();
 b15zdnd00an1n02x5 FILLER_230_825 ();
 b15zdnd00an1n01x5 FILLER_230_827 ();
 b15zdnd11an1n32x5 FILLER_230_844 ();
 b15zdnd00an1n01x5 FILLER_230_876 ();
 b15zdnd11an1n04x5 FILLER_230_886 ();
 b15zdnd11an1n64x5 FILLER_230_916 ();
 b15zdnd11an1n16x5 FILLER_230_980 ();
 b15zdnd11an1n08x5 FILLER_230_996 ();
 b15zdnd11an1n04x5 FILLER_230_1004 ();
 b15zdnd00an1n01x5 FILLER_230_1008 ();
 b15zdnd11an1n08x5 FILLER_230_1022 ();
 b15zdnd11an1n04x5 FILLER_230_1030 ();
 b15zdnd11an1n04x5 FILLER_230_1058 ();
 b15zdnd11an1n64x5 FILLER_230_1076 ();
 b15zdnd11an1n64x5 FILLER_230_1140 ();
 b15zdnd11an1n64x5 FILLER_230_1204 ();
 b15zdnd11an1n64x5 FILLER_230_1268 ();
 b15zdnd11an1n64x5 FILLER_230_1332 ();
 b15zdnd11an1n64x5 FILLER_230_1396 ();
 b15zdnd11an1n64x5 FILLER_230_1460 ();
 b15zdnd11an1n64x5 FILLER_230_1524 ();
 b15zdnd11an1n64x5 FILLER_230_1588 ();
 b15zdnd00an1n02x5 FILLER_230_1652 ();
 b15zdnd00an1n01x5 FILLER_230_1654 ();
 b15zdnd11an1n64x5 FILLER_230_1664 ();
 b15zdnd11an1n32x5 FILLER_230_1728 ();
 b15zdnd11an1n08x5 FILLER_230_1760 ();
 b15zdnd11an1n64x5 FILLER_230_1786 ();
 b15zdnd11an1n64x5 FILLER_230_1850 ();
 b15zdnd11an1n64x5 FILLER_230_1914 ();
 b15zdnd11an1n16x5 FILLER_230_1978 ();
 b15zdnd11an1n04x5 FILLER_230_1994 ();
 b15zdnd00an1n02x5 FILLER_230_1998 ();
 b15zdnd11an1n32x5 FILLER_230_2007 ();
 b15zdnd11an1n04x5 FILLER_230_2039 ();
 b15zdnd00an1n01x5 FILLER_230_2043 ();
 b15zdnd11an1n08x5 FILLER_230_2047 ();
 b15zdnd00an1n02x5 FILLER_230_2055 ();
 b15zdnd11an1n04x5 FILLER_230_2064 ();
 b15zdnd11an1n64x5 FILLER_230_2071 ();
 b15zdnd11an1n16x5 FILLER_230_2135 ();
 b15zdnd00an1n02x5 FILLER_230_2151 ();
 b15zdnd00an1n01x5 FILLER_230_2153 ();
 b15zdnd11an1n64x5 FILLER_230_2162 ();
 b15zdnd11an1n32x5 FILLER_230_2226 ();
 b15zdnd11an1n16x5 FILLER_230_2258 ();
 b15zdnd00an1n02x5 FILLER_230_2274 ();
 b15zdnd11an1n64x5 FILLER_231_0 ();
 b15zdnd11an1n64x5 FILLER_231_64 ();
 b15zdnd11an1n64x5 FILLER_231_128 ();
 b15zdnd11an1n64x5 FILLER_231_192 ();
 b15zdnd11an1n64x5 FILLER_231_256 ();
 b15zdnd11an1n64x5 FILLER_231_320 ();
 b15zdnd11an1n64x5 FILLER_231_384 ();
 b15zdnd11an1n64x5 FILLER_231_448 ();
 b15zdnd00an1n02x5 FILLER_231_512 ();
 b15zdnd11an1n08x5 FILLER_231_517 ();
 b15zdnd11an1n04x5 FILLER_231_525 ();
 b15zdnd00an1n02x5 FILLER_231_529 ();
 b15zdnd11an1n64x5 FILLER_231_552 ();
 b15zdnd11an1n64x5 FILLER_231_616 ();
 b15zdnd11an1n64x5 FILLER_231_680 ();
 b15zdnd11an1n32x5 FILLER_231_744 ();
 b15zdnd11an1n16x5 FILLER_231_776 ();
 b15zdnd11an1n04x5 FILLER_231_792 ();
 b15zdnd11an1n04x5 FILLER_231_806 ();
 b15zdnd11an1n16x5 FILLER_231_814 ();
 b15zdnd00an1n02x5 FILLER_231_830 ();
 b15zdnd11an1n64x5 FILLER_231_845 ();
 b15zdnd11an1n64x5 FILLER_231_918 ();
 b15zdnd11an1n64x5 FILLER_231_982 ();
 b15zdnd11an1n64x5 FILLER_231_1046 ();
 b15zdnd11an1n08x5 FILLER_231_1110 ();
 b15zdnd11an1n04x5 FILLER_231_1118 ();
 b15zdnd11an1n08x5 FILLER_231_1136 ();
 b15zdnd11an1n04x5 FILLER_231_1144 ();
 b15zdnd11an1n04x5 FILLER_231_1154 ();
 b15zdnd00an1n02x5 FILLER_231_1158 ();
 b15zdnd11an1n64x5 FILLER_231_1171 ();
 b15zdnd11an1n64x5 FILLER_231_1235 ();
 b15zdnd11an1n64x5 FILLER_231_1299 ();
 b15zdnd11an1n64x5 FILLER_231_1363 ();
 b15zdnd11an1n64x5 FILLER_231_1427 ();
 b15zdnd11an1n32x5 FILLER_231_1491 ();
 b15zdnd11an1n08x5 FILLER_231_1523 ();
 b15zdnd11an1n64x5 FILLER_231_1539 ();
 b15zdnd11an1n64x5 FILLER_231_1603 ();
 b15zdnd11an1n64x5 FILLER_231_1667 ();
 b15zdnd11an1n64x5 FILLER_231_1731 ();
 b15zdnd11an1n64x5 FILLER_231_1795 ();
 b15zdnd11an1n64x5 FILLER_231_1859 ();
 b15zdnd11an1n32x5 FILLER_231_1923 ();
 b15zdnd11an1n16x5 FILLER_231_1972 ();
 b15zdnd11an1n32x5 FILLER_231_1994 ();
 b15zdnd11an1n16x5 FILLER_231_2026 ();
 b15zdnd00an1n02x5 FILLER_231_2042 ();
 b15zdnd11an1n16x5 FILLER_231_2086 ();
 b15zdnd00an1n01x5 FILLER_231_2102 ();
 b15zdnd11an1n64x5 FILLER_231_2117 ();
 b15zdnd11an1n64x5 FILLER_231_2181 ();
 b15zdnd11an1n32x5 FILLER_231_2245 ();
 b15zdnd11an1n04x5 FILLER_231_2277 ();
 b15zdnd00an1n02x5 FILLER_231_2281 ();
 b15zdnd00an1n01x5 FILLER_231_2283 ();
 b15zdnd11an1n64x5 FILLER_232_8 ();
 b15zdnd11an1n64x5 FILLER_232_72 ();
 b15zdnd11an1n64x5 FILLER_232_136 ();
 b15zdnd11an1n64x5 FILLER_232_200 ();
 b15zdnd11an1n64x5 FILLER_232_264 ();
 b15zdnd11an1n32x5 FILLER_232_328 ();
 b15zdnd11an1n08x5 FILLER_232_360 ();
 b15zdnd00an1n02x5 FILLER_232_368 ();
 b15zdnd11an1n64x5 FILLER_232_373 ();
 b15zdnd11an1n64x5 FILLER_232_437 ();
 b15zdnd11an1n32x5 FILLER_232_501 ();
 b15zdnd11an1n08x5 FILLER_232_533 ();
 b15zdnd11an1n04x5 FILLER_232_541 ();
 b15zdnd00an1n01x5 FILLER_232_545 ();
 b15zdnd11an1n64x5 FILLER_232_550 ();
 b15zdnd11an1n64x5 FILLER_232_614 ();
 b15zdnd11an1n32x5 FILLER_232_678 ();
 b15zdnd11an1n08x5 FILLER_232_710 ();
 b15zdnd11an1n64x5 FILLER_232_726 ();
 b15zdnd11an1n64x5 FILLER_232_790 ();
 b15zdnd11an1n64x5 FILLER_232_854 ();
 b15zdnd11an1n32x5 FILLER_232_918 ();
 b15zdnd11an1n04x5 FILLER_232_950 ();
 b15zdnd00an1n01x5 FILLER_232_954 ();
 b15zdnd11an1n32x5 FILLER_232_965 ();
 b15zdnd11an1n04x5 FILLER_232_997 ();
 b15zdnd00an1n02x5 FILLER_232_1001 ();
 b15zdnd11an1n16x5 FILLER_232_1017 ();
 b15zdnd11an1n08x5 FILLER_232_1033 ();
 b15zdnd00an1n02x5 FILLER_232_1041 ();
 b15zdnd11an1n16x5 FILLER_232_1057 ();
 b15zdnd11an1n04x5 FILLER_232_1073 ();
 b15zdnd00an1n01x5 FILLER_232_1077 ();
 b15zdnd11an1n64x5 FILLER_232_1098 ();
 b15zdnd11an1n64x5 FILLER_232_1162 ();
 b15zdnd11an1n64x5 FILLER_232_1226 ();
 b15zdnd11an1n64x5 FILLER_232_1290 ();
 b15zdnd11an1n64x5 FILLER_232_1354 ();
 b15zdnd11an1n64x5 FILLER_232_1418 ();
 b15zdnd11an1n64x5 FILLER_232_1482 ();
 b15zdnd11an1n64x5 FILLER_232_1546 ();
 b15zdnd11an1n64x5 FILLER_232_1610 ();
 b15zdnd11an1n64x5 FILLER_232_1674 ();
 b15zdnd11an1n64x5 FILLER_232_1738 ();
 b15zdnd11an1n64x5 FILLER_232_1802 ();
 b15zdnd11an1n64x5 FILLER_232_1866 ();
 b15zdnd11an1n32x5 FILLER_232_1930 ();
 b15zdnd11an1n08x5 FILLER_232_1962 ();
 b15zdnd11an1n04x5 FILLER_232_1970 ();
 b15zdnd00an1n01x5 FILLER_232_1974 ();
 b15zdnd11an1n64x5 FILLER_232_1989 ();
 b15zdnd11an1n32x5 FILLER_232_2053 ();
 b15zdnd11an1n16x5 FILLER_232_2085 ();
 b15zdnd11an1n08x5 FILLER_232_2101 ();
 b15zdnd00an1n02x5 FILLER_232_2109 ();
 b15zdnd00an1n01x5 FILLER_232_2111 ();
 b15zdnd11an1n32x5 FILLER_232_2119 ();
 b15zdnd00an1n02x5 FILLER_232_2151 ();
 b15zdnd00an1n01x5 FILLER_232_2153 ();
 b15zdnd11an1n64x5 FILLER_232_2162 ();
 b15zdnd11an1n32x5 FILLER_232_2226 ();
 b15zdnd11an1n16x5 FILLER_232_2258 ();
 b15zdnd00an1n02x5 FILLER_232_2274 ();
 b15zdnd11an1n64x5 FILLER_233_0 ();
 b15zdnd11an1n64x5 FILLER_233_64 ();
 b15zdnd11an1n64x5 FILLER_233_128 ();
 b15zdnd11an1n64x5 FILLER_233_192 ();
 b15zdnd11an1n64x5 FILLER_233_256 ();
 b15zdnd11an1n16x5 FILLER_233_320 ();
 b15zdnd11an1n04x5 FILLER_233_336 ();
 b15zdnd00an1n02x5 FILLER_233_340 ();
 b15zdnd00an1n01x5 FILLER_233_342 ();
 b15zdnd11an1n64x5 FILLER_233_395 ();
 b15zdnd11an1n64x5 FILLER_233_459 ();
 b15zdnd11an1n64x5 FILLER_233_523 ();
 b15zdnd11an1n64x5 FILLER_233_587 ();
 b15zdnd11an1n64x5 FILLER_233_651 ();
 b15zdnd11an1n16x5 FILLER_233_715 ();
 b15zdnd00an1n02x5 FILLER_233_731 ();
 b15zdnd00an1n01x5 FILLER_233_733 ();
 b15zdnd11an1n64x5 FILLER_233_752 ();
 b15zdnd11an1n08x5 FILLER_233_816 ();
 b15zdnd11an1n04x5 FILLER_233_824 ();
 b15zdnd00an1n02x5 FILLER_233_828 ();
 b15zdnd00an1n01x5 FILLER_233_830 ();
 b15zdnd11an1n16x5 FILLER_233_841 ();
 b15zdnd11an1n08x5 FILLER_233_857 ();
 b15zdnd11an1n64x5 FILLER_233_868 ();
 b15zdnd11an1n64x5 FILLER_233_932 ();
 b15zdnd11an1n32x5 FILLER_233_996 ();
 b15zdnd11an1n16x5 FILLER_233_1028 ();
 b15zdnd11an1n04x5 FILLER_233_1044 ();
 b15zdnd00an1n01x5 FILLER_233_1048 ();
 b15zdnd11an1n16x5 FILLER_233_1056 ();
 b15zdnd11an1n04x5 FILLER_233_1072 ();
 b15zdnd00an1n01x5 FILLER_233_1076 ();
 b15zdnd11an1n64x5 FILLER_233_1088 ();
 b15zdnd11an1n08x5 FILLER_233_1152 ();
 b15zdnd11an1n04x5 FILLER_233_1160 ();
 b15zdnd11an1n04x5 FILLER_233_1190 ();
 b15zdnd00an1n02x5 FILLER_233_1194 ();
 b15zdnd00an1n01x5 FILLER_233_1196 ();
 b15zdnd11an1n08x5 FILLER_233_1217 ();
 b15zdnd00an1n02x5 FILLER_233_1225 ();
 b15zdnd00an1n01x5 FILLER_233_1227 ();
 b15zdnd11an1n04x5 FILLER_233_1236 ();
 b15zdnd11an1n32x5 FILLER_233_1260 ();
 b15zdnd11an1n64x5 FILLER_233_1312 ();
 b15zdnd11an1n64x5 FILLER_233_1376 ();
 b15zdnd11an1n64x5 FILLER_233_1440 ();
 b15zdnd11an1n08x5 FILLER_233_1504 ();
 b15zdnd00an1n02x5 FILLER_233_1512 ();
 b15zdnd11an1n64x5 FILLER_233_1518 ();
 b15zdnd11an1n64x5 FILLER_233_1582 ();
 b15zdnd11an1n64x5 FILLER_233_1646 ();
 b15zdnd11an1n64x5 FILLER_233_1710 ();
 b15zdnd11an1n16x5 FILLER_233_1774 ();
 b15zdnd11an1n08x5 FILLER_233_1790 ();
 b15zdnd00an1n02x5 FILLER_233_1798 ();
 b15zdnd11an1n32x5 FILLER_233_1815 ();
 b15zdnd11an1n16x5 FILLER_233_1847 ();
 b15zdnd11an1n08x5 FILLER_233_1863 ();
 b15zdnd00an1n02x5 FILLER_233_1871 ();
 b15zdnd11an1n04x5 FILLER_233_1884 ();
 b15zdnd11an1n64x5 FILLER_233_1898 ();
 b15zdnd11an1n64x5 FILLER_233_1962 ();
 b15zdnd11an1n64x5 FILLER_233_2026 ();
 b15zdnd11an1n64x5 FILLER_233_2090 ();
 b15zdnd11an1n64x5 FILLER_233_2154 ();
 b15zdnd11an1n64x5 FILLER_233_2218 ();
 b15zdnd00an1n02x5 FILLER_233_2282 ();
 b15zdnd11an1n64x5 FILLER_234_8 ();
 b15zdnd11an1n64x5 FILLER_234_72 ();
 b15zdnd11an1n64x5 FILLER_234_136 ();
 b15zdnd11an1n64x5 FILLER_234_200 ();
 b15zdnd11an1n32x5 FILLER_234_264 ();
 b15zdnd11an1n16x5 FILLER_234_296 ();
 b15zdnd11an1n08x5 FILLER_234_312 ();
 b15zdnd11an1n04x5 FILLER_234_323 ();
 b15zdnd11an1n04x5 FILLER_234_330 ();
 b15zdnd11an1n16x5 FILLER_234_337 ();
 b15zdnd11an1n04x5 FILLER_234_353 ();
 b15zdnd00an1n02x5 FILLER_234_357 ();
 b15zdnd11an1n64x5 FILLER_234_401 ();
 b15zdnd11an1n64x5 FILLER_234_465 ();
 b15zdnd11an1n64x5 FILLER_234_529 ();
 b15zdnd11an1n64x5 FILLER_234_593 ();
 b15zdnd11an1n32x5 FILLER_234_657 ();
 b15zdnd00an1n01x5 FILLER_234_689 ();
 b15zdnd11an1n16x5 FILLER_234_697 ();
 b15zdnd11an1n04x5 FILLER_234_713 ();
 b15zdnd00an1n01x5 FILLER_234_717 ();
 b15zdnd11an1n64x5 FILLER_234_726 ();
 b15zdnd11an1n32x5 FILLER_234_790 ();
 b15zdnd11an1n08x5 FILLER_234_822 ();
 b15zdnd00an1n01x5 FILLER_234_830 ();
 b15zdnd11an1n32x5 FILLER_234_834 ();
 b15zdnd00an1n02x5 FILLER_234_866 ();
 b15zdnd00an1n01x5 FILLER_234_868 ();
 b15zdnd11an1n64x5 FILLER_234_879 ();
 b15zdnd11an1n64x5 FILLER_234_943 ();
 b15zdnd11an1n16x5 FILLER_234_1007 ();
 b15zdnd11an1n08x5 FILLER_234_1023 ();
 b15zdnd11an1n04x5 FILLER_234_1031 ();
 b15zdnd00an1n01x5 FILLER_234_1035 ();
 b15zdnd11an1n64x5 FILLER_234_1056 ();
 b15zdnd11an1n32x5 FILLER_234_1120 ();
 b15zdnd11an1n08x5 FILLER_234_1152 ();
 b15zdnd11an1n04x5 FILLER_234_1160 ();
 b15zdnd11an1n32x5 FILLER_234_1171 ();
 b15zdnd11an1n04x5 FILLER_234_1203 ();
 b15zdnd11an1n04x5 FILLER_234_1221 ();
 b15zdnd11an1n16x5 FILLER_234_1245 ();
 b15zdnd11an1n04x5 FILLER_234_1261 ();
 b15zdnd00an1n02x5 FILLER_234_1265 ();
 b15zdnd11an1n16x5 FILLER_234_1281 ();
 b15zdnd11an1n64x5 FILLER_234_1307 ();
 b15zdnd11an1n64x5 FILLER_234_1371 ();
 b15zdnd11an1n64x5 FILLER_234_1435 ();
 b15zdnd11an1n64x5 FILLER_234_1499 ();
 b15zdnd11an1n64x5 FILLER_234_1563 ();
 b15zdnd11an1n64x5 FILLER_234_1627 ();
 b15zdnd11an1n64x5 FILLER_234_1691 ();
 b15zdnd11an1n32x5 FILLER_234_1755 ();
 b15zdnd11an1n16x5 FILLER_234_1787 ();
 b15zdnd11an1n08x5 FILLER_234_1803 ();
 b15zdnd00an1n02x5 FILLER_234_1811 ();
 b15zdnd00an1n01x5 FILLER_234_1813 ();
 b15zdnd11an1n32x5 FILLER_234_1832 ();
 b15zdnd11an1n16x5 FILLER_234_1864 ();
 b15zdnd11an1n08x5 FILLER_234_1880 ();
 b15zdnd11an1n04x5 FILLER_234_1888 ();
 b15zdnd00an1n02x5 FILLER_234_1892 ();
 b15zdnd11an1n64x5 FILLER_234_1898 ();
 b15zdnd11an1n64x5 FILLER_234_1962 ();
 b15zdnd11an1n64x5 FILLER_234_2026 ();
 b15zdnd11an1n64x5 FILLER_234_2090 ();
 b15zdnd11an1n32x5 FILLER_234_2162 ();
 b15zdnd11an1n08x5 FILLER_234_2194 ();
 b15zdnd11an1n04x5 FILLER_234_2202 ();
 b15zdnd11an1n32x5 FILLER_234_2213 ();
 b15zdnd11an1n16x5 FILLER_234_2245 ();
 b15zdnd11an1n08x5 FILLER_234_2261 ();
 b15zdnd11an1n04x5 FILLER_234_2269 ();
 b15zdnd00an1n02x5 FILLER_234_2273 ();
 b15zdnd00an1n01x5 FILLER_234_2275 ();
 b15zdnd11an1n64x5 FILLER_235_0 ();
 b15zdnd11an1n64x5 FILLER_235_64 ();
 b15zdnd11an1n64x5 FILLER_235_128 ();
 b15zdnd11an1n16x5 FILLER_235_192 ();
 b15zdnd11an1n08x5 FILLER_235_208 ();
 b15zdnd00an1n01x5 FILLER_235_216 ();
 b15zdnd11an1n64x5 FILLER_235_220 ();
 b15zdnd11an1n16x5 FILLER_235_284 ();
 b15zdnd11an1n08x5 FILLER_235_352 ();
 b15zdnd00an1n01x5 FILLER_235_360 ();
 b15zdnd11an1n04x5 FILLER_235_364 ();
 b15zdnd11an1n64x5 FILLER_235_371 ();
 b15zdnd11an1n64x5 FILLER_235_435 ();
 b15zdnd11an1n64x5 FILLER_235_499 ();
 b15zdnd11an1n64x5 FILLER_235_563 ();
 b15zdnd11an1n64x5 FILLER_235_627 ();
 b15zdnd11an1n64x5 FILLER_235_691 ();
 b15zdnd11an1n64x5 FILLER_235_755 ();
 b15zdnd11an1n64x5 FILLER_235_819 ();
 b15zdnd11an1n64x5 FILLER_235_883 ();
 b15zdnd11an1n64x5 FILLER_235_947 ();
 b15zdnd11an1n16x5 FILLER_235_1011 ();
 b15zdnd11an1n04x5 FILLER_235_1027 ();
 b15zdnd00an1n02x5 FILLER_235_1031 ();
 b15zdnd00an1n01x5 FILLER_235_1033 ();
 b15zdnd11an1n04x5 FILLER_235_1054 ();
 b15zdnd11an1n64x5 FILLER_235_1072 ();
 b15zdnd11an1n32x5 FILLER_235_1136 ();
 b15zdnd11an1n16x5 FILLER_235_1168 ();
 b15zdnd11an1n08x5 FILLER_235_1184 ();
 b15zdnd00an1n02x5 FILLER_235_1192 ();
 b15zdnd00an1n01x5 FILLER_235_1194 ();
 b15zdnd11an1n64x5 FILLER_235_1209 ();
 b15zdnd11an1n64x5 FILLER_235_1273 ();
 b15zdnd11an1n64x5 FILLER_235_1337 ();
 b15zdnd11an1n64x5 FILLER_235_1401 ();
 b15zdnd11an1n64x5 FILLER_235_1465 ();
 b15zdnd11an1n64x5 FILLER_235_1529 ();
 b15zdnd11an1n64x5 FILLER_235_1593 ();
 b15zdnd11an1n64x5 FILLER_235_1657 ();
 b15zdnd11an1n64x5 FILLER_235_1721 ();
 b15zdnd11an1n64x5 FILLER_235_1785 ();
 b15zdnd11an1n64x5 FILLER_235_1849 ();
 b15zdnd11an1n04x5 FILLER_235_1913 ();
 b15zdnd11an1n32x5 FILLER_235_1923 ();
 b15zdnd11an1n16x5 FILLER_235_1955 ();
 b15zdnd11an1n08x5 FILLER_235_1971 ();
 b15zdnd11an1n04x5 FILLER_235_1979 ();
 b15zdnd00an1n02x5 FILLER_235_1983 ();
 b15zdnd00an1n01x5 FILLER_235_1985 ();
 b15zdnd11an1n32x5 FILLER_235_1993 ();
 b15zdnd11an1n16x5 FILLER_235_2025 ();
 b15zdnd11an1n04x5 FILLER_235_2041 ();
 b15zdnd00an1n02x5 FILLER_235_2045 ();
 b15zdnd00an1n01x5 FILLER_235_2047 ();
 b15zdnd11an1n64x5 FILLER_235_2053 ();
 b15zdnd11an1n64x5 FILLER_235_2117 ();
 b15zdnd11an1n04x5 FILLER_235_2181 ();
 b15zdnd00an1n01x5 FILLER_235_2185 ();
 b15zdnd11an1n64x5 FILLER_235_2211 ();
 b15zdnd11an1n08x5 FILLER_235_2275 ();
 b15zdnd00an1n01x5 FILLER_235_2283 ();
 b15zdnd11an1n64x5 FILLER_236_8 ();
 b15zdnd11an1n64x5 FILLER_236_72 ();
 b15zdnd11an1n32x5 FILLER_236_136 ();
 b15zdnd11an1n16x5 FILLER_236_168 ();
 b15zdnd11an1n04x5 FILLER_236_184 ();
 b15zdnd00an1n02x5 FILLER_236_188 ();
 b15zdnd11an1n64x5 FILLER_236_242 ();
 b15zdnd11an1n32x5 FILLER_236_306 ();
 b15zdnd11an1n08x5 FILLER_236_338 ();
 b15zdnd11an1n04x5 FILLER_236_346 ();
 b15zdnd11an1n64x5 FILLER_236_392 ();
 b15zdnd11an1n64x5 FILLER_236_456 ();
 b15zdnd11an1n64x5 FILLER_236_520 ();
 b15zdnd11an1n64x5 FILLER_236_584 ();
 b15zdnd11an1n64x5 FILLER_236_648 ();
 b15zdnd11an1n04x5 FILLER_236_712 ();
 b15zdnd00an1n02x5 FILLER_236_716 ();
 b15zdnd11an1n64x5 FILLER_236_726 ();
 b15zdnd11an1n64x5 FILLER_236_790 ();
 b15zdnd11an1n08x5 FILLER_236_854 ();
 b15zdnd11an1n04x5 FILLER_236_862 ();
 b15zdnd00an1n01x5 FILLER_236_866 ();
 b15zdnd11an1n32x5 FILLER_236_898 ();
 b15zdnd11an1n08x5 FILLER_236_930 ();
 b15zdnd11an1n04x5 FILLER_236_938 ();
 b15zdnd00an1n02x5 FILLER_236_942 ();
 b15zdnd11an1n64x5 FILLER_236_947 ();
 b15zdnd11an1n08x5 FILLER_236_1011 ();
 b15zdnd11an1n64x5 FILLER_236_1022 ();
 b15zdnd11an1n64x5 FILLER_236_1086 ();
 b15zdnd11an1n08x5 FILLER_236_1150 ();
 b15zdnd00an1n02x5 FILLER_236_1158 ();
 b15zdnd11an1n64x5 FILLER_236_1171 ();
 b15zdnd11an1n64x5 FILLER_236_1235 ();
 b15zdnd11an1n64x5 FILLER_236_1299 ();
 b15zdnd11an1n64x5 FILLER_236_1363 ();
 b15zdnd11an1n16x5 FILLER_236_1427 ();
 b15zdnd11an1n04x5 FILLER_236_1443 ();
 b15zdnd00an1n02x5 FILLER_236_1447 ();
 b15zdnd00an1n01x5 FILLER_236_1449 ();
 b15zdnd11an1n04x5 FILLER_236_1457 ();
 b15zdnd00an1n02x5 FILLER_236_1461 ();
 b15zdnd11an1n64x5 FILLER_236_1466 ();
 b15zdnd11an1n64x5 FILLER_236_1530 ();
 b15zdnd11an1n32x5 FILLER_236_1594 ();
 b15zdnd11an1n16x5 FILLER_236_1626 ();
 b15zdnd11an1n04x5 FILLER_236_1642 ();
 b15zdnd00an1n02x5 FILLER_236_1646 ();
 b15zdnd11an1n64x5 FILLER_236_1700 ();
 b15zdnd11an1n64x5 FILLER_236_1764 ();
 b15zdnd11an1n32x5 FILLER_236_1828 ();
 b15zdnd11an1n08x5 FILLER_236_1860 ();
 b15zdnd11an1n04x5 FILLER_236_1868 ();
 b15zdnd00an1n02x5 FILLER_236_1872 ();
 b15zdnd00an1n01x5 FILLER_236_1874 ();
 b15zdnd11an1n08x5 FILLER_236_1917 ();
 b15zdnd00an1n02x5 FILLER_236_1925 ();
 b15zdnd11an1n64x5 FILLER_236_1954 ();
 b15zdnd11an1n64x5 FILLER_236_2018 ();
 b15zdnd11an1n64x5 FILLER_236_2082 ();
 b15zdnd11an1n08x5 FILLER_236_2146 ();
 b15zdnd11an1n64x5 FILLER_236_2162 ();
 b15zdnd11an1n32x5 FILLER_236_2226 ();
 b15zdnd11an1n16x5 FILLER_236_2258 ();
 b15zdnd00an1n02x5 FILLER_236_2274 ();
 b15zdnd11an1n64x5 FILLER_237_0 ();
 b15zdnd11an1n64x5 FILLER_237_64 ();
 b15zdnd11an1n64x5 FILLER_237_128 ();
 b15zdnd11an1n16x5 FILLER_237_192 ();
 b15zdnd11an1n04x5 FILLER_237_211 ();
 b15zdnd11an1n64x5 FILLER_237_218 ();
 b15zdnd11an1n32x5 FILLER_237_282 ();
 b15zdnd11an1n16x5 FILLER_237_314 ();
 b15zdnd00an1n01x5 FILLER_237_330 ();
 b15zdnd11an1n64x5 FILLER_237_362 ();
 b15zdnd11an1n64x5 FILLER_237_426 ();
 b15zdnd11an1n64x5 FILLER_237_490 ();
 b15zdnd11an1n16x5 FILLER_237_554 ();
 b15zdnd11an1n08x5 FILLER_237_570 ();
 b15zdnd11an1n64x5 FILLER_237_605 ();
 b15zdnd11an1n64x5 FILLER_237_669 ();
 b15zdnd11an1n64x5 FILLER_237_733 ();
 b15zdnd11an1n04x5 FILLER_237_797 ();
 b15zdnd00an1n02x5 FILLER_237_801 ();
 b15zdnd11an1n04x5 FILLER_237_823 ();
 b15zdnd11an1n16x5 FILLER_237_841 ();
 b15zdnd00an1n01x5 FILLER_237_857 ();
 b15zdnd11an1n04x5 FILLER_237_878 ();
 b15zdnd11an1n16x5 FILLER_237_900 ();
 b15zdnd00an1n01x5 FILLER_237_916 ();
 b15zdnd11an1n64x5 FILLER_237_969 ();
 b15zdnd11an1n64x5 FILLER_237_1033 ();
 b15zdnd11an1n32x5 FILLER_237_1097 ();
 b15zdnd11an1n16x5 FILLER_237_1129 ();
 b15zdnd00an1n02x5 FILLER_237_1145 ();
 b15zdnd11an1n16x5 FILLER_237_1154 ();
 b15zdnd11an1n08x5 FILLER_237_1170 ();
 b15zdnd11an1n04x5 FILLER_237_1178 ();
 b15zdnd11an1n64x5 FILLER_237_1193 ();
 b15zdnd11an1n64x5 FILLER_237_1257 ();
 b15zdnd11an1n64x5 FILLER_237_1321 ();
 b15zdnd11an1n32x5 FILLER_237_1385 ();
 b15zdnd11an1n16x5 FILLER_237_1417 ();
 b15zdnd11an1n04x5 FILLER_237_1433 ();
 b15zdnd00an1n01x5 FILLER_237_1437 ();
 b15zdnd11an1n32x5 FILLER_237_1490 ();
 b15zdnd11an1n16x5 FILLER_237_1522 ();
 b15zdnd11an1n08x5 FILLER_237_1538 ();
 b15zdnd11an1n04x5 FILLER_237_1546 ();
 b15zdnd00an1n02x5 FILLER_237_1550 ();
 b15zdnd11an1n64x5 FILLER_237_1560 ();
 b15zdnd11an1n16x5 FILLER_237_1624 ();
 b15zdnd11an1n08x5 FILLER_237_1640 ();
 b15zdnd11an1n04x5 FILLER_237_1648 ();
 b15zdnd00an1n02x5 FILLER_237_1652 ();
 b15zdnd11an1n64x5 FILLER_237_1706 ();
 b15zdnd11an1n64x5 FILLER_237_1770 ();
 b15zdnd11an1n64x5 FILLER_237_1834 ();
 b15zdnd11an1n04x5 FILLER_237_1898 ();
 b15zdnd11an1n16x5 FILLER_237_1905 ();
 b15zdnd11an1n08x5 FILLER_237_1921 ();
 b15zdnd11an1n04x5 FILLER_237_1929 ();
 b15zdnd00an1n02x5 FILLER_237_1933 ();
 b15zdnd11an1n64x5 FILLER_237_1938 ();
 b15zdnd11an1n64x5 FILLER_237_2002 ();
 b15zdnd11an1n64x5 FILLER_237_2066 ();
 b15zdnd11an1n64x5 FILLER_237_2130 ();
 b15zdnd11an1n64x5 FILLER_237_2194 ();
 b15zdnd11an1n16x5 FILLER_237_2258 ();
 b15zdnd11an1n08x5 FILLER_237_2274 ();
 b15zdnd00an1n02x5 FILLER_237_2282 ();
 b15zdnd11an1n08x5 FILLER_238_8 ();
 b15zdnd11an1n04x5 FILLER_238_16 ();
 b15zdnd00an1n02x5 FILLER_238_20 ();
 b15zdnd00an1n01x5 FILLER_238_22 ();
 b15zdnd11an1n64x5 FILLER_238_28 ();
 b15zdnd11an1n64x5 FILLER_238_92 ();
 b15zdnd11an1n64x5 FILLER_238_156 ();
 b15zdnd11an1n64x5 FILLER_238_220 ();
 b15zdnd11an1n64x5 FILLER_238_284 ();
 b15zdnd11an1n64x5 FILLER_238_348 ();
 b15zdnd11an1n64x5 FILLER_238_412 ();
 b15zdnd11an1n64x5 FILLER_238_476 ();
 b15zdnd11an1n32x5 FILLER_238_540 ();
 b15zdnd11an1n16x5 FILLER_238_572 ();
 b15zdnd11an1n08x5 FILLER_238_588 ();
 b15zdnd00an1n02x5 FILLER_238_596 ();
 b15zdnd11an1n16x5 FILLER_238_602 ();
 b15zdnd11an1n04x5 FILLER_238_618 ();
 b15zdnd00an1n02x5 FILLER_238_622 ();
 b15zdnd00an1n01x5 FILLER_238_624 ();
 b15zdnd11an1n64x5 FILLER_238_632 ();
 b15zdnd11an1n16x5 FILLER_238_696 ();
 b15zdnd11an1n04x5 FILLER_238_712 ();
 b15zdnd00an1n02x5 FILLER_238_716 ();
 b15zdnd11an1n64x5 FILLER_238_726 ();
 b15zdnd11an1n16x5 FILLER_238_790 ();
 b15zdnd11an1n08x5 FILLER_238_806 ();
 b15zdnd11an1n04x5 FILLER_238_814 ();
 b15zdnd00an1n02x5 FILLER_238_818 ();
 b15zdnd11an1n08x5 FILLER_238_862 ();
 b15zdnd11an1n04x5 FILLER_238_870 ();
 b15zdnd11an1n08x5 FILLER_238_888 ();
 b15zdnd00an1n02x5 FILLER_238_896 ();
 b15zdnd11an1n04x5 FILLER_238_940 ();
 b15zdnd11an1n64x5 FILLER_238_947 ();
 b15zdnd11an1n64x5 FILLER_238_1011 ();
 b15zdnd11an1n64x5 FILLER_238_1075 ();
 b15zdnd11an1n16x5 FILLER_238_1139 ();
 b15zdnd11an1n08x5 FILLER_238_1155 ();
 b15zdnd11an1n64x5 FILLER_238_1183 ();
 b15zdnd11an1n64x5 FILLER_238_1247 ();
 b15zdnd11an1n64x5 FILLER_238_1311 ();
 b15zdnd11an1n64x5 FILLER_238_1375 ();
 b15zdnd11an1n04x5 FILLER_238_1439 ();
 b15zdnd00an1n02x5 FILLER_238_1443 ();
 b15zdnd11an1n04x5 FILLER_238_1452 ();
 b15zdnd11an1n64x5 FILLER_238_1508 ();
 b15zdnd11an1n32x5 FILLER_238_1572 ();
 b15zdnd11an1n08x5 FILLER_238_1604 ();
 b15zdnd11an1n04x5 FILLER_238_1612 ();
 b15zdnd00an1n02x5 FILLER_238_1616 ();
 b15zdnd11an1n04x5 FILLER_238_1670 ();
 b15zdnd11an1n04x5 FILLER_238_1677 ();
 b15zdnd11an1n04x5 FILLER_238_1684 ();
 b15zdnd11an1n64x5 FILLER_238_1691 ();
 b15zdnd11an1n32x5 FILLER_238_1755 ();
 b15zdnd11an1n04x5 FILLER_238_1787 ();
 b15zdnd11an1n64x5 FILLER_238_1822 ();
 b15zdnd11an1n64x5 FILLER_238_1886 ();
 b15zdnd11an1n64x5 FILLER_238_1950 ();
 b15zdnd11an1n64x5 FILLER_238_2014 ();
 b15zdnd11an1n64x5 FILLER_238_2078 ();
 b15zdnd11an1n08x5 FILLER_238_2142 ();
 b15zdnd11an1n04x5 FILLER_238_2150 ();
 b15zdnd11an1n64x5 FILLER_238_2162 ();
 b15zdnd11an1n32x5 FILLER_238_2226 ();
 b15zdnd11an1n16x5 FILLER_238_2258 ();
 b15zdnd00an1n02x5 FILLER_238_2274 ();
 b15zdnd11an1n64x5 FILLER_239_0 ();
 b15zdnd11an1n64x5 FILLER_239_64 ();
 b15zdnd11an1n64x5 FILLER_239_128 ();
 b15zdnd11an1n64x5 FILLER_239_192 ();
 b15zdnd11an1n64x5 FILLER_239_256 ();
 b15zdnd11an1n64x5 FILLER_239_320 ();
 b15zdnd11an1n32x5 FILLER_239_384 ();
 b15zdnd11an1n16x5 FILLER_239_416 ();
 b15zdnd11an1n08x5 FILLER_239_432 ();
 b15zdnd11an1n64x5 FILLER_239_480 ();
 b15zdnd11an1n64x5 FILLER_239_544 ();
 b15zdnd11an1n32x5 FILLER_239_608 ();
 b15zdnd11an1n08x5 FILLER_239_640 ();
 b15zdnd11an1n04x5 FILLER_239_648 ();
 b15zdnd00an1n01x5 FILLER_239_652 ();
 b15zdnd11an1n64x5 FILLER_239_668 ();
 b15zdnd11an1n16x5 FILLER_239_732 ();
 b15zdnd11an1n08x5 FILLER_239_748 ();
 b15zdnd00an1n02x5 FILLER_239_756 ();
 b15zdnd11an1n32x5 FILLER_239_783 ();
 b15zdnd11an1n16x5 FILLER_239_815 ();
 b15zdnd11an1n08x5 FILLER_239_831 ();
 b15zdnd11an1n16x5 FILLER_239_842 ();
 b15zdnd00an1n01x5 FILLER_239_858 ();
 b15zdnd11an1n32x5 FILLER_239_901 ();
 b15zdnd00an1n02x5 FILLER_239_933 ();
 b15zdnd11an1n64x5 FILLER_239_938 ();
 b15zdnd11an1n64x5 FILLER_239_1002 ();
 b15zdnd11an1n32x5 FILLER_239_1066 ();
 b15zdnd11an1n04x5 FILLER_239_1098 ();
 b15zdnd00an1n02x5 FILLER_239_1102 ();
 b15zdnd11an1n32x5 FILLER_239_1111 ();
 b15zdnd11an1n16x5 FILLER_239_1143 ();
 b15zdnd11an1n08x5 FILLER_239_1159 ();
 b15zdnd00an1n02x5 FILLER_239_1167 ();
 b15zdnd00an1n01x5 FILLER_239_1169 ();
 b15zdnd11an1n64x5 FILLER_239_1182 ();
 b15zdnd11an1n08x5 FILLER_239_1246 ();
 b15zdnd00an1n02x5 FILLER_239_1254 ();
 b15zdnd00an1n01x5 FILLER_239_1256 ();
 b15zdnd11an1n04x5 FILLER_239_1261 ();
 b15zdnd00an1n01x5 FILLER_239_1265 ();
 b15zdnd11an1n64x5 FILLER_239_1280 ();
 b15zdnd11an1n64x5 FILLER_239_1344 ();
 b15zdnd11an1n32x5 FILLER_239_1408 ();
 b15zdnd11an1n16x5 FILLER_239_1440 ();
 b15zdnd11an1n04x5 FILLER_239_1456 ();
 b15zdnd00an1n01x5 FILLER_239_1460 ();
 b15zdnd11an1n04x5 FILLER_239_1464 ();
 b15zdnd11an1n04x5 FILLER_239_1471 ();
 b15zdnd11an1n04x5 FILLER_239_1478 ();
 b15zdnd11an1n64x5 FILLER_239_1485 ();
 b15zdnd11an1n64x5 FILLER_239_1549 ();
 b15zdnd11an1n04x5 FILLER_239_1613 ();
 b15zdnd00an1n02x5 FILLER_239_1617 ();
 b15zdnd00an1n01x5 FILLER_239_1619 ();
 b15zdnd11an1n04x5 FILLER_239_1672 ();
 b15zdnd00an1n01x5 FILLER_239_1676 ();
 b15zdnd11an1n04x5 FILLER_239_1680 ();
 b15zdnd11an1n64x5 FILLER_239_1687 ();
 b15zdnd11an1n64x5 FILLER_239_1751 ();
 b15zdnd11an1n64x5 FILLER_239_1815 ();
 b15zdnd11an1n64x5 FILLER_239_1879 ();
 b15zdnd11an1n64x5 FILLER_239_1943 ();
 b15zdnd11an1n64x5 FILLER_239_2007 ();
 b15zdnd11an1n64x5 FILLER_239_2071 ();
 b15zdnd11an1n32x5 FILLER_239_2135 ();
 b15zdnd11an1n16x5 FILLER_239_2167 ();
 b15zdnd11an1n64x5 FILLER_239_2189 ();
 b15zdnd11an1n16x5 FILLER_239_2253 ();
 b15zdnd11an1n08x5 FILLER_239_2269 ();
 b15zdnd11an1n04x5 FILLER_239_2277 ();
 b15zdnd00an1n02x5 FILLER_239_2281 ();
 b15zdnd00an1n01x5 FILLER_239_2283 ();
 b15zdnd11an1n64x5 FILLER_240_8 ();
 b15zdnd11an1n64x5 FILLER_240_72 ();
 b15zdnd11an1n64x5 FILLER_240_136 ();
 b15zdnd11an1n64x5 FILLER_240_200 ();
 b15zdnd11an1n32x5 FILLER_240_264 ();
 b15zdnd11an1n04x5 FILLER_240_296 ();
 b15zdnd00an1n02x5 FILLER_240_300 ();
 b15zdnd11an1n64x5 FILLER_240_344 ();
 b15zdnd11an1n32x5 FILLER_240_408 ();
 b15zdnd11an1n16x5 FILLER_240_440 ();
 b15zdnd11an1n08x5 FILLER_240_456 ();
 b15zdnd11an1n04x5 FILLER_240_464 ();
 b15zdnd00an1n02x5 FILLER_240_468 ();
 b15zdnd00an1n01x5 FILLER_240_470 ();
 b15zdnd11an1n04x5 FILLER_240_474 ();
 b15zdnd11an1n64x5 FILLER_240_481 ();
 b15zdnd11an1n64x5 FILLER_240_545 ();
 b15zdnd11an1n32x5 FILLER_240_609 ();
 b15zdnd11an1n16x5 FILLER_240_641 ();
 b15zdnd11an1n08x5 FILLER_240_657 ();
 b15zdnd11an1n04x5 FILLER_240_665 ();
 b15zdnd11an1n32x5 FILLER_240_672 ();
 b15zdnd11an1n08x5 FILLER_240_704 ();
 b15zdnd11an1n04x5 FILLER_240_712 ();
 b15zdnd00an1n02x5 FILLER_240_716 ();
 b15zdnd11an1n64x5 FILLER_240_726 ();
 b15zdnd11an1n64x5 FILLER_240_790 ();
 b15zdnd11an1n16x5 FILLER_240_854 ();
 b15zdnd00an1n02x5 FILLER_240_870 ();
 b15zdnd00an1n01x5 FILLER_240_872 ();
 b15zdnd11an1n64x5 FILLER_240_876 ();
 b15zdnd11an1n64x5 FILLER_240_940 ();
 b15zdnd11an1n64x5 FILLER_240_1004 ();
 b15zdnd11an1n64x5 FILLER_240_1068 ();
 b15zdnd11an1n64x5 FILLER_240_1132 ();
 b15zdnd11an1n32x5 FILLER_240_1196 ();
 b15zdnd11an1n08x5 FILLER_240_1228 ();
 b15zdnd00an1n02x5 FILLER_240_1236 ();
 b15zdnd11an1n64x5 FILLER_240_1245 ();
 b15zdnd11an1n64x5 FILLER_240_1309 ();
 b15zdnd11an1n32x5 FILLER_240_1373 ();
 b15zdnd11an1n64x5 FILLER_240_1414 ();
 b15zdnd11an1n04x5 FILLER_240_1478 ();
 b15zdnd11an1n64x5 FILLER_240_1485 ();
 b15zdnd11an1n64x5 FILLER_240_1549 ();
 b15zdnd11an1n16x5 FILLER_240_1613 ();
 b15zdnd11an1n04x5 FILLER_240_1629 ();
 b15zdnd00an1n02x5 FILLER_240_1633 ();
 b15zdnd00an1n01x5 FILLER_240_1635 ();
 b15zdnd11an1n04x5 FILLER_240_1639 ();
 b15zdnd11an1n08x5 FILLER_240_1646 ();
 b15zdnd11an1n04x5 FILLER_240_1661 ();
 b15zdnd11an1n64x5 FILLER_240_1707 ();
 b15zdnd11an1n64x5 FILLER_240_1771 ();
 b15zdnd11an1n64x5 FILLER_240_1835 ();
 b15zdnd11an1n32x5 FILLER_240_1899 ();
 b15zdnd11an1n16x5 FILLER_240_1931 ();
 b15zdnd00an1n01x5 FILLER_240_1947 ();
 b15zdnd11an1n64x5 FILLER_240_1954 ();
 b15zdnd11an1n64x5 FILLER_240_2018 ();
 b15zdnd11an1n64x5 FILLER_240_2082 ();
 b15zdnd11an1n08x5 FILLER_240_2146 ();
 b15zdnd11an1n64x5 FILLER_240_2162 ();
 b15zdnd11an1n32x5 FILLER_240_2226 ();
 b15zdnd11an1n16x5 FILLER_240_2258 ();
 b15zdnd00an1n02x5 FILLER_240_2274 ();
 b15zdnd11an1n64x5 FILLER_241_0 ();
 b15zdnd11an1n64x5 FILLER_241_64 ();
 b15zdnd11an1n64x5 FILLER_241_128 ();
 b15zdnd11an1n64x5 FILLER_241_192 ();
 b15zdnd11an1n32x5 FILLER_241_256 ();
 b15zdnd11an1n08x5 FILLER_241_288 ();
 b15zdnd11an1n04x5 FILLER_241_296 ();
 b15zdnd00an1n01x5 FILLER_241_300 ();
 b15zdnd11an1n64x5 FILLER_241_307 ();
 b15zdnd11an1n64x5 FILLER_241_371 ();
 b15zdnd11an1n64x5 FILLER_241_435 ();
 b15zdnd11an1n32x5 FILLER_241_499 ();
 b15zdnd11an1n16x5 FILLER_241_531 ();
 b15zdnd11an1n08x5 FILLER_241_547 ();
 b15zdnd00an1n02x5 FILLER_241_555 ();
 b15zdnd00an1n01x5 FILLER_241_557 ();
 b15zdnd11an1n04x5 FILLER_241_561 ();
 b15zdnd11an1n32x5 FILLER_241_607 ();
 b15zdnd11an1n16x5 FILLER_241_639 ();
 b15zdnd11an1n08x5 FILLER_241_655 ();
 b15zdnd11an1n04x5 FILLER_241_663 ();
 b15zdnd11an1n64x5 FILLER_241_688 ();
 b15zdnd11an1n64x5 FILLER_241_752 ();
 b15zdnd11an1n64x5 FILLER_241_816 ();
 b15zdnd11an1n64x5 FILLER_241_880 ();
 b15zdnd11an1n64x5 FILLER_241_944 ();
 b15zdnd11an1n64x5 FILLER_241_1008 ();
 b15zdnd11an1n64x5 FILLER_241_1072 ();
 b15zdnd11an1n64x5 FILLER_241_1136 ();
 b15zdnd11an1n16x5 FILLER_241_1200 ();
 b15zdnd00an1n02x5 FILLER_241_1216 ();
 b15zdnd11an1n32x5 FILLER_241_1257 ();
 b15zdnd11an1n16x5 FILLER_241_1289 ();
 b15zdnd11an1n08x5 FILLER_241_1305 ();
 b15zdnd00an1n02x5 FILLER_241_1313 ();
 b15zdnd11an1n64x5 FILLER_241_1342 ();
 b15zdnd11an1n64x5 FILLER_241_1406 ();
 b15zdnd11an1n64x5 FILLER_241_1470 ();
 b15zdnd11an1n64x5 FILLER_241_1534 ();
 b15zdnd11an1n32x5 FILLER_241_1598 ();
 b15zdnd11an1n08x5 FILLER_241_1630 ();
 b15zdnd11an1n08x5 FILLER_241_1641 ();
 b15zdnd00an1n01x5 FILLER_241_1649 ();
 b15zdnd11an1n04x5 FILLER_241_1653 ();
 b15zdnd11an1n16x5 FILLER_241_1660 ();
 b15zdnd11an1n04x5 FILLER_241_1676 ();
 b15zdnd11an1n64x5 FILLER_241_1683 ();
 b15zdnd11an1n64x5 FILLER_241_1747 ();
 b15zdnd11an1n64x5 FILLER_241_1811 ();
 b15zdnd11an1n64x5 FILLER_241_1875 ();
 b15zdnd11an1n64x5 FILLER_241_1939 ();
 b15zdnd11an1n64x5 FILLER_241_2003 ();
 b15zdnd11an1n64x5 FILLER_241_2067 ();
 b15zdnd11an1n16x5 FILLER_241_2131 ();
 b15zdnd11an1n04x5 FILLER_241_2147 ();
 b15zdnd11an1n64x5 FILLER_241_2161 ();
 b15zdnd11an1n32x5 FILLER_241_2225 ();
 b15zdnd11an1n16x5 FILLER_241_2257 ();
 b15zdnd11an1n08x5 FILLER_241_2273 ();
 b15zdnd00an1n02x5 FILLER_241_2281 ();
 b15zdnd00an1n01x5 FILLER_241_2283 ();
 b15zdnd11an1n64x5 FILLER_242_8 ();
 b15zdnd11an1n64x5 FILLER_242_72 ();
 b15zdnd11an1n64x5 FILLER_242_136 ();
 b15zdnd11an1n64x5 FILLER_242_200 ();
 b15zdnd11an1n64x5 FILLER_242_264 ();
 b15zdnd11an1n64x5 FILLER_242_328 ();
 b15zdnd11an1n64x5 FILLER_242_392 ();
 b15zdnd11an1n32x5 FILLER_242_456 ();
 b15zdnd11an1n04x5 FILLER_242_488 ();
 b15zdnd11an1n04x5 FILLER_242_495 ();
 b15zdnd00an1n02x5 FILLER_242_499 ();
 b15zdnd00an1n01x5 FILLER_242_501 ();
 b15zdnd11an1n16x5 FILLER_242_509 ();
 b15zdnd00an1n01x5 FILLER_242_525 ();
 b15zdnd11an1n04x5 FILLER_242_566 ();
 b15zdnd11an1n64x5 FILLER_242_574 ();
 b15zdnd11an1n64x5 FILLER_242_638 ();
 b15zdnd11an1n16x5 FILLER_242_702 ();
 b15zdnd11an1n64x5 FILLER_242_726 ();
 b15zdnd11an1n64x5 FILLER_242_790 ();
 b15zdnd11an1n64x5 FILLER_242_854 ();
 b15zdnd11an1n32x5 FILLER_242_918 ();
 b15zdnd11an1n08x5 FILLER_242_950 ();
 b15zdnd00an1n01x5 FILLER_242_958 ();
 b15zdnd11an1n04x5 FILLER_242_969 ();
 b15zdnd00an1n01x5 FILLER_242_973 ();
 b15zdnd11an1n08x5 FILLER_242_992 ();
 b15zdnd11an1n04x5 FILLER_242_1000 ();
 b15zdnd11an1n64x5 FILLER_242_1008 ();
 b15zdnd11an1n64x5 FILLER_242_1072 ();
 b15zdnd11an1n64x5 FILLER_242_1136 ();
 b15zdnd11an1n64x5 FILLER_242_1200 ();
 b15zdnd11an1n32x5 FILLER_242_1264 ();
 b15zdnd11an1n16x5 FILLER_242_1296 ();
 b15zdnd11an1n04x5 FILLER_242_1312 ();
 b15zdnd00an1n01x5 FILLER_242_1316 ();
 b15zdnd11an1n04x5 FILLER_242_1320 ();
 b15zdnd11an1n64x5 FILLER_242_1331 ();
 b15zdnd11an1n32x5 FILLER_242_1395 ();
 b15zdnd11an1n16x5 FILLER_242_1427 ();
 b15zdnd00an1n02x5 FILLER_242_1443 ();
 b15zdnd00an1n01x5 FILLER_242_1445 ();
 b15zdnd11an1n04x5 FILLER_242_1498 ();
 b15zdnd11an1n64x5 FILLER_242_1544 ();
 b15zdnd11an1n32x5 FILLER_242_1608 ();
 b15zdnd00an1n02x5 FILLER_242_1640 ();
 b15zdnd00an1n01x5 FILLER_242_1642 ();
 b15zdnd11an1n64x5 FILLER_242_1646 ();
 b15zdnd11an1n64x5 FILLER_242_1710 ();
 b15zdnd11an1n64x5 FILLER_242_1774 ();
 b15zdnd11an1n64x5 FILLER_242_1838 ();
 b15zdnd11an1n64x5 FILLER_242_1902 ();
 b15zdnd11an1n64x5 FILLER_242_1966 ();
 b15zdnd11an1n64x5 FILLER_242_2030 ();
 b15zdnd11an1n32x5 FILLER_242_2094 ();
 b15zdnd11an1n16x5 FILLER_242_2126 ();
 b15zdnd11an1n08x5 FILLER_242_2142 ();
 b15zdnd11an1n04x5 FILLER_242_2150 ();
 b15zdnd11an1n64x5 FILLER_242_2162 ();
 b15zdnd11an1n16x5 FILLER_242_2226 ();
 b15zdnd11an1n08x5 FILLER_242_2242 ();
 b15zdnd11an1n04x5 FILLER_242_2250 ();
 b15zdnd00an1n02x5 FILLER_242_2254 ();
 b15zdnd11an1n16x5 FILLER_242_2260 ();
 b15zdnd11an1n64x5 FILLER_243_0 ();
 b15zdnd11an1n64x5 FILLER_243_64 ();
 b15zdnd11an1n64x5 FILLER_243_128 ();
 b15zdnd11an1n64x5 FILLER_243_192 ();
 b15zdnd11an1n64x5 FILLER_243_256 ();
 b15zdnd11an1n64x5 FILLER_243_320 ();
 b15zdnd11an1n64x5 FILLER_243_384 ();
 b15zdnd11an1n16x5 FILLER_243_448 ();
 b15zdnd11an1n04x5 FILLER_243_464 ();
 b15zdnd00an1n01x5 FILLER_243_468 ();
 b15zdnd11an1n32x5 FILLER_243_521 ();
 b15zdnd11an1n04x5 FILLER_243_553 ();
 b15zdnd00an1n02x5 FILLER_243_557 ();
 b15zdnd11an1n64x5 FILLER_243_562 ();
 b15zdnd11an1n32x5 FILLER_243_626 ();
 b15zdnd00an1n02x5 FILLER_243_658 ();
 b15zdnd00an1n01x5 FILLER_243_660 ();
 b15zdnd11an1n64x5 FILLER_243_670 ();
 b15zdnd11an1n64x5 FILLER_243_734 ();
 b15zdnd11an1n64x5 FILLER_243_798 ();
 b15zdnd11an1n64x5 FILLER_243_862 ();
 b15zdnd11an1n32x5 FILLER_243_926 ();
 b15zdnd11an1n64x5 FILLER_243_972 ();
 b15zdnd11an1n16x5 FILLER_243_1036 ();
 b15zdnd00an1n02x5 FILLER_243_1052 ();
 b15zdnd11an1n16x5 FILLER_243_1094 ();
 b15zdnd00an1n02x5 FILLER_243_1110 ();
 b15zdnd11an1n64x5 FILLER_243_1134 ();
 b15zdnd11an1n64x5 FILLER_243_1198 ();
 b15zdnd11an1n64x5 FILLER_243_1262 ();
 b15zdnd00an1n02x5 FILLER_243_1326 ();
 b15zdnd11an1n04x5 FILLER_243_1331 ();
 b15zdnd11an1n04x5 FILLER_243_1338 ();
 b15zdnd11an1n64x5 FILLER_243_1345 ();
 b15zdnd11an1n32x5 FILLER_243_1409 ();
 b15zdnd11an1n16x5 FILLER_243_1441 ();
 b15zdnd11an1n08x5 FILLER_243_1457 ();
 b15zdnd00an1n01x5 FILLER_243_1465 ();
 b15zdnd11an1n64x5 FILLER_243_1469 ();
 b15zdnd11an1n64x5 FILLER_243_1533 ();
 b15zdnd11an1n64x5 FILLER_243_1597 ();
 b15zdnd11an1n64x5 FILLER_243_1661 ();
 b15zdnd11an1n64x5 FILLER_243_1725 ();
 b15zdnd11an1n64x5 FILLER_243_1789 ();
 b15zdnd11an1n64x5 FILLER_243_1853 ();
 b15zdnd11an1n64x5 FILLER_243_1917 ();
 b15zdnd11an1n64x5 FILLER_243_1981 ();
 b15zdnd11an1n64x5 FILLER_243_2045 ();
 b15zdnd11an1n64x5 FILLER_243_2109 ();
 b15zdnd11an1n64x5 FILLER_243_2173 ();
 b15zdnd11an1n04x5 FILLER_243_2237 ();
 b15zdnd00an1n02x5 FILLER_243_2241 ();
 b15zdnd00an1n01x5 FILLER_243_2243 ();
 b15zdnd11an1n32x5 FILLER_243_2248 ();
 b15zdnd11an1n04x5 FILLER_243_2280 ();
 b15zdnd11an1n64x5 FILLER_244_8 ();
 b15zdnd11an1n64x5 FILLER_244_72 ();
 b15zdnd11an1n64x5 FILLER_244_136 ();
 b15zdnd11an1n64x5 FILLER_244_200 ();
 b15zdnd11an1n32x5 FILLER_244_264 ();
 b15zdnd11an1n04x5 FILLER_244_296 ();
 b15zdnd00an1n01x5 FILLER_244_300 ();
 b15zdnd11an1n64x5 FILLER_244_304 ();
 b15zdnd11an1n64x5 FILLER_244_368 ();
 b15zdnd11an1n32x5 FILLER_244_432 ();
 b15zdnd11an1n16x5 FILLER_244_464 ();
 b15zdnd11an1n08x5 FILLER_244_480 ();
 b15zdnd00an1n01x5 FILLER_244_488 ();
 b15zdnd11an1n04x5 FILLER_244_492 ();
 b15zdnd11an1n64x5 FILLER_244_499 ();
 b15zdnd11an1n64x5 FILLER_244_563 ();
 b15zdnd11an1n64x5 FILLER_244_627 ();
 b15zdnd11an1n16x5 FILLER_244_691 ();
 b15zdnd11an1n08x5 FILLER_244_707 ();
 b15zdnd00an1n02x5 FILLER_244_715 ();
 b15zdnd00an1n01x5 FILLER_244_717 ();
 b15zdnd11an1n32x5 FILLER_244_726 ();
 b15zdnd11an1n08x5 FILLER_244_758 ();
 b15zdnd00an1n02x5 FILLER_244_766 ();
 b15zdnd00an1n01x5 FILLER_244_768 ();
 b15zdnd11an1n04x5 FILLER_244_811 ();
 b15zdnd11an1n64x5 FILLER_244_827 ();
 b15zdnd11an1n32x5 FILLER_244_891 ();
 b15zdnd11an1n16x5 FILLER_244_923 ();
 b15zdnd11an1n04x5 FILLER_244_939 ();
 b15zdnd00an1n02x5 FILLER_244_943 ();
 b15zdnd00an1n01x5 FILLER_244_945 ();
 b15zdnd11an1n08x5 FILLER_244_957 ();
 b15zdnd11an1n64x5 FILLER_244_991 ();
 b15zdnd11an1n16x5 FILLER_244_1055 ();
 b15zdnd00an1n02x5 FILLER_244_1071 ();
 b15zdnd00an1n01x5 FILLER_244_1073 ();
 b15zdnd11an1n08x5 FILLER_244_1080 ();
 b15zdnd00an1n01x5 FILLER_244_1088 ();
 b15zdnd11an1n64x5 FILLER_244_1092 ();
 b15zdnd11an1n64x5 FILLER_244_1156 ();
 b15zdnd11an1n08x5 FILLER_244_1220 ();
 b15zdnd11an1n04x5 FILLER_244_1228 ();
 b15zdnd00an1n01x5 FILLER_244_1232 ();
 b15zdnd11an1n64x5 FILLER_244_1244 ();
 b15zdnd00an1n02x5 FILLER_244_1308 ();
 b15zdnd11an1n08x5 FILLER_244_1362 ();
 b15zdnd11an1n04x5 FILLER_244_1370 ();
 b15zdnd00an1n02x5 FILLER_244_1374 ();
 b15zdnd11an1n16x5 FILLER_244_1383 ();
 b15zdnd11an1n08x5 FILLER_244_1399 ();
 b15zdnd00an1n01x5 FILLER_244_1407 ();
 b15zdnd11an1n32x5 FILLER_244_1417 ();
 b15zdnd11an1n16x5 FILLER_244_1449 ();
 b15zdnd00an1n02x5 FILLER_244_1465 ();
 b15zdnd11an1n04x5 FILLER_244_1470 ();
 b15zdnd11an1n32x5 FILLER_244_1477 ();
 b15zdnd11an1n08x5 FILLER_244_1509 ();
 b15zdnd00an1n02x5 FILLER_244_1517 ();
 b15zdnd00an1n01x5 FILLER_244_1519 ();
 b15zdnd11an1n04x5 FILLER_244_1527 ();
 b15zdnd11an1n64x5 FILLER_244_1539 ();
 b15zdnd11an1n64x5 FILLER_244_1603 ();
 b15zdnd11an1n64x5 FILLER_244_1667 ();
 b15zdnd11an1n64x5 FILLER_244_1731 ();
 b15zdnd11an1n64x5 FILLER_244_1795 ();
 b15zdnd11an1n64x5 FILLER_244_1859 ();
 b15zdnd11an1n64x5 FILLER_244_1923 ();
 b15zdnd11an1n64x5 FILLER_244_1987 ();
 b15zdnd11an1n64x5 FILLER_244_2051 ();
 b15zdnd11an1n32x5 FILLER_244_2115 ();
 b15zdnd11an1n04x5 FILLER_244_2147 ();
 b15zdnd00an1n02x5 FILLER_244_2151 ();
 b15zdnd00an1n01x5 FILLER_244_2153 ();
 b15zdnd11an1n64x5 FILLER_244_2162 ();
 b15zdnd11an1n32x5 FILLER_244_2226 ();
 b15zdnd11an1n16x5 FILLER_244_2258 ();
 b15zdnd00an1n02x5 FILLER_244_2274 ();
 b15zdnd11an1n64x5 FILLER_245_0 ();
 b15zdnd11an1n64x5 FILLER_245_64 ();
 b15zdnd11an1n64x5 FILLER_245_128 ();
 b15zdnd11an1n64x5 FILLER_245_192 ();
 b15zdnd11an1n64x5 FILLER_245_256 ();
 b15zdnd11an1n64x5 FILLER_245_320 ();
 b15zdnd11an1n64x5 FILLER_245_384 ();
 b15zdnd11an1n64x5 FILLER_245_448 ();
 b15zdnd11an1n64x5 FILLER_245_512 ();
 b15zdnd11an1n64x5 FILLER_245_576 ();
 b15zdnd11an1n64x5 FILLER_245_640 ();
 b15zdnd11an1n64x5 FILLER_245_704 ();
 b15zdnd11an1n64x5 FILLER_245_768 ();
 b15zdnd11an1n64x5 FILLER_245_832 ();
 b15zdnd11an1n32x5 FILLER_245_896 ();
 b15zdnd11an1n16x5 FILLER_245_928 ();
 b15zdnd11an1n04x5 FILLER_245_944 ();
 b15zdnd11an1n64x5 FILLER_245_975 ();
 b15zdnd11an1n32x5 FILLER_245_1039 ();
 b15zdnd11an1n16x5 FILLER_245_1071 ();
 b15zdnd00an1n01x5 FILLER_245_1087 ();
 b15zdnd11an1n64x5 FILLER_245_1091 ();
 b15zdnd11an1n32x5 FILLER_245_1155 ();
 b15zdnd11an1n04x5 FILLER_245_1187 ();
 b15zdnd00an1n02x5 FILLER_245_1191 ();
 b15zdnd00an1n01x5 FILLER_245_1193 ();
 b15zdnd11an1n64x5 FILLER_245_1205 ();
 b15zdnd11an1n32x5 FILLER_245_1269 ();
 b15zdnd11an1n08x5 FILLER_245_1301 ();
 b15zdnd11an1n16x5 FILLER_245_1361 ();
 b15zdnd11an1n32x5 FILLER_245_1386 ();
 b15zdnd11an1n16x5 FILLER_245_1418 ();
 b15zdnd11an1n08x5 FILLER_245_1434 ();
 b15zdnd11an1n04x5 FILLER_245_1442 ();
 b15zdnd00an1n02x5 FILLER_245_1446 ();
 b15zdnd00an1n01x5 FILLER_245_1448 ();
 b15zdnd11an1n08x5 FILLER_245_1469 ();
 b15zdnd11an1n04x5 FILLER_245_1477 ();
 b15zdnd00an1n01x5 FILLER_245_1481 ();
 b15zdnd11an1n64x5 FILLER_245_1490 ();
 b15zdnd11an1n64x5 FILLER_245_1554 ();
 b15zdnd11an1n64x5 FILLER_245_1618 ();
 b15zdnd11an1n64x5 FILLER_245_1682 ();
 b15zdnd11an1n64x5 FILLER_245_1746 ();
 b15zdnd11an1n64x5 FILLER_245_1810 ();
 b15zdnd11an1n32x5 FILLER_245_1874 ();
 b15zdnd11an1n08x5 FILLER_245_1906 ();
 b15zdnd11an1n04x5 FILLER_245_1914 ();
 b15zdnd00an1n02x5 FILLER_245_1918 ();
 b15zdnd00an1n01x5 FILLER_245_1920 ();
 b15zdnd11an1n64x5 FILLER_245_1973 ();
 b15zdnd11an1n64x5 FILLER_245_2037 ();
 b15zdnd11an1n64x5 FILLER_245_2101 ();
 b15zdnd11an1n64x5 FILLER_245_2165 ();
 b15zdnd11an1n32x5 FILLER_245_2229 ();
 b15zdnd11an1n16x5 FILLER_245_2261 ();
 b15zdnd11an1n04x5 FILLER_245_2277 ();
 b15zdnd00an1n02x5 FILLER_245_2281 ();
 b15zdnd00an1n01x5 FILLER_245_2283 ();
 b15zdnd11an1n64x5 FILLER_246_8 ();
 b15zdnd11an1n64x5 FILLER_246_72 ();
 b15zdnd11an1n64x5 FILLER_246_136 ();
 b15zdnd11an1n64x5 FILLER_246_200 ();
 b15zdnd11an1n64x5 FILLER_246_264 ();
 b15zdnd11an1n64x5 FILLER_246_328 ();
 b15zdnd11an1n64x5 FILLER_246_392 ();
 b15zdnd11an1n64x5 FILLER_246_456 ();
 b15zdnd11an1n64x5 FILLER_246_520 ();
 b15zdnd11an1n64x5 FILLER_246_584 ();
 b15zdnd11an1n08x5 FILLER_246_648 ();
 b15zdnd00an1n02x5 FILLER_246_656 ();
 b15zdnd00an1n01x5 FILLER_246_658 ();
 b15zdnd11an1n32x5 FILLER_246_664 ();
 b15zdnd11an1n16x5 FILLER_246_696 ();
 b15zdnd11an1n04x5 FILLER_246_712 ();
 b15zdnd00an1n02x5 FILLER_246_716 ();
 b15zdnd11an1n64x5 FILLER_246_726 ();
 b15zdnd11an1n64x5 FILLER_246_790 ();
 b15zdnd11an1n64x5 FILLER_246_854 ();
 b15zdnd11an1n64x5 FILLER_246_918 ();
 b15zdnd11an1n16x5 FILLER_246_982 ();
 b15zdnd11an1n04x5 FILLER_246_998 ();
 b15zdnd00an1n02x5 FILLER_246_1002 ();
 b15zdnd11an1n64x5 FILLER_246_1018 ();
 b15zdnd11an1n64x5 FILLER_246_1082 ();
 b15zdnd11an1n64x5 FILLER_246_1146 ();
 b15zdnd11an1n08x5 FILLER_246_1210 ();
 b15zdnd00an1n02x5 FILLER_246_1218 ();
 b15zdnd00an1n01x5 FILLER_246_1220 ();
 b15zdnd11an1n64x5 FILLER_246_1226 ();
 b15zdnd11an1n16x5 FILLER_246_1290 ();
 b15zdnd11an1n04x5 FILLER_246_1306 ();
 b15zdnd00an1n02x5 FILLER_246_1310 ();
 b15zdnd11an1n08x5 FILLER_246_1320 ();
 b15zdnd00an1n01x5 FILLER_246_1328 ();
 b15zdnd11an1n04x5 FILLER_246_1332 ();
 b15zdnd11an1n04x5 FILLER_246_1356 ();
 b15zdnd00an1n01x5 FILLER_246_1360 ();
 b15zdnd11an1n04x5 FILLER_246_1368 ();
 b15zdnd00an1n01x5 FILLER_246_1372 ();
 b15zdnd11an1n64x5 FILLER_246_1380 ();
 b15zdnd11an1n64x5 FILLER_246_1444 ();
 b15zdnd11an1n64x5 FILLER_246_1508 ();
 b15zdnd11an1n64x5 FILLER_246_1572 ();
 b15zdnd11an1n64x5 FILLER_246_1636 ();
 b15zdnd11an1n64x5 FILLER_246_1700 ();
 b15zdnd11an1n64x5 FILLER_246_1764 ();
 b15zdnd11an1n64x5 FILLER_246_1828 ();
 b15zdnd11an1n32x5 FILLER_246_1892 ();
 b15zdnd11an1n08x5 FILLER_246_1924 ();
 b15zdnd11an1n04x5 FILLER_246_1935 ();
 b15zdnd11an1n04x5 FILLER_246_1942 ();
 b15zdnd00an1n01x5 FILLER_246_1946 ();
 b15zdnd11an1n16x5 FILLER_246_1950 ();
 b15zdnd11an1n04x5 FILLER_246_1966 ();
 b15zdnd00an1n02x5 FILLER_246_1970 ();
 b15zdnd00an1n01x5 FILLER_246_1972 ();
 b15zdnd11an1n64x5 FILLER_246_1976 ();
 b15zdnd11an1n08x5 FILLER_246_2040 ();
 b15zdnd11an1n04x5 FILLER_246_2048 ();
 b15zdnd11an1n64x5 FILLER_246_2072 ();
 b15zdnd11an1n16x5 FILLER_246_2136 ();
 b15zdnd00an1n02x5 FILLER_246_2152 ();
 b15zdnd11an1n08x5 FILLER_246_2162 ();
 b15zdnd11an1n64x5 FILLER_246_2184 ();
 b15zdnd11an1n16x5 FILLER_246_2248 ();
 b15zdnd11an1n08x5 FILLER_246_2264 ();
 b15zdnd11an1n04x5 FILLER_246_2272 ();
 b15zdnd11an1n64x5 FILLER_247_0 ();
 b15zdnd11an1n64x5 FILLER_247_64 ();
 b15zdnd11an1n64x5 FILLER_247_128 ();
 b15zdnd11an1n64x5 FILLER_247_192 ();
 b15zdnd11an1n64x5 FILLER_247_256 ();
 b15zdnd11an1n64x5 FILLER_247_320 ();
 b15zdnd11an1n64x5 FILLER_247_384 ();
 b15zdnd11an1n64x5 FILLER_247_448 ();
 b15zdnd11an1n64x5 FILLER_247_512 ();
 b15zdnd11an1n64x5 FILLER_247_576 ();
 b15zdnd00an1n01x5 FILLER_247_640 ();
 b15zdnd11an1n04x5 FILLER_247_683 ();
 b15zdnd11an1n32x5 FILLER_247_695 ();
 b15zdnd11an1n16x5 FILLER_247_727 ();
 b15zdnd11an1n08x5 FILLER_247_743 ();
 b15zdnd11an1n04x5 FILLER_247_751 ();
 b15zdnd11an1n64x5 FILLER_247_758 ();
 b15zdnd11an1n64x5 FILLER_247_822 ();
 b15zdnd11an1n64x5 FILLER_247_886 ();
 b15zdnd11an1n64x5 FILLER_247_950 ();
 b15zdnd11an1n64x5 FILLER_247_1014 ();
 b15zdnd11an1n64x5 FILLER_247_1078 ();
 b15zdnd11an1n64x5 FILLER_247_1142 ();
 b15zdnd11an1n08x5 FILLER_247_1206 ();
 b15zdnd00an1n01x5 FILLER_247_1214 ();
 b15zdnd11an1n32x5 FILLER_247_1257 ();
 b15zdnd11an1n16x5 FILLER_247_1289 ();
 b15zdnd11an1n64x5 FILLER_247_1357 ();
 b15zdnd11an1n16x5 FILLER_247_1421 ();
 b15zdnd11an1n08x5 FILLER_247_1437 ();
 b15zdnd11an1n04x5 FILLER_247_1445 ();
 b15zdnd00an1n02x5 FILLER_247_1449 ();
 b15zdnd00an1n01x5 FILLER_247_1451 ();
 b15zdnd11an1n64x5 FILLER_247_1455 ();
 b15zdnd11an1n64x5 FILLER_247_1519 ();
 b15zdnd11an1n64x5 FILLER_247_1583 ();
 b15zdnd11an1n64x5 FILLER_247_1647 ();
 b15zdnd11an1n64x5 FILLER_247_1711 ();
 b15zdnd11an1n64x5 FILLER_247_1775 ();
 b15zdnd11an1n32x5 FILLER_247_1839 ();
 b15zdnd11an1n16x5 FILLER_247_1871 ();
 b15zdnd00an1n02x5 FILLER_247_1887 ();
 b15zdnd00an1n01x5 FILLER_247_1889 ();
 b15zdnd11an1n04x5 FILLER_247_1932 ();
 b15zdnd11an1n32x5 FILLER_247_1976 ();
 b15zdnd11an1n16x5 FILLER_247_2008 ();
 b15zdnd11an1n08x5 FILLER_247_2024 ();
 b15zdnd11an1n04x5 FILLER_247_2032 ();
 b15zdnd00an1n02x5 FILLER_247_2036 ();
 b15zdnd00an1n01x5 FILLER_247_2038 ();
 b15zdnd11an1n08x5 FILLER_247_2059 ();
 b15zdnd00an1n02x5 FILLER_247_2067 ();
 b15zdnd00an1n01x5 FILLER_247_2069 ();
 b15zdnd11an1n64x5 FILLER_247_2073 ();
 b15zdnd11an1n16x5 FILLER_247_2137 ();
 b15zdnd00an1n02x5 FILLER_247_2153 ();
 b15zdnd11an1n64x5 FILLER_247_2169 ();
 b15zdnd11an1n32x5 FILLER_247_2233 ();
 b15zdnd11an1n16x5 FILLER_247_2265 ();
 b15zdnd00an1n02x5 FILLER_247_2281 ();
 b15zdnd00an1n01x5 FILLER_247_2283 ();
 b15zdnd11an1n64x5 FILLER_248_8 ();
 b15zdnd11an1n64x5 FILLER_248_72 ();
 b15zdnd11an1n64x5 FILLER_248_136 ();
 b15zdnd11an1n64x5 FILLER_248_200 ();
 b15zdnd11an1n64x5 FILLER_248_264 ();
 b15zdnd11an1n64x5 FILLER_248_328 ();
 b15zdnd11an1n64x5 FILLER_248_392 ();
 b15zdnd11an1n64x5 FILLER_248_456 ();
 b15zdnd11an1n64x5 FILLER_248_520 ();
 b15zdnd11an1n64x5 FILLER_248_584 ();
 b15zdnd11an1n08x5 FILLER_248_648 ();
 b15zdnd11an1n04x5 FILLER_248_663 ();
 b15zdnd11an1n04x5 FILLER_248_671 ();
 b15zdnd11an1n08x5 FILLER_248_680 ();
 b15zdnd11an1n16x5 FILLER_248_694 ();
 b15zdnd11an1n08x5 FILLER_248_710 ();
 b15zdnd00an1n02x5 FILLER_248_726 ();
 b15zdnd11an1n64x5 FILLER_248_780 ();
 b15zdnd11an1n64x5 FILLER_248_844 ();
 b15zdnd11an1n64x5 FILLER_248_908 ();
 b15zdnd11an1n64x5 FILLER_248_972 ();
 b15zdnd11an1n32x5 FILLER_248_1036 ();
 b15zdnd11an1n08x5 FILLER_248_1068 ();
 b15zdnd11an1n04x5 FILLER_248_1076 ();
 b15zdnd00an1n02x5 FILLER_248_1080 ();
 b15zdnd11an1n64x5 FILLER_248_1096 ();
 b15zdnd11an1n16x5 FILLER_248_1160 ();
 b15zdnd11an1n08x5 FILLER_248_1176 ();
 b15zdnd11an1n04x5 FILLER_248_1184 ();
 b15zdnd11an1n04x5 FILLER_248_1228 ();
 b15zdnd11an1n64x5 FILLER_248_1235 ();
 b15zdnd11an1n16x5 FILLER_248_1299 ();
 b15zdnd11an1n08x5 FILLER_248_1315 ();
 b15zdnd11an1n04x5 FILLER_248_1323 ();
 b15zdnd11an1n04x5 FILLER_248_1330 ();
 b15zdnd11an1n04x5 FILLER_248_1337 ();
 b15zdnd11an1n08x5 FILLER_248_1344 ();
 b15zdnd00an1n02x5 FILLER_248_1352 ();
 b15zdnd00an1n01x5 FILLER_248_1354 ();
 b15zdnd11an1n64x5 FILLER_248_1362 ();
 b15zdnd11an1n16x5 FILLER_248_1426 ();
 b15zdnd11an1n04x5 FILLER_248_1445 ();
 b15zdnd00an1n02x5 FILLER_248_1449 ();
 b15zdnd11an1n64x5 FILLER_248_1454 ();
 b15zdnd11an1n64x5 FILLER_248_1518 ();
 b15zdnd11an1n64x5 FILLER_248_1582 ();
 b15zdnd11an1n64x5 FILLER_248_1646 ();
 b15zdnd11an1n64x5 FILLER_248_1710 ();
 b15zdnd11an1n64x5 FILLER_248_1774 ();
 b15zdnd11an1n32x5 FILLER_248_1838 ();
 b15zdnd11an1n04x5 FILLER_248_1870 ();
 b15zdnd11an1n32x5 FILLER_248_1926 ();
 b15zdnd11an1n08x5 FILLER_248_1958 ();
 b15zdnd00an1n02x5 FILLER_248_1966 ();
 b15zdnd11an1n64x5 FILLER_248_1971 ();
 b15zdnd11an1n08x5 FILLER_248_2035 ();
 b15zdnd00an1n01x5 FILLER_248_2043 ();
 b15zdnd11an1n04x5 FILLER_248_2096 ();
 b15zdnd11an1n16x5 FILLER_248_2131 ();
 b15zdnd11an1n04x5 FILLER_248_2147 ();
 b15zdnd00an1n02x5 FILLER_248_2151 ();
 b15zdnd00an1n01x5 FILLER_248_2153 ();
 b15zdnd11an1n64x5 FILLER_248_2162 ();
 b15zdnd11an1n32x5 FILLER_248_2226 ();
 b15zdnd11an1n16x5 FILLER_248_2258 ();
 b15zdnd00an1n02x5 FILLER_248_2274 ();
 b15zdnd11an1n64x5 FILLER_249_0 ();
 b15zdnd11an1n64x5 FILLER_249_64 ();
 b15zdnd11an1n64x5 FILLER_249_128 ();
 b15zdnd11an1n64x5 FILLER_249_192 ();
 b15zdnd11an1n32x5 FILLER_249_256 ();
 b15zdnd00an1n01x5 FILLER_249_288 ();
 b15zdnd11an1n64x5 FILLER_249_295 ();
 b15zdnd11an1n64x5 FILLER_249_359 ();
 b15zdnd11an1n64x5 FILLER_249_423 ();
 b15zdnd11an1n64x5 FILLER_249_487 ();
 b15zdnd11an1n64x5 FILLER_249_551 ();
 b15zdnd11an1n08x5 FILLER_249_615 ();
 b15zdnd11an1n16x5 FILLER_249_626 ();
 b15zdnd11an1n08x5 FILLER_249_642 ();
 b15zdnd11an1n04x5 FILLER_249_650 ();
 b15zdnd11an1n32x5 FILLER_249_696 ();
 b15zdnd11an1n16x5 FILLER_249_728 ();
 b15zdnd11an1n08x5 FILLER_249_744 ();
 b15zdnd00an1n01x5 FILLER_249_752 ();
 b15zdnd11an1n64x5 FILLER_249_756 ();
 b15zdnd11an1n08x5 FILLER_249_820 ();
 b15zdnd11an1n04x5 FILLER_249_828 ();
 b15zdnd11an1n64x5 FILLER_249_874 ();
 b15zdnd11an1n64x5 FILLER_249_938 ();
 b15zdnd11an1n64x5 FILLER_249_1002 ();
 b15zdnd11an1n08x5 FILLER_249_1088 ();
 b15zdnd11an1n04x5 FILLER_249_1096 ();
 b15zdnd11an1n16x5 FILLER_249_1121 ();
 b15zdnd11an1n08x5 FILLER_249_1137 ();
 b15zdnd11an1n04x5 FILLER_249_1145 ();
 b15zdnd11an1n32x5 FILLER_249_1169 ();
 b15zdnd11an1n16x5 FILLER_249_1201 ();
 b15zdnd11an1n04x5 FILLER_249_1217 ();
 b15zdnd00an1n02x5 FILLER_249_1221 ();
 b15zdnd00an1n01x5 FILLER_249_1223 ();
 b15zdnd11an1n64x5 FILLER_249_1227 ();
 b15zdnd11an1n32x5 FILLER_249_1291 ();
 b15zdnd11an1n04x5 FILLER_249_1323 ();
 b15zdnd00an1n02x5 FILLER_249_1327 ();
 b15zdnd00an1n01x5 FILLER_249_1329 ();
 b15zdnd11an1n04x5 FILLER_249_1333 ();
 b15zdnd11an1n64x5 FILLER_249_1340 ();
 b15zdnd11an1n16x5 FILLER_249_1404 ();
 b15zdnd11an1n04x5 FILLER_249_1420 ();
 b15zdnd00an1n02x5 FILLER_249_1424 ();
 b15zdnd11an1n64x5 FILLER_249_1478 ();
 b15zdnd11an1n64x5 FILLER_249_1542 ();
 b15zdnd11an1n64x5 FILLER_249_1606 ();
 b15zdnd11an1n32x5 FILLER_249_1670 ();
 b15zdnd11an1n16x5 FILLER_249_1702 ();
 b15zdnd11an1n08x5 FILLER_249_1718 ();
 b15zdnd00an1n01x5 FILLER_249_1726 ();
 b15zdnd11an1n32x5 FILLER_249_1735 ();
 b15zdnd11an1n16x5 FILLER_249_1767 ();
 b15zdnd11an1n08x5 FILLER_249_1783 ();
 b15zdnd00an1n02x5 FILLER_249_1791 ();
 b15zdnd00an1n01x5 FILLER_249_1793 ();
 b15zdnd11an1n64x5 FILLER_249_1806 ();
 b15zdnd11an1n16x5 FILLER_249_1870 ();
 b15zdnd11an1n04x5 FILLER_249_1886 ();
 b15zdnd00an1n02x5 FILLER_249_1890 ();
 b15zdnd11an1n04x5 FILLER_249_1895 ();
 b15zdnd11an1n64x5 FILLER_249_1902 ();
 b15zdnd11an1n64x5 FILLER_249_1966 ();
 b15zdnd11an1n32x5 FILLER_249_2030 ();
 b15zdnd11an1n04x5 FILLER_249_2065 ();
 b15zdnd11an1n64x5 FILLER_249_2072 ();
 b15zdnd11an1n64x5 FILLER_249_2136 ();
 b15zdnd11an1n64x5 FILLER_249_2200 ();
 b15zdnd11an1n16x5 FILLER_249_2264 ();
 b15zdnd11an1n04x5 FILLER_249_2280 ();
 b15zdnd11an1n64x5 FILLER_250_8 ();
 b15zdnd11an1n64x5 FILLER_250_72 ();
 b15zdnd11an1n64x5 FILLER_250_136 ();
 b15zdnd11an1n64x5 FILLER_250_200 ();
 b15zdnd11an1n64x5 FILLER_250_264 ();
 b15zdnd11an1n64x5 FILLER_250_328 ();
 b15zdnd11an1n64x5 FILLER_250_392 ();
 b15zdnd11an1n64x5 FILLER_250_456 ();
 b15zdnd11an1n64x5 FILLER_250_520 ();
 b15zdnd11an1n08x5 FILLER_250_584 ();
 b15zdnd11an1n04x5 FILLER_250_592 ();
 b15zdnd11an1n08x5 FILLER_250_648 ();
 b15zdnd00an1n02x5 FILLER_250_656 ();
 b15zdnd11an1n04x5 FILLER_250_663 ();
 b15zdnd11an1n08x5 FILLER_250_709 ();
 b15zdnd00an1n01x5 FILLER_250_717 ();
 b15zdnd11an1n16x5 FILLER_250_726 ();
 b15zdnd11an1n08x5 FILLER_250_742 ();
 b15zdnd00an1n02x5 FILLER_250_750 ();
 b15zdnd11an1n64x5 FILLER_250_755 ();
 b15zdnd11an1n32x5 FILLER_250_819 ();
 b15zdnd11an1n08x5 FILLER_250_851 ();
 b15zdnd11an1n04x5 FILLER_250_859 ();
 b15zdnd00an1n02x5 FILLER_250_863 ();
 b15zdnd11an1n64x5 FILLER_250_907 ();
 b15zdnd11an1n64x5 FILLER_250_971 ();
 b15zdnd00an1n02x5 FILLER_250_1035 ();
 b15zdnd11an1n32x5 FILLER_250_1041 ();
 b15zdnd11an1n16x5 FILLER_250_1073 ();
 b15zdnd11an1n08x5 FILLER_250_1089 ();
 b15zdnd11an1n04x5 FILLER_250_1097 ();
 b15zdnd11an1n08x5 FILLER_250_1111 ();
 b15zdnd11an1n04x5 FILLER_250_1119 ();
 b15zdnd00an1n02x5 FILLER_250_1123 ();
 b15zdnd00an1n01x5 FILLER_250_1125 ();
 b15zdnd11an1n64x5 FILLER_250_1137 ();
 b15zdnd11an1n64x5 FILLER_250_1201 ();
 b15zdnd11an1n64x5 FILLER_250_1265 ();
 b15zdnd11an1n64x5 FILLER_250_1329 ();
 b15zdnd11an1n16x5 FILLER_250_1393 ();
 b15zdnd11an1n08x5 FILLER_250_1416 ();
 b15zdnd11an1n04x5 FILLER_250_1424 ();
 b15zdnd11an1n64x5 FILLER_250_1480 ();
 b15zdnd11an1n64x5 FILLER_250_1544 ();
 b15zdnd11an1n64x5 FILLER_250_1608 ();
 b15zdnd11an1n32x5 FILLER_250_1672 ();
 b15zdnd00an1n01x5 FILLER_250_1704 ();
 b15zdnd11an1n64x5 FILLER_250_1713 ();
 b15zdnd11an1n08x5 FILLER_250_1777 ();
 b15zdnd00an1n02x5 FILLER_250_1785 ();
 b15zdnd00an1n01x5 FILLER_250_1787 ();
 b15zdnd11an1n64x5 FILLER_250_1812 ();
 b15zdnd11an1n16x5 FILLER_250_1876 ();
 b15zdnd11an1n08x5 FILLER_250_1892 ();
 b15zdnd11an1n64x5 FILLER_250_1903 ();
 b15zdnd11an1n64x5 FILLER_250_1967 ();
 b15zdnd11an1n64x5 FILLER_250_2031 ();
 b15zdnd11an1n32x5 FILLER_250_2095 ();
 b15zdnd11an1n16x5 FILLER_250_2127 ();
 b15zdnd11an1n08x5 FILLER_250_2143 ();
 b15zdnd00an1n02x5 FILLER_250_2151 ();
 b15zdnd00an1n01x5 FILLER_250_2153 ();
 b15zdnd11an1n64x5 FILLER_250_2162 ();
 b15zdnd11an1n32x5 FILLER_250_2226 ();
 b15zdnd11an1n16x5 FILLER_250_2258 ();
 b15zdnd00an1n02x5 FILLER_250_2274 ();
 b15zdnd11an1n64x5 FILLER_251_0 ();
 b15zdnd11an1n64x5 FILLER_251_64 ();
 b15zdnd11an1n64x5 FILLER_251_128 ();
 b15zdnd11an1n64x5 FILLER_251_192 ();
 b15zdnd11an1n32x5 FILLER_251_256 ();
 b15zdnd00an1n02x5 FILLER_251_288 ();
 b15zdnd00an1n01x5 FILLER_251_290 ();
 b15zdnd11an1n64x5 FILLER_251_295 ();
 b15zdnd11an1n64x5 FILLER_251_359 ();
 b15zdnd11an1n64x5 FILLER_251_423 ();
 b15zdnd11an1n64x5 FILLER_251_487 ();
 b15zdnd11an1n32x5 FILLER_251_551 ();
 b15zdnd11an1n16x5 FILLER_251_583 ();
 b15zdnd11an1n08x5 FILLER_251_599 ();
 b15zdnd11an1n04x5 FILLER_251_607 ();
 b15zdnd00an1n02x5 FILLER_251_611 ();
 b15zdnd00an1n01x5 FILLER_251_613 ();
 b15zdnd11an1n04x5 FILLER_251_617 ();
 b15zdnd11an1n16x5 FILLER_251_624 ();
 b15zdnd11an1n08x5 FILLER_251_640 ();
 b15zdnd11an1n04x5 FILLER_251_648 ();
 b15zdnd00an1n01x5 FILLER_251_652 ();
 b15zdnd11an1n64x5 FILLER_251_695 ();
 b15zdnd11an1n64x5 FILLER_251_759 ();
 b15zdnd11an1n32x5 FILLER_251_823 ();
 b15zdnd11an1n16x5 FILLER_251_855 ();
 b15zdnd00an1n01x5 FILLER_251_871 ();
 b15zdnd11an1n64x5 FILLER_251_914 ();
 b15zdnd11an1n64x5 FILLER_251_978 ();
 b15zdnd11an1n64x5 FILLER_251_1042 ();
 b15zdnd11an1n32x5 FILLER_251_1106 ();
 b15zdnd11an1n16x5 FILLER_251_1138 ();
 b15zdnd11an1n04x5 FILLER_251_1154 ();
 b15zdnd00an1n02x5 FILLER_251_1158 ();
 b15zdnd11an1n64x5 FILLER_251_1170 ();
 b15zdnd11an1n64x5 FILLER_251_1234 ();
 b15zdnd11an1n64x5 FILLER_251_1298 ();
 b15zdnd11an1n64x5 FILLER_251_1362 ();
 b15zdnd11an1n08x5 FILLER_251_1426 ();
 b15zdnd00an1n01x5 FILLER_251_1434 ();
 b15zdnd11an1n08x5 FILLER_251_1477 ();
 b15zdnd11an1n04x5 FILLER_251_1485 ();
 b15zdnd00an1n01x5 FILLER_251_1489 ();
 b15zdnd11an1n64x5 FILLER_251_1497 ();
 b15zdnd11an1n64x5 FILLER_251_1561 ();
 b15zdnd11an1n64x5 FILLER_251_1625 ();
 b15zdnd11an1n64x5 FILLER_251_1689 ();
 b15zdnd11an1n32x5 FILLER_251_1753 ();
 b15zdnd00an1n02x5 FILLER_251_1785 ();
 b15zdnd11an1n64x5 FILLER_251_1805 ();
 b15zdnd11an1n64x5 FILLER_251_1869 ();
 b15zdnd11an1n64x5 FILLER_251_1933 ();
 b15zdnd11an1n64x5 FILLER_251_1997 ();
 b15zdnd11an1n32x5 FILLER_251_2061 ();
 b15zdnd11an1n04x5 FILLER_251_2093 ();
 b15zdnd11an1n04x5 FILLER_251_2139 ();
 b15zdnd11an1n64x5 FILLER_251_2185 ();
 b15zdnd11an1n16x5 FILLER_251_2254 ();
 b15zdnd11an1n08x5 FILLER_251_2270 ();
 b15zdnd11an1n04x5 FILLER_251_2278 ();
 b15zdnd00an1n02x5 FILLER_251_2282 ();
 b15zdnd11an1n64x5 FILLER_252_8 ();
 b15zdnd11an1n64x5 FILLER_252_72 ();
 b15zdnd11an1n64x5 FILLER_252_136 ();
 b15zdnd11an1n64x5 FILLER_252_200 ();
 b15zdnd11an1n16x5 FILLER_252_264 ();
 b15zdnd11an1n64x5 FILLER_252_295 ();
 b15zdnd11an1n64x5 FILLER_252_359 ();
 b15zdnd11an1n64x5 FILLER_252_423 ();
 b15zdnd11an1n64x5 FILLER_252_487 ();
 b15zdnd11an1n64x5 FILLER_252_551 ();
 b15zdnd11an1n32x5 FILLER_252_615 ();
 b15zdnd11an1n08x5 FILLER_252_647 ();
 b15zdnd11an1n04x5 FILLER_252_655 ();
 b15zdnd00an1n01x5 FILLER_252_659 ();
 b15zdnd11an1n16x5 FILLER_252_663 ();
 b15zdnd11an1n04x5 FILLER_252_679 ();
 b15zdnd00an1n01x5 FILLER_252_683 ();
 b15zdnd11an1n16x5 FILLER_252_690 ();
 b15zdnd11an1n08x5 FILLER_252_706 ();
 b15zdnd11an1n04x5 FILLER_252_714 ();
 b15zdnd11an1n64x5 FILLER_252_726 ();
 b15zdnd11an1n64x5 FILLER_252_790 ();
 b15zdnd11an1n64x5 FILLER_252_854 ();
 b15zdnd11an1n64x5 FILLER_252_918 ();
 b15zdnd11an1n64x5 FILLER_252_982 ();
 b15zdnd11an1n32x5 FILLER_252_1046 ();
 b15zdnd11an1n16x5 FILLER_252_1078 ();
 b15zdnd11an1n08x5 FILLER_252_1094 ();
 b15zdnd11an1n04x5 FILLER_252_1102 ();
 b15zdnd11an1n16x5 FILLER_252_1126 ();
 b15zdnd11an1n04x5 FILLER_252_1142 ();
 b15zdnd00an1n02x5 FILLER_252_1146 ();
 b15zdnd11an1n64x5 FILLER_252_1162 ();
 b15zdnd11an1n64x5 FILLER_252_1226 ();
 b15zdnd11an1n64x5 FILLER_252_1290 ();
 b15zdnd11an1n64x5 FILLER_252_1354 ();
 b15zdnd11an1n16x5 FILLER_252_1418 ();
 b15zdnd11an1n04x5 FILLER_252_1434 ();
 b15zdnd00an1n01x5 FILLER_252_1438 ();
 b15zdnd11an1n04x5 FILLER_252_1446 ();
 b15zdnd00an1n01x5 FILLER_252_1450 ();
 b15zdnd11an1n04x5 FILLER_252_1454 ();
 b15zdnd11an1n64x5 FILLER_252_1461 ();
 b15zdnd11an1n64x5 FILLER_252_1525 ();
 b15zdnd11an1n16x5 FILLER_252_1589 ();
 b15zdnd11an1n08x5 FILLER_252_1605 ();
 b15zdnd00an1n01x5 FILLER_252_1613 ();
 b15zdnd11an1n32x5 FILLER_252_1636 ();
 b15zdnd11an1n16x5 FILLER_252_1668 ();
 b15zdnd11an1n04x5 FILLER_252_1684 ();
 b15zdnd00an1n01x5 FILLER_252_1688 ();
 b15zdnd11an1n64x5 FILLER_252_1693 ();
 b15zdnd11an1n16x5 FILLER_252_1757 ();
 b15zdnd11an1n08x5 FILLER_252_1773 ();
 b15zdnd11an1n04x5 FILLER_252_1781 ();
 b15zdnd00an1n01x5 FILLER_252_1785 ();
 b15zdnd11an1n64x5 FILLER_252_1801 ();
 b15zdnd11an1n64x5 FILLER_252_1865 ();
 b15zdnd11an1n64x5 FILLER_252_1929 ();
 b15zdnd11an1n64x5 FILLER_252_1993 ();
 b15zdnd11an1n64x5 FILLER_252_2057 ();
 b15zdnd11an1n32x5 FILLER_252_2121 ();
 b15zdnd00an1n01x5 FILLER_252_2153 ();
 b15zdnd11an1n64x5 FILLER_252_2162 ();
 b15zdnd11an1n32x5 FILLER_252_2226 ();
 b15zdnd11an1n16x5 FILLER_252_2258 ();
 b15zdnd00an1n02x5 FILLER_252_2274 ();
 b15zdnd11an1n64x5 FILLER_253_0 ();
 b15zdnd11an1n64x5 FILLER_253_64 ();
 b15zdnd11an1n64x5 FILLER_253_128 ();
 b15zdnd11an1n64x5 FILLER_253_192 ();
 b15zdnd11an1n32x5 FILLER_253_256 ();
 b15zdnd00an1n01x5 FILLER_253_288 ();
 b15zdnd11an1n64x5 FILLER_253_331 ();
 b15zdnd11an1n64x5 FILLER_253_395 ();
 b15zdnd11an1n64x5 FILLER_253_459 ();
 b15zdnd11an1n64x5 FILLER_253_523 ();
 b15zdnd11an1n64x5 FILLER_253_587 ();
 b15zdnd11an1n16x5 FILLER_253_651 ();
 b15zdnd11an1n08x5 FILLER_253_667 ();
 b15zdnd11an1n64x5 FILLER_253_678 ();
 b15zdnd11an1n64x5 FILLER_253_742 ();
 b15zdnd11an1n64x5 FILLER_253_806 ();
 b15zdnd11an1n64x5 FILLER_253_870 ();
 b15zdnd11an1n64x5 FILLER_253_934 ();
 b15zdnd11an1n64x5 FILLER_253_998 ();
 b15zdnd11an1n32x5 FILLER_253_1062 ();
 b15zdnd11an1n04x5 FILLER_253_1094 ();
 b15zdnd00an1n02x5 FILLER_253_1098 ();
 b15zdnd11an1n32x5 FILLER_253_1103 ();
 b15zdnd11an1n16x5 FILLER_253_1135 ();
 b15zdnd11an1n08x5 FILLER_253_1151 ();
 b15zdnd11an1n04x5 FILLER_253_1159 ();
 b15zdnd00an1n02x5 FILLER_253_1163 ();
 b15zdnd00an1n01x5 FILLER_253_1165 ();
 b15zdnd11an1n64x5 FILLER_253_1180 ();
 b15zdnd11an1n64x5 FILLER_253_1244 ();
 b15zdnd11an1n64x5 FILLER_253_1308 ();
 b15zdnd11an1n64x5 FILLER_253_1372 ();
 b15zdnd11an1n08x5 FILLER_253_1436 ();
 b15zdnd11an1n04x5 FILLER_253_1444 ();
 b15zdnd11an1n64x5 FILLER_253_1451 ();
 b15zdnd11an1n16x5 FILLER_253_1515 ();
 b15zdnd11an1n04x5 FILLER_253_1531 ();
 b15zdnd00an1n02x5 FILLER_253_1535 ();
 b15zdnd00an1n01x5 FILLER_253_1537 ();
 b15zdnd11an1n64x5 FILLER_253_1542 ();
 b15zdnd11an1n08x5 FILLER_253_1606 ();
 b15zdnd11an1n04x5 FILLER_253_1614 ();
 b15zdnd11an1n64x5 FILLER_253_1632 ();
 b15zdnd11an1n64x5 FILLER_253_1696 ();
 b15zdnd11an1n64x5 FILLER_253_1760 ();
 b15zdnd11an1n64x5 FILLER_253_1824 ();
 b15zdnd11an1n16x5 FILLER_253_1888 ();
 b15zdnd11an1n08x5 FILLER_253_1904 ();
 b15zdnd00an1n02x5 FILLER_253_1912 ();
 b15zdnd00an1n01x5 FILLER_253_1914 ();
 b15zdnd11an1n64x5 FILLER_253_1957 ();
 b15zdnd11an1n64x5 FILLER_253_2021 ();
 b15zdnd11an1n32x5 FILLER_253_2085 ();
 b15zdnd11an1n16x5 FILLER_253_2117 ();
 b15zdnd11an1n08x5 FILLER_253_2133 ();
 b15zdnd11an1n04x5 FILLER_253_2141 ();
 b15zdnd11an1n04x5 FILLER_253_2187 ();
 b15zdnd11an1n32x5 FILLER_253_2222 ();
 b15zdnd11an1n16x5 FILLER_253_2254 ();
 b15zdnd11an1n08x5 FILLER_253_2270 ();
 b15zdnd11an1n04x5 FILLER_253_2278 ();
 b15zdnd00an1n02x5 FILLER_253_2282 ();
 b15zdnd11an1n64x5 FILLER_254_8 ();
 b15zdnd11an1n64x5 FILLER_254_72 ();
 b15zdnd11an1n32x5 FILLER_254_136 ();
 b15zdnd11an1n08x5 FILLER_254_168 ();
 b15zdnd00an1n02x5 FILLER_254_176 ();
 b15zdnd00an1n01x5 FILLER_254_178 ();
 b15zdnd11an1n04x5 FILLER_254_182 ();
 b15zdnd11an1n04x5 FILLER_254_189 ();
 b15zdnd11an1n64x5 FILLER_254_196 ();
 b15zdnd11an1n16x5 FILLER_254_260 ();
 b15zdnd11an1n08x5 FILLER_254_276 ();
 b15zdnd00an1n02x5 FILLER_254_284 ();
 b15zdnd11an1n04x5 FILLER_254_292 ();
 b15zdnd11an1n64x5 FILLER_254_300 ();
 b15zdnd11an1n64x5 FILLER_254_364 ();
 b15zdnd11an1n64x5 FILLER_254_428 ();
 b15zdnd11an1n64x5 FILLER_254_492 ();
 b15zdnd11an1n64x5 FILLER_254_556 ();
 b15zdnd11an1n64x5 FILLER_254_620 ();
 b15zdnd11an1n32x5 FILLER_254_684 ();
 b15zdnd00an1n02x5 FILLER_254_716 ();
 b15zdnd11an1n64x5 FILLER_254_726 ();
 b15zdnd11an1n64x5 FILLER_254_790 ();
 b15zdnd11an1n64x5 FILLER_254_854 ();
 b15zdnd11an1n64x5 FILLER_254_918 ();
 b15zdnd11an1n64x5 FILLER_254_982 ();
 b15zdnd11an1n64x5 FILLER_254_1046 ();
 b15zdnd11an1n32x5 FILLER_254_1110 ();
 b15zdnd11an1n04x5 FILLER_254_1142 ();
 b15zdnd00an1n02x5 FILLER_254_1146 ();
 b15zdnd11an1n04x5 FILLER_254_1157 ();
 b15zdnd11an1n64x5 FILLER_254_1172 ();
 b15zdnd11an1n64x5 FILLER_254_1236 ();
 b15zdnd11an1n64x5 FILLER_254_1300 ();
 b15zdnd11an1n64x5 FILLER_254_1364 ();
 b15zdnd11an1n64x5 FILLER_254_1428 ();
 b15zdnd11an1n64x5 FILLER_254_1492 ();
 b15zdnd11an1n32x5 FILLER_254_1556 ();
 b15zdnd11an1n08x5 FILLER_254_1588 ();
 b15zdnd00an1n01x5 FILLER_254_1596 ();
 b15zdnd11an1n32x5 FILLER_254_1601 ();
 b15zdnd11an1n08x5 FILLER_254_1633 ();
 b15zdnd00an1n02x5 FILLER_254_1641 ();
 b15zdnd00an1n01x5 FILLER_254_1643 ();
 b15zdnd11an1n16x5 FILLER_254_1648 ();
 b15zdnd11an1n04x5 FILLER_254_1664 ();
 b15zdnd00an1n02x5 FILLER_254_1668 ();
 b15zdnd00an1n01x5 FILLER_254_1670 ();
 b15zdnd11an1n64x5 FILLER_254_1675 ();
 b15zdnd11an1n64x5 FILLER_254_1739 ();
 b15zdnd11an1n64x5 FILLER_254_1803 ();
 b15zdnd11an1n64x5 FILLER_254_1867 ();
 b15zdnd11an1n64x5 FILLER_254_1931 ();
 b15zdnd11an1n64x5 FILLER_254_1995 ();
 b15zdnd11an1n64x5 FILLER_254_2059 ();
 b15zdnd11an1n16x5 FILLER_254_2123 ();
 b15zdnd11an1n08x5 FILLER_254_2139 ();
 b15zdnd11an1n04x5 FILLER_254_2147 ();
 b15zdnd00an1n02x5 FILLER_254_2151 ();
 b15zdnd00an1n01x5 FILLER_254_2153 ();
 b15zdnd11an1n16x5 FILLER_254_2162 ();
 b15zdnd11an1n04x5 FILLER_254_2178 ();
 b15zdnd00an1n01x5 FILLER_254_2182 ();
 b15zdnd11an1n32x5 FILLER_254_2225 ();
 b15zdnd11an1n16x5 FILLER_254_2257 ();
 b15zdnd00an1n02x5 FILLER_254_2273 ();
 b15zdnd00an1n01x5 FILLER_254_2275 ();
 b15zdnd11an1n64x5 FILLER_255_0 ();
 b15zdnd11an1n64x5 FILLER_255_64 ();
 b15zdnd11an1n32x5 FILLER_255_128 ();
 b15zdnd11an1n16x5 FILLER_255_160 ();
 b15zdnd11an1n32x5 FILLER_255_218 ();
 b15zdnd11an1n16x5 FILLER_255_250 ();
 b15zdnd11an1n04x5 FILLER_255_266 ();
 b15zdnd00an1n02x5 FILLER_255_270 ();
 b15zdnd11an1n64x5 FILLER_255_314 ();
 b15zdnd11an1n32x5 FILLER_255_378 ();
 b15zdnd11an1n16x5 FILLER_255_410 ();
 b15zdnd11an1n04x5 FILLER_255_426 ();
 b15zdnd00an1n02x5 FILLER_255_430 ();
 b15zdnd00an1n01x5 FILLER_255_432 ();
 b15zdnd11an1n64x5 FILLER_255_436 ();
 b15zdnd11an1n64x5 FILLER_255_500 ();
 b15zdnd11an1n64x5 FILLER_255_564 ();
 b15zdnd11an1n64x5 FILLER_255_628 ();
 b15zdnd11an1n64x5 FILLER_255_692 ();
 b15zdnd11an1n64x5 FILLER_255_756 ();
 b15zdnd11an1n64x5 FILLER_255_820 ();
 b15zdnd11an1n64x5 FILLER_255_884 ();
 b15zdnd11an1n64x5 FILLER_255_948 ();
 b15zdnd11an1n08x5 FILLER_255_1012 ();
 b15zdnd11an1n04x5 FILLER_255_1020 ();
 b15zdnd11an1n64x5 FILLER_255_1028 ();
 b15zdnd11an1n64x5 FILLER_255_1092 ();
 b15zdnd11an1n64x5 FILLER_255_1176 ();
 b15zdnd11an1n32x5 FILLER_255_1240 ();
 b15zdnd11an1n08x5 FILLER_255_1272 ();
 b15zdnd00an1n02x5 FILLER_255_1280 ();
 b15zdnd11an1n64x5 FILLER_255_1306 ();
 b15zdnd11an1n64x5 FILLER_255_1370 ();
 b15zdnd11an1n64x5 FILLER_255_1434 ();
 b15zdnd00an1n01x5 FILLER_255_1498 ();
 b15zdnd11an1n64x5 FILLER_255_1503 ();
 b15zdnd11an1n64x5 FILLER_255_1567 ();
 b15zdnd11an1n32x5 FILLER_255_1631 ();
 b15zdnd11an1n08x5 FILLER_255_1663 ();
 b15zdnd00an1n02x5 FILLER_255_1671 ();
 b15zdnd00an1n01x5 FILLER_255_1673 ();
 b15zdnd11an1n64x5 FILLER_255_1680 ();
 b15zdnd11an1n32x5 FILLER_255_1744 ();
 b15zdnd11an1n16x5 FILLER_255_1776 ();
 b15zdnd11an1n08x5 FILLER_255_1792 ();
 b15zdnd00an1n01x5 FILLER_255_1800 ();
 b15zdnd11an1n64x5 FILLER_255_1843 ();
 b15zdnd11an1n64x5 FILLER_255_1907 ();
 b15zdnd11an1n64x5 FILLER_255_1971 ();
 b15zdnd11an1n64x5 FILLER_255_2035 ();
 b15zdnd11an1n64x5 FILLER_255_2099 ();
 b15zdnd11an1n64x5 FILLER_255_2163 ();
 b15zdnd11an1n32x5 FILLER_255_2227 ();
 b15zdnd11an1n16x5 FILLER_255_2259 ();
 b15zdnd11an1n08x5 FILLER_255_2275 ();
 b15zdnd00an1n01x5 FILLER_255_2283 ();
 b15zdnd11an1n64x5 FILLER_256_8 ();
 b15zdnd11an1n64x5 FILLER_256_72 ();
 b15zdnd11an1n16x5 FILLER_256_136 ();
 b15zdnd11an1n08x5 FILLER_256_152 ();
 b15zdnd11an1n32x5 FILLER_256_212 ();
 b15zdnd11an1n08x5 FILLER_256_244 ();
 b15zdnd11an1n04x5 FILLER_256_252 ();
 b15zdnd11an1n04x5 FILLER_256_259 ();
 b15zdnd00an1n02x5 FILLER_256_263 ();
 b15zdnd00an1n01x5 FILLER_256_265 ();
 b15zdnd11an1n04x5 FILLER_256_276 ();
 b15zdnd00an1n02x5 FILLER_256_280 ();
 b15zdnd11an1n04x5 FILLER_256_291 ();
 b15zdnd11an1n64x5 FILLER_256_302 ();
 b15zdnd11an1n32x5 FILLER_256_366 ();
 b15zdnd11an1n08x5 FILLER_256_398 ();
 b15zdnd11an1n64x5 FILLER_256_458 ();
 b15zdnd11an1n64x5 FILLER_256_522 ();
 b15zdnd11an1n64x5 FILLER_256_586 ();
 b15zdnd11an1n64x5 FILLER_256_650 ();
 b15zdnd11an1n04x5 FILLER_256_714 ();
 b15zdnd11an1n64x5 FILLER_256_726 ();
 b15zdnd11an1n64x5 FILLER_256_790 ();
 b15zdnd11an1n64x5 FILLER_256_854 ();
 b15zdnd11an1n64x5 FILLER_256_918 ();
 b15zdnd11an1n32x5 FILLER_256_982 ();
 b15zdnd00an1n02x5 FILLER_256_1014 ();
 b15zdnd00an1n01x5 FILLER_256_1016 ();
 b15zdnd11an1n64x5 FILLER_256_1027 ();
 b15zdnd11an1n64x5 FILLER_256_1091 ();
 b15zdnd11an1n64x5 FILLER_256_1155 ();
 b15zdnd11an1n64x5 FILLER_256_1219 ();
 b15zdnd11an1n64x5 FILLER_256_1283 ();
 b15zdnd11an1n64x5 FILLER_256_1347 ();
 b15zdnd11an1n64x5 FILLER_256_1411 ();
 b15zdnd11an1n64x5 FILLER_256_1475 ();
 b15zdnd11an1n16x5 FILLER_256_1539 ();
 b15zdnd11an1n04x5 FILLER_256_1555 ();
 b15zdnd00an1n02x5 FILLER_256_1559 ();
 b15zdnd11an1n64x5 FILLER_256_1584 ();
 b15zdnd11an1n64x5 FILLER_256_1648 ();
 b15zdnd11an1n64x5 FILLER_256_1712 ();
 b15zdnd11an1n08x5 FILLER_256_1776 ();
 b15zdnd00an1n01x5 FILLER_256_1784 ();
 b15zdnd11an1n64x5 FILLER_256_1837 ();
 b15zdnd11an1n64x5 FILLER_256_1901 ();
 b15zdnd11an1n64x5 FILLER_256_1965 ();
 b15zdnd11an1n64x5 FILLER_256_2029 ();
 b15zdnd11an1n16x5 FILLER_256_2093 ();
 b15zdnd11an1n08x5 FILLER_256_2109 ();
 b15zdnd11an1n04x5 FILLER_256_2117 ();
 b15zdnd00an1n01x5 FILLER_256_2121 ();
 b15zdnd11an1n16x5 FILLER_256_2136 ();
 b15zdnd00an1n02x5 FILLER_256_2152 ();
 b15zdnd11an1n64x5 FILLER_256_2162 ();
 b15zdnd11an1n32x5 FILLER_256_2226 ();
 b15zdnd11an1n16x5 FILLER_256_2258 ();
 b15zdnd00an1n02x5 FILLER_256_2274 ();
 b15zdnd11an1n64x5 FILLER_257_0 ();
 b15zdnd11an1n64x5 FILLER_257_64 ();
 b15zdnd11an1n64x5 FILLER_257_128 ();
 b15zdnd11an1n16x5 FILLER_257_192 ();
 b15zdnd00an1n02x5 FILLER_257_208 ();
 b15zdnd00an1n01x5 FILLER_257_210 ();
 b15zdnd11an1n04x5 FILLER_257_225 ();
 b15zdnd11an1n04x5 FILLER_257_281 ();
 b15zdnd11an1n64x5 FILLER_257_327 ();
 b15zdnd11an1n32x5 FILLER_257_391 ();
 b15zdnd00an1n01x5 FILLER_257_423 ();
 b15zdnd11an1n04x5 FILLER_257_427 ();
 b15zdnd11an1n08x5 FILLER_257_434 ();
 b15zdnd00an1n02x5 FILLER_257_442 ();
 b15zdnd00an1n01x5 FILLER_257_444 ();
 b15zdnd11an1n08x5 FILLER_257_448 ();
 b15zdnd00an1n02x5 FILLER_257_456 ();
 b15zdnd00an1n01x5 FILLER_257_458 ();
 b15zdnd11an1n64x5 FILLER_257_501 ();
 b15zdnd11an1n64x5 FILLER_257_565 ();
 b15zdnd11an1n64x5 FILLER_257_629 ();
 b15zdnd11an1n64x5 FILLER_257_693 ();
 b15zdnd11an1n64x5 FILLER_257_757 ();
 b15zdnd11an1n16x5 FILLER_257_821 ();
 b15zdnd00an1n02x5 FILLER_257_837 ();
 b15zdnd11an1n64x5 FILLER_257_842 ();
 b15zdnd11an1n64x5 FILLER_257_906 ();
 b15zdnd11an1n64x5 FILLER_257_970 ();
 b15zdnd11an1n64x5 FILLER_257_1034 ();
 b15zdnd11an1n64x5 FILLER_257_1098 ();
 b15zdnd11an1n64x5 FILLER_257_1162 ();
 b15zdnd11an1n64x5 FILLER_257_1226 ();
 b15zdnd11an1n64x5 FILLER_257_1290 ();
 b15zdnd11an1n64x5 FILLER_257_1354 ();
 b15zdnd11an1n64x5 FILLER_257_1418 ();
 b15zdnd11an1n64x5 FILLER_257_1482 ();
 b15zdnd11an1n64x5 FILLER_257_1546 ();
 b15zdnd11an1n64x5 FILLER_257_1610 ();
 b15zdnd11an1n64x5 FILLER_257_1674 ();
 b15zdnd11an1n32x5 FILLER_257_1738 ();
 b15zdnd11an1n08x5 FILLER_257_1770 ();
 b15zdnd00an1n01x5 FILLER_257_1778 ();
 b15zdnd11an1n04x5 FILLER_257_1818 ();
 b15zdnd11an1n64x5 FILLER_257_1829 ();
 b15zdnd11an1n32x5 FILLER_257_1893 ();
 b15zdnd11an1n08x5 FILLER_257_1925 ();
 b15zdnd11an1n04x5 FILLER_257_1933 ();
 b15zdnd00an1n02x5 FILLER_257_1937 ();
 b15zdnd00an1n01x5 FILLER_257_1939 ();
 b15zdnd11an1n32x5 FILLER_257_1982 ();
 b15zdnd11an1n16x5 FILLER_257_2014 ();
 b15zdnd00an1n02x5 FILLER_257_2030 ();
 b15zdnd00an1n01x5 FILLER_257_2032 ();
 b15zdnd11an1n04x5 FILLER_257_2036 ();
 b15zdnd11an1n64x5 FILLER_257_2043 ();
 b15zdnd11an1n32x5 FILLER_257_2107 ();
 b15zdnd11an1n16x5 FILLER_257_2139 ();
 b15zdnd11an1n08x5 FILLER_257_2155 ();
 b15zdnd11an1n04x5 FILLER_257_2163 ();
 b15zdnd11an1n64x5 FILLER_257_2176 ();
 b15zdnd00an1n02x5 FILLER_257_2240 ();
 b15zdnd11an1n08x5 FILLER_257_2246 ();
 b15zdnd11an1n08x5 FILLER_257_2258 ();
 b15zdnd11an1n04x5 FILLER_257_2266 ();
 b15zdnd11an1n08x5 FILLER_257_2274 ();
 b15zdnd00an1n02x5 FILLER_257_2282 ();
 b15zdnd11an1n64x5 FILLER_258_8 ();
 b15zdnd11an1n64x5 FILLER_258_72 ();
 b15zdnd11an1n64x5 FILLER_258_136 ();
 b15zdnd11an1n32x5 FILLER_258_200 ();
 b15zdnd11an1n08x5 FILLER_258_232 ();
 b15zdnd11an1n04x5 FILLER_258_240 ();
 b15zdnd00an1n02x5 FILLER_258_244 ();
 b15zdnd00an1n01x5 FILLER_258_246 ();
 b15zdnd11an1n04x5 FILLER_258_250 ();
 b15zdnd11an1n04x5 FILLER_258_257 ();
 b15zdnd00an1n01x5 FILLER_258_261 ();
 b15zdnd11an1n64x5 FILLER_258_304 ();
 b15zdnd11an1n32x5 FILLER_258_368 ();
 b15zdnd11an1n04x5 FILLER_258_400 ();
 b15zdnd00an1n01x5 FILLER_258_404 ();
 b15zdnd11an1n04x5 FILLER_258_416 ();
 b15zdnd11an1n64x5 FILLER_258_472 ();
 b15zdnd11an1n64x5 FILLER_258_536 ();
 b15zdnd11an1n64x5 FILLER_258_600 ();
 b15zdnd11an1n32x5 FILLER_258_664 ();
 b15zdnd11an1n16x5 FILLER_258_696 ();
 b15zdnd11an1n04x5 FILLER_258_712 ();
 b15zdnd00an1n02x5 FILLER_258_716 ();
 b15zdnd11an1n64x5 FILLER_258_726 ();
 b15zdnd11an1n16x5 FILLER_258_790 ();
 b15zdnd11an1n04x5 FILLER_258_806 ();
 b15zdnd00an1n02x5 FILLER_258_810 ();
 b15zdnd11an1n32x5 FILLER_258_864 ();
 b15zdnd11an1n16x5 FILLER_258_896 ();
 b15zdnd11an1n08x5 FILLER_258_912 ();
 b15zdnd11an1n16x5 FILLER_258_932 ();
 b15zdnd11an1n08x5 FILLER_258_948 ();
 b15zdnd11an1n04x5 FILLER_258_956 ();
 b15zdnd00an1n01x5 FILLER_258_960 ();
 b15zdnd11an1n32x5 FILLER_258_969 ();
 b15zdnd11an1n08x5 FILLER_258_1001 ();
 b15zdnd11an1n04x5 FILLER_258_1009 ();
 b15zdnd00an1n01x5 FILLER_258_1013 ();
 b15zdnd11an1n64x5 FILLER_258_1017 ();
 b15zdnd11an1n64x5 FILLER_258_1081 ();
 b15zdnd11an1n64x5 FILLER_258_1145 ();
 b15zdnd11an1n32x5 FILLER_258_1209 ();
 b15zdnd11an1n08x5 FILLER_258_1241 ();
 b15zdnd00an1n02x5 FILLER_258_1249 ();
 b15zdnd00an1n01x5 FILLER_258_1251 ();
 b15zdnd11an1n64x5 FILLER_258_1264 ();
 b15zdnd11an1n04x5 FILLER_258_1328 ();
 b15zdnd00an1n01x5 FILLER_258_1332 ();
 b15zdnd11an1n64x5 FILLER_258_1347 ();
 b15zdnd11an1n64x5 FILLER_258_1411 ();
 b15zdnd11an1n64x5 FILLER_258_1475 ();
 b15zdnd11an1n64x5 FILLER_258_1539 ();
 b15zdnd11an1n16x5 FILLER_258_1603 ();
 b15zdnd11an1n08x5 FILLER_258_1619 ();
 b15zdnd11an1n08x5 FILLER_258_1634 ();
 b15zdnd00an1n02x5 FILLER_258_1642 ();
 b15zdnd00an1n01x5 FILLER_258_1644 ();
 b15zdnd11an1n64x5 FILLER_258_1649 ();
 b15zdnd11an1n64x5 FILLER_258_1713 ();
 b15zdnd11an1n08x5 FILLER_258_1777 ();
 b15zdnd11an1n08x5 FILLER_258_1793 ();
 b15zdnd00an1n01x5 FILLER_258_1801 ();
 b15zdnd11an1n04x5 FILLER_258_1805 ();
 b15zdnd11an1n04x5 FILLER_258_1812 ();
 b15zdnd00an1n01x5 FILLER_258_1816 ();
 b15zdnd11an1n64x5 FILLER_258_1820 ();
 b15zdnd11an1n64x5 FILLER_258_1884 ();
 b15zdnd11an1n32x5 FILLER_258_1948 ();
 b15zdnd11an1n16x5 FILLER_258_1980 ();
 b15zdnd11an1n08x5 FILLER_258_1996 ();
 b15zdnd11an1n04x5 FILLER_258_2004 ();
 b15zdnd11an1n32x5 FILLER_258_2060 ();
 b15zdnd11an1n16x5 FILLER_258_2092 ();
 b15zdnd11an1n04x5 FILLER_258_2108 ();
 b15zdnd00an1n02x5 FILLER_258_2112 ();
 b15zdnd11an1n16x5 FILLER_258_2138 ();
 b15zdnd11an1n64x5 FILLER_258_2162 ();
 b15zdnd11an1n04x5 FILLER_258_2226 ();
 b15zdnd00an1n02x5 FILLER_258_2230 ();
 b15zdnd00an1n02x5 FILLER_258_2274 ();
 b15zdnd11an1n08x5 FILLER_259_0 ();
 b15zdnd00an1n01x5 FILLER_259_8 ();
 b15zdnd11an1n64x5 FILLER_259_13 ();
 b15zdnd11an1n64x5 FILLER_259_77 ();
 b15zdnd11an1n32x5 FILLER_259_141 ();
 b15zdnd11an1n16x5 FILLER_259_173 ();
 b15zdnd11an1n08x5 FILLER_259_189 ();
 b15zdnd11an1n04x5 FILLER_259_197 ();
 b15zdnd00an1n02x5 FILLER_259_201 ();
 b15zdnd00an1n01x5 FILLER_259_203 ();
 b15zdnd11an1n32x5 FILLER_259_218 ();
 b15zdnd00an1n01x5 FILLER_259_250 ();
 b15zdnd11an1n04x5 FILLER_259_293 ();
 b15zdnd11an1n64x5 FILLER_259_305 ();
 b15zdnd11an1n32x5 FILLER_259_369 ();
 b15zdnd11an1n16x5 FILLER_259_401 ();
 b15zdnd11an1n04x5 FILLER_259_417 ();
 b15zdnd11an1n08x5 FILLER_259_428 ();
 b15zdnd00an1n02x5 FILLER_259_436 ();
 b15zdnd11an1n04x5 FILLER_259_441 ();
 b15zdnd11an1n16x5 FILLER_259_448 ();
 b15zdnd11an1n04x5 FILLER_259_464 ();
 b15zdnd00an1n02x5 FILLER_259_468 ();
 b15zdnd11an1n32x5 FILLER_259_477 ();
 b15zdnd11an1n16x5 FILLER_259_509 ();
 b15zdnd11an1n08x5 FILLER_259_525 ();
 b15zdnd00an1n02x5 FILLER_259_533 ();
 b15zdnd00an1n01x5 FILLER_259_535 ();
 b15zdnd11an1n04x5 FILLER_259_539 ();
 b15zdnd11an1n16x5 FILLER_259_546 ();
 b15zdnd00an1n02x5 FILLER_259_562 ();
 b15zdnd11an1n64x5 FILLER_259_568 ();
 b15zdnd11an1n64x5 FILLER_259_632 ();
 b15zdnd11an1n64x5 FILLER_259_696 ();
 b15zdnd11an1n64x5 FILLER_259_760 ();
 b15zdnd11an1n04x5 FILLER_259_824 ();
 b15zdnd00an1n02x5 FILLER_259_828 ();
 b15zdnd11an1n04x5 FILLER_259_833 ();
 b15zdnd11an1n16x5 FILLER_259_840 ();
 b15zdnd11an1n04x5 FILLER_259_856 ();
 b15zdnd00an1n02x5 FILLER_259_860 ();
 b15zdnd11an1n64x5 FILLER_259_865 ();
 b15zdnd00an1n01x5 FILLER_259_929 ();
 b15zdnd11an1n16x5 FILLER_259_956 ();
 b15zdnd11an1n04x5 FILLER_259_972 ();
 b15zdnd11an1n04x5 FILLER_259_1016 ();
 b15zdnd11an1n64x5 FILLER_259_1034 ();
 b15zdnd11an1n64x5 FILLER_259_1098 ();
 b15zdnd11an1n32x5 FILLER_259_1162 ();
 b15zdnd11an1n16x5 FILLER_259_1194 ();
 b15zdnd11an1n08x5 FILLER_259_1210 ();
 b15zdnd00an1n02x5 FILLER_259_1218 ();
 b15zdnd11an1n04x5 FILLER_259_1223 ();
 b15zdnd11an1n32x5 FILLER_259_1230 ();
 b15zdnd11an1n16x5 FILLER_259_1262 ();
 b15zdnd11an1n08x5 FILLER_259_1278 ();
 b15zdnd00an1n02x5 FILLER_259_1286 ();
 b15zdnd00an1n01x5 FILLER_259_1288 ();
 b15zdnd11an1n16x5 FILLER_259_1309 ();
 b15zdnd00an1n01x5 FILLER_259_1325 ();
 b15zdnd11an1n64x5 FILLER_259_1337 ();
 b15zdnd11an1n64x5 FILLER_259_1401 ();
 b15zdnd11an1n64x5 FILLER_259_1465 ();
 b15zdnd11an1n64x5 FILLER_259_1529 ();
 b15zdnd11an1n16x5 FILLER_259_1593 ();
 b15zdnd11an1n08x5 FILLER_259_1609 ();
 b15zdnd11an1n04x5 FILLER_259_1617 ();
 b15zdnd00an1n02x5 FILLER_259_1621 ();
 b15zdnd11an1n64x5 FILLER_259_1631 ();
 b15zdnd11an1n64x5 FILLER_259_1695 ();
 b15zdnd11an1n64x5 FILLER_259_1759 ();
 b15zdnd11an1n64x5 FILLER_259_1823 ();
 b15zdnd11an1n64x5 FILLER_259_1887 ();
 b15zdnd11an1n64x5 FILLER_259_1951 ();
 b15zdnd11an1n16x5 FILLER_259_2015 ();
 b15zdnd00an1n02x5 FILLER_259_2031 ();
 b15zdnd11an1n64x5 FILLER_259_2036 ();
 b15zdnd11an1n64x5 FILLER_259_2100 ();
 b15zdnd11an1n64x5 FILLER_259_2164 ();
 b15zdnd11an1n08x5 FILLER_259_2228 ();
 b15zdnd11an1n04x5 FILLER_259_2236 ();
 b15zdnd00an1n02x5 FILLER_259_2282 ();
 b15zdnd11an1n64x5 FILLER_260_8 ();
 b15zdnd11an1n64x5 FILLER_260_72 ();
 b15zdnd11an1n64x5 FILLER_260_136 ();
 b15zdnd11an1n64x5 FILLER_260_200 ();
 b15zdnd11an1n08x5 FILLER_260_264 ();
 b15zdnd11an1n04x5 FILLER_260_272 ();
 b15zdnd00an1n02x5 FILLER_260_276 ();
 b15zdnd00an1n01x5 FILLER_260_278 ();
 b15zdnd11an1n64x5 FILLER_260_289 ();
 b15zdnd11an1n64x5 FILLER_260_353 ();
 b15zdnd11an1n32x5 FILLER_260_417 ();
 b15zdnd11an1n08x5 FILLER_260_449 ();
 b15zdnd00an1n01x5 FILLER_260_457 ();
 b15zdnd11an1n16x5 FILLER_260_489 ();
 b15zdnd11an1n08x5 FILLER_260_505 ();
 b15zdnd11an1n04x5 FILLER_260_513 ();
 b15zdnd00an1n01x5 FILLER_260_517 ();
 b15zdnd11an1n04x5 FILLER_260_570 ();
 b15zdnd11an1n64x5 FILLER_260_616 ();
 b15zdnd11an1n32x5 FILLER_260_680 ();
 b15zdnd11an1n04x5 FILLER_260_712 ();
 b15zdnd00an1n02x5 FILLER_260_716 ();
 b15zdnd11an1n64x5 FILLER_260_726 ();
 b15zdnd11an1n32x5 FILLER_260_790 ();
 b15zdnd11an1n08x5 FILLER_260_822 ();
 b15zdnd11an1n04x5 FILLER_260_830 ();
 b15zdnd00an1n01x5 FILLER_260_834 ();
 b15zdnd11an1n64x5 FILLER_260_887 ();
 b15zdnd11an1n08x5 FILLER_260_951 ();
 b15zdnd11an1n04x5 FILLER_260_959 ();
 b15zdnd11an1n16x5 FILLER_260_977 ();
 b15zdnd11an1n08x5 FILLER_260_993 ();
 b15zdnd11an1n04x5 FILLER_260_1001 ();
 b15zdnd00an1n02x5 FILLER_260_1005 ();
 b15zdnd00an1n01x5 FILLER_260_1007 ();
 b15zdnd11an1n08x5 FILLER_260_1011 ();
 b15zdnd11an1n16x5 FILLER_260_1032 ();
 b15zdnd11an1n04x5 FILLER_260_1048 ();
 b15zdnd00an1n02x5 FILLER_260_1052 ();
 b15zdnd11an1n16x5 FILLER_260_1070 ();
 b15zdnd11an1n08x5 FILLER_260_1086 ();
 b15zdnd00an1n01x5 FILLER_260_1094 ();
 b15zdnd11an1n64x5 FILLER_260_1107 ();
 b15zdnd11an1n16x5 FILLER_260_1171 ();
 b15zdnd11an1n08x5 FILLER_260_1187 ();
 b15zdnd11an1n16x5 FILLER_260_1247 ();
 b15zdnd11an1n08x5 FILLER_260_1263 ();
 b15zdnd11an1n04x5 FILLER_260_1271 ();
 b15zdnd00an1n02x5 FILLER_260_1275 ();
 b15zdnd00an1n01x5 FILLER_260_1277 ();
 b15zdnd11an1n64x5 FILLER_260_1289 ();
 b15zdnd11an1n16x5 FILLER_260_1353 ();
 b15zdnd11an1n04x5 FILLER_260_1369 ();
 b15zdnd00an1n01x5 FILLER_260_1373 ();
 b15zdnd11an1n64x5 FILLER_260_1386 ();
 b15zdnd11an1n64x5 FILLER_260_1450 ();
 b15zdnd11an1n64x5 FILLER_260_1514 ();
 b15zdnd11an1n08x5 FILLER_260_1578 ();
 b15zdnd00an1n02x5 FILLER_260_1586 ();
 b15zdnd00an1n01x5 FILLER_260_1588 ();
 b15zdnd11an1n16x5 FILLER_260_1598 ();
 b15zdnd11an1n08x5 FILLER_260_1614 ();
 b15zdnd00an1n02x5 FILLER_260_1622 ();
 b15zdnd11an1n16x5 FILLER_260_1635 ();
 b15zdnd11an1n08x5 FILLER_260_1651 ();
 b15zdnd11an1n04x5 FILLER_260_1659 ();
 b15zdnd11an1n16x5 FILLER_260_1670 ();
 b15zdnd11an1n04x5 FILLER_260_1686 ();
 b15zdnd00an1n02x5 FILLER_260_1690 ();
 b15zdnd11an1n04x5 FILLER_260_1731 ();
 b15zdnd11an1n64x5 FILLER_260_1742 ();
 b15zdnd11an1n64x5 FILLER_260_1806 ();
 b15zdnd11an1n64x5 FILLER_260_1870 ();
 b15zdnd11an1n64x5 FILLER_260_1934 ();
 b15zdnd11an1n64x5 FILLER_260_1998 ();
 b15zdnd11an1n64x5 FILLER_260_2062 ();
 b15zdnd11an1n16x5 FILLER_260_2126 ();
 b15zdnd11an1n08x5 FILLER_260_2142 ();
 b15zdnd11an1n04x5 FILLER_260_2150 ();
 b15zdnd11an1n64x5 FILLER_260_2162 ();
 b15zdnd11an1n32x5 FILLER_260_2226 ();
 b15zdnd11an1n16x5 FILLER_260_2258 ();
 b15zdnd00an1n02x5 FILLER_260_2274 ();
 b15zdnd11an1n64x5 FILLER_261_0 ();
 b15zdnd11an1n64x5 FILLER_261_64 ();
 b15zdnd11an1n64x5 FILLER_261_128 ();
 b15zdnd11an1n64x5 FILLER_261_192 ();
 b15zdnd11an1n64x5 FILLER_261_256 ();
 b15zdnd11an1n64x5 FILLER_261_320 ();
 b15zdnd11an1n64x5 FILLER_261_384 ();
 b15zdnd11an1n64x5 FILLER_261_448 ();
 b15zdnd11an1n32x5 FILLER_261_512 ();
 b15zdnd11an1n04x5 FILLER_261_544 ();
 b15zdnd11an1n64x5 FILLER_261_551 ();
 b15zdnd11an1n64x5 FILLER_261_615 ();
 b15zdnd11an1n16x5 FILLER_261_679 ();
 b15zdnd11an1n08x5 FILLER_261_695 ();
 b15zdnd00an1n02x5 FILLER_261_703 ();
 b15zdnd11an1n64x5 FILLER_261_733 ();
 b15zdnd11an1n32x5 FILLER_261_797 ();
 b15zdnd11an1n16x5 FILLER_261_829 ();
 b15zdnd11an1n08x5 FILLER_261_845 ();
 b15zdnd11an1n04x5 FILLER_261_856 ();
 b15zdnd11an1n64x5 FILLER_261_863 ();
 b15zdnd11an1n64x5 FILLER_261_927 ();
 b15zdnd11an1n16x5 FILLER_261_991 ();
 b15zdnd11an1n04x5 FILLER_261_1007 ();
 b15zdnd11an1n04x5 FILLER_261_1016 ();
 b15zdnd00an1n02x5 FILLER_261_1020 ();
 b15zdnd11an1n04x5 FILLER_261_1026 ();
 b15zdnd11an1n64x5 FILLER_261_1035 ();
 b15zdnd11an1n64x5 FILLER_261_1099 ();
 b15zdnd11an1n32x5 FILLER_261_1163 ();
 b15zdnd11an1n16x5 FILLER_261_1195 ();
 b15zdnd11an1n08x5 FILLER_261_1211 ();
 b15zdnd00an1n01x5 FILLER_261_1219 ();
 b15zdnd11an1n64x5 FILLER_261_1223 ();
 b15zdnd11an1n64x5 FILLER_261_1287 ();
 b15zdnd11an1n64x5 FILLER_261_1351 ();
 b15zdnd11an1n64x5 FILLER_261_1415 ();
 b15zdnd11an1n32x5 FILLER_261_1479 ();
 b15zdnd11an1n16x5 FILLER_261_1511 ();
 b15zdnd00an1n02x5 FILLER_261_1527 ();
 b15zdnd00an1n01x5 FILLER_261_1529 ();
 b15zdnd11an1n04x5 FILLER_261_1569 ();
 b15zdnd11an1n04x5 FILLER_261_1576 ();
 b15zdnd11an1n16x5 FILLER_261_1607 ();
 b15zdnd11an1n64x5 FILLER_261_1627 ();
 b15zdnd00an1n02x5 FILLER_261_1691 ();
 b15zdnd00an1n01x5 FILLER_261_1693 ();
 b15zdnd11an1n64x5 FILLER_261_1698 ();
 b15zdnd11an1n64x5 FILLER_261_1762 ();
 b15zdnd11an1n64x5 FILLER_261_1826 ();
 b15zdnd11an1n64x5 FILLER_261_1890 ();
 b15zdnd11an1n64x5 FILLER_261_1954 ();
 b15zdnd11an1n32x5 FILLER_261_2018 ();
 b15zdnd11an1n16x5 FILLER_261_2050 ();
 b15zdnd00an1n02x5 FILLER_261_2066 ();
 b15zdnd11an1n16x5 FILLER_261_2080 ();
 b15zdnd11an1n04x5 FILLER_261_2096 ();
 b15zdnd00an1n01x5 FILLER_261_2100 ();
 b15zdnd11an1n04x5 FILLER_261_2104 ();
 b15zdnd11an1n04x5 FILLER_261_2111 ();
 b15zdnd11an1n64x5 FILLER_261_2120 ();
 b15zdnd11an1n64x5 FILLER_261_2184 ();
 b15zdnd00an1n02x5 FILLER_261_2248 ();
 b15zdnd11an1n16x5 FILLER_261_2256 ();
 b15zdnd11an1n08x5 FILLER_261_2272 ();
 b15zdnd11an1n04x5 FILLER_261_2280 ();
 b15zdnd11an1n04x5 FILLER_262_8 ();
 b15zdnd00an1n02x5 FILLER_262_12 ();
 b15zdnd00an1n01x5 FILLER_262_14 ();
 b15zdnd11an1n64x5 FILLER_262_21 ();
 b15zdnd11an1n64x5 FILLER_262_85 ();
 b15zdnd11an1n64x5 FILLER_262_149 ();
 b15zdnd11an1n64x5 FILLER_262_213 ();
 b15zdnd11an1n64x5 FILLER_262_277 ();
 b15zdnd11an1n64x5 FILLER_262_341 ();
 b15zdnd11an1n64x5 FILLER_262_405 ();
 b15zdnd11an1n64x5 FILLER_262_469 ();
 b15zdnd11an1n04x5 FILLER_262_533 ();
 b15zdnd00an1n02x5 FILLER_262_537 ();
 b15zdnd00an1n01x5 FILLER_262_539 ();
 b15zdnd11an1n64x5 FILLER_262_546 ();
 b15zdnd11an1n64x5 FILLER_262_610 ();
 b15zdnd11an1n32x5 FILLER_262_674 ();
 b15zdnd11an1n08x5 FILLER_262_706 ();
 b15zdnd11an1n04x5 FILLER_262_714 ();
 b15zdnd00an1n02x5 FILLER_262_726 ();
 b15zdnd11an1n64x5 FILLER_262_731 ();
 b15zdnd11an1n64x5 FILLER_262_795 ();
 b15zdnd11an1n64x5 FILLER_262_859 ();
 b15zdnd11an1n32x5 FILLER_262_923 ();
 b15zdnd11an1n16x5 FILLER_262_955 ();
 b15zdnd11an1n08x5 FILLER_262_971 ();
 b15zdnd00an1n02x5 FILLER_262_979 ();
 b15zdnd00an1n01x5 FILLER_262_981 ();
 b15zdnd11an1n64x5 FILLER_262_1024 ();
 b15zdnd11an1n64x5 FILLER_262_1088 ();
 b15zdnd11an1n64x5 FILLER_262_1152 ();
 b15zdnd11an1n64x5 FILLER_262_1216 ();
 b15zdnd11an1n64x5 FILLER_262_1280 ();
 b15zdnd11an1n64x5 FILLER_262_1344 ();
 b15zdnd11an1n64x5 FILLER_262_1408 ();
 b15zdnd11an1n32x5 FILLER_262_1472 ();
 b15zdnd11an1n04x5 FILLER_262_1549 ();
 b15zdnd11an1n64x5 FILLER_262_1557 ();
 b15zdnd11an1n64x5 FILLER_262_1621 ();
 b15zdnd11an1n64x5 FILLER_262_1685 ();
 b15zdnd11an1n64x5 FILLER_262_1749 ();
 b15zdnd11an1n64x5 FILLER_262_1813 ();
 b15zdnd11an1n64x5 FILLER_262_1877 ();
 b15zdnd11an1n64x5 FILLER_262_1941 ();
 b15zdnd11an1n64x5 FILLER_262_2005 ();
 b15zdnd00an1n02x5 FILLER_262_2069 ();
 b15zdnd00an1n01x5 FILLER_262_2071 ();
 b15zdnd11an1n04x5 FILLER_262_2079 ();
 b15zdnd11an1n16x5 FILLER_262_2135 ();
 b15zdnd00an1n02x5 FILLER_262_2151 ();
 b15zdnd00an1n01x5 FILLER_262_2153 ();
 b15zdnd11an1n64x5 FILLER_262_2162 ();
 b15zdnd11an1n16x5 FILLER_262_2226 ();
 b15zdnd11an1n08x5 FILLER_262_2242 ();
 b15zdnd11an1n04x5 FILLER_262_2250 ();
 b15zdnd00an1n02x5 FILLER_262_2254 ();
 b15zdnd11an1n16x5 FILLER_262_2260 ();
 b15zdnd11an1n64x5 FILLER_263_0 ();
 b15zdnd11an1n64x5 FILLER_263_64 ();
 b15zdnd11an1n64x5 FILLER_263_128 ();
 b15zdnd11an1n64x5 FILLER_263_192 ();
 b15zdnd11an1n64x5 FILLER_263_256 ();
 b15zdnd11an1n64x5 FILLER_263_320 ();
 b15zdnd11an1n64x5 FILLER_263_384 ();
 b15zdnd11an1n64x5 FILLER_263_448 ();
 b15zdnd11an1n08x5 FILLER_263_512 ();
 b15zdnd11an1n04x5 FILLER_263_520 ();
 b15zdnd00an1n01x5 FILLER_263_524 ();
 b15zdnd11an1n64x5 FILLER_263_567 ();
 b15zdnd11an1n64x5 FILLER_263_631 ();
 b15zdnd11an1n32x5 FILLER_263_695 ();
 b15zdnd11an1n64x5 FILLER_263_730 ();
 b15zdnd11an1n64x5 FILLER_263_794 ();
 b15zdnd11an1n64x5 FILLER_263_858 ();
 b15zdnd11an1n16x5 FILLER_263_922 ();
 b15zdnd00an1n02x5 FILLER_263_938 ();
 b15zdnd11an1n64x5 FILLER_263_943 ();
 b15zdnd11an1n64x5 FILLER_263_1007 ();
 b15zdnd11an1n16x5 FILLER_263_1071 ();
 b15zdnd11an1n04x5 FILLER_263_1087 ();
 b15zdnd11an1n64x5 FILLER_263_1122 ();
 b15zdnd11an1n64x5 FILLER_263_1186 ();
 b15zdnd11an1n16x5 FILLER_263_1250 ();
 b15zdnd11an1n04x5 FILLER_263_1266 ();
 b15zdnd11an1n64x5 FILLER_263_1282 ();
 b15zdnd11an1n64x5 FILLER_263_1346 ();
 b15zdnd11an1n64x5 FILLER_263_1410 ();
 b15zdnd11an1n64x5 FILLER_263_1474 ();
 b15zdnd11an1n64x5 FILLER_263_1538 ();
 b15zdnd11an1n64x5 FILLER_263_1602 ();
 b15zdnd11an1n64x5 FILLER_263_1666 ();
 b15zdnd11an1n64x5 FILLER_263_1730 ();
 b15zdnd11an1n64x5 FILLER_263_1794 ();
 b15zdnd11an1n64x5 FILLER_263_1858 ();
 b15zdnd11an1n32x5 FILLER_263_1922 ();
 b15zdnd00an1n02x5 FILLER_263_1954 ();
 b15zdnd00an1n01x5 FILLER_263_1956 ();
 b15zdnd11an1n64x5 FILLER_263_1972 ();
 b15zdnd11an1n16x5 FILLER_263_2036 ();
 b15zdnd11an1n04x5 FILLER_263_2052 ();
 b15zdnd00an1n02x5 FILLER_263_2056 ();
 b15zdnd11an1n32x5 FILLER_263_2064 ();
 b15zdnd11an1n08x5 FILLER_263_2096 ();
 b15zdnd11an1n04x5 FILLER_263_2104 ();
 b15zdnd11an1n04x5 FILLER_263_2111 ();
 b15zdnd11an1n32x5 FILLER_263_2120 ();
 b15zdnd00an1n02x5 FILLER_263_2152 ();
 b15zdnd11an1n64x5 FILLER_263_2160 ();
 b15zdnd11an1n32x5 FILLER_263_2224 ();
 b15zdnd11an1n16x5 FILLER_263_2256 ();
 b15zdnd11an1n08x5 FILLER_263_2272 ();
 b15zdnd11an1n04x5 FILLER_263_2280 ();
 b15zdnd11an1n64x5 FILLER_264_8 ();
 b15zdnd11an1n64x5 FILLER_264_72 ();
 b15zdnd11an1n64x5 FILLER_264_136 ();
 b15zdnd11an1n64x5 FILLER_264_200 ();
 b15zdnd11an1n64x5 FILLER_264_264 ();
 b15zdnd11an1n64x5 FILLER_264_328 ();
 b15zdnd11an1n64x5 FILLER_264_392 ();
 b15zdnd11an1n32x5 FILLER_264_456 ();
 b15zdnd11an1n08x5 FILLER_264_488 ();
 b15zdnd00an1n02x5 FILLER_264_496 ();
 b15zdnd00an1n01x5 FILLER_264_498 ();
 b15zdnd11an1n08x5 FILLER_264_504 ();
 b15zdnd00an1n02x5 FILLER_264_512 ();
 b15zdnd11an1n64x5 FILLER_264_519 ();
 b15zdnd11an1n64x5 FILLER_264_583 ();
 b15zdnd11an1n64x5 FILLER_264_647 ();
 b15zdnd11an1n04x5 FILLER_264_711 ();
 b15zdnd00an1n02x5 FILLER_264_715 ();
 b15zdnd00an1n01x5 FILLER_264_717 ();
 b15zdnd11an1n64x5 FILLER_264_726 ();
 b15zdnd11an1n64x5 FILLER_264_790 ();
 b15zdnd11an1n64x5 FILLER_264_854 ();
 b15zdnd11an1n04x5 FILLER_264_918 ();
 b15zdnd11an1n64x5 FILLER_264_974 ();
 b15zdnd11an1n64x5 FILLER_264_1038 ();
 b15zdnd11an1n64x5 FILLER_264_1102 ();
 b15zdnd11an1n64x5 FILLER_264_1166 ();
 b15zdnd11an1n64x5 FILLER_264_1230 ();
 b15zdnd11an1n64x5 FILLER_264_1294 ();
 b15zdnd11an1n64x5 FILLER_264_1358 ();
 b15zdnd11an1n64x5 FILLER_264_1422 ();
 b15zdnd11an1n64x5 FILLER_264_1486 ();
 b15zdnd11an1n64x5 FILLER_264_1550 ();
 b15zdnd11an1n64x5 FILLER_264_1614 ();
 b15zdnd11an1n64x5 FILLER_264_1678 ();
 b15zdnd11an1n64x5 FILLER_264_1742 ();
 b15zdnd11an1n64x5 FILLER_264_1806 ();
 b15zdnd11an1n64x5 FILLER_264_1870 ();
 b15zdnd11an1n08x5 FILLER_264_1934 ();
 b15zdnd00an1n01x5 FILLER_264_1942 ();
 b15zdnd11an1n04x5 FILLER_264_1946 ();
 b15zdnd11an1n16x5 FILLER_264_1953 ();
 b15zdnd00an1n01x5 FILLER_264_1969 ();
 b15zdnd11an1n64x5 FILLER_264_2012 ();
 b15zdnd11an1n64x5 FILLER_264_2076 ();
 b15zdnd11an1n08x5 FILLER_264_2140 ();
 b15zdnd11an1n04x5 FILLER_264_2148 ();
 b15zdnd00an1n02x5 FILLER_264_2152 ();
 b15zdnd11an1n64x5 FILLER_264_2162 ();
 b15zdnd11an1n32x5 FILLER_264_2226 ();
 b15zdnd11an1n16x5 FILLER_264_2258 ();
 b15zdnd00an1n02x5 FILLER_264_2274 ();
 b15zdnd11an1n64x5 FILLER_265_0 ();
 b15zdnd11an1n64x5 FILLER_265_64 ();
 b15zdnd11an1n64x5 FILLER_265_128 ();
 b15zdnd11an1n64x5 FILLER_265_192 ();
 b15zdnd11an1n64x5 FILLER_265_256 ();
 b15zdnd11an1n64x5 FILLER_265_320 ();
 b15zdnd11an1n64x5 FILLER_265_384 ();
 b15zdnd11an1n64x5 FILLER_265_448 ();
 b15zdnd11an1n04x5 FILLER_265_512 ();
 b15zdnd00an1n02x5 FILLER_265_516 ();
 b15zdnd00an1n01x5 FILLER_265_518 ();
 b15zdnd11an1n64x5 FILLER_265_561 ();
 b15zdnd11an1n64x5 FILLER_265_625 ();
 b15zdnd11an1n64x5 FILLER_265_689 ();
 b15zdnd11an1n64x5 FILLER_265_753 ();
 b15zdnd11an1n64x5 FILLER_265_817 ();
 b15zdnd11an1n32x5 FILLER_265_881 ();
 b15zdnd11an1n08x5 FILLER_265_913 ();
 b15zdnd00an1n02x5 FILLER_265_921 ();
 b15zdnd00an1n01x5 FILLER_265_923 ();
 b15zdnd11an1n16x5 FILLER_265_927 ();
 b15zdnd11an1n04x5 FILLER_265_943 ();
 b15zdnd11an1n64x5 FILLER_265_950 ();
 b15zdnd11an1n04x5 FILLER_265_1025 ();
 b15zdnd11an1n64x5 FILLER_265_1032 ();
 b15zdnd11an1n64x5 FILLER_265_1096 ();
 b15zdnd11an1n64x5 FILLER_265_1160 ();
 b15zdnd11an1n64x5 FILLER_265_1224 ();
 b15zdnd11an1n64x5 FILLER_265_1288 ();
 b15zdnd11an1n64x5 FILLER_265_1352 ();
 b15zdnd11an1n64x5 FILLER_265_1416 ();
 b15zdnd11an1n32x5 FILLER_265_1480 ();
 b15zdnd11an1n08x5 FILLER_265_1512 ();
 b15zdnd00an1n01x5 FILLER_265_1520 ();
 b15zdnd11an1n64x5 FILLER_265_1532 ();
 b15zdnd11an1n64x5 FILLER_265_1596 ();
 b15zdnd11an1n64x5 FILLER_265_1660 ();
 b15zdnd11an1n64x5 FILLER_265_1724 ();
 b15zdnd11an1n64x5 FILLER_265_1788 ();
 b15zdnd11an1n64x5 FILLER_265_1852 ();
 b15zdnd11an1n08x5 FILLER_265_1916 ();
 b15zdnd00an1n01x5 FILLER_265_1924 ();
 b15zdnd11an1n64x5 FILLER_265_1977 ();
 b15zdnd11an1n64x5 FILLER_265_2041 ();
 b15zdnd11an1n16x5 FILLER_265_2105 ();
 b15zdnd11an1n64x5 FILLER_265_2130 ();
 b15zdnd11an1n64x5 FILLER_265_2194 ();
 b15zdnd11an1n16x5 FILLER_265_2258 ();
 b15zdnd11an1n08x5 FILLER_265_2274 ();
 b15zdnd00an1n02x5 FILLER_265_2282 ();
 b15zdnd11an1n64x5 FILLER_266_8 ();
 b15zdnd11an1n64x5 FILLER_266_72 ();
 b15zdnd11an1n64x5 FILLER_266_136 ();
 b15zdnd11an1n64x5 FILLER_266_200 ();
 b15zdnd11an1n64x5 FILLER_266_264 ();
 b15zdnd11an1n64x5 FILLER_266_328 ();
 b15zdnd11an1n64x5 FILLER_266_392 ();
 b15zdnd11an1n64x5 FILLER_266_456 ();
 b15zdnd11an1n64x5 FILLER_266_520 ();
 b15zdnd11an1n64x5 FILLER_266_584 ();
 b15zdnd11an1n64x5 FILLER_266_648 ();
 b15zdnd11an1n04x5 FILLER_266_712 ();
 b15zdnd00an1n02x5 FILLER_266_716 ();
 b15zdnd11an1n16x5 FILLER_266_726 ();
 b15zdnd11an1n64x5 FILLER_266_745 ();
 b15zdnd11an1n64x5 FILLER_266_809 ();
 b15zdnd11an1n64x5 FILLER_266_873 ();
 b15zdnd11an1n64x5 FILLER_266_937 ();
 b15zdnd11an1n64x5 FILLER_266_1001 ();
 b15zdnd11an1n32x5 FILLER_266_1065 ();
 b15zdnd11an1n04x5 FILLER_266_1097 ();
 b15zdnd11an1n64x5 FILLER_266_1127 ();
 b15zdnd11an1n64x5 FILLER_266_1191 ();
 b15zdnd11an1n64x5 FILLER_266_1255 ();
 b15zdnd11an1n64x5 FILLER_266_1319 ();
 b15zdnd11an1n64x5 FILLER_266_1383 ();
 b15zdnd11an1n64x5 FILLER_266_1447 ();
 b15zdnd11an1n64x5 FILLER_266_1511 ();
 b15zdnd11an1n64x5 FILLER_266_1575 ();
 b15zdnd11an1n64x5 FILLER_266_1639 ();
 b15zdnd11an1n64x5 FILLER_266_1703 ();
 b15zdnd11an1n64x5 FILLER_266_1767 ();
 b15zdnd11an1n64x5 FILLER_266_1831 ();
 b15zdnd11an1n32x5 FILLER_266_1895 ();
 b15zdnd00an1n01x5 FILLER_266_1927 ();
 b15zdnd11an1n64x5 FILLER_266_1970 ();
 b15zdnd11an1n64x5 FILLER_266_2034 ();
 b15zdnd11an1n32x5 FILLER_266_2098 ();
 b15zdnd11an1n16x5 FILLER_266_2130 ();
 b15zdnd11an1n08x5 FILLER_266_2146 ();
 b15zdnd11an1n64x5 FILLER_266_2162 ();
 b15zdnd11an1n32x5 FILLER_266_2226 ();
 b15zdnd11an1n16x5 FILLER_266_2258 ();
 b15zdnd00an1n02x5 FILLER_266_2274 ();
 b15zdnd11an1n64x5 FILLER_267_0 ();
 b15zdnd11an1n64x5 FILLER_267_64 ();
 b15zdnd11an1n64x5 FILLER_267_128 ();
 b15zdnd11an1n64x5 FILLER_267_192 ();
 b15zdnd11an1n16x5 FILLER_267_256 ();
 b15zdnd11an1n08x5 FILLER_267_272 ();
 b15zdnd00an1n02x5 FILLER_267_280 ();
 b15zdnd00an1n01x5 FILLER_267_282 ();
 b15zdnd11an1n64x5 FILLER_267_325 ();
 b15zdnd11an1n64x5 FILLER_267_389 ();
 b15zdnd11an1n64x5 FILLER_267_453 ();
 b15zdnd11an1n64x5 FILLER_267_517 ();
 b15zdnd11an1n64x5 FILLER_267_581 ();
 b15zdnd11an1n64x5 FILLER_267_645 ();
 b15zdnd11an1n16x5 FILLER_267_709 ();
 b15zdnd11an1n04x5 FILLER_267_725 ();
 b15zdnd11an1n64x5 FILLER_267_750 ();
 b15zdnd11an1n16x5 FILLER_267_814 ();
 b15zdnd00an1n01x5 FILLER_267_830 ();
 b15zdnd11an1n64x5 FILLER_267_875 ();
 b15zdnd11an1n64x5 FILLER_267_939 ();
 b15zdnd11an1n64x5 FILLER_267_1003 ();
 b15zdnd11an1n64x5 FILLER_267_1067 ();
 b15zdnd11an1n16x5 FILLER_267_1131 ();
 b15zdnd11an1n04x5 FILLER_267_1147 ();
 b15zdnd00an1n02x5 FILLER_267_1151 ();
 b15zdnd11an1n64x5 FILLER_267_1156 ();
 b15zdnd11an1n64x5 FILLER_267_1220 ();
 b15zdnd11an1n16x5 FILLER_267_1284 ();
 b15zdnd11an1n04x5 FILLER_267_1300 ();
 b15zdnd11an1n04x5 FILLER_267_1316 ();
 b15zdnd11an1n04x5 FILLER_267_1323 ();
 b15zdnd11an1n64x5 FILLER_267_1330 ();
 b15zdnd11an1n64x5 FILLER_267_1394 ();
 b15zdnd11an1n16x5 FILLER_267_1458 ();
 b15zdnd11an1n08x5 FILLER_267_1474 ();
 b15zdnd11an1n04x5 FILLER_267_1482 ();
 b15zdnd00an1n01x5 FILLER_267_1486 ();
 b15zdnd11an1n64x5 FILLER_267_1490 ();
 b15zdnd11an1n64x5 FILLER_267_1554 ();
 b15zdnd11an1n64x5 FILLER_267_1618 ();
 b15zdnd11an1n64x5 FILLER_267_1682 ();
 b15zdnd11an1n64x5 FILLER_267_1746 ();
 b15zdnd11an1n64x5 FILLER_267_1810 ();
 b15zdnd11an1n32x5 FILLER_267_1874 ();
 b15zdnd11an1n16x5 FILLER_267_1906 ();
 b15zdnd00an1n02x5 FILLER_267_1922 ();
 b15zdnd11an1n04x5 FILLER_267_1930 ();
 b15zdnd00an1n02x5 FILLER_267_1934 ();
 b15zdnd00an1n01x5 FILLER_267_1936 ();
 b15zdnd11an1n64x5 FILLER_267_1979 ();
 b15zdnd11an1n64x5 FILLER_267_2043 ();
 b15zdnd11an1n32x5 FILLER_267_2107 ();
 b15zdnd11an1n16x5 FILLER_267_2139 ();
 b15zdnd11an1n64x5 FILLER_267_2164 ();
 b15zdnd11an1n32x5 FILLER_267_2228 ();
 b15zdnd11an1n16x5 FILLER_267_2260 ();
 b15zdnd11an1n08x5 FILLER_267_2276 ();
 b15zdnd11an1n04x5 FILLER_268_8 ();
 b15zdnd00an1n02x5 FILLER_268_12 ();
 b15zdnd11an1n64x5 FILLER_268_18 ();
 b15zdnd11an1n64x5 FILLER_268_82 ();
 b15zdnd11an1n64x5 FILLER_268_146 ();
 b15zdnd11an1n64x5 FILLER_268_210 ();
 b15zdnd11an1n64x5 FILLER_268_274 ();
 b15zdnd11an1n64x5 FILLER_268_338 ();
 b15zdnd11an1n64x5 FILLER_268_402 ();
 b15zdnd11an1n08x5 FILLER_268_466 ();
 b15zdnd11an1n04x5 FILLER_268_474 ();
 b15zdnd11an1n64x5 FILLER_268_496 ();
 b15zdnd11an1n64x5 FILLER_268_560 ();
 b15zdnd11an1n64x5 FILLER_268_624 ();
 b15zdnd11an1n16x5 FILLER_268_688 ();
 b15zdnd11an1n08x5 FILLER_268_704 ();
 b15zdnd11an1n04x5 FILLER_268_712 ();
 b15zdnd00an1n02x5 FILLER_268_716 ();
 b15zdnd11an1n04x5 FILLER_268_726 ();
 b15zdnd11an1n64x5 FILLER_268_734 ();
 b15zdnd11an1n32x5 FILLER_268_798 ();
 b15zdnd11an1n16x5 FILLER_268_830 ();
 b15zdnd11an1n04x5 FILLER_268_846 ();
 b15zdnd00an1n01x5 FILLER_268_850 ();
 b15zdnd11an1n04x5 FILLER_268_854 ();
 b15zdnd11an1n64x5 FILLER_268_861 ();
 b15zdnd11an1n32x5 FILLER_268_925 ();
 b15zdnd11an1n16x5 FILLER_268_957 ();
 b15zdnd11an1n08x5 FILLER_268_973 ();
 b15zdnd11an1n04x5 FILLER_268_981 ();
 b15zdnd00an1n02x5 FILLER_268_985 ();
 b15zdnd11an1n64x5 FILLER_268_1010 ();
 b15zdnd11an1n32x5 FILLER_268_1074 ();
 b15zdnd11an1n16x5 FILLER_268_1106 ();
 b15zdnd11an1n08x5 FILLER_268_1122 ();
 b15zdnd00an1n02x5 FILLER_268_1130 ();
 b15zdnd11an1n16x5 FILLER_268_1184 ();
 b15zdnd11an1n64x5 FILLER_268_1220 ();
 b15zdnd00an1n02x5 FILLER_268_1284 ();
 b15zdnd11an1n32x5 FILLER_268_1326 ();
 b15zdnd11an1n16x5 FILLER_268_1358 ();
 b15zdnd11an1n04x5 FILLER_268_1374 ();
 b15zdnd00an1n02x5 FILLER_268_1378 ();
 b15zdnd00an1n01x5 FILLER_268_1380 ();
 b15zdnd11an1n64x5 FILLER_268_1389 ();
 b15zdnd11an1n32x5 FILLER_268_1453 ();
 b15zdnd00an1n01x5 FILLER_268_1485 ();
 b15zdnd11an1n04x5 FILLER_268_1489 ();
 b15zdnd11an1n64x5 FILLER_268_1496 ();
 b15zdnd11an1n64x5 FILLER_268_1560 ();
 b15zdnd11an1n64x5 FILLER_268_1624 ();
 b15zdnd11an1n64x5 FILLER_268_1688 ();
 b15zdnd11an1n64x5 FILLER_268_1752 ();
 b15zdnd11an1n64x5 FILLER_268_1816 ();
 b15zdnd11an1n32x5 FILLER_268_1880 ();
 b15zdnd11an1n08x5 FILLER_268_1912 ();
 b15zdnd11an1n04x5 FILLER_268_1920 ();
 b15zdnd00an1n02x5 FILLER_268_1924 ();
 b15zdnd00an1n01x5 FILLER_268_1926 ();
 b15zdnd11an1n16x5 FILLER_268_1930 ();
 b15zdnd11an1n04x5 FILLER_268_1946 ();
 b15zdnd11an1n64x5 FILLER_268_1953 ();
 b15zdnd11an1n64x5 FILLER_268_2017 ();
 b15zdnd11an1n64x5 FILLER_268_2081 ();
 b15zdnd11an1n08x5 FILLER_268_2145 ();
 b15zdnd00an1n01x5 FILLER_268_2153 ();
 b15zdnd11an1n64x5 FILLER_268_2162 ();
 b15zdnd11an1n32x5 FILLER_268_2226 ();
 b15zdnd11an1n16x5 FILLER_268_2258 ();
 b15zdnd00an1n02x5 FILLER_268_2274 ();
 b15zdnd11an1n64x5 FILLER_269_0 ();
 b15zdnd11an1n64x5 FILLER_269_64 ();
 b15zdnd11an1n64x5 FILLER_269_128 ();
 b15zdnd11an1n64x5 FILLER_269_192 ();
 b15zdnd11an1n64x5 FILLER_269_256 ();
 b15zdnd11an1n64x5 FILLER_269_320 ();
 b15zdnd11an1n64x5 FILLER_269_384 ();
 b15zdnd11an1n32x5 FILLER_269_448 ();
 b15zdnd11an1n08x5 FILLER_269_480 ();
 b15zdnd00an1n01x5 FILLER_269_488 ();
 b15zdnd11an1n04x5 FILLER_269_492 ();
 b15zdnd00an1n02x5 FILLER_269_496 ();
 b15zdnd11an1n64x5 FILLER_269_511 ();
 b15zdnd11an1n64x5 FILLER_269_575 ();
 b15zdnd11an1n64x5 FILLER_269_639 ();
 b15zdnd11an1n16x5 FILLER_269_703 ();
 b15zdnd11an1n04x5 FILLER_269_719 ();
 b15zdnd00an1n02x5 FILLER_269_723 ();
 b15zdnd00an1n01x5 FILLER_269_725 ();
 b15zdnd11an1n64x5 FILLER_269_744 ();
 b15zdnd11an1n32x5 FILLER_269_808 ();
 b15zdnd11an1n08x5 FILLER_269_840 ();
 b15zdnd00an1n02x5 FILLER_269_848 ();
 b15zdnd11an1n16x5 FILLER_269_853 ();
 b15zdnd11an1n64x5 FILLER_269_911 ();
 b15zdnd11an1n16x5 FILLER_269_975 ();
 b15zdnd00an1n02x5 FILLER_269_991 ();
 b15zdnd11an1n64x5 FILLER_269_1010 ();
 b15zdnd11an1n32x5 FILLER_269_1074 ();
 b15zdnd00an1n01x5 FILLER_269_1106 ();
 b15zdnd11an1n04x5 FILLER_269_1114 ();
 b15zdnd00an1n02x5 FILLER_269_1118 ();
 b15zdnd00an1n01x5 FILLER_269_1120 ();
 b15zdnd11an1n64x5 FILLER_269_1163 ();
 b15zdnd11an1n64x5 FILLER_269_1227 ();
 b15zdnd11an1n32x5 FILLER_269_1291 ();
 b15zdnd11an1n08x5 FILLER_269_1323 ();
 b15zdnd11an1n04x5 FILLER_269_1331 ();
 b15zdnd00an1n02x5 FILLER_269_1335 ();
 b15zdnd00an1n01x5 FILLER_269_1337 ();
 b15zdnd11an1n08x5 FILLER_269_1380 ();
 b15zdnd11an1n04x5 FILLER_269_1388 ();
 b15zdnd00an1n01x5 FILLER_269_1392 ();
 b15zdnd11an1n32x5 FILLER_269_1420 ();
 b15zdnd11an1n08x5 FILLER_269_1452 ();
 b15zdnd00an1n01x5 FILLER_269_1460 ();
 b15zdnd11an1n64x5 FILLER_269_1513 ();
 b15zdnd11an1n64x5 FILLER_269_1577 ();
 b15zdnd11an1n04x5 FILLER_269_1641 ();
 b15zdnd00an1n02x5 FILLER_269_1645 ();
 b15zdnd11an1n64x5 FILLER_269_1650 ();
 b15zdnd11an1n64x5 FILLER_269_1714 ();
 b15zdnd11an1n64x5 FILLER_269_1778 ();
 b15zdnd11an1n64x5 FILLER_269_1842 ();
 b15zdnd11an1n64x5 FILLER_269_1906 ();
 b15zdnd11an1n64x5 FILLER_269_1970 ();
 b15zdnd11an1n64x5 FILLER_269_2034 ();
 b15zdnd11an1n64x5 FILLER_269_2098 ();
 b15zdnd11an1n64x5 FILLER_269_2162 ();
 b15zdnd11an1n32x5 FILLER_269_2226 ();
 b15zdnd11an1n16x5 FILLER_269_2258 ();
 b15zdnd11an1n08x5 FILLER_269_2274 ();
 b15zdnd00an1n02x5 FILLER_269_2282 ();
 b15zdnd11an1n64x5 FILLER_270_8 ();
 b15zdnd11an1n64x5 FILLER_270_72 ();
 b15zdnd11an1n64x5 FILLER_270_136 ();
 b15zdnd11an1n64x5 FILLER_270_200 ();
 b15zdnd11an1n64x5 FILLER_270_264 ();
 b15zdnd11an1n64x5 FILLER_270_328 ();
 b15zdnd11an1n64x5 FILLER_270_392 ();
 b15zdnd11an1n16x5 FILLER_270_456 ();
 b15zdnd11an1n08x5 FILLER_270_472 ();
 b15zdnd11an1n04x5 FILLER_270_480 ();
 b15zdnd00an1n02x5 FILLER_270_484 ();
 b15zdnd00an1n01x5 FILLER_270_486 ();
 b15zdnd11an1n04x5 FILLER_270_492 ();
 b15zdnd11an1n64x5 FILLER_270_512 ();
 b15zdnd11an1n64x5 FILLER_270_576 ();
 b15zdnd11an1n64x5 FILLER_270_640 ();
 b15zdnd11an1n08x5 FILLER_270_704 ();
 b15zdnd11an1n04x5 FILLER_270_712 ();
 b15zdnd00an1n02x5 FILLER_270_716 ();
 b15zdnd11an1n64x5 FILLER_270_726 ();
 b15zdnd11an1n64x5 FILLER_270_790 ();
 b15zdnd11an1n64x5 FILLER_270_854 ();
 b15zdnd11an1n64x5 FILLER_270_918 ();
 b15zdnd11an1n64x5 FILLER_270_982 ();
 b15zdnd11an1n64x5 FILLER_270_1046 ();
 b15zdnd11an1n32x5 FILLER_270_1110 ();
 b15zdnd11an1n04x5 FILLER_270_1142 ();
 b15zdnd11an1n04x5 FILLER_270_1149 ();
 b15zdnd11an1n64x5 FILLER_270_1156 ();
 b15zdnd11an1n64x5 FILLER_270_1220 ();
 b15zdnd11an1n64x5 FILLER_270_1284 ();
 b15zdnd11an1n64x5 FILLER_270_1348 ();
 b15zdnd11an1n32x5 FILLER_270_1412 ();
 b15zdnd11an1n16x5 FILLER_270_1444 ();
 b15zdnd11an1n04x5 FILLER_270_1460 ();
 b15zdnd11an1n08x5 FILLER_270_1482 ();
 b15zdnd00an1n01x5 FILLER_270_1490 ();
 b15zdnd11an1n64x5 FILLER_270_1533 ();
 b15zdnd11an1n32x5 FILLER_270_1597 ();
 b15zdnd11an1n08x5 FILLER_270_1629 ();
 b15zdnd11an1n04x5 FILLER_270_1637 ();
 b15zdnd11an1n04x5 FILLER_270_1644 ();
 b15zdnd11an1n64x5 FILLER_270_1651 ();
 b15zdnd11an1n64x5 FILLER_270_1715 ();
 b15zdnd11an1n64x5 FILLER_270_1779 ();
 b15zdnd11an1n64x5 FILLER_270_1843 ();
 b15zdnd11an1n08x5 FILLER_270_1907 ();
 b15zdnd11an1n04x5 FILLER_270_1915 ();
 b15zdnd00an1n01x5 FILLER_270_1919 ();
 b15zdnd11an1n64x5 FILLER_270_1926 ();
 b15zdnd11an1n64x5 FILLER_270_1990 ();
 b15zdnd11an1n64x5 FILLER_270_2054 ();
 b15zdnd11an1n32x5 FILLER_270_2118 ();
 b15zdnd11an1n04x5 FILLER_270_2150 ();
 b15zdnd11an1n64x5 FILLER_270_2162 ();
 b15zdnd11an1n32x5 FILLER_270_2226 ();
 b15zdnd11an1n16x5 FILLER_270_2258 ();
 b15zdnd00an1n02x5 FILLER_270_2274 ();
 b15zdnd11an1n16x5 FILLER_271_0 ();
 b15zdnd11an1n08x5 FILLER_271_16 ();
 b15zdnd11an1n04x5 FILLER_271_24 ();
 b15zdnd00an1n01x5 FILLER_271_28 ();
 b15zdnd11an1n64x5 FILLER_271_33 ();
 b15zdnd11an1n64x5 FILLER_271_97 ();
 b15zdnd11an1n64x5 FILLER_271_161 ();
 b15zdnd11an1n64x5 FILLER_271_225 ();
 b15zdnd11an1n64x5 FILLER_271_289 ();
 b15zdnd11an1n64x5 FILLER_271_353 ();
 b15zdnd11an1n64x5 FILLER_271_417 ();
 b15zdnd11an1n64x5 FILLER_271_481 ();
 b15zdnd11an1n64x5 FILLER_271_545 ();
 b15zdnd11an1n08x5 FILLER_271_609 ();
 b15zdnd11an1n04x5 FILLER_271_617 ();
 b15zdnd00an1n02x5 FILLER_271_621 ();
 b15zdnd11an1n64x5 FILLER_271_626 ();
 b15zdnd11an1n32x5 FILLER_271_690 ();
 b15zdnd11an1n16x5 FILLER_271_722 ();
 b15zdnd00an1n01x5 FILLER_271_738 ();
 b15zdnd11an1n64x5 FILLER_271_745 ();
 b15zdnd11an1n64x5 FILLER_271_809 ();
 b15zdnd11an1n64x5 FILLER_271_873 ();
 b15zdnd11an1n32x5 FILLER_271_937 ();
 b15zdnd11an1n16x5 FILLER_271_969 ();
 b15zdnd00an1n02x5 FILLER_271_985 ();
 b15zdnd11an1n04x5 FILLER_271_994 ();
 b15zdnd11an1n08x5 FILLER_271_1012 ();
 b15zdnd11an1n32x5 FILLER_271_1046 ();
 b15zdnd11an1n16x5 FILLER_271_1078 ();
 b15zdnd11an1n64x5 FILLER_271_1104 ();
 b15zdnd11an1n64x5 FILLER_271_1168 ();
 b15zdnd11an1n64x5 FILLER_271_1232 ();
 b15zdnd00an1n01x5 FILLER_271_1296 ();
 b15zdnd11an1n64x5 FILLER_271_1325 ();
 b15zdnd11an1n64x5 FILLER_271_1389 ();
 b15zdnd11an1n08x5 FILLER_271_1453 ();
 b15zdnd11an1n04x5 FILLER_271_1461 ();
 b15zdnd00an1n02x5 FILLER_271_1465 ();
 b15zdnd11an1n32x5 FILLER_271_1509 ();
 b15zdnd11an1n08x5 FILLER_271_1541 ();
 b15zdnd00an1n01x5 FILLER_271_1549 ();
 b15zdnd11an1n16x5 FILLER_271_1592 ();
 b15zdnd11an1n08x5 FILLER_271_1608 ();
 b15zdnd11an1n04x5 FILLER_271_1616 ();
 b15zdnd00an1n02x5 FILLER_271_1620 ();
 b15zdnd00an1n01x5 FILLER_271_1622 ();
 b15zdnd11an1n64x5 FILLER_271_1675 ();
 b15zdnd11an1n64x5 FILLER_271_1739 ();
 b15zdnd11an1n64x5 FILLER_271_1803 ();
 b15zdnd11an1n64x5 FILLER_271_1867 ();
 b15zdnd11an1n64x5 FILLER_271_1931 ();
 b15zdnd11an1n64x5 FILLER_271_1995 ();
 b15zdnd11an1n64x5 FILLER_271_2059 ();
 b15zdnd11an1n64x5 FILLER_271_2123 ();
 b15zdnd11an1n64x5 FILLER_271_2187 ();
 b15zdnd11an1n32x5 FILLER_271_2251 ();
 b15zdnd00an1n01x5 FILLER_271_2283 ();
 b15zdnd11an1n64x5 FILLER_272_8 ();
 b15zdnd11an1n64x5 FILLER_272_72 ();
 b15zdnd11an1n64x5 FILLER_272_136 ();
 b15zdnd11an1n64x5 FILLER_272_200 ();
 b15zdnd11an1n64x5 FILLER_272_264 ();
 b15zdnd11an1n64x5 FILLER_272_328 ();
 b15zdnd11an1n64x5 FILLER_272_392 ();
 b15zdnd11an1n32x5 FILLER_272_456 ();
 b15zdnd11an1n64x5 FILLER_272_499 ();
 b15zdnd11an1n32x5 FILLER_272_563 ();
 b15zdnd00an1n01x5 FILLER_272_595 ();
 b15zdnd11an1n64x5 FILLER_272_648 ();
 b15zdnd11an1n04x5 FILLER_272_712 ();
 b15zdnd00an1n02x5 FILLER_272_716 ();
 b15zdnd11an1n64x5 FILLER_272_726 ();
 b15zdnd11an1n64x5 FILLER_272_790 ();
 b15zdnd11an1n64x5 FILLER_272_854 ();
 b15zdnd11an1n64x5 FILLER_272_918 ();
 b15zdnd00an1n02x5 FILLER_272_982 ();
 b15zdnd11an1n64x5 FILLER_272_1000 ();
 b15zdnd11an1n64x5 FILLER_272_1064 ();
 b15zdnd11an1n64x5 FILLER_272_1128 ();
 b15zdnd11an1n64x5 FILLER_272_1192 ();
 b15zdnd11an1n64x5 FILLER_272_1256 ();
 b15zdnd11an1n32x5 FILLER_272_1320 ();
 b15zdnd11an1n16x5 FILLER_272_1352 ();
 b15zdnd11an1n08x5 FILLER_272_1368 ();
 b15zdnd00an1n01x5 FILLER_272_1376 ();
 b15zdnd11an1n08x5 FILLER_272_1380 ();
 b15zdnd00an1n02x5 FILLER_272_1388 ();
 b15zdnd00an1n01x5 FILLER_272_1390 ();
 b15zdnd11an1n08x5 FILLER_272_1395 ();
 b15zdnd00an1n02x5 FILLER_272_1403 ();
 b15zdnd00an1n01x5 FILLER_272_1405 ();
 b15zdnd11an1n32x5 FILLER_272_1420 ();
 b15zdnd11an1n08x5 FILLER_272_1455 ();
 b15zdnd11an1n04x5 FILLER_272_1463 ();
 b15zdnd11an1n64x5 FILLER_272_1509 ();
 b15zdnd11an1n64x5 FILLER_272_1573 ();
 b15zdnd11an1n64x5 FILLER_272_1637 ();
 b15zdnd11an1n64x5 FILLER_272_1701 ();
 b15zdnd11an1n64x5 FILLER_272_1765 ();
 b15zdnd11an1n64x5 FILLER_272_1829 ();
 b15zdnd11an1n64x5 FILLER_272_1893 ();
 b15zdnd11an1n64x5 FILLER_272_1957 ();
 b15zdnd11an1n64x5 FILLER_272_2021 ();
 b15zdnd11an1n32x5 FILLER_272_2085 ();
 b15zdnd00an1n02x5 FILLER_272_2117 ();
 b15zdnd00an1n01x5 FILLER_272_2119 ();
 b15zdnd11an1n16x5 FILLER_272_2123 ();
 b15zdnd11an1n08x5 FILLER_272_2139 ();
 b15zdnd11an1n04x5 FILLER_272_2147 ();
 b15zdnd00an1n02x5 FILLER_272_2151 ();
 b15zdnd00an1n01x5 FILLER_272_2153 ();
 b15zdnd11an1n64x5 FILLER_272_2162 ();
 b15zdnd11an1n32x5 FILLER_272_2226 ();
 b15zdnd11an1n16x5 FILLER_272_2258 ();
 b15zdnd00an1n02x5 FILLER_272_2274 ();
 b15zdnd11an1n64x5 FILLER_273_0 ();
 b15zdnd11an1n64x5 FILLER_273_64 ();
 b15zdnd11an1n64x5 FILLER_273_128 ();
 b15zdnd11an1n64x5 FILLER_273_192 ();
 b15zdnd11an1n64x5 FILLER_273_256 ();
 b15zdnd11an1n64x5 FILLER_273_320 ();
 b15zdnd11an1n64x5 FILLER_273_384 ();
 b15zdnd11an1n64x5 FILLER_273_448 ();
 b15zdnd11an1n64x5 FILLER_273_512 ();
 b15zdnd11an1n32x5 FILLER_273_576 ();
 b15zdnd11an1n04x5 FILLER_273_608 ();
 b15zdnd00an1n02x5 FILLER_273_612 ();
 b15zdnd11an1n04x5 FILLER_273_617 ();
 b15zdnd11an1n64x5 FILLER_273_624 ();
 b15zdnd11an1n64x5 FILLER_273_688 ();
 b15zdnd11an1n64x5 FILLER_273_752 ();
 b15zdnd11an1n64x5 FILLER_273_816 ();
 b15zdnd11an1n64x5 FILLER_273_880 ();
 b15zdnd11an1n64x5 FILLER_273_944 ();
 b15zdnd11an1n64x5 FILLER_273_1008 ();
 b15zdnd11an1n64x5 FILLER_273_1072 ();
 b15zdnd11an1n16x5 FILLER_273_1136 ();
 b15zdnd11an1n08x5 FILLER_273_1152 ();
 b15zdnd11an1n04x5 FILLER_273_1160 ();
 b15zdnd00an1n02x5 FILLER_273_1164 ();
 b15zdnd00an1n01x5 FILLER_273_1166 ();
 b15zdnd11an1n64x5 FILLER_273_1209 ();
 b15zdnd11an1n32x5 FILLER_273_1273 ();
 b15zdnd11an1n16x5 FILLER_273_1330 ();
 b15zdnd11an1n08x5 FILLER_273_1346 ();
 b15zdnd11an1n04x5 FILLER_273_1354 ();
 b15zdnd00an1n01x5 FILLER_273_1358 ();
 b15zdnd11an1n08x5 FILLER_273_1363 ();
 b15zdnd11an1n04x5 FILLER_273_1371 ();
 b15zdnd11an1n64x5 FILLER_273_1385 ();
 b15zdnd00an1n02x5 FILLER_273_1449 ();
 b15zdnd00an1n01x5 FILLER_273_1451 ();
 b15zdnd11an1n08x5 FILLER_273_1459 ();
 b15zdnd00an1n02x5 FILLER_273_1467 ();
 b15zdnd00an1n01x5 FILLER_273_1469 ();
 b15zdnd11an1n64x5 FILLER_273_1476 ();
 b15zdnd11an1n64x5 FILLER_273_1540 ();
 b15zdnd11an1n32x5 FILLER_273_1604 ();
 b15zdnd11an1n16x5 FILLER_273_1636 ();
 b15zdnd11an1n08x5 FILLER_273_1652 ();
 b15zdnd00an1n02x5 FILLER_273_1660 ();
 b15zdnd00an1n01x5 FILLER_273_1662 ();
 b15zdnd11an1n64x5 FILLER_273_1683 ();
 b15zdnd11an1n16x5 FILLER_273_1747 ();
 b15zdnd11an1n04x5 FILLER_273_1766 ();
 b15zdnd11an1n64x5 FILLER_273_1773 ();
 b15zdnd11an1n32x5 FILLER_273_1837 ();
 b15zdnd11an1n16x5 FILLER_273_1869 ();
 b15zdnd11an1n04x5 FILLER_273_1885 ();
 b15zdnd00an1n02x5 FILLER_273_1889 ();
 b15zdnd11an1n04x5 FILLER_273_1897 ();
 b15zdnd11an1n04x5 FILLER_273_1908 ();
 b15zdnd11an1n04x5 FILLER_273_1916 ();
 b15zdnd11an1n64x5 FILLER_273_1924 ();
 b15zdnd11an1n32x5 FILLER_273_1988 ();
 b15zdnd00an1n01x5 FILLER_273_2020 ();
 b15zdnd11an1n32x5 FILLER_273_2073 ();
 b15zdnd11an1n08x5 FILLER_273_2105 ();
 b15zdnd00an1n02x5 FILLER_273_2113 ();
 b15zdnd00an1n01x5 FILLER_273_2115 ();
 b15zdnd11an1n64x5 FILLER_273_2125 ();
 b15zdnd11an1n64x5 FILLER_273_2189 ();
 b15zdnd11an1n16x5 FILLER_273_2253 ();
 b15zdnd11an1n08x5 FILLER_273_2269 ();
 b15zdnd11an1n04x5 FILLER_273_2277 ();
 b15zdnd00an1n02x5 FILLER_273_2281 ();
 b15zdnd00an1n01x5 FILLER_273_2283 ();
 b15zdnd11an1n64x5 FILLER_274_8 ();
 b15zdnd11an1n64x5 FILLER_274_72 ();
 b15zdnd11an1n64x5 FILLER_274_136 ();
 b15zdnd11an1n32x5 FILLER_274_200 ();
 b15zdnd11an1n16x5 FILLER_274_232 ();
 b15zdnd11an1n08x5 FILLER_274_248 ();
 b15zdnd11an1n04x5 FILLER_274_256 ();
 b15zdnd11an1n64x5 FILLER_274_263 ();
 b15zdnd11an1n64x5 FILLER_274_327 ();
 b15zdnd11an1n64x5 FILLER_274_391 ();
 b15zdnd11an1n64x5 FILLER_274_455 ();
 b15zdnd11an1n64x5 FILLER_274_519 ();
 b15zdnd11an1n32x5 FILLER_274_583 ();
 b15zdnd00an1n01x5 FILLER_274_615 ();
 b15zdnd11an1n04x5 FILLER_274_619 ();
 b15zdnd11an1n32x5 FILLER_274_665 ();
 b15zdnd11an1n16x5 FILLER_274_697 ();
 b15zdnd11an1n04x5 FILLER_274_713 ();
 b15zdnd00an1n01x5 FILLER_274_717 ();
 b15zdnd11an1n64x5 FILLER_274_726 ();
 b15zdnd11an1n64x5 FILLER_274_790 ();
 b15zdnd11an1n64x5 FILLER_274_854 ();
 b15zdnd11an1n64x5 FILLER_274_918 ();
 b15zdnd00an1n02x5 FILLER_274_982 ();
 b15zdnd11an1n04x5 FILLER_274_992 ();
 b15zdnd00an1n02x5 FILLER_274_996 ();
 b15zdnd11an1n64x5 FILLER_274_1022 ();
 b15zdnd11an1n16x5 FILLER_274_1086 ();
 b15zdnd11an1n08x5 FILLER_274_1102 ();
 b15zdnd11an1n04x5 FILLER_274_1110 ();
 b15zdnd00an1n02x5 FILLER_274_1114 ();
 b15zdnd00an1n01x5 FILLER_274_1116 ();
 b15zdnd11an1n16x5 FILLER_274_1126 ();
 b15zdnd11an1n04x5 FILLER_274_1142 ();
 b15zdnd00an1n02x5 FILLER_274_1146 ();
 b15zdnd00an1n01x5 FILLER_274_1148 ();
 b15zdnd11an1n64x5 FILLER_274_1169 ();
 b15zdnd11an1n64x5 FILLER_274_1233 ();
 b15zdnd11an1n64x5 FILLER_274_1297 ();
 b15zdnd11an1n64x5 FILLER_274_1361 ();
 b15zdnd11an1n32x5 FILLER_274_1425 ();
 b15zdnd11an1n08x5 FILLER_274_1457 ();
 b15zdnd11an1n64x5 FILLER_274_1507 ();
 b15zdnd11an1n32x5 FILLER_274_1571 ();
 b15zdnd11an1n16x5 FILLER_274_1603 ();
 b15zdnd11an1n08x5 FILLER_274_1619 ();
 b15zdnd11an1n04x5 FILLER_274_1627 ();
 b15zdnd11an1n64x5 FILLER_274_1673 ();
 b15zdnd00an1n01x5 FILLER_274_1737 ();
 b15zdnd11an1n64x5 FILLER_274_1790 ();
 b15zdnd11an1n16x5 FILLER_274_1854 ();
 b15zdnd11an1n08x5 FILLER_274_1912 ();
 b15zdnd11an1n16x5 FILLER_274_1962 ();
 b15zdnd11an1n08x5 FILLER_274_1978 ();
 b15zdnd00an1n02x5 FILLER_274_1986 ();
 b15zdnd00an1n01x5 FILLER_274_1988 ();
 b15zdnd11an1n08x5 FILLER_274_2031 ();
 b15zdnd11an1n04x5 FILLER_274_2039 ();
 b15zdnd11an1n04x5 FILLER_274_2046 ();
 b15zdnd11an1n64x5 FILLER_274_2053 ();
 b15zdnd11an1n32x5 FILLER_274_2117 ();
 b15zdnd11an1n04x5 FILLER_274_2149 ();
 b15zdnd00an1n01x5 FILLER_274_2153 ();
 b15zdnd11an1n64x5 FILLER_274_2162 ();
 b15zdnd11an1n32x5 FILLER_274_2226 ();
 b15zdnd11an1n16x5 FILLER_274_2258 ();
 b15zdnd00an1n02x5 FILLER_274_2274 ();
 b15zdnd11an1n64x5 FILLER_275_0 ();
 b15zdnd11an1n64x5 FILLER_275_64 ();
 b15zdnd11an1n64x5 FILLER_275_128 ();
 b15zdnd11an1n32x5 FILLER_275_192 ();
 b15zdnd11an1n08x5 FILLER_275_224 ();
 b15zdnd00an1n01x5 FILLER_275_232 ();
 b15zdnd11an1n64x5 FILLER_275_285 ();
 b15zdnd11an1n64x5 FILLER_275_349 ();
 b15zdnd11an1n64x5 FILLER_275_413 ();
 b15zdnd11an1n64x5 FILLER_275_477 ();
 b15zdnd11an1n64x5 FILLER_275_541 ();
 b15zdnd11an1n04x5 FILLER_275_605 ();
 b15zdnd11an1n04x5 FILLER_275_613 ();
 b15zdnd11an1n64x5 FILLER_275_622 ();
 b15zdnd11an1n64x5 FILLER_275_686 ();
 b15zdnd11an1n64x5 FILLER_275_750 ();
 b15zdnd11an1n64x5 FILLER_275_814 ();
 b15zdnd11an1n64x5 FILLER_275_878 ();
 b15zdnd11an1n32x5 FILLER_275_942 ();
 b15zdnd11an1n08x5 FILLER_275_974 ();
 b15zdnd11an1n04x5 FILLER_275_982 ();
 b15zdnd00an1n01x5 FILLER_275_986 ();
 b15zdnd11an1n64x5 FILLER_275_1011 ();
 b15zdnd11an1n32x5 FILLER_275_1075 ();
 b15zdnd11an1n08x5 FILLER_275_1107 ();
 b15zdnd11an1n04x5 FILLER_275_1126 ();
 b15zdnd11an1n32x5 FILLER_275_1156 ();
 b15zdnd11an1n16x5 FILLER_275_1188 ();
 b15zdnd11an1n08x5 FILLER_275_1204 ();
 b15zdnd11an1n04x5 FILLER_275_1212 ();
 b15zdnd00an1n02x5 FILLER_275_1216 ();
 b15zdnd11an1n64x5 FILLER_275_1260 ();
 b15zdnd11an1n64x5 FILLER_275_1324 ();
 b15zdnd11an1n64x5 FILLER_275_1388 ();
 b15zdnd11an1n08x5 FILLER_275_1452 ();
 b15zdnd11an1n64x5 FILLER_275_1502 ();
 b15zdnd11an1n64x5 FILLER_275_1566 ();
 b15zdnd11an1n64x5 FILLER_275_1630 ();
 b15zdnd11an1n64x5 FILLER_275_1694 ();
 b15zdnd11an1n04x5 FILLER_275_1758 ();
 b15zdnd00an1n02x5 FILLER_275_1762 ();
 b15zdnd11an1n64x5 FILLER_275_1767 ();
 b15zdnd11an1n04x5 FILLER_275_1831 ();
 b15zdnd11an1n04x5 FILLER_275_1887 ();
 b15zdnd00an1n01x5 FILLER_275_1891 ();
 b15zdnd11an1n64x5 FILLER_275_1934 ();
 b15zdnd11an1n32x5 FILLER_275_1998 ();
 b15zdnd11an1n16x5 FILLER_275_2030 ();
 b15zdnd11an1n64x5 FILLER_275_2049 ();
 b15zdnd11an1n08x5 FILLER_275_2113 ();
 b15zdnd00an1n02x5 FILLER_275_2121 ();
 b15zdnd00an1n01x5 FILLER_275_2123 ();
 b15zdnd11an1n64x5 FILLER_275_2127 ();
 b15zdnd11an1n64x5 FILLER_275_2191 ();
 b15zdnd11an1n16x5 FILLER_275_2255 ();
 b15zdnd11an1n08x5 FILLER_275_2271 ();
 b15zdnd11an1n04x5 FILLER_275_2279 ();
 b15zdnd00an1n01x5 FILLER_275_2283 ();
 b15zdnd11an1n64x5 FILLER_276_8 ();
 b15zdnd11an1n64x5 FILLER_276_72 ();
 b15zdnd11an1n64x5 FILLER_276_136 ();
 b15zdnd11an1n32x5 FILLER_276_200 ();
 b15zdnd11an1n16x5 FILLER_276_232 ();
 b15zdnd00an1n02x5 FILLER_276_248 ();
 b15zdnd00an1n01x5 FILLER_276_250 ();
 b15zdnd11an1n04x5 FILLER_276_254 ();
 b15zdnd11an1n64x5 FILLER_276_261 ();
 b15zdnd11an1n64x5 FILLER_276_325 ();
 b15zdnd11an1n64x5 FILLER_276_389 ();
 b15zdnd11an1n32x5 FILLER_276_453 ();
 b15zdnd11an1n08x5 FILLER_276_485 ();
 b15zdnd11an1n04x5 FILLER_276_493 ();
 b15zdnd11an1n64x5 FILLER_276_504 ();
 b15zdnd11an1n32x5 FILLER_276_568 ();
 b15zdnd11an1n08x5 FILLER_276_600 ();
 b15zdnd11an1n64x5 FILLER_276_650 ();
 b15zdnd11an1n04x5 FILLER_276_714 ();
 b15zdnd11an1n64x5 FILLER_276_726 ();
 b15zdnd11an1n64x5 FILLER_276_790 ();
 b15zdnd11an1n16x5 FILLER_276_854 ();
 b15zdnd11an1n08x5 FILLER_276_870 ();
 b15zdnd11an1n04x5 FILLER_276_878 ();
 b15zdnd00an1n02x5 FILLER_276_882 ();
 b15zdnd00an1n01x5 FILLER_276_884 ();
 b15zdnd11an1n16x5 FILLER_276_905 ();
 b15zdnd11an1n04x5 FILLER_276_921 ();
 b15zdnd11an1n32x5 FILLER_276_956 ();
 b15zdnd11an1n08x5 FILLER_276_988 ();
 b15zdnd11an1n64x5 FILLER_276_1012 ();
 b15zdnd11an1n16x5 FILLER_276_1076 ();
 b15zdnd11an1n04x5 FILLER_276_1092 ();
 b15zdnd00an1n01x5 FILLER_276_1096 ();
 b15zdnd11an1n04x5 FILLER_276_1121 ();
 b15zdnd11an1n08x5 FILLER_276_1136 ();
 b15zdnd11an1n04x5 FILLER_276_1144 ();
 b15zdnd00an1n02x5 FILLER_276_1148 ();
 b15zdnd11an1n32x5 FILLER_276_1157 ();
 b15zdnd11an1n08x5 FILLER_276_1189 ();
 b15zdnd11an1n04x5 FILLER_276_1197 ();
 b15zdnd11an1n64x5 FILLER_276_1221 ();
 b15zdnd11an1n64x5 FILLER_276_1285 ();
 b15zdnd11an1n64x5 FILLER_276_1349 ();
 b15zdnd11an1n32x5 FILLER_276_1413 ();
 b15zdnd11an1n04x5 FILLER_276_1445 ();
 b15zdnd00an1n02x5 FILLER_276_1449 ();
 b15zdnd00an1n01x5 FILLER_276_1451 ();
 b15zdnd11an1n64x5 FILLER_276_1456 ();
 b15zdnd11an1n64x5 FILLER_276_1520 ();
 b15zdnd11an1n08x5 FILLER_276_1584 ();
 b15zdnd00an1n02x5 FILLER_276_1592 ();
 b15zdnd11an1n04x5 FILLER_276_1597 ();
 b15zdnd11an1n64x5 FILLER_276_1604 ();
 b15zdnd11an1n64x5 FILLER_276_1668 ();
 b15zdnd11an1n64x5 FILLER_276_1759 ();
 b15zdnd11an1n16x5 FILLER_276_1823 ();
 b15zdnd11an1n08x5 FILLER_276_1839 ();
 b15zdnd11an1n04x5 FILLER_276_1847 ();
 b15zdnd00an1n02x5 FILLER_276_1851 ();
 b15zdnd11an1n04x5 FILLER_276_1856 ();
 b15zdnd11an1n04x5 FILLER_276_1863 ();
 b15zdnd11an1n16x5 FILLER_276_1870 ();
 b15zdnd11an1n04x5 FILLER_276_1886 ();
 b15zdnd00an1n01x5 FILLER_276_1890 ();
 b15zdnd11an1n08x5 FILLER_276_1904 ();
 b15zdnd00an1n02x5 FILLER_276_1912 ();
 b15zdnd00an1n01x5 FILLER_276_1914 ();
 b15zdnd11an1n04x5 FILLER_276_1924 ();
 b15zdnd11an1n64x5 FILLER_276_1935 ();
 b15zdnd11an1n64x5 FILLER_276_1999 ();
 b15zdnd11an1n04x5 FILLER_276_2063 ();
 b15zdnd00an1n02x5 FILLER_276_2067 ();
 b15zdnd11an1n32x5 FILLER_276_2111 ();
 b15zdnd11an1n08x5 FILLER_276_2143 ();
 b15zdnd00an1n02x5 FILLER_276_2151 ();
 b15zdnd00an1n01x5 FILLER_276_2153 ();
 b15zdnd11an1n64x5 FILLER_276_2162 ();
 b15zdnd11an1n32x5 FILLER_276_2226 ();
 b15zdnd11an1n16x5 FILLER_276_2258 ();
 b15zdnd00an1n02x5 FILLER_276_2274 ();
 b15zdnd11an1n64x5 FILLER_277_0 ();
 b15zdnd11an1n64x5 FILLER_277_64 ();
 b15zdnd11an1n64x5 FILLER_277_128 ();
 b15zdnd11an1n64x5 FILLER_277_192 ();
 b15zdnd11an1n64x5 FILLER_277_256 ();
 b15zdnd11an1n64x5 FILLER_277_320 ();
 b15zdnd11an1n16x5 FILLER_277_384 ();
 b15zdnd11an1n08x5 FILLER_277_400 ();
 b15zdnd11an1n64x5 FILLER_277_411 ();
 b15zdnd11an1n16x5 FILLER_277_475 ();
 b15zdnd11an1n08x5 FILLER_277_491 ();
 b15zdnd11an1n04x5 FILLER_277_499 ();
 b15zdnd11an1n64x5 FILLER_277_507 ();
 b15zdnd11an1n16x5 FILLER_277_571 ();
 b15zdnd11an1n08x5 FILLER_277_587 ();
 b15zdnd00an1n01x5 FILLER_277_595 ();
 b15zdnd11an1n04x5 FILLER_277_600 ();
 b15zdnd11an1n64x5 FILLER_277_646 ();
 b15zdnd11an1n64x5 FILLER_277_710 ();
 b15zdnd11an1n64x5 FILLER_277_774 ();
 b15zdnd11an1n32x5 FILLER_277_838 ();
 b15zdnd11an1n08x5 FILLER_277_870 ();
 b15zdnd00an1n02x5 FILLER_277_878 ();
 b15zdnd11an1n32x5 FILLER_277_887 ();
 b15zdnd11an1n08x5 FILLER_277_919 ();
 b15zdnd11an1n64x5 FILLER_277_953 ();
 b15zdnd11an1n64x5 FILLER_277_1017 ();
 b15zdnd11an1n32x5 FILLER_277_1081 ();
 b15zdnd11an1n04x5 FILLER_277_1127 ();
 b15zdnd11an1n08x5 FILLER_277_1136 ();
 b15zdnd11an1n04x5 FILLER_277_1144 ();
 b15zdnd00an1n02x5 FILLER_277_1148 ();
 b15zdnd11an1n64x5 FILLER_277_1176 ();
 b15zdnd11an1n64x5 FILLER_277_1240 ();
 b15zdnd11an1n32x5 FILLER_277_1304 ();
 b15zdnd11an1n16x5 FILLER_277_1336 ();
 b15zdnd00an1n02x5 FILLER_277_1352 ();
 b15zdnd00an1n01x5 FILLER_277_1354 ();
 b15zdnd11an1n64x5 FILLER_277_1358 ();
 b15zdnd11an1n64x5 FILLER_277_1422 ();
 b15zdnd11an1n64x5 FILLER_277_1486 ();
 b15zdnd11an1n16x5 FILLER_277_1550 ();
 b15zdnd00an1n02x5 FILLER_277_1566 ();
 b15zdnd00an1n01x5 FILLER_277_1568 ();
 b15zdnd11an1n64x5 FILLER_277_1621 ();
 b15zdnd11an1n32x5 FILLER_277_1685 ();
 b15zdnd11an1n16x5 FILLER_277_1717 ();
 b15zdnd11an1n08x5 FILLER_277_1733 ();
 b15zdnd11an1n04x5 FILLER_277_1741 ();
 b15zdnd00an1n02x5 FILLER_277_1745 ();
 b15zdnd00an1n01x5 FILLER_277_1747 ();
 b15zdnd11an1n08x5 FILLER_277_1756 ();
 b15zdnd11an1n04x5 FILLER_277_1764 ();
 b15zdnd00an1n02x5 FILLER_277_1768 ();
 b15zdnd00an1n01x5 FILLER_277_1770 ();
 b15zdnd11an1n64x5 FILLER_277_1775 ();
 b15zdnd11an1n32x5 FILLER_277_1839 ();
 b15zdnd11an1n16x5 FILLER_277_1871 ();
 b15zdnd11an1n08x5 FILLER_277_1887 ();
 b15zdnd00an1n01x5 FILLER_277_1895 ();
 b15zdnd11an1n04x5 FILLER_277_1904 ();
 b15zdnd00an1n01x5 FILLER_277_1908 ();
 b15zdnd11an1n64x5 FILLER_277_1916 ();
 b15zdnd11an1n64x5 FILLER_277_1980 ();
 b15zdnd11an1n64x5 FILLER_277_2044 ();
 b15zdnd11an1n16x5 FILLER_277_2108 ();
 b15zdnd11an1n08x5 FILLER_277_2124 ();
 b15zdnd11an1n04x5 FILLER_277_2132 ();
 b15zdnd11an1n64x5 FILLER_277_2143 ();
 b15zdnd11an1n64x5 FILLER_277_2207 ();
 b15zdnd11an1n08x5 FILLER_277_2271 ();
 b15zdnd11an1n04x5 FILLER_277_2279 ();
 b15zdnd00an1n01x5 FILLER_277_2283 ();
 b15zdnd11an1n64x5 FILLER_278_8 ();
 b15zdnd11an1n64x5 FILLER_278_72 ();
 b15zdnd11an1n64x5 FILLER_278_136 ();
 b15zdnd11an1n64x5 FILLER_278_200 ();
 b15zdnd11an1n32x5 FILLER_278_264 ();
 b15zdnd11an1n08x5 FILLER_278_296 ();
 b15zdnd00an1n01x5 FILLER_278_304 ();
 b15zdnd11an1n16x5 FILLER_278_347 ();
 b15zdnd11an1n08x5 FILLER_278_363 ();
 b15zdnd11an1n04x5 FILLER_278_374 ();
 b15zdnd11an1n08x5 FILLER_278_420 ();
 b15zdnd00an1n01x5 FILLER_278_428 ();
 b15zdnd11an1n64x5 FILLER_278_436 ();
 b15zdnd11an1n64x5 FILLER_278_500 ();
 b15zdnd00an1n02x5 FILLER_278_564 ();
 b15zdnd00an1n01x5 FILLER_278_566 ();
 b15zdnd11an1n08x5 FILLER_278_574 ();
 b15zdnd11an1n04x5 FILLER_278_582 ();
 b15zdnd00an1n02x5 FILLER_278_586 ();
 b15zdnd11an1n08x5 FILLER_278_594 ();
 b15zdnd00an1n01x5 FILLER_278_602 ();
 b15zdnd11an1n04x5 FILLER_278_609 ();
 b15zdnd11an1n64x5 FILLER_278_623 ();
 b15zdnd11an1n16x5 FILLER_278_687 ();
 b15zdnd11an1n08x5 FILLER_278_703 ();
 b15zdnd11an1n04x5 FILLER_278_711 ();
 b15zdnd00an1n02x5 FILLER_278_715 ();
 b15zdnd00an1n01x5 FILLER_278_717 ();
 b15zdnd11an1n64x5 FILLER_278_726 ();
 b15zdnd11an1n64x5 FILLER_278_790 ();
 b15zdnd11an1n64x5 FILLER_278_854 ();
 b15zdnd00an1n02x5 FILLER_278_918 ();
 b15zdnd11an1n64x5 FILLER_278_946 ();
 b15zdnd11an1n32x5 FILLER_278_1010 ();
 b15zdnd11an1n16x5 FILLER_278_1042 ();
 b15zdnd00an1n02x5 FILLER_278_1058 ();
 b15zdnd00an1n01x5 FILLER_278_1060 ();
 b15zdnd11an1n64x5 FILLER_278_1069 ();
 b15zdnd11an1n16x5 FILLER_278_1165 ();
 b15zdnd11an1n04x5 FILLER_278_1181 ();
 b15zdnd00an1n02x5 FILLER_278_1185 ();
 b15zdnd11an1n08x5 FILLER_278_1204 ();
 b15zdnd11an1n04x5 FILLER_278_1212 ();
 b15zdnd00an1n02x5 FILLER_278_1216 ();
 b15zdnd00an1n01x5 FILLER_278_1218 ();
 b15zdnd11an1n64x5 FILLER_278_1239 ();
 b15zdnd11an1n32x5 FILLER_278_1303 ();
 b15zdnd11an1n04x5 FILLER_278_1375 ();
 b15zdnd11an1n64x5 FILLER_278_1382 ();
 b15zdnd11an1n64x5 FILLER_278_1446 ();
 b15zdnd11an1n08x5 FILLER_278_1510 ();
 b15zdnd11an1n04x5 FILLER_278_1518 ();
 b15zdnd11an1n16x5 FILLER_278_1564 ();
 b15zdnd11an1n08x5 FILLER_278_1580 ();
 b15zdnd11an1n04x5 FILLER_278_1588 ();
 b15zdnd00an1n02x5 FILLER_278_1592 ();
 b15zdnd00an1n01x5 FILLER_278_1594 ();
 b15zdnd11an1n64x5 FILLER_278_1598 ();
 b15zdnd11an1n64x5 FILLER_278_1662 ();
 b15zdnd11an1n16x5 FILLER_278_1726 ();
 b15zdnd11an1n04x5 FILLER_278_1742 ();
 b15zdnd00an1n01x5 FILLER_278_1746 ();
 b15zdnd11an1n64x5 FILLER_278_1750 ();
 b15zdnd11an1n64x5 FILLER_278_1814 ();
 b15zdnd11an1n64x5 FILLER_278_1878 ();
 b15zdnd11an1n64x5 FILLER_278_1942 ();
 b15zdnd11an1n64x5 FILLER_278_2006 ();
 b15zdnd11an1n32x5 FILLER_278_2070 ();
 b15zdnd11an1n08x5 FILLER_278_2102 ();
 b15zdnd11an1n04x5 FILLER_278_2110 ();
 b15zdnd11an1n04x5 FILLER_278_2118 ();
 b15zdnd11an1n04x5 FILLER_278_2129 ();
 b15zdnd11an1n08x5 FILLER_278_2145 ();
 b15zdnd00an1n01x5 FILLER_278_2153 ();
 b15zdnd11an1n64x5 FILLER_278_2162 ();
 b15zdnd11an1n16x5 FILLER_278_2226 ();
 b15zdnd11an1n08x5 FILLER_278_2242 ();
 b15zdnd00an1n02x5 FILLER_278_2250 ();
 b15zdnd11an1n16x5 FILLER_278_2258 ();
 b15zdnd00an1n02x5 FILLER_278_2274 ();
 b15zdnd11an1n64x5 FILLER_279_0 ();
 b15zdnd00an1n01x5 FILLER_279_64 ();
 b15zdnd11an1n64x5 FILLER_279_110 ();
 b15zdnd11an1n64x5 FILLER_279_174 ();
 b15zdnd11an1n64x5 FILLER_279_238 ();
 b15zdnd11an1n32x5 FILLER_279_302 ();
 b15zdnd11an1n08x5 FILLER_279_334 ();
 b15zdnd00an1n02x5 FILLER_279_342 ();
 b15zdnd00an1n01x5 FILLER_279_344 ();
 b15zdnd11an1n04x5 FILLER_279_397 ();
 b15zdnd00an1n01x5 FILLER_279_401 ();
 b15zdnd11an1n04x5 FILLER_279_407 ();
 b15zdnd11an1n64x5 FILLER_279_453 ();
 b15zdnd11an1n32x5 FILLER_279_517 ();
 b15zdnd11an1n04x5 FILLER_279_549 ();
 b15zdnd00an1n02x5 FILLER_279_553 ();
 b15zdnd00an1n01x5 FILLER_279_555 ();
 b15zdnd11an1n04x5 FILLER_279_561 ();
 b15zdnd11an1n16x5 FILLER_279_607 ();
 b15zdnd11an1n08x5 FILLER_279_623 ();
 b15zdnd11an1n64x5 FILLER_279_638 ();
 b15zdnd11an1n64x5 FILLER_279_702 ();
 b15zdnd11an1n64x5 FILLER_279_766 ();
 b15zdnd11an1n64x5 FILLER_279_830 ();
 b15zdnd11an1n08x5 FILLER_279_894 ();
 b15zdnd00an1n02x5 FILLER_279_902 ();
 b15zdnd00an1n01x5 FILLER_279_904 ();
 b15zdnd11an1n16x5 FILLER_279_925 ();
 b15zdnd11an1n08x5 FILLER_279_941 ();
 b15zdnd00an1n01x5 FILLER_279_949 ();
 b15zdnd11an1n04x5 FILLER_279_976 ();
 b15zdnd11an1n64x5 FILLER_279_1000 ();
 b15zdnd11an1n64x5 FILLER_279_1064 ();
 b15zdnd11an1n16x5 FILLER_279_1128 ();
 b15zdnd00an1n02x5 FILLER_279_1144 ();
 b15zdnd11an1n08x5 FILLER_279_1188 ();
 b15zdnd11an1n04x5 FILLER_279_1196 ();
 b15zdnd00an1n02x5 FILLER_279_1200 ();
 b15zdnd11an1n64x5 FILLER_279_1216 ();
 b15zdnd11an1n64x5 FILLER_279_1280 ();
 b15zdnd11an1n64x5 FILLER_279_1344 ();
 b15zdnd11an1n16x5 FILLER_279_1408 ();
 b15zdnd00an1n02x5 FILLER_279_1424 ();
 b15zdnd00an1n01x5 FILLER_279_1426 ();
 b15zdnd11an1n64x5 FILLER_279_1431 ();
 b15zdnd11an1n64x5 FILLER_279_1495 ();
 b15zdnd11an1n64x5 FILLER_279_1559 ();
 b15zdnd11an1n64x5 FILLER_279_1623 ();
 b15zdnd11an1n32x5 FILLER_279_1687 ();
 b15zdnd11an1n04x5 FILLER_279_1719 ();
 b15zdnd00an1n02x5 FILLER_279_1723 ();
 b15zdnd11an1n64x5 FILLER_279_1777 ();
 b15zdnd11an1n64x5 FILLER_279_1841 ();
 b15zdnd11an1n64x5 FILLER_279_1905 ();
 b15zdnd11an1n64x5 FILLER_279_1969 ();
 b15zdnd11an1n64x5 FILLER_279_2033 ();
 b15zdnd11an1n16x5 FILLER_279_2097 ();
 b15zdnd00an1n01x5 FILLER_279_2113 ();
 b15zdnd11an1n04x5 FILLER_279_2120 ();
 b15zdnd11an1n04x5 FILLER_279_2129 ();
 b15zdnd11an1n64x5 FILLER_279_2175 ();
 b15zdnd11an1n32x5 FILLER_279_2239 ();
 b15zdnd11an1n08x5 FILLER_279_2271 ();
 b15zdnd11an1n04x5 FILLER_279_2279 ();
 b15zdnd00an1n01x5 FILLER_279_2283 ();
 b15zdnd11an1n64x5 FILLER_280_8 ();
 b15zdnd11an1n64x5 FILLER_280_72 ();
 b15zdnd11an1n64x5 FILLER_280_136 ();
 b15zdnd11an1n64x5 FILLER_280_200 ();
 b15zdnd11an1n64x5 FILLER_280_264 ();
 b15zdnd11an1n32x5 FILLER_280_328 ();
 b15zdnd00an1n02x5 FILLER_280_360 ();
 b15zdnd00an1n01x5 FILLER_280_362 ();
 b15zdnd11an1n04x5 FILLER_280_366 ();
 b15zdnd11an1n16x5 FILLER_280_373 ();
 b15zdnd11an1n08x5 FILLER_280_389 ();
 b15zdnd11an1n64x5 FILLER_280_439 ();
 b15zdnd11an1n64x5 FILLER_280_503 ();
 b15zdnd11an1n04x5 FILLER_280_571 ();
 b15zdnd11an1n64x5 FILLER_280_617 ();
 b15zdnd11an1n32x5 FILLER_280_681 ();
 b15zdnd11an1n04x5 FILLER_280_713 ();
 b15zdnd00an1n01x5 FILLER_280_717 ();
 b15zdnd11an1n32x5 FILLER_280_726 ();
 b15zdnd11an1n08x5 FILLER_280_758 ();
 b15zdnd11an1n04x5 FILLER_280_766 ();
 b15zdnd00an1n02x5 FILLER_280_770 ();
 b15zdnd00an1n01x5 FILLER_280_772 ();
 b15zdnd11an1n64x5 FILLER_280_776 ();
 b15zdnd11an1n64x5 FILLER_280_840 ();
 b15zdnd11an1n64x5 FILLER_280_904 ();
 b15zdnd11an1n64x5 FILLER_280_968 ();
 b15zdnd11an1n64x5 FILLER_280_1032 ();
 b15zdnd11an1n32x5 FILLER_280_1096 ();
 b15zdnd11an1n16x5 FILLER_280_1128 ();
 b15zdnd11an1n08x5 FILLER_280_1144 ();
 b15zdnd11an1n04x5 FILLER_280_1152 ();
 b15zdnd00an1n01x5 FILLER_280_1156 ();
 b15zdnd11an1n64x5 FILLER_280_1209 ();
 b15zdnd11an1n64x5 FILLER_280_1273 ();
 b15zdnd11an1n64x5 FILLER_280_1337 ();
 b15zdnd11an1n32x5 FILLER_280_1401 ();
 b15zdnd11an1n16x5 FILLER_280_1433 ();
 b15zdnd11an1n04x5 FILLER_280_1458 ();
 b15zdnd11an1n64x5 FILLER_280_1468 ();
 b15zdnd11an1n64x5 FILLER_280_1532 ();
 b15zdnd11an1n64x5 FILLER_280_1596 ();
 b15zdnd11an1n64x5 FILLER_280_1660 ();
 b15zdnd11an1n16x5 FILLER_280_1724 ();
 b15zdnd00an1n01x5 FILLER_280_1740 ();
 b15zdnd11an1n64x5 FILLER_280_1783 ();
 b15zdnd11an1n32x5 FILLER_280_1847 ();
 b15zdnd11an1n16x5 FILLER_280_1879 ();
 b15zdnd11an1n08x5 FILLER_280_1895 ();
 b15zdnd11an1n04x5 FILLER_280_1903 ();
 b15zdnd00an1n01x5 FILLER_280_1907 ();
 b15zdnd11an1n64x5 FILLER_280_1916 ();
 b15zdnd11an1n64x5 FILLER_280_1980 ();
 b15zdnd11an1n64x5 FILLER_280_2044 ();
 b15zdnd11an1n08x5 FILLER_280_2108 ();
 b15zdnd11an1n04x5 FILLER_280_2116 ();
 b15zdnd00an1n02x5 FILLER_280_2120 ();
 b15zdnd00an1n01x5 FILLER_280_2122 ();
 b15zdnd11an1n16x5 FILLER_280_2134 ();
 b15zdnd11an1n04x5 FILLER_280_2150 ();
 b15zdnd11an1n64x5 FILLER_280_2162 ();
 b15zdnd11an1n32x5 FILLER_280_2226 ();
 b15zdnd11an1n16x5 FILLER_280_2258 ();
 b15zdnd00an1n02x5 FILLER_280_2274 ();
 b15zdnd11an1n64x5 FILLER_281_0 ();
 b15zdnd11an1n64x5 FILLER_281_64 ();
 b15zdnd11an1n64x5 FILLER_281_128 ();
 b15zdnd11an1n64x5 FILLER_281_192 ();
 b15zdnd11an1n64x5 FILLER_281_256 ();
 b15zdnd11an1n64x5 FILLER_281_320 ();
 b15zdnd00an1n02x5 FILLER_281_384 ();
 b15zdnd00an1n01x5 FILLER_281_386 ();
 b15zdnd11an1n16x5 FILLER_281_405 ();
 b15zdnd00an1n02x5 FILLER_281_421 ();
 b15zdnd00an1n01x5 FILLER_281_423 ();
 b15zdnd11an1n64x5 FILLER_281_428 ();
 b15zdnd11an1n32x5 FILLER_281_492 ();
 b15zdnd11an1n08x5 FILLER_281_524 ();
 b15zdnd11an1n04x5 FILLER_281_532 ();
 b15zdnd00an1n02x5 FILLER_281_536 ();
 b15zdnd11an1n04x5 FILLER_281_590 ();
 b15zdnd11an1n64x5 FILLER_281_599 ();
 b15zdnd11an1n64x5 FILLER_281_663 ();
 b15zdnd00an1n02x5 FILLER_281_727 ();
 b15zdnd11an1n32x5 FILLER_281_733 ();
 b15zdnd00an1n02x5 FILLER_281_765 ();
 b15zdnd11an1n04x5 FILLER_281_770 ();
 b15zdnd11an1n04x5 FILLER_281_777 ();
 b15zdnd11an1n64x5 FILLER_281_784 ();
 b15zdnd11an1n64x5 FILLER_281_848 ();
 b15zdnd11an1n32x5 FILLER_281_912 ();
 b15zdnd11an1n16x5 FILLER_281_944 ();
 b15zdnd11an1n04x5 FILLER_281_960 ();
 b15zdnd11an1n32x5 FILLER_281_976 ();
 b15zdnd11an1n04x5 FILLER_281_1008 ();
 b15zdnd00an1n01x5 FILLER_281_1012 ();
 b15zdnd11an1n04x5 FILLER_281_1036 ();
 b15zdnd11an1n64x5 FILLER_281_1052 ();
 b15zdnd11an1n16x5 FILLER_281_1116 ();
 b15zdnd11an1n08x5 FILLER_281_1132 ();
 b15zdnd00an1n01x5 FILLER_281_1140 ();
 b15zdnd11an1n16x5 FILLER_281_1149 ();
 b15zdnd11an1n08x5 FILLER_281_1165 ();
 b15zdnd11an1n04x5 FILLER_281_1173 ();
 b15zdnd00an1n02x5 FILLER_281_1177 ();
 b15zdnd00an1n01x5 FILLER_281_1179 ();
 b15zdnd11an1n04x5 FILLER_281_1183 ();
 b15zdnd11an1n64x5 FILLER_281_1190 ();
 b15zdnd11an1n64x5 FILLER_281_1254 ();
 b15zdnd11an1n64x5 FILLER_281_1318 ();
 b15zdnd11an1n64x5 FILLER_281_1382 ();
 b15zdnd11an1n08x5 FILLER_281_1446 ();
 b15zdnd11an1n04x5 FILLER_281_1458 ();
 b15zdnd00an1n02x5 FILLER_281_1462 ();
 b15zdnd11an1n64x5 FILLER_281_1475 ();
 b15zdnd11an1n64x5 FILLER_281_1539 ();
 b15zdnd11an1n64x5 FILLER_281_1603 ();
 b15zdnd11an1n64x5 FILLER_281_1667 ();
 b15zdnd11an1n16x5 FILLER_281_1731 ();
 b15zdnd00an1n02x5 FILLER_281_1747 ();
 b15zdnd00an1n01x5 FILLER_281_1749 ();
 b15zdnd11an1n04x5 FILLER_281_1753 ();
 b15zdnd11an1n64x5 FILLER_281_1760 ();
 b15zdnd11an1n64x5 FILLER_281_1824 ();
 b15zdnd11an1n64x5 FILLER_281_1888 ();
 b15zdnd11an1n32x5 FILLER_281_1952 ();
 b15zdnd11an1n16x5 FILLER_281_1984 ();
 b15zdnd00an1n01x5 FILLER_281_2000 ();
 b15zdnd11an1n64x5 FILLER_281_2040 ();
 b15zdnd11an1n08x5 FILLER_281_2104 ();
 b15zdnd11an1n04x5 FILLER_281_2112 ();
 b15zdnd00an1n01x5 FILLER_281_2116 ();
 b15zdnd11an1n64x5 FILLER_281_2130 ();
 b15zdnd11an1n64x5 FILLER_281_2194 ();
 b15zdnd11an1n16x5 FILLER_281_2258 ();
 b15zdnd11an1n08x5 FILLER_281_2274 ();
 b15zdnd00an1n02x5 FILLER_281_2282 ();
 b15zdnd11an1n64x5 FILLER_282_8 ();
 b15zdnd11an1n64x5 FILLER_282_72 ();
 b15zdnd11an1n64x5 FILLER_282_136 ();
 b15zdnd11an1n64x5 FILLER_282_200 ();
 b15zdnd11an1n64x5 FILLER_282_264 ();
 b15zdnd11an1n64x5 FILLER_282_328 ();
 b15zdnd11an1n16x5 FILLER_282_392 ();
 b15zdnd00an1n02x5 FILLER_282_408 ();
 b15zdnd00an1n01x5 FILLER_282_410 ();
 b15zdnd11an1n64x5 FILLER_282_415 ();
 b15zdnd11an1n64x5 FILLER_282_479 ();
 b15zdnd11an1n04x5 FILLER_282_543 ();
 b15zdnd00an1n01x5 FILLER_282_547 ();
 b15zdnd11an1n04x5 FILLER_282_551 ();
 b15zdnd11an1n64x5 FILLER_282_597 ();
 b15zdnd11an1n32x5 FILLER_282_661 ();
 b15zdnd11an1n16x5 FILLER_282_693 ();
 b15zdnd11an1n08x5 FILLER_282_709 ();
 b15zdnd00an1n01x5 FILLER_282_717 ();
 b15zdnd11an1n16x5 FILLER_282_726 ();
 b15zdnd11an1n04x5 FILLER_282_742 ();
 b15zdnd00an1n01x5 FILLER_282_746 ();
 b15zdnd11an1n32x5 FILLER_282_799 ();
 b15zdnd11an1n16x5 FILLER_282_831 ();
 b15zdnd11an1n04x5 FILLER_282_847 ();
 b15zdnd00an1n02x5 FILLER_282_851 ();
 b15zdnd11an1n64x5 FILLER_282_856 ();
 b15zdnd11an1n08x5 FILLER_282_920 ();
 b15zdnd11an1n04x5 FILLER_282_928 ();
 b15zdnd00an1n02x5 FILLER_282_932 ();
 b15zdnd11an1n64x5 FILLER_282_939 ();
 b15zdnd11an1n64x5 FILLER_282_1003 ();
 b15zdnd11an1n64x5 FILLER_282_1067 ();
 b15zdnd11an1n16x5 FILLER_282_1131 ();
 b15zdnd11an1n08x5 FILLER_282_1147 ();
 b15zdnd11an1n04x5 FILLER_282_1155 ();
 b15zdnd00an1n02x5 FILLER_282_1159 ();
 b15zdnd00an1n01x5 FILLER_282_1161 ();
 b15zdnd11an1n04x5 FILLER_282_1168 ();
 b15zdnd00an1n02x5 FILLER_282_1172 ();
 b15zdnd00an1n01x5 FILLER_282_1174 ();
 b15zdnd11an1n64x5 FILLER_282_1217 ();
 b15zdnd11an1n64x5 FILLER_282_1281 ();
 b15zdnd11an1n64x5 FILLER_282_1345 ();
 b15zdnd11an1n64x5 FILLER_282_1409 ();
 b15zdnd11an1n64x5 FILLER_282_1473 ();
 b15zdnd11an1n64x5 FILLER_282_1537 ();
 b15zdnd11an1n64x5 FILLER_282_1601 ();
 b15zdnd11an1n64x5 FILLER_282_1665 ();
 b15zdnd11an1n64x5 FILLER_282_1729 ();
 b15zdnd11an1n64x5 FILLER_282_1793 ();
 b15zdnd11an1n64x5 FILLER_282_1857 ();
 b15zdnd11an1n04x5 FILLER_282_1921 ();
 b15zdnd00an1n01x5 FILLER_282_1925 ();
 b15zdnd11an1n32x5 FILLER_282_1968 ();
 b15zdnd11an1n04x5 FILLER_282_2000 ();
 b15zdnd11an1n64x5 FILLER_282_2015 ();
 b15zdnd11an1n64x5 FILLER_282_2079 ();
 b15zdnd11an1n08x5 FILLER_282_2143 ();
 b15zdnd00an1n02x5 FILLER_282_2151 ();
 b15zdnd00an1n01x5 FILLER_282_2153 ();
 b15zdnd11an1n64x5 FILLER_282_2162 ();
 b15zdnd11an1n32x5 FILLER_282_2226 ();
 b15zdnd11an1n16x5 FILLER_282_2258 ();
 b15zdnd00an1n02x5 FILLER_282_2274 ();
 b15zdnd11an1n64x5 FILLER_283_0 ();
 b15zdnd11an1n64x5 FILLER_283_64 ();
 b15zdnd11an1n64x5 FILLER_283_128 ();
 b15zdnd11an1n64x5 FILLER_283_192 ();
 b15zdnd11an1n64x5 FILLER_283_256 ();
 b15zdnd11an1n64x5 FILLER_283_320 ();
 b15zdnd11an1n16x5 FILLER_283_384 ();
 b15zdnd00an1n01x5 FILLER_283_400 ();
 b15zdnd11an1n04x5 FILLER_283_407 ();
 b15zdnd00an1n01x5 FILLER_283_411 ();
 b15zdnd11an1n64x5 FILLER_283_424 ();
 b15zdnd11an1n32x5 FILLER_283_488 ();
 b15zdnd11an1n08x5 FILLER_283_520 ();
 b15zdnd11an1n04x5 FILLER_283_528 ();
 b15zdnd00an1n02x5 FILLER_283_532 ();
 b15zdnd11an1n64x5 FILLER_283_576 ();
 b15zdnd11an1n64x5 FILLER_283_640 ();
 b15zdnd11an1n32x5 FILLER_283_704 ();
 b15zdnd11an1n08x5 FILLER_283_736 ();
 b15zdnd11an1n04x5 FILLER_283_744 ();
 b15zdnd11an1n04x5 FILLER_283_754 ();
 b15zdnd00an1n01x5 FILLER_283_758 ();
 b15zdnd11an1n04x5 FILLER_283_764 ();
 b15zdnd11an1n04x5 FILLER_283_810 ();
 b15zdnd11an1n04x5 FILLER_283_854 ();
 b15zdnd00an1n02x5 FILLER_283_858 ();
 b15zdnd11an1n64x5 FILLER_283_863 ();
 b15zdnd11an1n64x5 FILLER_283_927 ();
 b15zdnd11an1n64x5 FILLER_283_991 ();
 b15zdnd11an1n64x5 FILLER_283_1055 ();
 b15zdnd11an1n16x5 FILLER_283_1119 ();
 b15zdnd11an1n04x5 FILLER_283_1135 ();
 b15zdnd00an1n02x5 FILLER_283_1139 ();
 b15zdnd00an1n01x5 FILLER_283_1141 ();
 b15zdnd11an1n08x5 FILLER_283_1167 ();
 b15zdnd11an1n04x5 FILLER_283_1175 ();
 b15zdnd00an1n01x5 FILLER_283_1179 ();
 b15zdnd11an1n64x5 FILLER_283_1183 ();
 b15zdnd11an1n64x5 FILLER_283_1247 ();
 b15zdnd11an1n64x5 FILLER_283_1311 ();
 b15zdnd11an1n64x5 FILLER_283_1375 ();
 b15zdnd11an1n08x5 FILLER_283_1439 ();
 b15zdnd11an1n04x5 FILLER_283_1447 ();
 b15zdnd11an1n64x5 FILLER_283_1456 ();
 b15zdnd11an1n32x5 FILLER_283_1520 ();
 b15zdnd11an1n16x5 FILLER_283_1552 ();
 b15zdnd00an1n02x5 FILLER_283_1568 ();
 b15zdnd00an1n01x5 FILLER_283_1570 ();
 b15zdnd11an1n64x5 FILLER_283_1580 ();
 b15zdnd11an1n64x5 FILLER_283_1644 ();
 b15zdnd11an1n32x5 FILLER_283_1708 ();
 b15zdnd11an1n16x5 FILLER_283_1740 ();
 b15zdnd11an1n04x5 FILLER_283_1756 ();
 b15zdnd00an1n02x5 FILLER_283_1760 ();
 b15zdnd11an1n64x5 FILLER_283_1804 ();
 b15zdnd11an1n64x5 FILLER_283_1868 ();
 b15zdnd11an1n04x5 FILLER_283_1932 ();
 b15zdnd00an1n01x5 FILLER_283_1936 ();
 b15zdnd11an1n64x5 FILLER_283_1979 ();
 b15zdnd11an1n64x5 FILLER_283_2043 ();
 b15zdnd11an1n04x5 FILLER_283_2107 ();
 b15zdnd11an1n64x5 FILLER_283_2153 ();
 b15zdnd11an1n64x5 FILLER_283_2217 ();
 b15zdnd00an1n02x5 FILLER_283_2281 ();
 b15zdnd00an1n01x5 FILLER_283_2283 ();
 b15zdnd11an1n64x5 FILLER_284_8 ();
 b15zdnd11an1n64x5 FILLER_284_72 ();
 b15zdnd11an1n64x5 FILLER_284_136 ();
 b15zdnd11an1n64x5 FILLER_284_200 ();
 b15zdnd11an1n64x5 FILLER_284_264 ();
 b15zdnd11an1n64x5 FILLER_284_328 ();
 b15zdnd00an1n02x5 FILLER_284_392 ();
 b15zdnd11an1n04x5 FILLER_284_400 ();
 b15zdnd11an1n64x5 FILLER_284_446 ();
 b15zdnd11an1n32x5 FILLER_284_510 ();
 b15zdnd11an1n16x5 FILLER_284_542 ();
 b15zdnd00an1n02x5 FILLER_284_558 ();
 b15zdnd00an1n01x5 FILLER_284_560 ();
 b15zdnd11an1n04x5 FILLER_284_564 ();
 b15zdnd11an1n64x5 FILLER_284_571 ();
 b15zdnd11an1n64x5 FILLER_284_635 ();
 b15zdnd11an1n16x5 FILLER_284_699 ();
 b15zdnd00an1n02x5 FILLER_284_715 ();
 b15zdnd00an1n01x5 FILLER_284_717 ();
 b15zdnd11an1n16x5 FILLER_284_726 ();
 b15zdnd00an1n02x5 FILLER_284_742 ();
 b15zdnd11an1n64x5 FILLER_284_786 ();
 b15zdnd11an1n64x5 FILLER_284_850 ();
 b15zdnd11an1n64x5 FILLER_284_914 ();
 b15zdnd11an1n16x5 FILLER_284_978 ();
 b15zdnd11an1n04x5 FILLER_284_994 ();
 b15zdnd00an1n01x5 FILLER_284_998 ();
 b15zdnd11an1n64x5 FILLER_284_1022 ();
 b15zdnd11an1n64x5 FILLER_284_1086 ();
 b15zdnd11an1n64x5 FILLER_284_1150 ();
 b15zdnd11an1n64x5 FILLER_284_1214 ();
 b15zdnd11an1n64x5 FILLER_284_1278 ();
 b15zdnd11an1n64x5 FILLER_284_1342 ();
 b15zdnd11an1n16x5 FILLER_284_1406 ();
 b15zdnd11an1n08x5 FILLER_284_1422 ();
 b15zdnd11an1n04x5 FILLER_284_1450 ();
 b15zdnd11an1n64x5 FILLER_284_1464 ();
 b15zdnd11an1n64x5 FILLER_284_1528 ();
 b15zdnd11an1n32x5 FILLER_284_1592 ();
 b15zdnd11an1n16x5 FILLER_284_1624 ();
 b15zdnd11an1n04x5 FILLER_284_1640 ();
 b15zdnd00an1n02x5 FILLER_284_1644 ();
 b15zdnd00an1n01x5 FILLER_284_1646 ();
 b15zdnd11an1n04x5 FILLER_284_1650 ();
 b15zdnd11an1n64x5 FILLER_284_1657 ();
 b15zdnd11an1n64x5 FILLER_284_1721 ();
 b15zdnd11an1n64x5 FILLER_284_1785 ();
 b15zdnd11an1n64x5 FILLER_284_1849 ();
 b15zdnd11an1n16x5 FILLER_284_1913 ();
 b15zdnd00an1n02x5 FILLER_284_1929 ();
 b15zdnd11an1n64x5 FILLER_284_1940 ();
 b15zdnd11an1n64x5 FILLER_284_2004 ();
 b15zdnd11an1n16x5 FILLER_284_2068 ();
 b15zdnd11an1n04x5 FILLER_284_2084 ();
 b15zdnd00an1n01x5 FILLER_284_2088 ();
 b15zdnd11an1n16x5 FILLER_284_2131 ();
 b15zdnd11an1n04x5 FILLER_284_2147 ();
 b15zdnd00an1n02x5 FILLER_284_2151 ();
 b15zdnd00an1n01x5 FILLER_284_2153 ();
 b15zdnd11an1n64x5 FILLER_284_2162 ();
 b15zdnd11an1n32x5 FILLER_284_2226 ();
 b15zdnd11an1n16x5 FILLER_284_2258 ();
 b15zdnd00an1n02x5 FILLER_284_2274 ();
 b15zdnd11an1n64x5 FILLER_285_0 ();
 b15zdnd11an1n64x5 FILLER_285_64 ();
 b15zdnd11an1n64x5 FILLER_285_128 ();
 b15zdnd11an1n64x5 FILLER_285_192 ();
 b15zdnd11an1n64x5 FILLER_285_256 ();
 b15zdnd11an1n64x5 FILLER_285_320 ();
 b15zdnd11an1n16x5 FILLER_285_384 ();
 b15zdnd11an1n04x5 FILLER_285_400 ();
 b15zdnd00an1n02x5 FILLER_285_404 ();
 b15zdnd00an1n01x5 FILLER_285_406 ();
 b15zdnd11an1n04x5 FILLER_285_420 ();
 b15zdnd11an1n64x5 FILLER_285_431 ();
 b15zdnd11an1n64x5 FILLER_285_495 ();
 b15zdnd11an1n64x5 FILLER_285_559 ();
 b15zdnd11an1n64x5 FILLER_285_623 ();
 b15zdnd11an1n32x5 FILLER_285_687 ();
 b15zdnd11an1n08x5 FILLER_285_719 ();
 b15zdnd11an1n04x5 FILLER_285_727 ();
 b15zdnd00an1n02x5 FILLER_285_731 ();
 b15zdnd00an1n01x5 FILLER_285_733 ();
 b15zdnd11an1n08x5 FILLER_285_740 ();
 b15zdnd11an1n04x5 FILLER_285_748 ();
 b15zdnd00an1n02x5 FILLER_285_752 ();
 b15zdnd11an1n64x5 FILLER_285_796 ();
 b15zdnd11an1n64x5 FILLER_285_860 ();
 b15zdnd11an1n64x5 FILLER_285_924 ();
 b15zdnd11an1n64x5 FILLER_285_988 ();
 b15zdnd00an1n02x5 FILLER_285_1052 ();
 b15zdnd00an1n01x5 FILLER_285_1054 ();
 b15zdnd11an1n08x5 FILLER_285_1059 ();
 b15zdnd11an1n04x5 FILLER_285_1067 ();
 b15zdnd00an1n02x5 FILLER_285_1071 ();
 b15zdnd00an1n01x5 FILLER_285_1073 ();
 b15zdnd11an1n16x5 FILLER_285_1105 ();
 b15zdnd11an1n08x5 FILLER_285_1121 ();
 b15zdnd11an1n04x5 FILLER_285_1129 ();
 b15zdnd00an1n02x5 FILLER_285_1133 ();
 b15zdnd11an1n64x5 FILLER_285_1156 ();
 b15zdnd11an1n64x5 FILLER_285_1220 ();
 b15zdnd11an1n64x5 FILLER_285_1284 ();
 b15zdnd11an1n64x5 FILLER_285_1348 ();
 b15zdnd11an1n08x5 FILLER_285_1412 ();
 b15zdnd11an1n04x5 FILLER_285_1420 ();
 b15zdnd00an1n02x5 FILLER_285_1424 ();
 b15zdnd11an1n64x5 FILLER_285_1438 ();
 b15zdnd11an1n64x5 FILLER_285_1502 ();
 b15zdnd11an1n32x5 FILLER_285_1566 ();
 b15zdnd11an1n16x5 FILLER_285_1598 ();
 b15zdnd00an1n01x5 FILLER_285_1614 ();
 b15zdnd11an1n64x5 FILLER_285_1655 ();
 b15zdnd11an1n64x5 FILLER_285_1719 ();
 b15zdnd11an1n64x5 FILLER_285_1783 ();
 b15zdnd11an1n64x5 FILLER_285_1847 ();
 b15zdnd11an1n64x5 FILLER_285_1911 ();
 b15zdnd11an1n64x5 FILLER_285_1975 ();
 b15zdnd11an1n04x5 FILLER_285_2039 ();
 b15zdnd00an1n02x5 FILLER_285_2043 ();
 b15zdnd11an1n08x5 FILLER_285_2048 ();
 b15zdnd00an1n02x5 FILLER_285_2056 ();
 b15zdnd00an1n01x5 FILLER_285_2058 ();
 b15zdnd11an1n16x5 FILLER_285_2062 ();
 b15zdnd11an1n04x5 FILLER_285_2078 ();
 b15zdnd00an1n01x5 FILLER_285_2082 ();
 b15zdnd11an1n64x5 FILLER_285_2089 ();
 b15zdnd11an1n64x5 FILLER_285_2153 ();
 b15zdnd11an1n64x5 FILLER_285_2217 ();
 b15zdnd00an1n02x5 FILLER_285_2281 ();
 b15zdnd00an1n01x5 FILLER_285_2283 ();
 b15zdnd11an1n64x5 FILLER_286_8 ();
 b15zdnd11an1n64x5 FILLER_286_72 ();
 b15zdnd11an1n64x5 FILLER_286_136 ();
 b15zdnd11an1n64x5 FILLER_286_200 ();
 b15zdnd11an1n64x5 FILLER_286_264 ();
 b15zdnd11an1n64x5 FILLER_286_328 ();
 b15zdnd11an1n16x5 FILLER_286_392 ();
 b15zdnd11an1n04x5 FILLER_286_408 ();
 b15zdnd11an1n64x5 FILLER_286_422 ();
 b15zdnd11an1n64x5 FILLER_286_486 ();
 b15zdnd11an1n64x5 FILLER_286_550 ();
 b15zdnd11an1n64x5 FILLER_286_614 ();
 b15zdnd11an1n32x5 FILLER_286_678 ();
 b15zdnd11an1n08x5 FILLER_286_710 ();
 b15zdnd11an1n04x5 FILLER_286_726 ();
 b15zdnd11an1n64x5 FILLER_286_743 ();
 b15zdnd11an1n64x5 FILLER_286_807 ();
 b15zdnd11an1n64x5 FILLER_286_871 ();
 b15zdnd11an1n64x5 FILLER_286_935 ();
 b15zdnd11an1n64x5 FILLER_286_999 ();
 b15zdnd11an1n64x5 FILLER_286_1063 ();
 b15zdnd11an1n64x5 FILLER_286_1127 ();
 b15zdnd11an1n64x5 FILLER_286_1191 ();
 b15zdnd11an1n64x5 FILLER_286_1255 ();
 b15zdnd11an1n64x5 FILLER_286_1319 ();
 b15zdnd11an1n64x5 FILLER_286_1383 ();
 b15zdnd11an1n08x5 FILLER_286_1447 ();
 b15zdnd00an1n02x5 FILLER_286_1455 ();
 b15zdnd00an1n01x5 FILLER_286_1457 ();
 b15zdnd11an1n64x5 FILLER_286_1466 ();
 b15zdnd11an1n64x5 FILLER_286_1530 ();
 b15zdnd11an1n64x5 FILLER_286_1594 ();
 b15zdnd11an1n64x5 FILLER_286_1658 ();
 b15zdnd11an1n64x5 FILLER_286_1722 ();
 b15zdnd11an1n16x5 FILLER_286_1786 ();
 b15zdnd11an1n64x5 FILLER_286_1805 ();
 b15zdnd11an1n64x5 FILLER_286_1869 ();
 b15zdnd11an1n64x5 FILLER_286_1933 ();
 b15zdnd11an1n32x5 FILLER_286_1997 ();
 b15zdnd00an1n02x5 FILLER_286_2029 ();
 b15zdnd11an1n64x5 FILLER_286_2083 ();
 b15zdnd11an1n04x5 FILLER_286_2147 ();
 b15zdnd00an1n02x5 FILLER_286_2151 ();
 b15zdnd00an1n01x5 FILLER_286_2153 ();
 b15zdnd11an1n64x5 FILLER_286_2162 ();
 b15zdnd11an1n32x5 FILLER_286_2226 ();
 b15zdnd11an1n16x5 FILLER_286_2258 ();
 b15zdnd00an1n02x5 FILLER_286_2274 ();
 b15zdnd11an1n64x5 FILLER_287_0 ();
 b15zdnd11an1n64x5 FILLER_287_64 ();
 b15zdnd11an1n64x5 FILLER_287_128 ();
 b15zdnd11an1n64x5 FILLER_287_192 ();
 b15zdnd11an1n64x5 FILLER_287_256 ();
 b15zdnd11an1n64x5 FILLER_287_320 ();
 b15zdnd11an1n16x5 FILLER_287_384 ();
 b15zdnd11an1n08x5 FILLER_287_400 ();
 b15zdnd00an1n01x5 FILLER_287_408 ();
 b15zdnd11an1n64x5 FILLER_287_423 ();
 b15zdnd11an1n64x5 FILLER_287_487 ();
 b15zdnd11an1n64x5 FILLER_287_551 ();
 b15zdnd11an1n64x5 FILLER_287_615 ();
 b15zdnd11an1n32x5 FILLER_287_679 ();
 b15zdnd11an1n16x5 FILLER_287_711 ();
 b15zdnd11an1n04x5 FILLER_287_727 ();
 b15zdnd00an1n01x5 FILLER_287_731 ();
 b15zdnd11an1n04x5 FILLER_287_738 ();
 b15zdnd00an1n01x5 FILLER_287_742 ();
 b15zdnd11an1n64x5 FILLER_287_785 ();
 b15zdnd11an1n64x5 FILLER_287_849 ();
 b15zdnd11an1n32x5 FILLER_287_913 ();
 b15zdnd11an1n16x5 FILLER_287_945 ();
 b15zdnd11an1n08x5 FILLER_287_961 ();
 b15zdnd00an1n02x5 FILLER_287_969 ();
 b15zdnd00an1n01x5 FILLER_287_971 ();
 b15zdnd11an1n64x5 FILLER_287_975 ();
 b15zdnd11an1n64x5 FILLER_287_1039 ();
 b15zdnd11an1n32x5 FILLER_287_1103 ();
 b15zdnd11an1n08x5 FILLER_287_1135 ();
 b15zdnd11an1n04x5 FILLER_287_1143 ();
 b15zdnd00an1n01x5 FILLER_287_1147 ();
 b15zdnd11an1n32x5 FILLER_287_1152 ();
 b15zdnd11an1n04x5 FILLER_287_1184 ();
 b15zdnd00an1n02x5 FILLER_287_1188 ();
 b15zdnd00an1n01x5 FILLER_287_1190 ();
 b15zdnd11an1n64x5 FILLER_287_1194 ();
 b15zdnd11an1n64x5 FILLER_287_1258 ();
 b15zdnd11an1n64x5 FILLER_287_1322 ();
 b15zdnd11an1n64x5 FILLER_287_1386 ();
 b15zdnd00an1n02x5 FILLER_287_1450 ();
 b15zdnd00an1n01x5 FILLER_287_1452 ();
 b15zdnd11an1n64x5 FILLER_287_1463 ();
 b15zdnd11an1n64x5 FILLER_287_1527 ();
 b15zdnd11an1n64x5 FILLER_287_1591 ();
 b15zdnd11an1n64x5 FILLER_287_1655 ();
 b15zdnd11an1n08x5 FILLER_287_1719 ();
 b15zdnd11an1n04x5 FILLER_287_1727 ();
 b15zdnd11an1n04x5 FILLER_287_1762 ();
 b15zdnd11an1n64x5 FILLER_287_1806 ();
 b15zdnd11an1n32x5 FILLER_287_1870 ();
 b15zdnd11an1n16x5 FILLER_287_1902 ();
 b15zdnd11an1n04x5 FILLER_287_1921 ();
 b15zdnd11an1n64x5 FILLER_287_1928 ();
 b15zdnd11an1n64x5 FILLER_287_1992 ();
 b15zdnd11an1n64x5 FILLER_287_2059 ();
 b15zdnd11an1n64x5 FILLER_287_2123 ();
 b15zdnd11an1n64x5 FILLER_287_2187 ();
 b15zdnd11an1n32x5 FILLER_287_2251 ();
 b15zdnd00an1n01x5 FILLER_287_2283 ();
 b15zdnd11an1n64x5 FILLER_288_8 ();
 b15zdnd11an1n64x5 FILLER_288_72 ();
 b15zdnd11an1n64x5 FILLER_288_136 ();
 b15zdnd11an1n64x5 FILLER_288_200 ();
 b15zdnd11an1n64x5 FILLER_288_264 ();
 b15zdnd11an1n64x5 FILLER_288_328 ();
 b15zdnd11an1n64x5 FILLER_288_392 ();
 b15zdnd11an1n64x5 FILLER_288_456 ();
 b15zdnd11an1n64x5 FILLER_288_520 ();
 b15zdnd11an1n64x5 FILLER_288_584 ();
 b15zdnd11an1n64x5 FILLER_288_648 ();
 b15zdnd11an1n04x5 FILLER_288_712 ();
 b15zdnd00an1n02x5 FILLER_288_716 ();
 b15zdnd11an1n64x5 FILLER_288_726 ();
 b15zdnd11an1n64x5 FILLER_288_790 ();
 b15zdnd11an1n64x5 FILLER_288_854 ();
 b15zdnd11an1n16x5 FILLER_288_918 ();
 b15zdnd11an1n04x5 FILLER_288_934 ();
 b15zdnd00an1n02x5 FILLER_288_938 ();
 b15zdnd00an1n01x5 FILLER_288_940 ();
 b15zdnd11an1n16x5 FILLER_288_983 ();
 b15zdnd11an1n04x5 FILLER_288_999 ();
 b15zdnd00an1n02x5 FILLER_288_1003 ();
 b15zdnd00an1n01x5 FILLER_288_1005 ();
 b15zdnd11an1n64x5 FILLER_288_1026 ();
 b15zdnd11an1n64x5 FILLER_288_1090 ();
 b15zdnd11an1n32x5 FILLER_288_1154 ();
 b15zdnd00an1n02x5 FILLER_288_1186 ();
 b15zdnd00an1n01x5 FILLER_288_1188 ();
 b15zdnd11an1n04x5 FILLER_288_1192 ();
 b15zdnd11an1n64x5 FILLER_288_1199 ();
 b15zdnd11an1n64x5 FILLER_288_1263 ();
 b15zdnd11an1n64x5 FILLER_288_1327 ();
 b15zdnd11an1n64x5 FILLER_288_1391 ();
 b15zdnd11an1n64x5 FILLER_288_1455 ();
 b15zdnd11an1n64x5 FILLER_288_1519 ();
 b15zdnd11an1n64x5 FILLER_288_1583 ();
 b15zdnd11an1n64x5 FILLER_288_1647 ();
 b15zdnd11an1n64x5 FILLER_288_1711 ();
 b15zdnd11an1n16x5 FILLER_288_1775 ();
 b15zdnd11an1n08x5 FILLER_288_1791 ();
 b15zdnd11an1n04x5 FILLER_288_1799 ();
 b15zdnd00an1n01x5 FILLER_288_1803 ();
 b15zdnd11an1n64x5 FILLER_288_1807 ();
 b15zdnd11an1n16x5 FILLER_288_1871 ();
 b15zdnd11an1n08x5 FILLER_288_1887 ();
 b15zdnd11an1n04x5 FILLER_288_1895 ();
 b15zdnd00an1n01x5 FILLER_288_1899 ();
 b15zdnd11an1n64x5 FILLER_288_1952 ();
 b15zdnd11an1n64x5 FILLER_288_2016 ();
 b15zdnd11an1n64x5 FILLER_288_2080 ();
 b15zdnd11an1n08x5 FILLER_288_2144 ();
 b15zdnd00an1n02x5 FILLER_288_2152 ();
 b15zdnd11an1n64x5 FILLER_288_2162 ();
 b15zdnd11an1n32x5 FILLER_288_2226 ();
 b15zdnd11an1n16x5 FILLER_288_2258 ();
 b15zdnd00an1n02x5 FILLER_288_2274 ();
 b15zdnd11an1n64x5 FILLER_289_0 ();
 b15zdnd11an1n64x5 FILLER_289_64 ();
 b15zdnd11an1n64x5 FILLER_289_128 ();
 b15zdnd11an1n64x5 FILLER_289_192 ();
 b15zdnd11an1n64x5 FILLER_289_256 ();
 b15zdnd11an1n64x5 FILLER_289_320 ();
 b15zdnd11an1n16x5 FILLER_289_384 ();
 b15zdnd11an1n08x5 FILLER_289_400 ();
 b15zdnd11an1n04x5 FILLER_289_408 ();
 b15zdnd00an1n02x5 FILLER_289_412 ();
 b15zdnd00an1n01x5 FILLER_289_414 ();
 b15zdnd11an1n64x5 FILLER_289_422 ();
 b15zdnd11an1n64x5 FILLER_289_486 ();
 b15zdnd11an1n16x5 FILLER_289_550 ();
 b15zdnd11an1n08x5 FILLER_289_566 ();
 b15zdnd00an1n02x5 FILLER_289_574 ();
 b15zdnd11an1n64x5 FILLER_289_618 ();
 b15zdnd11an1n16x5 FILLER_289_682 ();
 b15zdnd11an1n04x5 FILLER_289_698 ();
 b15zdnd00an1n02x5 FILLER_289_702 ();
 b15zdnd11an1n64x5 FILLER_289_707 ();
 b15zdnd11an1n64x5 FILLER_289_771 ();
 b15zdnd11an1n64x5 FILLER_289_835 ();
 b15zdnd11an1n32x5 FILLER_289_899 ();
 b15zdnd00an1n02x5 FILLER_289_931 ();
 b15zdnd00an1n01x5 FILLER_289_933 ();
 b15zdnd11an1n04x5 FILLER_289_941 ();
 b15zdnd11an1n64x5 FILLER_289_997 ();
 b15zdnd11an1n64x5 FILLER_289_1061 ();
 b15zdnd11an1n32x5 FILLER_289_1125 ();
 b15zdnd11an1n08x5 FILLER_289_1157 ();
 b15zdnd11an1n04x5 FILLER_289_1165 ();
 b15zdnd00an1n02x5 FILLER_289_1169 ();
 b15zdnd11an1n64x5 FILLER_289_1223 ();
 b15zdnd11an1n64x5 FILLER_289_1287 ();
 b15zdnd11an1n64x5 FILLER_289_1351 ();
 b15zdnd11an1n32x5 FILLER_289_1415 ();
 b15zdnd11an1n08x5 FILLER_289_1447 ();
 b15zdnd11an1n32x5 FILLER_289_1470 ();
 b15zdnd00an1n02x5 FILLER_289_1502 ();
 b15zdnd00an1n01x5 FILLER_289_1504 ();
 b15zdnd11an1n16x5 FILLER_289_1526 ();
 b15zdnd00an1n02x5 FILLER_289_1542 ();
 b15zdnd00an1n01x5 FILLER_289_1544 ();
 b15zdnd11an1n04x5 FILLER_289_1548 ();
 b15zdnd11an1n64x5 FILLER_289_1555 ();
 b15zdnd11an1n64x5 FILLER_289_1619 ();
 b15zdnd11an1n64x5 FILLER_289_1683 ();
 b15zdnd11an1n64x5 FILLER_289_1747 ();
 b15zdnd11an1n64x5 FILLER_289_1811 ();
 b15zdnd11an1n32x5 FILLER_289_1875 ();
 b15zdnd11an1n16x5 FILLER_289_1907 ();
 b15zdnd00an1n02x5 FILLER_289_1923 ();
 b15zdnd00an1n01x5 FILLER_289_1925 ();
 b15zdnd11an1n64x5 FILLER_289_1929 ();
 b15zdnd11an1n64x5 FILLER_289_1993 ();
 b15zdnd11an1n64x5 FILLER_289_2057 ();
 b15zdnd11an1n64x5 FILLER_289_2121 ();
 b15zdnd11an1n64x5 FILLER_289_2185 ();
 b15zdnd11an1n32x5 FILLER_289_2249 ();
 b15zdnd00an1n02x5 FILLER_289_2281 ();
 b15zdnd00an1n01x5 FILLER_289_2283 ();
 b15zdnd11an1n64x5 FILLER_290_8 ();
 b15zdnd11an1n64x5 FILLER_290_72 ();
 b15zdnd11an1n64x5 FILLER_290_136 ();
 b15zdnd11an1n64x5 FILLER_290_200 ();
 b15zdnd11an1n64x5 FILLER_290_264 ();
 b15zdnd11an1n32x5 FILLER_290_328 ();
 b15zdnd11an1n16x5 FILLER_290_360 ();
 b15zdnd11an1n08x5 FILLER_290_376 ();
 b15zdnd11an1n04x5 FILLER_290_384 ();
 b15zdnd00an1n02x5 FILLER_290_388 ();
 b15zdnd11an1n64x5 FILLER_290_432 ();
 b15zdnd11an1n64x5 FILLER_290_496 ();
 b15zdnd11an1n64x5 FILLER_290_560 ();
 b15zdnd11an1n64x5 FILLER_290_624 ();
 b15zdnd11an1n08x5 FILLER_290_688 ();
 b15zdnd11an1n04x5 FILLER_290_696 ();
 b15zdnd00an1n02x5 FILLER_290_700 ();
 b15zdnd00an1n01x5 FILLER_290_702 ();
 b15zdnd00an1n02x5 FILLER_290_716 ();
 b15zdnd11an1n64x5 FILLER_290_726 ();
 b15zdnd11an1n64x5 FILLER_290_790 ();
 b15zdnd11an1n64x5 FILLER_290_854 ();
 b15zdnd11an1n32x5 FILLER_290_918 ();
 b15zdnd11an1n08x5 FILLER_290_950 ();
 b15zdnd11an1n04x5 FILLER_290_958 ();
 b15zdnd11an1n04x5 FILLER_290_965 ();
 b15zdnd00an1n01x5 FILLER_290_969 ();
 b15zdnd11an1n64x5 FILLER_290_973 ();
 b15zdnd11an1n64x5 FILLER_290_1037 ();
 b15zdnd11an1n64x5 FILLER_290_1101 ();
 b15zdnd11an1n16x5 FILLER_290_1165 ();
 b15zdnd11an1n04x5 FILLER_290_1181 ();
 b15zdnd11an1n04x5 FILLER_290_1216 ();
 b15zdnd11an1n64x5 FILLER_290_1246 ();
 b15zdnd11an1n64x5 FILLER_290_1310 ();
 b15zdnd11an1n64x5 FILLER_290_1374 ();
 b15zdnd11an1n08x5 FILLER_290_1438 ();
 b15zdnd11an1n04x5 FILLER_290_1446 ();
 b15zdnd11an1n32x5 FILLER_290_1455 ();
 b15zdnd11an1n16x5 FILLER_290_1487 ();
 b15zdnd00an1n02x5 FILLER_290_1503 ();
 b15zdnd11an1n04x5 FILLER_290_1509 ();
 b15zdnd11an1n64x5 FILLER_290_1553 ();
 b15zdnd11an1n64x5 FILLER_290_1617 ();
 b15zdnd11an1n64x5 FILLER_290_1681 ();
 b15zdnd11an1n64x5 FILLER_290_1745 ();
 b15zdnd11an1n64x5 FILLER_290_1809 ();
 b15zdnd11an1n64x5 FILLER_290_1873 ();
 b15zdnd11an1n64x5 FILLER_290_1937 ();
 b15zdnd11an1n64x5 FILLER_290_2001 ();
 b15zdnd11an1n64x5 FILLER_290_2065 ();
 b15zdnd11an1n16x5 FILLER_290_2129 ();
 b15zdnd11an1n08x5 FILLER_290_2145 ();
 b15zdnd00an1n01x5 FILLER_290_2153 ();
 b15zdnd11an1n64x5 FILLER_290_2162 ();
 b15zdnd11an1n32x5 FILLER_290_2226 ();
 b15zdnd11an1n16x5 FILLER_290_2258 ();
 b15zdnd00an1n02x5 FILLER_290_2274 ();
 b15zdnd11an1n64x5 FILLER_291_0 ();
 b15zdnd11an1n64x5 FILLER_291_64 ();
 b15zdnd11an1n64x5 FILLER_291_128 ();
 b15zdnd11an1n64x5 FILLER_291_192 ();
 b15zdnd11an1n32x5 FILLER_291_256 ();
 b15zdnd11an1n16x5 FILLER_291_288 ();
 b15zdnd00an1n01x5 FILLER_291_304 ();
 b15zdnd11an1n64x5 FILLER_291_314 ();
 b15zdnd11an1n16x5 FILLER_291_378 ();
 b15zdnd11an1n04x5 FILLER_291_394 ();
 b15zdnd00an1n02x5 FILLER_291_398 ();
 b15zdnd00an1n01x5 FILLER_291_400 ();
 b15zdnd11an1n64x5 FILLER_291_443 ();
 b15zdnd11an1n64x5 FILLER_291_507 ();
 b15zdnd11an1n64x5 FILLER_291_571 ();
 b15zdnd11an1n64x5 FILLER_291_635 ();
 b15zdnd11an1n08x5 FILLER_291_699 ();
 b15zdnd00an1n02x5 FILLER_291_707 ();
 b15zdnd11an1n08x5 FILLER_291_713 ();
 b15zdnd11an1n04x5 FILLER_291_721 ();
 b15zdnd00an1n01x5 FILLER_291_725 ();
 b15zdnd11an1n04x5 FILLER_291_735 ();
 b15zdnd11an1n64x5 FILLER_291_748 ();
 b15zdnd11an1n32x5 FILLER_291_812 ();
 b15zdnd11an1n04x5 FILLER_291_844 ();
 b15zdnd00an1n02x5 FILLER_291_848 ();
 b15zdnd11an1n64x5 FILLER_291_902 ();
 b15zdnd11an1n32x5 FILLER_291_966 ();
 b15zdnd11an1n16x5 FILLER_291_998 ();
 b15zdnd00an1n02x5 FILLER_291_1014 ();
 b15zdnd11an1n04x5 FILLER_291_1039 ();
 b15zdnd11an1n64x5 FILLER_291_1059 ();
 b15zdnd11an1n64x5 FILLER_291_1123 ();
 b15zdnd11an1n64x5 FILLER_291_1187 ();
 b15zdnd11an1n64x5 FILLER_291_1251 ();
 b15zdnd11an1n64x5 FILLER_291_1315 ();
 b15zdnd11an1n64x5 FILLER_291_1379 ();
 b15zdnd11an1n08x5 FILLER_291_1443 ();
 b15zdnd00an1n02x5 FILLER_291_1451 ();
 b15zdnd11an1n64x5 FILLER_291_1495 ();
 b15zdnd11an1n32x5 FILLER_291_1559 ();
 b15zdnd11an1n16x5 FILLER_291_1591 ();
 b15zdnd11an1n04x5 FILLER_291_1607 ();
 b15zdnd00an1n01x5 FILLER_291_1611 ();
 b15zdnd11an1n64x5 FILLER_291_1654 ();
 b15zdnd11an1n64x5 FILLER_291_1718 ();
 b15zdnd11an1n64x5 FILLER_291_1782 ();
 b15zdnd11an1n64x5 FILLER_291_1846 ();
 b15zdnd11an1n64x5 FILLER_291_1910 ();
 b15zdnd11an1n64x5 FILLER_291_1974 ();
 b15zdnd11an1n64x5 FILLER_291_2038 ();
 b15zdnd11an1n64x5 FILLER_291_2102 ();
 b15zdnd11an1n64x5 FILLER_291_2166 ();
 b15zdnd11an1n32x5 FILLER_291_2230 ();
 b15zdnd11an1n16x5 FILLER_291_2262 ();
 b15zdnd11an1n04x5 FILLER_291_2278 ();
 b15zdnd00an1n02x5 FILLER_291_2282 ();
 b15zdnd11an1n64x5 FILLER_292_8 ();
 b15zdnd11an1n64x5 FILLER_292_72 ();
 b15zdnd11an1n64x5 FILLER_292_136 ();
 b15zdnd11an1n16x5 FILLER_292_200 ();
 b15zdnd11an1n08x5 FILLER_292_216 ();
 b15zdnd11an1n04x5 FILLER_292_224 ();
 b15zdnd00an1n02x5 FILLER_292_228 ();
 b15zdnd00an1n01x5 FILLER_292_230 ();
 b15zdnd11an1n64x5 FILLER_292_273 ();
 b15zdnd11an1n64x5 FILLER_292_337 ();
 b15zdnd11an1n64x5 FILLER_292_401 ();
 b15zdnd11an1n64x5 FILLER_292_465 ();
 b15zdnd11an1n64x5 FILLER_292_529 ();
 b15zdnd11an1n64x5 FILLER_292_593 ();
 b15zdnd11an1n32x5 FILLER_292_657 ();
 b15zdnd11an1n08x5 FILLER_292_689 ();
 b15zdnd11an1n04x5 FILLER_292_697 ();
 b15zdnd00an1n02x5 FILLER_292_701 ();
 b15zdnd11an1n08x5 FILLER_292_707 ();
 b15zdnd00an1n02x5 FILLER_292_715 ();
 b15zdnd00an1n01x5 FILLER_292_717 ();
 b15zdnd11an1n64x5 FILLER_292_726 ();
 b15zdnd11an1n08x5 FILLER_292_790 ();
 b15zdnd11an1n04x5 FILLER_292_798 ();
 b15zdnd11an1n16x5 FILLER_292_844 ();
 b15zdnd11an1n08x5 FILLER_292_860 ();
 b15zdnd00an1n02x5 FILLER_292_868 ();
 b15zdnd11an1n04x5 FILLER_292_873 ();
 b15zdnd11an1n64x5 FILLER_292_880 ();
 b15zdnd11an1n64x5 FILLER_292_944 ();
 b15zdnd11an1n08x5 FILLER_292_1008 ();
 b15zdnd00an1n02x5 FILLER_292_1016 ();
 b15zdnd00an1n01x5 FILLER_292_1018 ();
 b15zdnd11an1n64x5 FILLER_292_1042 ();
 b15zdnd11an1n64x5 FILLER_292_1106 ();
 b15zdnd11an1n64x5 FILLER_292_1170 ();
 b15zdnd11an1n64x5 FILLER_292_1234 ();
 b15zdnd11an1n64x5 FILLER_292_1298 ();
 b15zdnd11an1n64x5 FILLER_292_1362 ();
 b15zdnd11an1n32x5 FILLER_292_1426 ();
 b15zdnd11an1n16x5 FILLER_292_1458 ();
 b15zdnd00an1n02x5 FILLER_292_1474 ();
 b15zdnd00an1n01x5 FILLER_292_1476 ();
 b15zdnd11an1n64x5 FILLER_292_1519 ();
 b15zdnd11an1n64x5 FILLER_292_1583 ();
 b15zdnd11an1n64x5 FILLER_292_1647 ();
 b15zdnd11an1n64x5 FILLER_292_1711 ();
 b15zdnd11an1n64x5 FILLER_292_1775 ();
 b15zdnd11an1n64x5 FILLER_292_1839 ();
 b15zdnd11an1n32x5 FILLER_292_1903 ();
 b15zdnd11an1n16x5 FILLER_292_1935 ();
 b15zdnd00an1n01x5 FILLER_292_1951 ();
 b15zdnd11an1n64x5 FILLER_292_1994 ();
 b15zdnd11an1n64x5 FILLER_292_2058 ();
 b15zdnd11an1n32x5 FILLER_292_2122 ();
 b15zdnd11an1n64x5 FILLER_292_2162 ();
 b15zdnd11an1n32x5 FILLER_292_2226 ();
 b15zdnd11an1n16x5 FILLER_292_2258 ();
 b15zdnd00an1n02x5 FILLER_292_2274 ();
 b15zdnd11an1n16x5 FILLER_293_0 ();
 b15zdnd11an1n04x5 FILLER_293_16 ();
 b15zdnd11an1n64x5 FILLER_293_28 ();
 b15zdnd11an1n64x5 FILLER_293_92 ();
 b15zdnd11an1n64x5 FILLER_293_156 ();
 b15zdnd11an1n64x5 FILLER_293_220 ();
 b15zdnd11an1n64x5 FILLER_293_284 ();
 b15zdnd11an1n64x5 FILLER_293_348 ();
 b15zdnd11an1n64x5 FILLER_293_412 ();
 b15zdnd11an1n64x5 FILLER_293_476 ();
 b15zdnd11an1n64x5 FILLER_293_540 ();
 b15zdnd11an1n64x5 FILLER_293_604 ();
 b15zdnd11an1n64x5 FILLER_293_668 ();
 b15zdnd11an1n64x5 FILLER_293_732 ();
 b15zdnd11an1n64x5 FILLER_293_796 ();
 b15zdnd11an1n16x5 FILLER_293_860 ();
 b15zdnd11an1n64x5 FILLER_293_879 ();
 b15zdnd11an1n16x5 FILLER_293_943 ();
 b15zdnd00an1n02x5 FILLER_293_959 ();
 b15zdnd00an1n01x5 FILLER_293_961 ();
 b15zdnd11an1n64x5 FILLER_293_968 ();
 b15zdnd11an1n16x5 FILLER_293_1032 ();
 b15zdnd11an1n04x5 FILLER_293_1048 ();
 b15zdnd00an1n02x5 FILLER_293_1052 ();
 b15zdnd11an1n64x5 FILLER_293_1077 ();
 b15zdnd11an1n64x5 FILLER_293_1141 ();
 b15zdnd00an1n02x5 FILLER_293_1205 ();
 b15zdnd00an1n01x5 FILLER_293_1207 ();
 b15zdnd11an1n64x5 FILLER_293_1236 ();
 b15zdnd00an1n01x5 FILLER_293_1300 ();
 b15zdnd11an1n08x5 FILLER_293_1304 ();
 b15zdnd00an1n02x5 FILLER_293_1312 ();
 b15zdnd00an1n01x5 FILLER_293_1314 ();
 b15zdnd11an1n64x5 FILLER_293_1324 ();
 b15zdnd11an1n64x5 FILLER_293_1388 ();
 b15zdnd11an1n64x5 FILLER_293_1452 ();
 b15zdnd11an1n64x5 FILLER_293_1516 ();
 b15zdnd11an1n16x5 FILLER_293_1580 ();
 b15zdnd11an1n08x5 FILLER_293_1596 ();
 b15zdnd11an1n04x5 FILLER_293_1604 ();
 b15zdnd00an1n02x5 FILLER_293_1608 ();
 b15zdnd00an1n01x5 FILLER_293_1610 ();
 b15zdnd11an1n64x5 FILLER_293_1653 ();
 b15zdnd11an1n64x5 FILLER_293_1717 ();
 b15zdnd11an1n64x5 FILLER_293_1781 ();
 b15zdnd11an1n64x5 FILLER_293_1845 ();
 b15zdnd11an1n64x5 FILLER_293_1909 ();
 b15zdnd11an1n64x5 FILLER_293_1973 ();
 b15zdnd11an1n64x5 FILLER_293_2037 ();
 b15zdnd11an1n64x5 FILLER_293_2101 ();
 b15zdnd11an1n64x5 FILLER_293_2165 ();
 b15zdnd11an1n32x5 FILLER_293_2229 ();
 b15zdnd11an1n16x5 FILLER_293_2261 ();
 b15zdnd11an1n04x5 FILLER_293_2277 ();
 b15zdnd00an1n02x5 FILLER_293_2281 ();
 b15zdnd00an1n01x5 FILLER_293_2283 ();
 b15zdnd11an1n64x5 FILLER_294_8 ();
 b15zdnd11an1n64x5 FILLER_294_72 ();
 b15zdnd11an1n64x5 FILLER_294_136 ();
 b15zdnd11an1n64x5 FILLER_294_200 ();
 b15zdnd11an1n64x5 FILLER_294_264 ();
 b15zdnd11an1n64x5 FILLER_294_328 ();
 b15zdnd11an1n64x5 FILLER_294_392 ();
 b15zdnd11an1n64x5 FILLER_294_456 ();
 b15zdnd11an1n64x5 FILLER_294_520 ();
 b15zdnd11an1n64x5 FILLER_294_584 ();
 b15zdnd11an1n64x5 FILLER_294_648 ();
 b15zdnd11an1n04x5 FILLER_294_712 ();
 b15zdnd00an1n02x5 FILLER_294_716 ();
 b15zdnd11an1n64x5 FILLER_294_726 ();
 b15zdnd11an1n64x5 FILLER_294_790 ();
 b15zdnd11an1n64x5 FILLER_294_854 ();
 b15zdnd11an1n64x5 FILLER_294_918 ();
 b15zdnd11an1n16x5 FILLER_294_982 ();
 b15zdnd11an1n08x5 FILLER_294_998 ();
 b15zdnd11an1n04x5 FILLER_294_1006 ();
 b15zdnd11an1n16x5 FILLER_294_1018 ();
 b15zdnd11an1n08x5 FILLER_294_1034 ();
 b15zdnd00an1n02x5 FILLER_294_1042 ();
 b15zdnd00an1n01x5 FILLER_294_1044 ();
 b15zdnd11an1n64x5 FILLER_294_1087 ();
 b15zdnd11an1n64x5 FILLER_294_1151 ();
 b15zdnd11an1n64x5 FILLER_294_1215 ();
 b15zdnd11an1n08x5 FILLER_294_1279 ();
 b15zdnd11an1n04x5 FILLER_294_1287 ();
 b15zdnd00an1n02x5 FILLER_294_1291 ();
 b15zdnd00an1n01x5 FILLER_294_1293 ();
 b15zdnd11an1n04x5 FILLER_294_1297 ();
 b15zdnd11an1n04x5 FILLER_294_1306 ();
 b15zdnd11an1n04x5 FILLER_294_1318 ();
 b15zdnd11an1n64x5 FILLER_294_1364 ();
 b15zdnd11an1n64x5 FILLER_294_1428 ();
 b15zdnd11an1n64x5 FILLER_294_1492 ();
 b15zdnd11an1n64x5 FILLER_294_1556 ();
 b15zdnd11an1n64x5 FILLER_294_1620 ();
 b15zdnd11an1n64x5 FILLER_294_1684 ();
 b15zdnd11an1n64x5 FILLER_294_1748 ();
 b15zdnd11an1n64x5 FILLER_294_1812 ();
 b15zdnd11an1n64x5 FILLER_294_1876 ();
 b15zdnd11an1n32x5 FILLER_294_1940 ();
 b15zdnd11an1n04x5 FILLER_294_1972 ();
 b15zdnd00an1n02x5 FILLER_294_1976 ();
 b15zdnd11an1n64x5 FILLER_294_2018 ();
 b15zdnd11an1n64x5 FILLER_294_2082 ();
 b15zdnd11an1n08x5 FILLER_294_2146 ();
 b15zdnd11an1n64x5 FILLER_294_2162 ();
 b15zdnd11an1n32x5 FILLER_294_2226 ();
 b15zdnd11an1n16x5 FILLER_294_2258 ();
 b15zdnd00an1n02x5 FILLER_294_2274 ();
 b15zdnd11an1n64x5 FILLER_295_0 ();
 b15zdnd11an1n64x5 FILLER_295_64 ();
 b15zdnd11an1n64x5 FILLER_295_128 ();
 b15zdnd11an1n64x5 FILLER_295_192 ();
 b15zdnd11an1n64x5 FILLER_295_256 ();
 b15zdnd11an1n64x5 FILLER_295_320 ();
 b15zdnd11an1n64x5 FILLER_295_384 ();
 b15zdnd11an1n64x5 FILLER_295_448 ();
 b15zdnd11an1n64x5 FILLER_295_512 ();
 b15zdnd11an1n32x5 FILLER_295_576 ();
 b15zdnd11an1n16x5 FILLER_295_608 ();
 b15zdnd11an1n08x5 FILLER_295_624 ();
 b15zdnd11an1n04x5 FILLER_295_632 ();
 b15zdnd00an1n02x5 FILLER_295_636 ();
 b15zdnd00an1n01x5 FILLER_295_638 ();
 b15zdnd11an1n32x5 FILLER_295_642 ();
 b15zdnd11an1n08x5 FILLER_295_674 ();
 b15zdnd11an1n04x5 FILLER_295_682 ();
 b15zdnd00an1n02x5 FILLER_295_686 ();
 b15zdnd00an1n01x5 FILLER_295_688 ();
 b15zdnd11an1n64x5 FILLER_295_731 ();
 b15zdnd11an1n64x5 FILLER_295_795 ();
 b15zdnd11an1n64x5 FILLER_295_859 ();
 b15zdnd11an1n64x5 FILLER_295_923 ();
 b15zdnd11an1n32x5 FILLER_295_987 ();
 b15zdnd11an1n04x5 FILLER_295_1019 ();
 b15zdnd00an1n02x5 FILLER_295_1023 ();
 b15zdnd11an1n16x5 FILLER_295_1048 ();
 b15zdnd00an1n02x5 FILLER_295_1064 ();
 b15zdnd11an1n64x5 FILLER_295_1086 ();
 b15zdnd11an1n64x5 FILLER_295_1150 ();
 b15zdnd11an1n64x5 FILLER_295_1214 ();
 b15zdnd11an1n08x5 FILLER_295_1278 ();
 b15zdnd11an1n04x5 FILLER_295_1289 ();
 b15zdnd11an1n64x5 FILLER_295_1335 ();
 b15zdnd11an1n16x5 FILLER_295_1399 ();
 b15zdnd11an1n08x5 FILLER_295_1415 ();
 b15zdnd11an1n04x5 FILLER_295_1423 ();
 b15zdnd11an1n04x5 FILLER_295_1466 ();
 b15zdnd00an1n01x5 FILLER_295_1470 ();
 b15zdnd11an1n04x5 FILLER_295_1474 ();
 b15zdnd11an1n64x5 FILLER_295_1481 ();
 b15zdnd11an1n64x5 FILLER_295_1545 ();
 b15zdnd11an1n64x5 FILLER_295_1609 ();
 b15zdnd11an1n64x5 FILLER_295_1673 ();
 b15zdnd11an1n64x5 FILLER_295_1737 ();
 b15zdnd11an1n64x5 FILLER_295_1801 ();
 b15zdnd11an1n64x5 FILLER_295_1865 ();
 b15zdnd11an1n64x5 FILLER_295_1929 ();
 b15zdnd11an1n04x5 FILLER_295_1993 ();
 b15zdnd00an1n02x5 FILLER_295_1997 ();
 b15zdnd00an1n01x5 FILLER_295_1999 ();
 b15zdnd11an1n04x5 FILLER_295_2007 ();
 b15zdnd00an1n02x5 FILLER_295_2011 ();
 b15zdnd00an1n01x5 FILLER_295_2013 ();
 b15zdnd11an1n64x5 FILLER_295_2017 ();
 b15zdnd11an1n64x5 FILLER_295_2081 ();
 b15zdnd11an1n64x5 FILLER_295_2145 ();
 b15zdnd11an1n64x5 FILLER_295_2209 ();
 b15zdnd11an1n08x5 FILLER_295_2273 ();
 b15zdnd00an1n02x5 FILLER_295_2281 ();
 b15zdnd00an1n01x5 FILLER_295_2283 ();
 b15zdnd11an1n64x5 FILLER_296_8 ();
 b15zdnd11an1n64x5 FILLER_296_72 ();
 b15zdnd11an1n64x5 FILLER_296_136 ();
 b15zdnd11an1n64x5 FILLER_296_200 ();
 b15zdnd11an1n64x5 FILLER_296_264 ();
 b15zdnd11an1n32x5 FILLER_296_328 ();
 b15zdnd11an1n04x5 FILLER_296_360 ();
 b15zdnd00an1n02x5 FILLER_296_364 ();
 b15zdnd00an1n01x5 FILLER_296_366 ();
 b15zdnd11an1n32x5 FILLER_296_370 ();
 b15zdnd11an1n16x5 FILLER_296_402 ();
 b15zdnd00an1n01x5 FILLER_296_418 ();
 b15zdnd11an1n64x5 FILLER_296_461 ();
 b15zdnd11an1n64x5 FILLER_296_525 ();
 b15zdnd11an1n08x5 FILLER_296_589 ();
 b15zdnd11an1n04x5 FILLER_296_597 ();
 b15zdnd00an1n02x5 FILLER_296_601 ();
 b15zdnd11an1n64x5 FILLER_296_643 ();
 b15zdnd11an1n08x5 FILLER_296_707 ();
 b15zdnd00an1n02x5 FILLER_296_715 ();
 b15zdnd00an1n01x5 FILLER_296_717 ();
 b15zdnd11an1n32x5 FILLER_296_726 ();
 b15zdnd11an1n16x5 FILLER_296_758 ();
 b15zdnd00an1n02x5 FILLER_296_774 ();
 b15zdnd00an1n01x5 FILLER_296_776 ();
 b15zdnd11an1n64x5 FILLER_296_816 ();
 b15zdnd11an1n64x5 FILLER_296_880 ();
 b15zdnd11an1n32x5 FILLER_296_944 ();
 b15zdnd11an1n08x5 FILLER_296_976 ();
 b15zdnd11an1n04x5 FILLER_296_984 ();
 b15zdnd11an1n64x5 FILLER_296_996 ();
 b15zdnd11an1n08x5 FILLER_296_1060 ();
 b15zdnd11an1n04x5 FILLER_296_1068 ();
 b15zdnd00an1n01x5 FILLER_296_1072 ();
 b15zdnd11an1n16x5 FILLER_296_1084 ();
 b15zdnd00an1n01x5 FILLER_296_1100 ();
 b15zdnd11an1n64x5 FILLER_296_1111 ();
 b15zdnd11an1n64x5 FILLER_296_1175 ();
 b15zdnd11an1n32x5 FILLER_296_1239 ();
 b15zdnd11an1n04x5 FILLER_296_1271 ();
 b15zdnd11an1n04x5 FILLER_296_1327 ();
 b15zdnd11an1n64x5 FILLER_296_1373 ();
 b15zdnd11an1n08x5 FILLER_296_1437 ();
 b15zdnd00an1n01x5 FILLER_296_1445 ();
 b15zdnd11an1n64x5 FILLER_296_1498 ();
 b15zdnd11an1n64x5 FILLER_296_1562 ();
 b15zdnd11an1n64x5 FILLER_296_1626 ();
 b15zdnd11an1n64x5 FILLER_296_1690 ();
 b15zdnd11an1n64x5 FILLER_296_1754 ();
 b15zdnd11an1n64x5 FILLER_296_1818 ();
 b15zdnd11an1n64x5 FILLER_296_1882 ();
 b15zdnd11an1n64x5 FILLER_296_1946 ();
 b15zdnd11an1n04x5 FILLER_296_2010 ();
 b15zdnd00an1n01x5 FILLER_296_2014 ();
 b15zdnd11an1n64x5 FILLER_296_2018 ();
 b15zdnd11an1n64x5 FILLER_296_2082 ();
 b15zdnd11an1n08x5 FILLER_296_2146 ();
 b15zdnd11an1n64x5 FILLER_296_2162 ();
 b15zdnd11an1n32x5 FILLER_296_2226 ();
 b15zdnd11an1n16x5 FILLER_296_2258 ();
 b15zdnd00an1n02x5 FILLER_296_2274 ();
 b15zdnd11an1n64x5 FILLER_297_0 ();
 b15zdnd11an1n64x5 FILLER_297_64 ();
 b15zdnd11an1n64x5 FILLER_297_128 ();
 b15zdnd11an1n64x5 FILLER_297_192 ();
 b15zdnd11an1n64x5 FILLER_297_256 ();
 b15zdnd11an1n16x5 FILLER_297_320 ();
 b15zdnd11an1n08x5 FILLER_297_336 ();
 b15zdnd11an1n64x5 FILLER_297_396 ();
 b15zdnd11an1n64x5 FILLER_297_460 ();
 b15zdnd11an1n64x5 FILLER_297_524 ();
 b15zdnd11an1n32x5 FILLER_297_588 ();
 b15zdnd11an1n16x5 FILLER_297_620 ();
 b15zdnd11an1n04x5 FILLER_297_636 ();
 b15zdnd11an1n64x5 FILLER_297_643 ();
 b15zdnd11an1n64x5 FILLER_297_707 ();
 b15zdnd11an1n08x5 FILLER_297_771 ();
 b15zdnd11an1n04x5 FILLER_297_779 ();
 b15zdnd00an1n02x5 FILLER_297_783 ();
 b15zdnd00an1n01x5 FILLER_297_785 ();
 b15zdnd11an1n64x5 FILLER_297_794 ();
 b15zdnd11an1n08x5 FILLER_297_858 ();
 b15zdnd11an1n04x5 FILLER_297_866 ();
 b15zdnd00an1n01x5 FILLER_297_870 ();
 b15zdnd11an1n64x5 FILLER_297_913 ();
 b15zdnd11an1n64x5 FILLER_297_977 ();
 b15zdnd11an1n32x5 FILLER_297_1041 ();
 b15zdnd11an1n04x5 FILLER_297_1073 ();
 b15zdnd00an1n02x5 FILLER_297_1077 ();
 b15zdnd11an1n04x5 FILLER_297_1086 ();
 b15zdnd11an1n64x5 FILLER_297_1099 ();
 b15zdnd11an1n64x5 FILLER_297_1163 ();
 b15zdnd11an1n64x5 FILLER_297_1227 ();
 b15zdnd11an1n08x5 FILLER_297_1291 ();
 b15zdnd00an1n02x5 FILLER_297_1299 ();
 b15zdnd00an1n01x5 FILLER_297_1301 ();
 b15zdnd11an1n32x5 FILLER_297_1344 ();
 b15zdnd11an1n04x5 FILLER_297_1376 ();
 b15zdnd11an1n32x5 FILLER_297_1408 ();
 b15zdnd11an1n16x5 FILLER_297_1440 ();
 b15zdnd00an1n02x5 FILLER_297_1456 ();
 b15zdnd11an1n04x5 FILLER_297_1466 ();
 b15zdnd00an1n02x5 FILLER_297_1470 ();
 b15zdnd11an1n64x5 FILLER_297_1475 ();
 b15zdnd11an1n16x5 FILLER_297_1539 ();
 b15zdnd11an1n08x5 FILLER_297_1555 ();
 b15zdnd00an1n01x5 FILLER_297_1563 ();
 b15zdnd11an1n64x5 FILLER_297_1616 ();
 b15zdnd11an1n64x5 FILLER_297_1680 ();
 b15zdnd11an1n64x5 FILLER_297_1744 ();
 b15zdnd11an1n64x5 FILLER_297_1808 ();
 b15zdnd11an1n64x5 FILLER_297_1872 ();
 b15zdnd11an1n64x5 FILLER_297_1936 ();
 b15zdnd11an1n64x5 FILLER_297_2000 ();
 b15zdnd11an1n64x5 FILLER_297_2064 ();
 b15zdnd11an1n64x5 FILLER_297_2128 ();
 b15zdnd11an1n64x5 FILLER_297_2192 ();
 b15zdnd11an1n16x5 FILLER_297_2256 ();
 b15zdnd11an1n08x5 FILLER_297_2272 ();
 b15zdnd11an1n04x5 FILLER_297_2280 ();
 b15zdnd11an1n64x5 FILLER_298_8 ();
 b15zdnd11an1n64x5 FILLER_298_72 ();
 b15zdnd11an1n64x5 FILLER_298_136 ();
 b15zdnd11an1n64x5 FILLER_298_200 ();
 b15zdnd11an1n64x5 FILLER_298_264 ();
 b15zdnd11an1n32x5 FILLER_298_328 ();
 b15zdnd00an1n02x5 FILLER_298_360 ();
 b15zdnd00an1n01x5 FILLER_298_362 ();
 b15zdnd11an1n04x5 FILLER_298_366 ();
 b15zdnd11an1n64x5 FILLER_298_373 ();
 b15zdnd11an1n64x5 FILLER_298_437 ();
 b15zdnd11an1n16x5 FILLER_298_501 ();
 b15zdnd11an1n08x5 FILLER_298_517 ();
 b15zdnd11an1n04x5 FILLER_298_525 ();
 b15zdnd00an1n01x5 FILLER_298_529 ();
 b15zdnd11an1n04x5 FILLER_298_533 ();
 b15zdnd00an1n01x5 FILLER_298_537 ();
 b15zdnd11an1n64x5 FILLER_298_569 ();
 b15zdnd11an1n08x5 FILLER_298_633 ();
 b15zdnd00an1n02x5 FILLER_298_641 ();
 b15zdnd00an1n01x5 FILLER_298_643 ();
 b15zdnd11an1n16x5 FILLER_298_696 ();
 b15zdnd11an1n04x5 FILLER_298_712 ();
 b15zdnd00an1n02x5 FILLER_298_716 ();
 b15zdnd11an1n32x5 FILLER_298_726 ();
 b15zdnd11an1n16x5 FILLER_298_758 ();
 b15zdnd11an1n08x5 FILLER_298_774 ();
 b15zdnd11an1n04x5 FILLER_298_782 ();
 b15zdnd11an1n32x5 FILLER_298_828 ();
 b15zdnd11an1n04x5 FILLER_298_860 ();
 b15zdnd11an1n64x5 FILLER_298_906 ();
 b15zdnd11an1n64x5 FILLER_298_970 ();
 b15zdnd11an1n64x5 FILLER_298_1034 ();
 b15zdnd11an1n64x5 FILLER_298_1098 ();
 b15zdnd11an1n64x5 FILLER_298_1162 ();
 b15zdnd11an1n64x5 FILLER_298_1226 ();
 b15zdnd11an1n08x5 FILLER_298_1290 ();
 b15zdnd00an1n01x5 FILLER_298_1298 ();
 b15zdnd11an1n04x5 FILLER_298_1307 ();
 b15zdnd11an1n64x5 FILLER_298_1317 ();
 b15zdnd11an1n64x5 FILLER_298_1381 ();
 b15zdnd11an1n64x5 FILLER_298_1445 ();
 b15zdnd11an1n64x5 FILLER_298_1509 ();
 b15zdnd11an1n08x5 FILLER_298_1573 ();
 b15zdnd00an1n01x5 FILLER_298_1581 ();
 b15zdnd11an1n04x5 FILLER_298_1585 ();
 b15zdnd11an1n04x5 FILLER_298_1592 ();
 b15zdnd11an1n64x5 FILLER_298_1599 ();
 b15zdnd11an1n32x5 FILLER_298_1663 ();
 b15zdnd11an1n16x5 FILLER_298_1695 ();
 b15zdnd00an1n02x5 FILLER_298_1711 ();
 b15zdnd00an1n01x5 FILLER_298_1713 ();
 b15zdnd11an1n04x5 FILLER_298_1717 ();
 b15zdnd11an1n64x5 FILLER_298_1746 ();
 b15zdnd11an1n64x5 FILLER_298_1810 ();
 b15zdnd11an1n64x5 FILLER_298_1874 ();
 b15zdnd11an1n64x5 FILLER_298_1938 ();
 b15zdnd11an1n32x5 FILLER_298_2002 ();
 b15zdnd11an1n64x5 FILLER_298_2037 ();
 b15zdnd11an1n32x5 FILLER_298_2101 ();
 b15zdnd11an1n16x5 FILLER_298_2133 ();
 b15zdnd11an1n04x5 FILLER_298_2149 ();
 b15zdnd00an1n01x5 FILLER_298_2153 ();
 b15zdnd11an1n64x5 FILLER_298_2162 ();
 b15zdnd11an1n32x5 FILLER_298_2226 ();
 b15zdnd11an1n16x5 FILLER_298_2258 ();
 b15zdnd00an1n02x5 FILLER_298_2274 ();
 b15zdnd11an1n64x5 FILLER_299_0 ();
 b15zdnd11an1n64x5 FILLER_299_64 ();
 b15zdnd11an1n64x5 FILLER_299_128 ();
 b15zdnd11an1n64x5 FILLER_299_192 ();
 b15zdnd11an1n64x5 FILLER_299_256 ();
 b15zdnd11an1n64x5 FILLER_299_320 ();
 b15zdnd11an1n64x5 FILLER_299_384 ();
 b15zdnd11an1n64x5 FILLER_299_448 ();
 b15zdnd11an1n08x5 FILLER_299_512 ();
 b15zdnd00an1n02x5 FILLER_299_520 ();
 b15zdnd00an1n01x5 FILLER_299_522 ();
 b15zdnd11an1n64x5 FILLER_299_565 ();
 b15zdnd11an1n32x5 FILLER_299_629 ();
 b15zdnd11an1n04x5 FILLER_299_661 ();
 b15zdnd00an1n02x5 FILLER_299_665 ();
 b15zdnd11an1n64x5 FILLER_299_670 ();
 b15zdnd11an1n64x5 FILLER_299_734 ();
 b15zdnd11an1n32x5 FILLER_299_798 ();
 b15zdnd11an1n16x5 FILLER_299_830 ();
 b15zdnd11an1n08x5 FILLER_299_846 ();
 b15zdnd11an1n04x5 FILLER_299_854 ();
 b15zdnd00an1n02x5 FILLER_299_858 ();
 b15zdnd00an1n01x5 FILLER_299_860 ();
 b15zdnd11an1n64x5 FILLER_299_875 ();
 b15zdnd11an1n64x5 FILLER_299_939 ();
 b15zdnd00an1n02x5 FILLER_299_1003 ();
 b15zdnd00an1n01x5 FILLER_299_1005 ();
 b15zdnd11an1n32x5 FILLER_299_1013 ();
 b15zdnd11an1n16x5 FILLER_299_1045 ();
 b15zdnd11an1n08x5 FILLER_299_1061 ();
 b15zdnd00an1n01x5 FILLER_299_1069 ();
 b15zdnd11an1n64x5 FILLER_299_1093 ();
 b15zdnd11an1n64x5 FILLER_299_1157 ();
 b15zdnd11an1n64x5 FILLER_299_1221 ();
 b15zdnd11an1n16x5 FILLER_299_1285 ();
 b15zdnd11an1n04x5 FILLER_299_1301 ();
 b15zdnd11an1n04x5 FILLER_299_1311 ();
 b15zdnd11an1n64x5 FILLER_299_1319 ();
 b15zdnd11an1n64x5 FILLER_299_1383 ();
 b15zdnd11an1n64x5 FILLER_299_1447 ();
 b15zdnd11an1n64x5 FILLER_299_1511 ();
 b15zdnd11an1n64x5 FILLER_299_1575 ();
 b15zdnd11an1n64x5 FILLER_299_1639 ();
 b15zdnd11an1n04x5 FILLER_299_1703 ();
 b15zdnd00an1n02x5 FILLER_299_1707 ();
 b15zdnd00an1n01x5 FILLER_299_1709 ();
 b15zdnd11an1n04x5 FILLER_299_1713 ();
 b15zdnd11an1n16x5 FILLER_299_1720 ();
 b15zdnd11an1n04x5 FILLER_299_1736 ();
 b15zdnd00an1n01x5 FILLER_299_1740 ();
 b15zdnd11an1n64x5 FILLER_299_1783 ();
 b15zdnd11an1n64x5 FILLER_299_1847 ();
 b15zdnd11an1n64x5 FILLER_299_1911 ();
 b15zdnd11an1n32x5 FILLER_299_1975 ();
 b15zdnd11an1n16x5 FILLER_299_2007 ();
 b15zdnd11an1n08x5 FILLER_299_2023 ();
 b15zdnd00an1n01x5 FILLER_299_2031 ();
 b15zdnd11an1n04x5 FILLER_299_2035 ();
 b15zdnd11an1n08x5 FILLER_299_2042 ();
 b15zdnd11an1n04x5 FILLER_299_2050 ();
 b15zdnd00an1n02x5 FILLER_299_2054 ();
 b15zdnd00an1n01x5 FILLER_299_2056 ();
 b15zdnd11an1n64x5 FILLER_299_2060 ();
 b15zdnd11an1n64x5 FILLER_299_2124 ();
 b15zdnd11an1n64x5 FILLER_299_2188 ();
 b15zdnd11an1n32x5 FILLER_299_2252 ();
 b15zdnd11an1n64x5 FILLER_300_8 ();
 b15zdnd11an1n64x5 FILLER_300_72 ();
 b15zdnd11an1n64x5 FILLER_300_136 ();
 b15zdnd11an1n64x5 FILLER_300_200 ();
 b15zdnd11an1n64x5 FILLER_300_264 ();
 b15zdnd11an1n64x5 FILLER_300_328 ();
 b15zdnd11an1n64x5 FILLER_300_392 ();
 b15zdnd11an1n32x5 FILLER_300_456 ();
 b15zdnd11an1n08x5 FILLER_300_488 ();
 b15zdnd11an1n04x5 FILLER_300_496 ();
 b15zdnd00an1n02x5 FILLER_300_500 ();
 b15zdnd00an1n01x5 FILLER_300_502 ();
 b15zdnd11an1n64x5 FILLER_300_555 ();
 b15zdnd11an1n32x5 FILLER_300_619 ();
 b15zdnd11an1n16x5 FILLER_300_651 ();
 b15zdnd11an1n04x5 FILLER_300_667 ();
 b15zdnd00an1n01x5 FILLER_300_671 ();
 b15zdnd11an1n32x5 FILLER_300_675 ();
 b15zdnd11an1n08x5 FILLER_300_707 ();
 b15zdnd00an1n02x5 FILLER_300_715 ();
 b15zdnd00an1n01x5 FILLER_300_717 ();
 b15zdnd11an1n64x5 FILLER_300_726 ();
 b15zdnd11an1n64x5 FILLER_300_790 ();
 b15zdnd11an1n64x5 FILLER_300_854 ();
 b15zdnd11an1n64x5 FILLER_300_918 ();
 b15zdnd11an1n16x5 FILLER_300_982 ();
 b15zdnd00an1n01x5 FILLER_300_998 ();
 b15zdnd11an1n64x5 FILLER_300_1041 ();
 b15zdnd11an1n64x5 FILLER_300_1105 ();
 b15zdnd11an1n64x5 FILLER_300_1169 ();
 b15zdnd11an1n64x5 FILLER_300_1233 ();
 b15zdnd11an1n04x5 FILLER_300_1297 ();
 b15zdnd00an1n01x5 FILLER_300_1301 ();
 b15zdnd11an1n64x5 FILLER_300_1312 ();
 b15zdnd11an1n64x5 FILLER_300_1376 ();
 b15zdnd11an1n64x5 FILLER_300_1440 ();
 b15zdnd11an1n64x5 FILLER_300_1504 ();
 b15zdnd11an1n64x5 FILLER_300_1568 ();
 b15zdnd11an1n32x5 FILLER_300_1632 ();
 b15zdnd11an1n16x5 FILLER_300_1664 ();
 b15zdnd11an1n08x5 FILLER_300_1680 ();
 b15zdnd11an1n04x5 FILLER_300_1688 ();
 b15zdnd11an1n64x5 FILLER_300_1744 ();
 b15zdnd11an1n64x5 FILLER_300_1808 ();
 b15zdnd11an1n64x5 FILLER_300_1872 ();
 b15zdnd11an1n32x5 FILLER_300_1936 ();
 b15zdnd11an1n16x5 FILLER_300_1968 ();
 b15zdnd11an1n04x5 FILLER_300_1984 ();
 b15zdnd11an1n16x5 FILLER_300_1995 ();
 b15zdnd00an1n02x5 FILLER_300_2011 ();
 b15zdnd00an1n01x5 FILLER_300_2013 ();
 b15zdnd11an1n64x5 FILLER_300_2066 ();
 b15zdnd11an1n16x5 FILLER_300_2130 ();
 b15zdnd11an1n08x5 FILLER_300_2146 ();
 b15zdnd11an1n64x5 FILLER_300_2162 ();
 b15zdnd11an1n32x5 FILLER_300_2226 ();
 b15zdnd11an1n16x5 FILLER_300_2258 ();
 b15zdnd00an1n02x5 FILLER_300_2274 ();
 b15zdnd11an1n16x5 FILLER_301_0 ();
 b15zdnd11an1n08x5 FILLER_301_16 ();
 b15zdnd11an1n04x5 FILLER_301_24 ();
 b15zdnd00an1n02x5 FILLER_301_28 ();
 b15zdnd11an1n64x5 FILLER_301_34 ();
 b15zdnd11an1n64x5 FILLER_301_98 ();
 b15zdnd11an1n64x5 FILLER_301_162 ();
 b15zdnd11an1n64x5 FILLER_301_226 ();
 b15zdnd11an1n64x5 FILLER_301_290 ();
 b15zdnd11an1n64x5 FILLER_301_354 ();
 b15zdnd11an1n64x5 FILLER_301_418 ();
 b15zdnd11an1n32x5 FILLER_301_482 ();
 b15zdnd11an1n04x5 FILLER_301_514 ();
 b15zdnd00an1n02x5 FILLER_301_518 ();
 b15zdnd00an1n01x5 FILLER_301_520 ();
 b15zdnd11an1n04x5 FILLER_301_524 ();
 b15zdnd11an1n64x5 FILLER_301_531 ();
 b15zdnd11an1n32x5 FILLER_301_595 ();
 b15zdnd11an1n16x5 FILLER_301_627 ();
 b15zdnd11an1n08x5 FILLER_301_643 ();
 b15zdnd11an1n04x5 FILLER_301_651 ();
 b15zdnd00an1n01x5 FILLER_301_655 ();
 b15zdnd11an1n16x5 FILLER_301_659 ();
 b15zdnd11an1n04x5 FILLER_301_675 ();
 b15zdnd00an1n02x5 FILLER_301_679 ();
 b15zdnd11an1n64x5 FILLER_301_707 ();
 b15zdnd11an1n64x5 FILLER_301_771 ();
 b15zdnd11an1n16x5 FILLER_301_835 ();
 b15zdnd00an1n02x5 FILLER_301_851 ();
 b15zdnd11an1n64x5 FILLER_301_863 ();
 b15zdnd11an1n32x5 FILLER_301_927 ();
 b15zdnd11an1n16x5 FILLER_301_959 ();
 b15zdnd11an1n04x5 FILLER_301_975 ();
 b15zdnd00an1n02x5 FILLER_301_979 ();
 b15zdnd00an1n01x5 FILLER_301_981 ();
 b15zdnd11an1n64x5 FILLER_301_992 ();
 b15zdnd11an1n64x5 FILLER_301_1056 ();
 b15zdnd11an1n64x5 FILLER_301_1120 ();
 b15zdnd11an1n64x5 FILLER_301_1184 ();
 b15zdnd11an1n64x5 FILLER_301_1248 ();
 b15zdnd00an1n02x5 FILLER_301_1312 ();
 b15zdnd00an1n01x5 FILLER_301_1314 ();
 b15zdnd11an1n64x5 FILLER_301_1319 ();
 b15zdnd11an1n64x5 FILLER_301_1383 ();
 b15zdnd11an1n64x5 FILLER_301_1447 ();
 b15zdnd11an1n64x5 FILLER_301_1511 ();
 b15zdnd11an1n16x5 FILLER_301_1575 ();
 b15zdnd11an1n08x5 FILLER_301_1591 ();
 b15zdnd11an1n04x5 FILLER_301_1599 ();
 b15zdnd11an1n32x5 FILLER_301_1645 ();
 b15zdnd11an1n16x5 FILLER_301_1677 ();
 b15zdnd00an1n01x5 FILLER_301_1693 ();
 b15zdnd11an1n64x5 FILLER_301_1714 ();
 b15zdnd11an1n64x5 FILLER_301_1778 ();
 b15zdnd11an1n64x5 FILLER_301_1842 ();
 b15zdnd11an1n64x5 FILLER_301_1906 ();
 b15zdnd11an1n32x5 FILLER_301_1970 ();
 b15zdnd11an1n16x5 FILLER_301_2002 ();
 b15zdnd11an1n08x5 FILLER_301_2018 ();
 b15zdnd11an1n04x5 FILLER_301_2026 ();
 b15zdnd11an1n64x5 FILLER_301_2082 ();
 b15zdnd11an1n64x5 FILLER_301_2146 ();
 b15zdnd11an1n64x5 FILLER_301_2210 ();
 b15zdnd11an1n08x5 FILLER_301_2274 ();
 b15zdnd00an1n02x5 FILLER_301_2282 ();
 b15zdnd00an1n02x5 FILLER_302_8 ();
 b15zdnd00an1n01x5 FILLER_302_10 ();
 b15zdnd11an1n64x5 FILLER_302_53 ();
 b15zdnd11an1n64x5 FILLER_302_117 ();
 b15zdnd11an1n32x5 FILLER_302_181 ();
 b15zdnd11an1n04x5 FILLER_302_213 ();
 b15zdnd00an1n02x5 FILLER_302_217 ();
 b15zdnd00an1n01x5 FILLER_302_219 ();
 b15zdnd11an1n08x5 FILLER_302_240 ();
 b15zdnd11an1n64x5 FILLER_302_251 ();
 b15zdnd11an1n64x5 FILLER_302_315 ();
 b15zdnd11an1n64x5 FILLER_302_379 ();
 b15zdnd11an1n64x5 FILLER_302_443 ();
 b15zdnd11an1n64x5 FILLER_302_507 ();
 b15zdnd11an1n64x5 FILLER_302_571 ();
 b15zdnd11an1n64x5 FILLER_302_635 ();
 b15zdnd11an1n16x5 FILLER_302_699 ();
 b15zdnd00an1n02x5 FILLER_302_715 ();
 b15zdnd00an1n01x5 FILLER_302_717 ();
 b15zdnd11an1n32x5 FILLER_302_726 ();
 b15zdnd11an1n16x5 FILLER_302_758 ();
 b15zdnd11an1n04x5 FILLER_302_774 ();
 b15zdnd11an1n64x5 FILLER_302_782 ();
 b15zdnd11an1n08x5 FILLER_302_846 ();
 b15zdnd11an1n64x5 FILLER_302_859 ();
 b15zdnd11an1n64x5 FILLER_302_923 ();
 b15zdnd11an1n64x5 FILLER_302_987 ();
 b15zdnd11an1n64x5 FILLER_302_1051 ();
 b15zdnd11an1n04x5 FILLER_302_1115 ();
 b15zdnd00an1n02x5 FILLER_302_1119 ();
 b15zdnd00an1n01x5 FILLER_302_1121 ();
 b15zdnd11an1n64x5 FILLER_302_1138 ();
 b15zdnd11an1n64x5 FILLER_302_1202 ();
 b15zdnd11an1n64x5 FILLER_302_1266 ();
 b15zdnd11an1n64x5 FILLER_302_1330 ();
 b15zdnd11an1n64x5 FILLER_302_1394 ();
 b15zdnd11an1n16x5 FILLER_302_1458 ();
 b15zdnd11an1n08x5 FILLER_302_1474 ();
 b15zdnd11an1n04x5 FILLER_302_1482 ();
 b15zdnd00an1n02x5 FILLER_302_1486 ();
 b15zdnd11an1n64x5 FILLER_302_1497 ();
 b15zdnd11an1n32x5 FILLER_302_1561 ();
 b15zdnd11an1n16x5 FILLER_302_1593 ();
 b15zdnd11an1n04x5 FILLER_302_1609 ();
 b15zdnd00an1n01x5 FILLER_302_1613 ();
 b15zdnd11an1n64x5 FILLER_302_1656 ();
 b15zdnd11an1n32x5 FILLER_302_1720 ();
 b15zdnd11an1n16x5 FILLER_302_1752 ();
 b15zdnd11an1n08x5 FILLER_302_1768 ();
 b15zdnd11an1n04x5 FILLER_302_1779 ();
 b15zdnd11an1n08x5 FILLER_302_1786 ();
 b15zdnd00an1n02x5 FILLER_302_1794 ();
 b15zdnd00an1n01x5 FILLER_302_1796 ();
 b15zdnd11an1n32x5 FILLER_302_1822 ();
 b15zdnd11an1n16x5 FILLER_302_1854 ();
 b15zdnd00an1n02x5 FILLER_302_1870 ();
 b15zdnd00an1n01x5 FILLER_302_1872 ();
 b15zdnd11an1n64x5 FILLER_302_1880 ();
 b15zdnd11an1n64x5 FILLER_302_1944 ();
 b15zdnd11an1n16x5 FILLER_302_2008 ();
 b15zdnd11an1n08x5 FILLER_302_2024 ();
 b15zdnd00an1n01x5 FILLER_302_2032 ();
 b15zdnd11an1n64x5 FILLER_302_2075 ();
 b15zdnd11an1n08x5 FILLER_302_2139 ();
 b15zdnd11an1n04x5 FILLER_302_2147 ();
 b15zdnd00an1n02x5 FILLER_302_2151 ();
 b15zdnd00an1n01x5 FILLER_302_2153 ();
 b15zdnd11an1n64x5 FILLER_302_2162 ();
 b15zdnd11an1n32x5 FILLER_302_2226 ();
 b15zdnd11an1n16x5 FILLER_302_2258 ();
 b15zdnd00an1n02x5 FILLER_302_2274 ();
 b15zdnd11an1n16x5 FILLER_303_0 ();
 b15zdnd11an1n08x5 FILLER_303_16 ();
 b15zdnd11an1n04x5 FILLER_303_24 ();
 b15zdnd00an1n01x5 FILLER_303_28 ();
 b15zdnd11an1n64x5 FILLER_303_33 ();
 b15zdnd11an1n64x5 FILLER_303_97 ();
 b15zdnd11an1n64x5 FILLER_303_161 ();
 b15zdnd00an1n01x5 FILLER_303_225 ();
 b15zdnd11an1n04x5 FILLER_303_258 ();
 b15zdnd11an1n64x5 FILLER_303_265 ();
 b15zdnd11an1n64x5 FILLER_303_329 ();
 b15zdnd11an1n64x5 FILLER_303_393 ();
 b15zdnd11an1n64x5 FILLER_303_457 ();
 b15zdnd11an1n64x5 FILLER_303_521 ();
 b15zdnd11an1n64x5 FILLER_303_585 ();
 b15zdnd11an1n64x5 FILLER_303_649 ();
 b15zdnd11an1n16x5 FILLER_303_713 ();
 b15zdnd11an1n08x5 FILLER_303_729 ();
 b15zdnd00an1n02x5 FILLER_303_737 ();
 b15zdnd00an1n01x5 FILLER_303_739 ();
 b15zdnd11an1n64x5 FILLER_303_780 ();
 b15zdnd11an1n64x5 FILLER_303_844 ();
 b15zdnd11an1n64x5 FILLER_303_908 ();
 b15zdnd11an1n64x5 FILLER_303_972 ();
 b15zdnd11an1n64x5 FILLER_303_1036 ();
 b15zdnd11an1n64x5 FILLER_303_1100 ();
 b15zdnd11an1n64x5 FILLER_303_1164 ();
 b15zdnd11an1n64x5 FILLER_303_1228 ();
 b15zdnd11an1n08x5 FILLER_303_1292 ();
 b15zdnd11an1n04x5 FILLER_303_1300 ();
 b15zdnd00an1n01x5 FILLER_303_1304 ();
 b15zdnd11an1n64x5 FILLER_303_1347 ();
 b15zdnd11an1n32x5 FILLER_303_1411 ();
 b15zdnd11an1n04x5 FILLER_303_1443 ();
 b15zdnd00an1n01x5 FILLER_303_1447 ();
 b15zdnd11an1n64x5 FILLER_303_1452 ();
 b15zdnd11an1n64x5 FILLER_303_1516 ();
 b15zdnd11an1n16x5 FILLER_303_1580 ();
 b15zdnd00an1n02x5 FILLER_303_1596 ();
 b15zdnd11an1n64x5 FILLER_303_1640 ();
 b15zdnd11an1n32x5 FILLER_303_1704 ();
 b15zdnd11an1n16x5 FILLER_303_1736 ();
 b15zdnd11an1n04x5 FILLER_303_1752 ();
 b15zdnd00an1n02x5 FILLER_303_1756 ();
 b15zdnd11an1n04x5 FILLER_303_1810 ();
 b15zdnd11an1n64x5 FILLER_303_1856 ();
 b15zdnd11an1n64x5 FILLER_303_1920 ();
 b15zdnd11an1n64x5 FILLER_303_1984 ();
 b15zdnd11an1n04x5 FILLER_303_2051 ();
 b15zdnd11an1n64x5 FILLER_303_2058 ();
 b15zdnd11an1n64x5 FILLER_303_2122 ();
 b15zdnd11an1n64x5 FILLER_303_2186 ();
 b15zdnd11an1n32x5 FILLER_303_2250 ();
 b15zdnd00an1n02x5 FILLER_303_2282 ();
 b15zdnd00an1n02x5 FILLER_304_8 ();
 b15zdnd11an1n64x5 FILLER_304_52 ();
 b15zdnd11an1n16x5 FILLER_304_116 ();
 b15zdnd11an1n04x5 FILLER_304_132 ();
 b15zdnd00an1n02x5 FILLER_304_136 ();
 b15zdnd00an1n01x5 FILLER_304_138 ();
 b15zdnd11an1n16x5 FILLER_304_181 ();
 b15zdnd11an1n08x5 FILLER_304_197 ();
 b15zdnd11an1n04x5 FILLER_304_205 ();
 b15zdnd00an1n02x5 FILLER_304_209 ();
 b15zdnd00an1n01x5 FILLER_304_211 ();
 b15zdnd11an1n64x5 FILLER_304_254 ();
 b15zdnd11an1n04x5 FILLER_304_318 ();
 b15zdnd00an1n01x5 FILLER_304_322 ();
 b15zdnd11an1n64x5 FILLER_304_326 ();
 b15zdnd11an1n16x5 FILLER_304_390 ();
 b15zdnd11an1n08x5 FILLER_304_406 ();
 b15zdnd00an1n02x5 FILLER_304_414 ();
 b15zdnd00an1n01x5 FILLER_304_416 ();
 b15zdnd11an1n64x5 FILLER_304_420 ();
 b15zdnd11an1n64x5 FILLER_304_484 ();
 b15zdnd11an1n64x5 FILLER_304_548 ();
 b15zdnd11an1n64x5 FILLER_304_612 ();
 b15zdnd11an1n32x5 FILLER_304_676 ();
 b15zdnd11an1n08x5 FILLER_304_708 ();
 b15zdnd00an1n02x5 FILLER_304_716 ();
 b15zdnd11an1n32x5 FILLER_304_726 ();
 b15zdnd11an1n08x5 FILLER_304_758 ();
 b15zdnd00an1n02x5 FILLER_304_766 ();
 b15zdnd00an1n01x5 FILLER_304_768 ();
 b15zdnd11an1n04x5 FILLER_304_772 ();
 b15zdnd11an1n64x5 FILLER_304_779 ();
 b15zdnd11an1n08x5 FILLER_304_843 ();
 b15zdnd00an1n01x5 FILLER_304_851 ();
 b15zdnd11an1n64x5 FILLER_304_862 ();
 b15zdnd11an1n64x5 FILLER_304_926 ();
 b15zdnd11an1n16x5 FILLER_304_990 ();
 b15zdnd11an1n04x5 FILLER_304_1006 ();
 b15zdnd00an1n02x5 FILLER_304_1010 ();
 b15zdnd00an1n01x5 FILLER_304_1012 ();
 b15zdnd11an1n64x5 FILLER_304_1020 ();
 b15zdnd11an1n32x5 FILLER_304_1084 ();
 b15zdnd11an1n16x5 FILLER_304_1116 ();
 b15zdnd11an1n08x5 FILLER_304_1132 ();
 b15zdnd11an1n04x5 FILLER_304_1140 ();
 b15zdnd11an1n64x5 FILLER_304_1158 ();
 b15zdnd11an1n64x5 FILLER_304_1222 ();
 b15zdnd11an1n16x5 FILLER_304_1286 ();
 b15zdnd00an1n01x5 FILLER_304_1302 ();
 b15zdnd11an1n04x5 FILLER_304_1318 ();
 b15zdnd11an1n64x5 FILLER_304_1325 ();
 b15zdnd11an1n64x5 FILLER_304_1389 ();
 b15zdnd11an1n64x5 FILLER_304_1453 ();
 b15zdnd11an1n64x5 FILLER_304_1517 ();
 b15zdnd11an1n16x5 FILLER_304_1581 ();
 b15zdnd00an1n02x5 FILLER_304_1597 ();
 b15zdnd00an1n01x5 FILLER_304_1599 ();
 b15zdnd11an1n08x5 FILLER_304_1610 ();
 b15zdnd00an1n01x5 FILLER_304_1618 ();
 b15zdnd11an1n64x5 FILLER_304_1626 ();
 b15zdnd11an1n64x5 FILLER_304_1690 ();
 b15zdnd11an1n16x5 FILLER_304_1754 ();
 b15zdnd11an1n08x5 FILLER_304_1770 ();
 b15zdnd11an1n04x5 FILLER_304_1778 ();
 b15zdnd00an1n01x5 FILLER_304_1782 ();
 b15zdnd11an1n32x5 FILLER_304_1786 ();
 b15zdnd00an1n02x5 FILLER_304_1818 ();
 b15zdnd11an1n16x5 FILLER_304_1862 ();
 b15zdnd00an1n01x5 FILLER_304_1878 ();
 b15zdnd11an1n08x5 FILLER_304_1882 ();
 b15zdnd11an1n04x5 FILLER_304_1890 ();
 b15zdnd00an1n02x5 FILLER_304_1894 ();
 b15zdnd00an1n01x5 FILLER_304_1896 ();
 b15zdnd11an1n64x5 FILLER_304_1907 ();
 b15zdnd11an1n32x5 FILLER_304_1971 ();
 b15zdnd11an1n04x5 FILLER_304_2003 ();
 b15zdnd00an1n02x5 FILLER_304_2007 ();
 b15zdnd11an1n64x5 FILLER_304_2013 ();
 b15zdnd11an1n64x5 FILLER_304_2077 ();
 b15zdnd11an1n08x5 FILLER_304_2141 ();
 b15zdnd11an1n04x5 FILLER_304_2149 ();
 b15zdnd00an1n01x5 FILLER_304_2153 ();
 b15zdnd11an1n64x5 FILLER_304_2162 ();
 b15zdnd11an1n32x5 FILLER_304_2226 ();
 b15zdnd11an1n16x5 FILLER_304_2258 ();
 b15zdnd00an1n02x5 FILLER_304_2274 ();
 b15zdnd11an1n16x5 FILLER_305_0 ();
 b15zdnd00an1n01x5 FILLER_305_16 ();
 b15zdnd11an1n64x5 FILLER_305_22 ();
 b15zdnd11an1n16x5 FILLER_305_86 ();
 b15zdnd11an1n08x5 FILLER_305_102 ();
 b15zdnd11an1n04x5 FILLER_305_110 ();
 b15zdnd11an1n64x5 FILLER_305_156 ();
 b15zdnd11an1n08x5 FILLER_305_220 ();
 b15zdnd00an1n02x5 FILLER_305_228 ();
 b15zdnd00an1n01x5 FILLER_305_230 ();
 b15zdnd11an1n16x5 FILLER_305_273 ();
 b15zdnd11an1n08x5 FILLER_305_289 ();
 b15zdnd11an1n04x5 FILLER_305_297 ();
 b15zdnd00an1n02x5 FILLER_305_301 ();
 b15zdnd11an1n32x5 FILLER_305_345 ();
 b15zdnd11an1n08x5 FILLER_305_377 ();
 b15zdnd11an1n04x5 FILLER_305_385 ();
 b15zdnd00an1n01x5 FILLER_305_389 ();
 b15zdnd11an1n64x5 FILLER_305_442 ();
 b15zdnd11an1n64x5 FILLER_305_506 ();
 b15zdnd11an1n64x5 FILLER_305_570 ();
 b15zdnd11an1n64x5 FILLER_305_634 ();
 b15zdnd11an1n64x5 FILLER_305_698 ();
 b15zdnd11an1n64x5 FILLER_305_762 ();
 b15zdnd11an1n32x5 FILLER_305_826 ();
 b15zdnd00an1n01x5 FILLER_305_858 ();
 b15zdnd11an1n64x5 FILLER_305_901 ();
 b15zdnd11an1n16x5 FILLER_305_965 ();
 b15zdnd11an1n04x5 FILLER_305_981 ();
 b15zdnd11an1n32x5 FILLER_305_1037 ();
 b15zdnd11an1n08x5 FILLER_305_1069 ();
 b15zdnd11an1n04x5 FILLER_305_1122 ();
 b15zdnd11an1n04x5 FILLER_305_1146 ();
 b15zdnd00an1n02x5 FILLER_305_1150 ();
 b15zdnd11an1n64x5 FILLER_305_1159 ();
 b15zdnd11an1n32x5 FILLER_305_1223 ();
 b15zdnd00an1n01x5 FILLER_305_1255 ();
 b15zdnd11an1n16x5 FILLER_305_1276 ();
 b15zdnd00an1n02x5 FILLER_305_1292 ();
 b15zdnd11an1n64x5 FILLER_305_1336 ();
 b15zdnd11an1n64x5 FILLER_305_1400 ();
 b15zdnd11an1n64x5 FILLER_305_1464 ();
 b15zdnd11an1n64x5 FILLER_305_1528 ();
 b15zdnd11an1n16x5 FILLER_305_1592 ();
 b15zdnd11an1n04x5 FILLER_305_1614 ();
 b15zdnd00an1n01x5 FILLER_305_1618 ();
 b15zdnd11an1n04x5 FILLER_305_1623 ();
 b15zdnd00an1n01x5 FILLER_305_1627 ();
 b15zdnd11an1n04x5 FILLER_305_1631 ();
 b15zdnd00an1n01x5 FILLER_305_1635 ();
 b15zdnd11an1n64x5 FILLER_305_1641 ();
 b15zdnd11an1n64x5 FILLER_305_1705 ();
 b15zdnd11an1n64x5 FILLER_305_1769 ();
 b15zdnd11an1n16x5 FILLER_305_1833 ();
 b15zdnd11an1n08x5 FILLER_305_1849 ();
 b15zdnd00an1n02x5 FILLER_305_1857 ();
 b15zdnd11an1n08x5 FILLER_305_1864 ();
 b15zdnd00an1n02x5 FILLER_305_1872 ();
 b15zdnd00an1n01x5 FILLER_305_1874 ();
 b15zdnd11an1n08x5 FILLER_305_1879 ();
 b15zdnd00an1n01x5 FILLER_305_1887 ();
 b15zdnd11an1n04x5 FILLER_305_1902 ();
 b15zdnd11an1n04x5 FILLER_305_1909 ();
 b15zdnd11an1n64x5 FILLER_305_1916 ();
 b15zdnd11an1n64x5 FILLER_305_1980 ();
 b15zdnd11an1n64x5 FILLER_305_2044 ();
 b15zdnd11an1n64x5 FILLER_305_2108 ();
 b15zdnd11an1n64x5 FILLER_305_2172 ();
 b15zdnd11an1n32x5 FILLER_305_2236 ();
 b15zdnd11an1n16x5 FILLER_305_2268 ();
 b15zdnd11an1n64x5 FILLER_306_8 ();
 b15zdnd11an1n64x5 FILLER_306_72 ();
 b15zdnd11an1n16x5 FILLER_306_136 ();
 b15zdnd11an1n08x5 FILLER_306_152 ();
 b15zdnd11an1n04x5 FILLER_306_160 ();
 b15zdnd11an1n16x5 FILLER_306_206 ();
 b15zdnd11an1n08x5 FILLER_306_222 ();
 b15zdnd11an1n16x5 FILLER_306_272 ();
 b15zdnd11an1n04x5 FILLER_306_288 ();
 b15zdnd00an1n02x5 FILLER_306_292 ();
 b15zdnd00an1n01x5 FILLER_306_294 ();
 b15zdnd11an1n64x5 FILLER_306_327 ();
 b15zdnd11an1n16x5 FILLER_306_391 ();
 b15zdnd00an1n01x5 FILLER_306_407 ();
 b15zdnd11an1n04x5 FILLER_306_411 ();
 b15zdnd11an1n64x5 FILLER_306_418 ();
 b15zdnd11an1n64x5 FILLER_306_482 ();
 b15zdnd11an1n64x5 FILLER_306_546 ();
 b15zdnd11an1n64x5 FILLER_306_610 ();
 b15zdnd11an1n32x5 FILLER_306_674 ();
 b15zdnd11an1n08x5 FILLER_306_706 ();
 b15zdnd11an1n04x5 FILLER_306_714 ();
 b15zdnd11an1n64x5 FILLER_306_726 ();
 b15zdnd11an1n32x5 FILLER_306_790 ();
 b15zdnd11an1n16x5 FILLER_306_822 ();
 b15zdnd11an1n08x5 FILLER_306_838 ();
 b15zdnd11an1n04x5 FILLER_306_846 ();
 b15zdnd00an1n02x5 FILLER_306_850 ();
 b15zdnd11an1n64x5 FILLER_306_855 ();
 b15zdnd11an1n64x5 FILLER_306_919 ();
 b15zdnd11an1n16x5 FILLER_306_983 ();
 b15zdnd11an1n04x5 FILLER_306_999 ();
 b15zdnd00an1n02x5 FILLER_306_1003 ();
 b15zdnd11an1n04x5 FILLER_306_1008 ();
 b15zdnd11an1n64x5 FILLER_306_1015 ();
 b15zdnd11an1n64x5 FILLER_306_1079 ();
 b15zdnd11an1n64x5 FILLER_306_1143 ();
 b15zdnd11an1n64x5 FILLER_306_1207 ();
 b15zdnd11an1n32x5 FILLER_306_1271 ();
 b15zdnd11an1n04x5 FILLER_306_1303 ();
 b15zdnd11an1n04x5 FILLER_306_1313 ();
 b15zdnd00an1n02x5 FILLER_306_1317 ();
 b15zdnd00an1n01x5 FILLER_306_1319 ();
 b15zdnd11an1n64x5 FILLER_306_1362 ();
 b15zdnd11an1n64x5 FILLER_306_1426 ();
 b15zdnd11an1n64x5 FILLER_306_1490 ();
 b15zdnd11an1n32x5 FILLER_306_1554 ();
 b15zdnd11an1n16x5 FILLER_306_1586 ();
 b15zdnd11an1n04x5 FILLER_306_1602 ();
 b15zdnd00an1n02x5 FILLER_306_1606 ();
 b15zdnd11an1n64x5 FILLER_306_1614 ();
 b15zdnd11an1n64x5 FILLER_306_1678 ();
 b15zdnd11an1n64x5 FILLER_306_1742 ();
 b15zdnd11an1n32x5 FILLER_306_1806 ();
 b15zdnd11an1n16x5 FILLER_306_1838 ();
 b15zdnd11an1n04x5 FILLER_306_1854 ();
 b15zdnd00an1n01x5 FILLER_306_1858 ();
 b15zdnd11an1n64x5 FILLER_306_1911 ();
 b15zdnd11an1n64x5 FILLER_306_1975 ();
 b15zdnd11an1n64x5 FILLER_306_2039 ();
 b15zdnd11an1n32x5 FILLER_306_2103 ();
 b15zdnd11an1n16x5 FILLER_306_2135 ();
 b15zdnd00an1n02x5 FILLER_306_2151 ();
 b15zdnd00an1n01x5 FILLER_306_2153 ();
 b15zdnd11an1n64x5 FILLER_306_2162 ();
 b15zdnd11an1n32x5 FILLER_306_2226 ();
 b15zdnd11an1n16x5 FILLER_306_2258 ();
 b15zdnd00an1n02x5 FILLER_306_2274 ();
 b15zdnd11an1n64x5 FILLER_307_0 ();
 b15zdnd11an1n64x5 FILLER_307_64 ();
 b15zdnd11an1n64x5 FILLER_307_128 ();
 b15zdnd11an1n08x5 FILLER_307_192 ();
 b15zdnd11an1n04x5 FILLER_307_200 ();
 b15zdnd00an1n02x5 FILLER_307_204 ();
 b15zdnd00an1n01x5 FILLER_307_206 ();
 b15zdnd11an1n04x5 FILLER_307_239 ();
 b15zdnd11an1n64x5 FILLER_307_246 ();
 b15zdnd11an1n08x5 FILLER_307_310 ();
 b15zdnd11an1n04x5 FILLER_307_318 ();
 b15zdnd00an1n02x5 FILLER_307_322 ();
 b15zdnd11an1n64x5 FILLER_307_327 ();
 b15zdnd11an1n64x5 FILLER_307_391 ();
 b15zdnd11an1n64x5 FILLER_307_455 ();
 b15zdnd11an1n64x5 FILLER_307_519 ();
 b15zdnd11an1n64x5 FILLER_307_583 ();
 b15zdnd11an1n64x5 FILLER_307_647 ();
 b15zdnd11an1n64x5 FILLER_307_711 ();
 b15zdnd11an1n64x5 FILLER_307_775 ();
 b15zdnd11an1n08x5 FILLER_307_839 ();
 b15zdnd11an1n64x5 FILLER_307_860 ();
 b15zdnd11an1n64x5 FILLER_307_924 ();
 b15zdnd11an1n16x5 FILLER_307_988 ();
 b15zdnd11an1n04x5 FILLER_307_1004 ();
 b15zdnd00an1n02x5 FILLER_307_1008 ();
 b15zdnd11an1n64x5 FILLER_307_1013 ();
 b15zdnd11an1n64x5 FILLER_307_1077 ();
 b15zdnd11an1n64x5 FILLER_307_1141 ();
 b15zdnd11an1n64x5 FILLER_307_1205 ();
 b15zdnd11an1n32x5 FILLER_307_1269 ();
 b15zdnd00an1n02x5 FILLER_307_1301 ();
 b15zdnd00an1n01x5 FILLER_307_1303 ();
 b15zdnd11an1n64x5 FILLER_307_1346 ();
 b15zdnd11an1n64x5 FILLER_307_1410 ();
 b15zdnd11an1n64x5 FILLER_307_1474 ();
 b15zdnd11an1n64x5 FILLER_307_1538 ();
 b15zdnd11an1n04x5 FILLER_307_1605 ();
 b15zdnd11an1n64x5 FILLER_307_1619 ();
 b15zdnd11an1n64x5 FILLER_307_1683 ();
 b15zdnd11an1n64x5 FILLER_307_1747 ();
 b15zdnd11an1n32x5 FILLER_307_1811 ();
 b15zdnd11an1n16x5 FILLER_307_1843 ();
 b15zdnd11an1n16x5 FILLER_307_1862 ();
 b15zdnd00an1n01x5 FILLER_307_1878 ();
 b15zdnd11an1n08x5 FILLER_307_1885 ();
 b15zdnd00an1n01x5 FILLER_307_1893 ();
 b15zdnd11an1n04x5 FILLER_307_1904 ();
 b15zdnd11an1n64x5 FILLER_307_1913 ();
 b15zdnd11an1n64x5 FILLER_307_1977 ();
 b15zdnd11an1n64x5 FILLER_307_2041 ();
 b15zdnd11an1n64x5 FILLER_307_2105 ();
 b15zdnd11an1n64x5 FILLER_307_2169 ();
 b15zdnd11an1n32x5 FILLER_307_2233 ();
 b15zdnd11an1n16x5 FILLER_307_2265 ();
 b15zdnd00an1n02x5 FILLER_307_2281 ();
 b15zdnd00an1n01x5 FILLER_307_2283 ();
 b15zdnd11an1n64x5 FILLER_308_8 ();
 b15zdnd11an1n64x5 FILLER_308_72 ();
 b15zdnd11an1n32x5 FILLER_308_136 ();
 b15zdnd11an1n16x5 FILLER_308_168 ();
 b15zdnd00an1n02x5 FILLER_308_184 ();
 b15zdnd11an1n32x5 FILLER_308_189 ();
 b15zdnd11an1n08x5 FILLER_308_221 ();
 b15zdnd00an1n02x5 FILLER_308_229 ();
 b15zdnd11an1n64x5 FILLER_308_234 ();
 b15zdnd11an1n64x5 FILLER_308_298 ();
 b15zdnd11an1n64x5 FILLER_308_362 ();
 b15zdnd11an1n64x5 FILLER_308_426 ();
 b15zdnd11an1n64x5 FILLER_308_490 ();
 b15zdnd11an1n64x5 FILLER_308_554 ();
 b15zdnd11an1n64x5 FILLER_308_618 ();
 b15zdnd11an1n32x5 FILLER_308_682 ();
 b15zdnd11an1n04x5 FILLER_308_714 ();
 b15zdnd11an1n64x5 FILLER_308_726 ();
 b15zdnd11an1n32x5 FILLER_308_790 ();
 b15zdnd11an1n16x5 FILLER_308_822 ();
 b15zdnd11an1n04x5 FILLER_308_838 ();
 b15zdnd11an1n04x5 FILLER_308_847 ();
 b15zdnd11an1n04x5 FILLER_308_863 ();
 b15zdnd11an1n64x5 FILLER_308_871 ();
 b15zdnd11an1n64x5 FILLER_308_935 ();
 b15zdnd11an1n64x5 FILLER_308_999 ();
 b15zdnd11an1n32x5 FILLER_308_1063 ();
 b15zdnd11an1n16x5 FILLER_308_1095 ();
 b15zdnd00an1n01x5 FILLER_308_1111 ();
 b15zdnd11an1n64x5 FILLER_308_1115 ();
 b15zdnd11an1n64x5 FILLER_308_1179 ();
 b15zdnd11an1n32x5 FILLER_308_1243 ();
 b15zdnd11an1n08x5 FILLER_308_1275 ();
 b15zdnd00an1n02x5 FILLER_308_1283 ();
 b15zdnd11an1n16x5 FILLER_308_1288 ();
 b15zdnd11an1n04x5 FILLER_308_1307 ();
 b15zdnd11an1n64x5 FILLER_308_1353 ();
 b15zdnd11an1n32x5 FILLER_308_1417 ();
 b15zdnd11an1n08x5 FILLER_308_1449 ();
 b15zdnd11an1n64x5 FILLER_308_1465 ();
 b15zdnd11an1n64x5 FILLER_308_1529 ();
 b15zdnd11an1n08x5 FILLER_308_1593 ();
 b15zdnd11an1n04x5 FILLER_308_1601 ();
 b15zdnd00an1n02x5 FILLER_308_1605 ();
 b15zdnd00an1n01x5 FILLER_308_1607 ();
 b15zdnd11an1n64x5 FILLER_308_1617 ();
 b15zdnd11an1n64x5 FILLER_308_1681 ();
 b15zdnd11an1n64x5 FILLER_308_1745 ();
 b15zdnd11an1n64x5 FILLER_308_1809 ();
 b15zdnd11an1n08x5 FILLER_308_1873 ();
 b15zdnd00an1n02x5 FILLER_308_1881 ();
 b15zdnd00an1n01x5 FILLER_308_1883 ();
 b15zdnd11an1n04x5 FILLER_308_1887 ();
 b15zdnd00an1n02x5 FILLER_308_1891 ();
 b15zdnd00an1n01x5 FILLER_308_1893 ();
 b15zdnd11an1n64x5 FILLER_308_1904 ();
 b15zdnd11an1n64x5 FILLER_308_1968 ();
 b15zdnd11an1n64x5 FILLER_308_2032 ();
 b15zdnd11an1n32x5 FILLER_308_2096 ();
 b15zdnd11an1n16x5 FILLER_308_2128 ();
 b15zdnd11an1n08x5 FILLER_308_2144 ();
 b15zdnd00an1n02x5 FILLER_308_2152 ();
 b15zdnd11an1n64x5 FILLER_308_2162 ();
 b15zdnd11an1n32x5 FILLER_308_2226 ();
 b15zdnd11an1n16x5 FILLER_308_2258 ();
 b15zdnd00an1n02x5 FILLER_308_2274 ();
 b15zdnd11an1n64x5 FILLER_309_0 ();
 b15zdnd11an1n64x5 FILLER_309_64 ();
 b15zdnd11an1n16x5 FILLER_309_128 ();
 b15zdnd11an1n08x5 FILLER_309_144 ();
 b15zdnd11an1n04x5 FILLER_309_152 ();
 b15zdnd00an1n02x5 FILLER_309_156 ();
 b15zdnd00an1n01x5 FILLER_309_158 ();
 b15zdnd11an1n64x5 FILLER_309_211 ();
 b15zdnd11an1n64x5 FILLER_309_275 ();
 b15zdnd11an1n64x5 FILLER_309_339 ();
 b15zdnd11an1n64x5 FILLER_309_403 ();
 b15zdnd11an1n64x5 FILLER_309_467 ();
 b15zdnd11an1n64x5 FILLER_309_531 ();
 b15zdnd11an1n64x5 FILLER_309_595 ();
 b15zdnd11an1n64x5 FILLER_309_659 ();
 b15zdnd11an1n64x5 FILLER_309_723 ();
 b15zdnd11an1n32x5 FILLER_309_787 ();
 b15zdnd11an1n16x5 FILLER_309_819 ();
 b15zdnd00an1n02x5 FILLER_309_835 ();
 b15zdnd11an1n64x5 FILLER_309_879 ();
 b15zdnd11an1n64x5 FILLER_309_943 ();
 b15zdnd11an1n32x5 FILLER_309_1007 ();
 b15zdnd11an1n16x5 FILLER_309_1039 ();
 b15zdnd11an1n04x5 FILLER_309_1055 ();
 b15zdnd00an1n02x5 FILLER_309_1059 ();
 b15zdnd11an1n16x5 FILLER_309_1069 ();
 b15zdnd11an1n64x5 FILLER_309_1137 ();
 b15zdnd11an1n64x5 FILLER_309_1201 ();
 b15zdnd11an1n16x5 FILLER_309_1265 ();
 b15zdnd11an1n64x5 FILLER_309_1333 ();
 b15zdnd11an1n64x5 FILLER_309_1397 ();
 b15zdnd11an1n64x5 FILLER_309_1461 ();
 b15zdnd11an1n64x5 FILLER_309_1525 ();
 b15zdnd11an1n08x5 FILLER_309_1589 ();
 b15zdnd11an1n04x5 FILLER_309_1597 ();
 b15zdnd11an1n64x5 FILLER_309_1614 ();
 b15zdnd11an1n64x5 FILLER_309_1678 ();
 b15zdnd11an1n64x5 FILLER_309_1742 ();
 b15zdnd11an1n64x5 FILLER_309_1806 ();
 b15zdnd11an1n16x5 FILLER_309_1870 ();
 b15zdnd11an1n04x5 FILLER_309_1886 ();
 b15zdnd00an1n01x5 FILLER_309_1890 ();
 b15zdnd11an1n64x5 FILLER_309_1901 ();
 b15zdnd11an1n64x5 FILLER_309_1965 ();
 b15zdnd11an1n64x5 FILLER_309_2029 ();
 b15zdnd11an1n64x5 FILLER_309_2093 ();
 b15zdnd11an1n64x5 FILLER_309_2157 ();
 b15zdnd11an1n32x5 FILLER_309_2221 ();
 b15zdnd11an1n16x5 FILLER_309_2253 ();
 b15zdnd11an1n08x5 FILLER_309_2269 ();
 b15zdnd11an1n04x5 FILLER_309_2277 ();
 b15zdnd00an1n02x5 FILLER_309_2281 ();
 b15zdnd00an1n01x5 FILLER_309_2283 ();
 b15zdnd11an1n64x5 FILLER_310_8 ();
 b15zdnd11an1n64x5 FILLER_310_72 ();
 b15zdnd11an1n32x5 FILLER_310_136 ();
 b15zdnd11an1n16x5 FILLER_310_168 ();
 b15zdnd11an1n64x5 FILLER_310_187 ();
 b15zdnd11an1n64x5 FILLER_310_251 ();
 b15zdnd11an1n64x5 FILLER_310_315 ();
 b15zdnd11an1n64x5 FILLER_310_379 ();
 b15zdnd11an1n64x5 FILLER_310_443 ();
 b15zdnd11an1n64x5 FILLER_310_507 ();
 b15zdnd11an1n64x5 FILLER_310_571 ();
 b15zdnd11an1n64x5 FILLER_310_635 ();
 b15zdnd11an1n16x5 FILLER_310_699 ();
 b15zdnd00an1n02x5 FILLER_310_715 ();
 b15zdnd00an1n01x5 FILLER_310_717 ();
 b15zdnd11an1n64x5 FILLER_310_726 ();
 b15zdnd11an1n32x5 FILLER_310_790 ();
 b15zdnd11an1n16x5 FILLER_310_822 ();
 b15zdnd11an1n04x5 FILLER_310_838 ();
 b15zdnd11an1n04x5 FILLER_310_845 ();
 b15zdnd11an1n64x5 FILLER_310_891 ();
 b15zdnd11an1n64x5 FILLER_310_955 ();
 b15zdnd11an1n64x5 FILLER_310_1019 ();
 b15zdnd11an1n16x5 FILLER_310_1083 ();
 b15zdnd11an1n04x5 FILLER_310_1099 ();
 b15zdnd11an1n04x5 FILLER_310_1106 ();
 b15zdnd11an1n32x5 FILLER_310_1113 ();
 b15zdnd00an1n02x5 FILLER_310_1145 ();
 b15zdnd00an1n01x5 FILLER_310_1147 ();
 b15zdnd11an1n64x5 FILLER_310_1155 ();
 b15zdnd11an1n64x5 FILLER_310_1219 ();
 b15zdnd11an1n64x5 FILLER_310_1283 ();
 b15zdnd11an1n64x5 FILLER_310_1347 ();
 b15zdnd11an1n64x5 FILLER_310_1411 ();
 b15zdnd11an1n64x5 FILLER_310_1475 ();
 b15zdnd11an1n32x5 FILLER_310_1539 ();
 b15zdnd11an1n16x5 FILLER_310_1571 ();
 b15zdnd11an1n08x5 FILLER_310_1587 ();
 b15zdnd11an1n04x5 FILLER_310_1595 ();
 b15zdnd00an1n02x5 FILLER_310_1599 ();
 b15zdnd00an1n01x5 FILLER_310_1601 ();
 b15zdnd11an1n64x5 FILLER_310_1607 ();
 b15zdnd11an1n64x5 FILLER_310_1671 ();
 b15zdnd11an1n64x5 FILLER_310_1735 ();
 b15zdnd11an1n64x5 FILLER_310_1799 ();
 b15zdnd11an1n64x5 FILLER_310_1863 ();
 b15zdnd11an1n64x5 FILLER_310_1927 ();
 b15zdnd11an1n64x5 FILLER_310_1991 ();
 b15zdnd11an1n64x5 FILLER_310_2055 ();
 b15zdnd11an1n32x5 FILLER_310_2119 ();
 b15zdnd00an1n02x5 FILLER_310_2151 ();
 b15zdnd00an1n01x5 FILLER_310_2153 ();
 b15zdnd11an1n64x5 FILLER_310_2162 ();
 b15zdnd11an1n32x5 FILLER_310_2226 ();
 b15zdnd11an1n16x5 FILLER_310_2258 ();
 b15zdnd00an1n02x5 FILLER_310_2274 ();
 b15zdnd11an1n64x5 FILLER_311_0 ();
 b15zdnd11an1n64x5 FILLER_311_64 ();
 b15zdnd11an1n32x5 FILLER_311_128 ();
 b15zdnd11an1n16x5 FILLER_311_160 ();
 b15zdnd11an1n04x5 FILLER_311_176 ();
 b15zdnd00an1n02x5 FILLER_311_180 ();
 b15zdnd00an1n01x5 FILLER_311_182 ();
 b15zdnd11an1n64x5 FILLER_311_186 ();
 b15zdnd11an1n64x5 FILLER_311_250 ();
 b15zdnd11an1n32x5 FILLER_311_314 ();
 b15zdnd11an1n16x5 FILLER_311_346 ();
 b15zdnd11an1n08x5 FILLER_311_362 ();
 b15zdnd00an1n02x5 FILLER_311_370 ();
 b15zdnd00an1n01x5 FILLER_311_372 ();
 b15zdnd11an1n16x5 FILLER_311_379 ();
 b15zdnd11an1n08x5 FILLER_311_395 ();
 b15zdnd11an1n04x5 FILLER_311_403 ();
 b15zdnd11an1n64x5 FILLER_311_411 ();
 b15zdnd11an1n64x5 FILLER_311_475 ();
 b15zdnd11an1n64x5 FILLER_311_539 ();
 b15zdnd11an1n64x5 FILLER_311_603 ();
 b15zdnd11an1n64x5 FILLER_311_667 ();
 b15zdnd11an1n08x5 FILLER_311_731 ();
 b15zdnd11an1n64x5 FILLER_311_744 ();
 b15zdnd11an1n16x5 FILLER_311_808 ();
 b15zdnd11an1n08x5 FILLER_311_824 ();
 b15zdnd11an1n04x5 FILLER_311_832 ();
 b15zdnd11an1n04x5 FILLER_311_839 ();
 b15zdnd11an1n04x5 FILLER_311_848 ();
 b15zdnd11an1n08x5 FILLER_311_858 ();
 b15zdnd11an1n64x5 FILLER_311_908 ();
 b15zdnd11an1n16x5 FILLER_311_977 ();
 b15zdnd11an1n64x5 FILLER_311_1016 ();
 b15zdnd11an1n64x5 FILLER_311_1080 ();
 b15zdnd00an1n01x5 FILLER_311_1144 ();
 b15zdnd11an1n64x5 FILLER_311_1157 ();
 b15zdnd11an1n64x5 FILLER_311_1221 ();
 b15zdnd11an1n08x5 FILLER_311_1285 ();
 b15zdnd11an1n64x5 FILLER_311_1296 ();
 b15zdnd11an1n16x5 FILLER_311_1360 ();
 b15zdnd11an1n64x5 FILLER_311_1387 ();
 b15zdnd11an1n32x5 FILLER_311_1451 ();
 b15zdnd11an1n08x5 FILLER_311_1483 ();
 b15zdnd11an1n04x5 FILLER_311_1491 ();
 b15zdnd00an1n02x5 FILLER_311_1495 ();
 b15zdnd00an1n01x5 FILLER_311_1497 ();
 b15zdnd11an1n04x5 FILLER_311_1501 ();
 b15zdnd11an1n64x5 FILLER_311_1508 ();
 b15zdnd11an1n64x5 FILLER_311_1572 ();
 b15zdnd11an1n64x5 FILLER_311_1636 ();
 b15zdnd11an1n64x5 FILLER_311_1700 ();
 b15zdnd11an1n64x5 FILLER_311_1764 ();
 b15zdnd11an1n64x5 FILLER_311_1828 ();
 b15zdnd11an1n64x5 FILLER_311_1892 ();
 b15zdnd11an1n64x5 FILLER_311_1956 ();
 b15zdnd11an1n64x5 FILLER_311_2020 ();
 b15zdnd11an1n64x5 FILLER_311_2084 ();
 b15zdnd11an1n64x5 FILLER_311_2148 ();
 b15zdnd11an1n64x5 FILLER_311_2212 ();
 b15zdnd11an1n08x5 FILLER_311_2276 ();
 b15zdnd11an1n64x5 FILLER_312_8 ();
 b15zdnd11an1n64x5 FILLER_312_72 ();
 b15zdnd11an1n64x5 FILLER_312_136 ();
 b15zdnd11an1n64x5 FILLER_312_200 ();
 b15zdnd11an1n64x5 FILLER_312_264 ();
 b15zdnd11an1n64x5 FILLER_312_328 ();
 b15zdnd11an1n64x5 FILLER_312_392 ();
 b15zdnd11an1n64x5 FILLER_312_456 ();
 b15zdnd11an1n64x5 FILLER_312_520 ();
 b15zdnd11an1n64x5 FILLER_312_584 ();
 b15zdnd11an1n32x5 FILLER_312_648 ();
 b15zdnd11an1n16x5 FILLER_312_680 ();
 b15zdnd11an1n08x5 FILLER_312_696 ();
 b15zdnd00an1n01x5 FILLER_312_704 ();
 b15zdnd11an1n08x5 FILLER_312_708 ();
 b15zdnd00an1n02x5 FILLER_312_716 ();
 b15zdnd11an1n08x5 FILLER_312_726 ();
 b15zdnd11an1n04x5 FILLER_312_734 ();
 b15zdnd00an1n01x5 FILLER_312_738 ();
 b15zdnd11an1n64x5 FILLER_312_746 ();
 b15zdnd11an1n16x5 FILLER_312_810 ();
 b15zdnd11an1n64x5 FILLER_312_878 ();
 b15zdnd11an1n16x5 FILLER_312_942 ();
 b15zdnd11an1n04x5 FILLER_312_958 ();
 b15zdnd00an1n02x5 FILLER_312_962 ();
 b15zdnd00an1n01x5 FILLER_312_964 ();
 b15zdnd11an1n04x5 FILLER_312_979 ();
 b15zdnd11an1n64x5 FILLER_312_995 ();
 b15zdnd11an1n64x5 FILLER_312_1059 ();
 b15zdnd11an1n64x5 FILLER_312_1123 ();
 b15zdnd11an1n64x5 FILLER_312_1187 ();
 b15zdnd11an1n64x5 FILLER_312_1251 ();
 b15zdnd11an1n64x5 FILLER_312_1315 ();
 b15zdnd11an1n64x5 FILLER_312_1379 ();
 b15zdnd11an1n16x5 FILLER_312_1443 ();
 b15zdnd11an1n04x5 FILLER_312_1459 ();
 b15zdnd00an1n02x5 FILLER_312_1463 ();
 b15zdnd00an1n01x5 FILLER_312_1465 ();
 b15zdnd11an1n64x5 FILLER_312_1506 ();
 b15zdnd11an1n64x5 FILLER_312_1570 ();
 b15zdnd11an1n64x5 FILLER_312_1634 ();
 b15zdnd11an1n32x5 FILLER_312_1698 ();
 b15zdnd00an1n02x5 FILLER_312_1730 ();
 b15zdnd11an1n04x5 FILLER_312_1735 ();
 b15zdnd11an1n64x5 FILLER_312_1742 ();
 b15zdnd11an1n64x5 FILLER_312_1806 ();
 b15zdnd11an1n64x5 FILLER_312_1870 ();
 b15zdnd11an1n64x5 FILLER_312_1934 ();
 b15zdnd11an1n64x5 FILLER_312_1998 ();
 b15zdnd11an1n64x5 FILLER_312_2062 ();
 b15zdnd11an1n16x5 FILLER_312_2126 ();
 b15zdnd11an1n08x5 FILLER_312_2142 ();
 b15zdnd11an1n04x5 FILLER_312_2150 ();
 b15zdnd11an1n64x5 FILLER_312_2162 ();
 b15zdnd11an1n32x5 FILLER_312_2226 ();
 b15zdnd11an1n16x5 FILLER_312_2258 ();
 b15zdnd00an1n02x5 FILLER_312_2274 ();
 b15zdnd11an1n64x5 FILLER_313_0 ();
 b15zdnd11an1n64x5 FILLER_313_64 ();
 b15zdnd11an1n64x5 FILLER_313_128 ();
 b15zdnd11an1n64x5 FILLER_313_192 ();
 b15zdnd11an1n64x5 FILLER_313_256 ();
 b15zdnd11an1n64x5 FILLER_313_320 ();
 b15zdnd11an1n64x5 FILLER_313_384 ();
 b15zdnd11an1n64x5 FILLER_313_448 ();
 b15zdnd11an1n64x5 FILLER_313_512 ();
 b15zdnd11an1n64x5 FILLER_313_576 ();
 b15zdnd11an1n32x5 FILLER_313_640 ();
 b15zdnd11an1n04x5 FILLER_313_672 ();
 b15zdnd00an1n02x5 FILLER_313_676 ();
 b15zdnd11an1n64x5 FILLER_313_730 ();
 b15zdnd11an1n32x5 FILLER_313_794 ();
 b15zdnd11an1n16x5 FILLER_313_826 ();
 b15zdnd11an1n04x5 FILLER_313_842 ();
 b15zdnd11an1n04x5 FILLER_313_849 ();
 b15zdnd11an1n64x5 FILLER_313_856 ();
 b15zdnd11an1n64x5 FILLER_313_920 ();
 b15zdnd11an1n04x5 FILLER_313_984 ();
 b15zdnd00an1n02x5 FILLER_313_988 ();
 b15zdnd00an1n01x5 FILLER_313_990 ();
 b15zdnd11an1n64x5 FILLER_313_1014 ();
 b15zdnd11an1n64x5 FILLER_313_1078 ();
 b15zdnd11an1n08x5 FILLER_313_1142 ();
 b15zdnd11an1n04x5 FILLER_313_1150 ();
 b15zdnd11an1n64x5 FILLER_313_1174 ();
 b15zdnd11an1n64x5 FILLER_313_1238 ();
 b15zdnd11an1n64x5 FILLER_313_1302 ();
 b15zdnd11an1n32x5 FILLER_313_1366 ();
 b15zdnd11an1n16x5 FILLER_313_1398 ();
 b15zdnd11an1n04x5 FILLER_313_1414 ();
 b15zdnd00an1n02x5 FILLER_313_1418 ();
 b15zdnd11an1n04x5 FILLER_313_1440 ();
 b15zdnd11an1n64x5 FILLER_313_1459 ();
 b15zdnd11an1n64x5 FILLER_313_1523 ();
 b15zdnd11an1n64x5 FILLER_313_1587 ();
 b15zdnd11an1n64x5 FILLER_313_1651 ();
 b15zdnd11an1n08x5 FILLER_313_1715 ();
 b15zdnd11an1n04x5 FILLER_313_1723 ();
 b15zdnd00an1n02x5 FILLER_313_1727 ();
 b15zdnd00an1n01x5 FILLER_313_1729 ();
 b15zdnd11an1n64x5 FILLER_313_1772 ();
 b15zdnd11an1n64x5 FILLER_313_1836 ();
 b15zdnd11an1n64x5 FILLER_313_1900 ();
 b15zdnd11an1n64x5 FILLER_313_1964 ();
 b15zdnd11an1n64x5 FILLER_313_2028 ();
 b15zdnd11an1n64x5 FILLER_313_2092 ();
 b15zdnd11an1n64x5 FILLER_313_2156 ();
 b15zdnd11an1n64x5 FILLER_313_2220 ();
 b15zdnd11an1n64x5 FILLER_314_8 ();
 b15zdnd11an1n64x5 FILLER_314_72 ();
 b15zdnd11an1n32x5 FILLER_314_136 ();
 b15zdnd00an1n02x5 FILLER_314_168 ();
 b15zdnd11an1n64x5 FILLER_314_212 ();
 b15zdnd11an1n64x5 FILLER_314_276 ();
 b15zdnd11an1n64x5 FILLER_314_340 ();
 b15zdnd11an1n64x5 FILLER_314_404 ();
 b15zdnd11an1n64x5 FILLER_314_468 ();
 b15zdnd11an1n64x5 FILLER_314_532 ();
 b15zdnd11an1n64x5 FILLER_314_596 ();
 b15zdnd11an1n32x5 FILLER_314_660 ();
 b15zdnd11an1n04x5 FILLER_314_692 ();
 b15zdnd11an1n04x5 FILLER_314_699 ();
 b15zdnd11an1n08x5 FILLER_314_706 ();
 b15zdnd11an1n04x5 FILLER_314_714 ();
 b15zdnd11an1n64x5 FILLER_314_726 ();
 b15zdnd11an1n64x5 FILLER_314_790 ();
 b15zdnd11an1n64x5 FILLER_314_854 ();
 b15zdnd11an1n64x5 FILLER_314_918 ();
 b15zdnd00an1n01x5 FILLER_314_982 ();
 b15zdnd11an1n64x5 FILLER_314_999 ();
 b15zdnd11an1n64x5 FILLER_314_1063 ();
 b15zdnd11an1n64x5 FILLER_314_1127 ();
 b15zdnd11an1n64x5 FILLER_314_1191 ();
 b15zdnd11an1n64x5 FILLER_314_1255 ();
 b15zdnd11an1n64x5 FILLER_314_1319 ();
 b15zdnd11an1n64x5 FILLER_314_1383 ();
 b15zdnd11an1n64x5 FILLER_314_1447 ();
 b15zdnd11an1n64x5 FILLER_314_1511 ();
 b15zdnd11an1n64x5 FILLER_314_1575 ();
 b15zdnd11an1n64x5 FILLER_314_1639 ();
 b15zdnd11an1n08x5 FILLER_314_1703 ();
 b15zdnd00an1n02x5 FILLER_314_1711 ();
 b15zdnd00an1n01x5 FILLER_314_1713 ();
 b15zdnd11an1n64x5 FILLER_314_1766 ();
 b15zdnd11an1n64x5 FILLER_314_1830 ();
 b15zdnd11an1n64x5 FILLER_314_1894 ();
 b15zdnd11an1n64x5 FILLER_314_1958 ();
 b15zdnd11an1n64x5 FILLER_314_2022 ();
 b15zdnd11an1n64x5 FILLER_314_2086 ();
 b15zdnd11an1n04x5 FILLER_314_2150 ();
 b15zdnd11an1n64x5 FILLER_314_2162 ();
 b15zdnd11an1n32x5 FILLER_314_2226 ();
 b15zdnd11an1n16x5 FILLER_314_2258 ();
 b15zdnd00an1n02x5 FILLER_314_2274 ();
 b15zdnd11an1n64x5 FILLER_315_0 ();
 b15zdnd11an1n64x5 FILLER_315_64 ();
 b15zdnd11an1n64x5 FILLER_315_128 ();
 b15zdnd11an1n64x5 FILLER_315_192 ();
 b15zdnd11an1n64x5 FILLER_315_256 ();
 b15zdnd11an1n64x5 FILLER_315_320 ();
 b15zdnd11an1n64x5 FILLER_315_384 ();
 b15zdnd11an1n64x5 FILLER_315_448 ();
 b15zdnd11an1n64x5 FILLER_315_512 ();
 b15zdnd11an1n64x5 FILLER_315_576 ();
 b15zdnd11an1n08x5 FILLER_315_640 ();
 b15zdnd00an1n02x5 FILLER_315_648 ();
 b15zdnd00an1n01x5 FILLER_315_650 ();
 b15zdnd11an1n32x5 FILLER_315_654 ();
 b15zdnd11an1n08x5 FILLER_315_686 ();
 b15zdnd11an1n64x5 FILLER_315_736 ();
 b15zdnd11an1n16x5 FILLER_315_800 ();
 b15zdnd11an1n08x5 FILLER_315_816 ();
 b15zdnd11an1n04x5 FILLER_315_824 ();
 b15zdnd00an1n02x5 FILLER_315_828 ();
 b15zdnd11an1n64x5 FILLER_315_848 ();
 b15zdnd11an1n64x5 FILLER_315_912 ();
 b15zdnd11an1n64x5 FILLER_315_976 ();
 b15zdnd11an1n64x5 FILLER_315_1040 ();
 b15zdnd11an1n64x5 FILLER_315_1104 ();
 b15zdnd11an1n08x5 FILLER_315_1168 ();
 b15zdnd11an1n64x5 FILLER_315_1184 ();
 b15zdnd11an1n64x5 FILLER_315_1248 ();
 b15zdnd11an1n64x5 FILLER_315_1312 ();
 b15zdnd11an1n64x5 FILLER_315_1376 ();
 b15zdnd11an1n64x5 FILLER_315_1440 ();
 b15zdnd11an1n64x5 FILLER_315_1504 ();
 b15zdnd11an1n64x5 FILLER_315_1568 ();
 b15zdnd11an1n64x5 FILLER_315_1632 ();
 b15zdnd11an1n32x5 FILLER_315_1696 ();
 b15zdnd11an1n08x5 FILLER_315_1728 ();
 b15zdnd00an1n02x5 FILLER_315_1736 ();
 b15zdnd00an1n01x5 FILLER_315_1738 ();
 b15zdnd11an1n64x5 FILLER_315_1742 ();
 b15zdnd11an1n64x5 FILLER_315_1806 ();
 b15zdnd11an1n64x5 FILLER_315_1870 ();
 b15zdnd11an1n32x5 FILLER_315_1934 ();
 b15zdnd11an1n16x5 FILLER_315_1966 ();
 b15zdnd11an1n04x5 FILLER_315_1982 ();
 b15zdnd00an1n02x5 FILLER_315_1986 ();
 b15zdnd00an1n01x5 FILLER_315_1988 ();
 b15zdnd11an1n04x5 FILLER_315_2029 ();
 b15zdnd11an1n64x5 FILLER_315_2036 ();
 b15zdnd11an1n64x5 FILLER_315_2100 ();
 b15zdnd11an1n64x5 FILLER_315_2164 ();
 b15zdnd11an1n32x5 FILLER_315_2228 ();
 b15zdnd11an1n16x5 FILLER_315_2260 ();
 b15zdnd11an1n08x5 FILLER_315_2276 ();
 b15zdnd11an1n64x5 FILLER_316_8 ();
 b15zdnd11an1n64x5 FILLER_316_72 ();
 b15zdnd11an1n64x5 FILLER_316_136 ();
 b15zdnd11an1n64x5 FILLER_316_200 ();
 b15zdnd11an1n64x5 FILLER_316_264 ();
 b15zdnd11an1n64x5 FILLER_316_328 ();
 b15zdnd11an1n64x5 FILLER_316_392 ();
 b15zdnd11an1n64x5 FILLER_316_456 ();
 b15zdnd11an1n64x5 FILLER_316_520 ();
 b15zdnd11an1n32x5 FILLER_316_584 ();
 b15zdnd11an1n08x5 FILLER_316_616 ();
 b15zdnd11an1n32x5 FILLER_316_676 ();
 b15zdnd11an1n08x5 FILLER_316_708 ();
 b15zdnd00an1n02x5 FILLER_316_716 ();
 b15zdnd11an1n32x5 FILLER_316_726 ();
 b15zdnd11an1n64x5 FILLER_316_800 ();
 b15zdnd11an1n64x5 FILLER_316_864 ();
 b15zdnd11an1n64x5 FILLER_316_928 ();
 b15zdnd11an1n32x5 FILLER_316_992 ();
 b15zdnd00an1n01x5 FILLER_316_1024 ();
 b15zdnd11an1n64x5 FILLER_316_1031 ();
 b15zdnd11an1n64x5 FILLER_316_1095 ();
 b15zdnd11an1n04x5 FILLER_316_1159 ();
 b15zdnd11an1n32x5 FILLER_316_1173 ();
 b15zdnd11an1n08x5 FILLER_316_1205 ();
 b15zdnd00an1n01x5 FILLER_316_1213 ();
 b15zdnd11an1n64x5 FILLER_316_1225 ();
 b15zdnd11an1n64x5 FILLER_316_1289 ();
 b15zdnd11an1n64x5 FILLER_316_1353 ();
 b15zdnd11an1n64x5 FILLER_316_1417 ();
 b15zdnd11an1n64x5 FILLER_316_1481 ();
 b15zdnd11an1n64x5 FILLER_316_1545 ();
 b15zdnd11an1n64x5 FILLER_316_1609 ();
 b15zdnd11an1n64x5 FILLER_316_1673 ();
 b15zdnd11an1n64x5 FILLER_316_1737 ();
 b15zdnd11an1n64x5 FILLER_316_1801 ();
 b15zdnd11an1n64x5 FILLER_316_1865 ();
 b15zdnd11an1n64x5 FILLER_316_1929 ();
 b15zdnd11an1n32x5 FILLER_316_1993 ();
 b15zdnd11an1n64x5 FILLER_316_2028 ();
 b15zdnd11an1n32x5 FILLER_316_2092 ();
 b15zdnd11an1n16x5 FILLER_316_2124 ();
 b15zdnd11an1n08x5 FILLER_316_2140 ();
 b15zdnd11an1n04x5 FILLER_316_2148 ();
 b15zdnd00an1n02x5 FILLER_316_2152 ();
 b15zdnd11an1n64x5 FILLER_316_2162 ();
 b15zdnd11an1n16x5 FILLER_316_2226 ();
 b15zdnd11an1n08x5 FILLER_316_2242 ();
 b15zdnd00an1n02x5 FILLER_316_2250 ();
 b15zdnd11an1n16x5 FILLER_316_2258 ();
 b15zdnd00an1n02x5 FILLER_316_2274 ();
 b15zdnd11an1n64x5 FILLER_317_0 ();
 b15zdnd11an1n64x5 FILLER_317_64 ();
 b15zdnd11an1n64x5 FILLER_317_128 ();
 b15zdnd11an1n64x5 FILLER_317_192 ();
 b15zdnd11an1n16x5 FILLER_317_256 ();
 b15zdnd00an1n01x5 FILLER_317_272 ();
 b15zdnd11an1n64x5 FILLER_317_276 ();
 b15zdnd11an1n64x5 FILLER_317_340 ();
 b15zdnd11an1n64x5 FILLER_317_404 ();
 b15zdnd11an1n64x5 FILLER_317_468 ();
 b15zdnd11an1n64x5 FILLER_317_532 ();
 b15zdnd11an1n16x5 FILLER_317_596 ();
 b15zdnd11an1n08x5 FILLER_317_612 ();
 b15zdnd11an1n04x5 FILLER_317_620 ();
 b15zdnd00an1n01x5 FILLER_317_624 ();
 b15zdnd11an1n08x5 FILLER_317_630 ();
 b15zdnd11an1n04x5 FILLER_317_638 ();
 b15zdnd11an1n04x5 FILLER_317_645 ();
 b15zdnd11an1n64x5 FILLER_317_652 ();
 b15zdnd11an1n64x5 FILLER_317_716 ();
 b15zdnd11an1n64x5 FILLER_317_780 ();
 b15zdnd11an1n64x5 FILLER_317_844 ();
 b15zdnd11an1n64x5 FILLER_317_908 ();
 b15zdnd11an1n64x5 FILLER_317_972 ();
 b15zdnd11an1n64x5 FILLER_317_1036 ();
 b15zdnd11an1n64x5 FILLER_317_1100 ();
 b15zdnd11an1n64x5 FILLER_317_1164 ();
 b15zdnd11an1n64x5 FILLER_317_1228 ();
 b15zdnd11an1n32x5 FILLER_317_1292 ();
 b15zdnd11an1n16x5 FILLER_317_1324 ();
 b15zdnd11an1n08x5 FILLER_317_1340 ();
 b15zdnd00an1n01x5 FILLER_317_1348 ();
 b15zdnd11an1n04x5 FILLER_317_1352 ();
 b15zdnd11an1n64x5 FILLER_317_1359 ();
 b15zdnd11an1n64x5 FILLER_317_1423 ();
 b15zdnd11an1n64x5 FILLER_317_1487 ();
 b15zdnd11an1n64x5 FILLER_317_1551 ();
 b15zdnd11an1n64x5 FILLER_317_1615 ();
 b15zdnd11an1n64x5 FILLER_317_1679 ();
 b15zdnd11an1n64x5 FILLER_317_1743 ();
 b15zdnd11an1n64x5 FILLER_317_1807 ();
 b15zdnd11an1n64x5 FILLER_317_1871 ();
 b15zdnd11an1n64x5 FILLER_317_1935 ();
 b15zdnd11an1n64x5 FILLER_317_1999 ();
 b15zdnd11an1n64x5 FILLER_317_2063 ();
 b15zdnd11an1n64x5 FILLER_317_2127 ();
 b15zdnd11an1n64x5 FILLER_317_2191 ();
 b15zdnd11an1n16x5 FILLER_317_2255 ();
 b15zdnd11an1n08x5 FILLER_317_2271 ();
 b15zdnd11an1n04x5 FILLER_317_2279 ();
 b15zdnd00an1n01x5 FILLER_317_2283 ();
 b15zdnd11an1n64x5 FILLER_318_8 ();
 b15zdnd11an1n64x5 FILLER_318_72 ();
 b15zdnd11an1n32x5 FILLER_318_136 ();
 b15zdnd11an1n08x5 FILLER_318_168 ();
 b15zdnd11an1n32x5 FILLER_318_180 ();
 b15zdnd11an1n16x5 FILLER_318_212 ();
 b15zdnd11an1n08x5 FILLER_318_228 ();
 b15zdnd11an1n04x5 FILLER_318_236 ();
 b15zdnd00an1n01x5 FILLER_318_240 ();
 b15zdnd11an1n64x5 FILLER_318_281 ();
 b15zdnd11an1n64x5 FILLER_318_345 ();
 b15zdnd11an1n64x5 FILLER_318_409 ();
 b15zdnd11an1n64x5 FILLER_318_473 ();
 b15zdnd11an1n64x5 FILLER_318_537 ();
 b15zdnd11an1n16x5 FILLER_318_601 ();
 b15zdnd11an1n08x5 FILLER_318_617 ();
 b15zdnd00an1n01x5 FILLER_318_625 ();
 b15zdnd11an1n32x5 FILLER_318_668 ();
 b15zdnd11an1n16x5 FILLER_318_700 ();
 b15zdnd00an1n02x5 FILLER_318_716 ();
 b15zdnd11an1n64x5 FILLER_318_726 ();
 b15zdnd11an1n64x5 FILLER_318_790 ();
 b15zdnd11an1n64x5 FILLER_318_854 ();
 b15zdnd11an1n64x5 FILLER_318_918 ();
 b15zdnd11an1n64x5 FILLER_318_982 ();
 b15zdnd11an1n64x5 FILLER_318_1046 ();
 b15zdnd11an1n32x5 FILLER_318_1110 ();
 b15zdnd11an1n16x5 FILLER_318_1142 ();
 b15zdnd11an1n08x5 FILLER_318_1158 ();
 b15zdnd11an1n32x5 FILLER_318_1175 ();
 b15zdnd00an1n01x5 FILLER_318_1207 ();
 b15zdnd11an1n64x5 FILLER_318_1215 ();
 b15zdnd11an1n32x5 FILLER_318_1279 ();
 b15zdnd11an1n16x5 FILLER_318_1311 ();
 b15zdnd11an1n04x5 FILLER_318_1327 ();
 b15zdnd11an1n64x5 FILLER_318_1383 ();
 b15zdnd11an1n64x5 FILLER_318_1447 ();
 b15zdnd11an1n64x5 FILLER_318_1511 ();
 b15zdnd11an1n64x5 FILLER_318_1575 ();
 b15zdnd11an1n64x5 FILLER_318_1639 ();
 b15zdnd11an1n64x5 FILLER_318_1703 ();
 b15zdnd11an1n64x5 FILLER_318_1767 ();
 b15zdnd11an1n64x5 FILLER_318_1831 ();
 b15zdnd11an1n64x5 FILLER_318_1895 ();
 b15zdnd11an1n64x5 FILLER_318_1959 ();
 b15zdnd11an1n32x5 FILLER_318_2023 ();
 b15zdnd11an1n08x5 FILLER_318_2055 ();
 b15zdnd11an1n04x5 FILLER_318_2063 ();
 b15zdnd00an1n02x5 FILLER_318_2067 ();
 b15zdnd11an1n64x5 FILLER_318_2073 ();
 b15zdnd11an1n16x5 FILLER_318_2137 ();
 b15zdnd00an1n01x5 FILLER_318_2153 ();
 b15zdnd11an1n64x5 FILLER_318_2162 ();
 b15zdnd11an1n16x5 FILLER_318_2226 ();
 b15zdnd11an1n08x5 FILLER_318_2242 ();
 b15zdnd11an1n04x5 FILLER_318_2250 ();
 b15zdnd00an1n01x5 FILLER_318_2254 ();
 b15zdnd11an1n16x5 FILLER_318_2260 ();
 b15zdnd11an1n64x5 FILLER_319_0 ();
 b15zdnd11an1n64x5 FILLER_319_64 ();
 b15zdnd11an1n32x5 FILLER_319_128 ();
 b15zdnd11an1n08x5 FILLER_319_160 ();
 b15zdnd11an1n04x5 FILLER_319_168 ();
 b15zdnd00an1n02x5 FILLER_319_172 ();
 b15zdnd11an1n64x5 FILLER_319_181 ();
 b15zdnd11an1n32x5 FILLER_319_245 ();
 b15zdnd00an1n02x5 FILLER_319_277 ();
 b15zdnd11an1n64x5 FILLER_319_282 ();
 b15zdnd11an1n64x5 FILLER_319_346 ();
 b15zdnd11an1n64x5 FILLER_319_410 ();
 b15zdnd11an1n64x5 FILLER_319_474 ();
 b15zdnd11an1n32x5 FILLER_319_538 ();
 b15zdnd11an1n16x5 FILLER_319_570 ();
 b15zdnd11an1n08x5 FILLER_319_586 ();
 b15zdnd11an1n04x5 FILLER_319_594 ();
 b15zdnd00an1n01x5 FILLER_319_598 ();
 b15zdnd11an1n04x5 FILLER_319_602 ();
 b15zdnd11an1n64x5 FILLER_319_615 ();
 b15zdnd11an1n64x5 FILLER_319_679 ();
 b15zdnd11an1n64x5 FILLER_319_743 ();
 b15zdnd11an1n64x5 FILLER_319_807 ();
 b15zdnd11an1n64x5 FILLER_319_871 ();
 b15zdnd11an1n32x5 FILLER_319_935 ();
 b15zdnd11an1n16x5 FILLER_319_967 ();
 b15zdnd11an1n08x5 FILLER_319_983 ();
 b15zdnd11an1n04x5 FILLER_319_991 ();
 b15zdnd00an1n02x5 FILLER_319_995 ();
 b15zdnd00an1n01x5 FILLER_319_997 ();
 b15zdnd11an1n64x5 FILLER_319_1005 ();
 b15zdnd11an1n64x5 FILLER_319_1069 ();
 b15zdnd11an1n64x5 FILLER_319_1133 ();
 b15zdnd11an1n16x5 FILLER_319_1197 ();
 b15zdnd00an1n01x5 FILLER_319_1213 ();
 b15zdnd11an1n64x5 FILLER_319_1217 ();
 b15zdnd11an1n64x5 FILLER_319_1281 ();
 b15zdnd11an1n08x5 FILLER_319_1345 ();
 b15zdnd11an1n04x5 FILLER_319_1353 ();
 b15zdnd11an1n64x5 FILLER_319_1360 ();
 b15zdnd11an1n32x5 FILLER_319_1424 ();
 b15zdnd11an1n04x5 FILLER_319_1456 ();
 b15zdnd00an1n01x5 FILLER_319_1460 ();
 b15zdnd11an1n64x5 FILLER_319_1513 ();
 b15zdnd11an1n64x5 FILLER_319_1577 ();
 b15zdnd11an1n64x5 FILLER_319_1641 ();
 b15zdnd11an1n64x5 FILLER_319_1705 ();
 b15zdnd11an1n64x5 FILLER_319_1769 ();
 b15zdnd11an1n64x5 FILLER_319_1833 ();
 b15zdnd11an1n64x5 FILLER_319_1897 ();
 b15zdnd11an1n64x5 FILLER_319_1961 ();
 b15zdnd11an1n32x5 FILLER_319_2025 ();
 b15zdnd11an1n04x5 FILLER_319_2057 ();
 b15zdnd00an1n02x5 FILLER_319_2061 ();
 b15zdnd11an1n64x5 FILLER_319_2073 ();
 b15zdnd11an1n64x5 FILLER_319_2137 ();
 b15zdnd11an1n64x5 FILLER_319_2201 ();
 b15zdnd11an1n16x5 FILLER_319_2265 ();
 b15zdnd00an1n02x5 FILLER_319_2281 ();
 b15zdnd00an1n01x5 FILLER_319_2283 ();
 b15zdnd11an1n64x5 FILLER_320_8 ();
 b15zdnd11an1n64x5 FILLER_320_72 ();
 b15zdnd11an1n64x5 FILLER_320_136 ();
 b15zdnd11an1n08x5 FILLER_320_200 ();
 b15zdnd00an1n02x5 FILLER_320_208 ();
 b15zdnd00an1n01x5 FILLER_320_210 ();
 b15zdnd11an1n64x5 FILLER_320_253 ();
 b15zdnd11an1n64x5 FILLER_320_317 ();
 b15zdnd11an1n64x5 FILLER_320_381 ();
 b15zdnd11an1n32x5 FILLER_320_445 ();
 b15zdnd11an1n16x5 FILLER_320_477 ();
 b15zdnd00an1n02x5 FILLER_320_493 ();
 b15zdnd00an1n01x5 FILLER_320_495 ();
 b15zdnd11an1n04x5 FILLER_320_501 ();
 b15zdnd11an1n32x5 FILLER_320_516 ();
 b15zdnd11an1n16x5 FILLER_320_548 ();
 b15zdnd11an1n08x5 FILLER_320_564 ();
 b15zdnd11an1n04x5 FILLER_320_572 ();
 b15zdnd11an1n64x5 FILLER_320_628 ();
 b15zdnd11an1n16x5 FILLER_320_692 ();
 b15zdnd11an1n08x5 FILLER_320_708 ();
 b15zdnd00an1n02x5 FILLER_320_716 ();
 b15zdnd11an1n64x5 FILLER_320_726 ();
 b15zdnd11an1n64x5 FILLER_320_790 ();
 b15zdnd11an1n64x5 FILLER_320_854 ();
 b15zdnd11an1n64x5 FILLER_320_918 ();
 b15zdnd11an1n64x5 FILLER_320_982 ();
 b15zdnd11an1n16x5 FILLER_320_1046 ();
 b15zdnd11an1n08x5 FILLER_320_1062 ();
 b15zdnd11an1n04x5 FILLER_320_1070 ();
 b15zdnd00an1n01x5 FILLER_320_1074 ();
 b15zdnd11an1n04x5 FILLER_320_1085 ();
 b15zdnd11an1n64x5 FILLER_320_1101 ();
 b15zdnd11an1n64x5 FILLER_320_1165 ();
 b15zdnd11an1n64x5 FILLER_320_1229 ();
 b15zdnd11an1n64x5 FILLER_320_1293 ();
 b15zdnd11an1n64x5 FILLER_320_1357 ();
 b15zdnd11an1n32x5 FILLER_320_1421 ();
 b15zdnd11an1n16x5 FILLER_320_1453 ();
 b15zdnd11an1n08x5 FILLER_320_1469 ();
 b15zdnd11an1n04x5 FILLER_320_1480 ();
 b15zdnd11an1n64x5 FILLER_320_1487 ();
 b15zdnd11an1n64x5 FILLER_320_1551 ();
 b15zdnd11an1n64x5 FILLER_320_1615 ();
 b15zdnd11an1n64x5 FILLER_320_1679 ();
 b15zdnd11an1n32x5 FILLER_320_1743 ();
 b15zdnd11an1n08x5 FILLER_320_1775 ();
 b15zdnd11an1n64x5 FILLER_320_1789 ();
 b15zdnd11an1n64x5 FILLER_320_1853 ();
 b15zdnd11an1n64x5 FILLER_320_1917 ();
 b15zdnd11an1n64x5 FILLER_320_1981 ();
 b15zdnd11an1n64x5 FILLER_320_2045 ();
 b15zdnd11an1n32x5 FILLER_320_2109 ();
 b15zdnd11an1n08x5 FILLER_320_2141 ();
 b15zdnd11an1n04x5 FILLER_320_2149 ();
 b15zdnd00an1n01x5 FILLER_320_2153 ();
 b15zdnd11an1n64x5 FILLER_320_2162 ();
 b15zdnd11an1n32x5 FILLER_320_2226 ();
 b15zdnd11an1n16x5 FILLER_320_2258 ();
 b15zdnd00an1n02x5 FILLER_320_2274 ();
 b15zdnd11an1n64x5 FILLER_321_0 ();
 b15zdnd11an1n64x5 FILLER_321_64 ();
 b15zdnd11an1n64x5 FILLER_321_128 ();
 b15zdnd11an1n64x5 FILLER_321_192 ();
 b15zdnd11an1n64x5 FILLER_321_256 ();
 b15zdnd11an1n16x5 FILLER_321_320 ();
 b15zdnd11an1n08x5 FILLER_321_336 ();
 b15zdnd00an1n01x5 FILLER_321_344 ();
 b15zdnd11an1n64x5 FILLER_321_348 ();
 b15zdnd11an1n32x5 FILLER_321_412 ();
 b15zdnd11an1n16x5 FILLER_321_444 ();
 b15zdnd11an1n08x5 FILLER_321_460 ();
 b15zdnd11an1n04x5 FILLER_321_468 ();
 b15zdnd00an1n02x5 FILLER_321_472 ();
 b15zdnd00an1n01x5 FILLER_321_474 ();
 b15zdnd11an1n16x5 FILLER_321_486 ();
 b15zdnd11an1n64x5 FILLER_321_511 ();
 b15zdnd11an1n16x5 FILLER_321_575 ();
 b15zdnd11an1n04x5 FILLER_321_591 ();
 b15zdnd00an1n01x5 FILLER_321_595 ();
 b15zdnd11an1n04x5 FILLER_321_599 ();
 b15zdnd11an1n64x5 FILLER_321_606 ();
 b15zdnd11an1n64x5 FILLER_321_670 ();
 b15zdnd11an1n64x5 FILLER_321_734 ();
 b15zdnd11an1n64x5 FILLER_321_798 ();
 b15zdnd11an1n64x5 FILLER_321_862 ();
 b15zdnd11an1n64x5 FILLER_321_926 ();
 b15zdnd11an1n32x5 FILLER_321_990 ();
 b15zdnd11an1n08x5 FILLER_321_1022 ();
 b15zdnd11an1n04x5 FILLER_321_1030 ();
 b15zdnd00an1n02x5 FILLER_321_1034 ();
 b15zdnd11an1n64x5 FILLER_321_1078 ();
 b15zdnd11an1n04x5 FILLER_321_1142 ();
 b15zdnd00an1n02x5 FILLER_321_1146 ();
 b15zdnd00an1n01x5 FILLER_321_1148 ();
 b15zdnd11an1n64x5 FILLER_321_1167 ();
 b15zdnd11an1n08x5 FILLER_321_1231 ();
 b15zdnd11an1n64x5 FILLER_321_1249 ();
 b15zdnd11an1n64x5 FILLER_321_1313 ();
 b15zdnd11an1n64x5 FILLER_321_1377 ();
 b15zdnd11an1n16x5 FILLER_321_1441 ();
 b15zdnd11an1n08x5 FILLER_321_1457 ();
 b15zdnd11an1n04x5 FILLER_321_1465 ();
 b15zdnd00an1n01x5 FILLER_321_1469 ();
 b15zdnd11an1n64x5 FILLER_321_1473 ();
 b15zdnd11an1n32x5 FILLER_321_1537 ();
 b15zdnd11an1n08x5 FILLER_321_1569 ();
 b15zdnd11an1n04x5 FILLER_321_1577 ();
 b15zdnd00an1n02x5 FILLER_321_1581 ();
 b15zdnd00an1n01x5 FILLER_321_1583 ();
 b15zdnd11an1n64x5 FILLER_321_1595 ();
 b15zdnd11an1n64x5 FILLER_321_1659 ();
 b15zdnd11an1n64x5 FILLER_321_1723 ();
 b15zdnd11an1n64x5 FILLER_321_1787 ();
 b15zdnd11an1n16x5 FILLER_321_1851 ();
 b15zdnd11an1n64x5 FILLER_321_1874 ();
 b15zdnd11an1n64x5 FILLER_321_1938 ();
 b15zdnd11an1n64x5 FILLER_321_2002 ();
 b15zdnd11an1n64x5 FILLER_321_2066 ();
 b15zdnd11an1n64x5 FILLER_321_2130 ();
 b15zdnd11an1n64x5 FILLER_321_2194 ();
 b15zdnd11an1n16x5 FILLER_321_2258 ();
 b15zdnd11an1n08x5 FILLER_321_2274 ();
 b15zdnd00an1n02x5 FILLER_321_2282 ();
 b15zdnd11an1n64x5 FILLER_322_8 ();
 b15zdnd11an1n64x5 FILLER_322_72 ();
 b15zdnd11an1n64x5 FILLER_322_136 ();
 b15zdnd11an1n64x5 FILLER_322_200 ();
 b15zdnd11an1n16x5 FILLER_322_264 ();
 b15zdnd11an1n04x5 FILLER_322_280 ();
 b15zdnd00an1n02x5 FILLER_322_284 ();
 b15zdnd11an1n64x5 FILLER_322_292 ();
 b15zdnd11an1n64x5 FILLER_322_356 ();
 b15zdnd11an1n64x5 FILLER_322_420 ();
 b15zdnd11an1n04x5 FILLER_322_490 ();
 b15zdnd11an1n64x5 FILLER_322_502 ();
 b15zdnd11an1n64x5 FILLER_322_566 ();
 b15zdnd11an1n64x5 FILLER_322_630 ();
 b15zdnd11an1n16x5 FILLER_322_694 ();
 b15zdnd11an1n08x5 FILLER_322_710 ();
 b15zdnd11an1n64x5 FILLER_322_726 ();
 b15zdnd11an1n64x5 FILLER_322_790 ();
 b15zdnd11an1n64x5 FILLER_322_854 ();
 b15zdnd11an1n64x5 FILLER_322_918 ();
 b15zdnd11an1n64x5 FILLER_322_982 ();
 b15zdnd11an1n32x5 FILLER_322_1046 ();
 b15zdnd11an1n16x5 FILLER_322_1109 ();
 b15zdnd11an1n08x5 FILLER_322_1125 ();
 b15zdnd00an1n02x5 FILLER_322_1133 ();
 b15zdnd11an1n64x5 FILLER_322_1150 ();
 b15zdnd11an1n64x5 FILLER_322_1214 ();
 b15zdnd11an1n64x5 FILLER_322_1278 ();
 b15zdnd11an1n64x5 FILLER_322_1342 ();
 b15zdnd11an1n64x5 FILLER_322_1406 ();
 b15zdnd11an1n64x5 FILLER_322_1470 ();
 b15zdnd11an1n32x5 FILLER_322_1534 ();
 b15zdnd11an1n16x5 FILLER_322_1566 ();
 b15zdnd11an1n08x5 FILLER_322_1582 ();
 b15zdnd00an1n02x5 FILLER_322_1590 ();
 b15zdnd11an1n16x5 FILLER_322_1602 ();
 b15zdnd11an1n08x5 FILLER_322_1618 ();
 b15zdnd00an1n01x5 FILLER_322_1626 ();
 b15zdnd11an1n04x5 FILLER_322_1630 ();
 b15zdnd11an1n64x5 FILLER_322_1637 ();
 b15zdnd11an1n64x5 FILLER_322_1701 ();
 b15zdnd11an1n64x5 FILLER_322_1765 ();
 b15zdnd11an1n32x5 FILLER_322_1829 ();
 b15zdnd11an1n16x5 FILLER_322_1861 ();
 b15zdnd11an1n08x5 FILLER_322_1877 ();
 b15zdnd11an1n64x5 FILLER_322_1910 ();
 b15zdnd11an1n64x5 FILLER_322_1974 ();
 b15zdnd11an1n16x5 FILLER_322_2038 ();
 b15zdnd00an1n01x5 FILLER_322_2054 ();
 b15zdnd11an1n64x5 FILLER_322_2067 ();
 b15zdnd11an1n16x5 FILLER_322_2131 ();
 b15zdnd11an1n04x5 FILLER_322_2147 ();
 b15zdnd00an1n02x5 FILLER_322_2151 ();
 b15zdnd00an1n01x5 FILLER_322_2153 ();
 b15zdnd11an1n64x5 FILLER_322_2162 ();
 b15zdnd11an1n32x5 FILLER_322_2226 ();
 b15zdnd11an1n16x5 FILLER_322_2258 ();
 b15zdnd00an1n02x5 FILLER_322_2274 ();
 b15zdnd11an1n64x5 FILLER_323_0 ();
 b15zdnd11an1n64x5 FILLER_323_64 ();
 b15zdnd11an1n64x5 FILLER_323_128 ();
 b15zdnd11an1n64x5 FILLER_323_192 ();
 b15zdnd11an1n16x5 FILLER_323_256 ();
 b15zdnd11an1n04x5 FILLER_323_272 ();
 b15zdnd00an1n02x5 FILLER_323_276 ();
 b15zdnd00an1n01x5 FILLER_323_278 ();
 b15zdnd11an1n04x5 FILLER_323_285 ();
 b15zdnd11an1n04x5 FILLER_323_304 ();
 b15zdnd11an1n64x5 FILLER_323_320 ();
 b15zdnd11an1n08x5 FILLER_323_384 ();
 b15zdnd11an1n04x5 FILLER_323_392 ();
 b15zdnd00an1n02x5 FILLER_323_396 ();
 b15zdnd11an1n64x5 FILLER_323_401 ();
 b15zdnd11an1n08x5 FILLER_323_465 ();
 b15zdnd00an1n01x5 FILLER_323_473 ();
 b15zdnd11an1n04x5 FILLER_323_483 ();
 b15zdnd11an1n16x5 FILLER_323_491 ();
 b15zdnd11an1n64x5 FILLER_323_511 ();
 b15zdnd11an1n64x5 FILLER_323_575 ();
 b15zdnd11an1n64x5 FILLER_323_639 ();
 b15zdnd11an1n04x5 FILLER_323_703 ();
 b15zdnd00an1n02x5 FILLER_323_707 ();
 b15zdnd00an1n01x5 FILLER_323_709 ();
 b15zdnd11an1n64x5 FILLER_323_752 ();
 b15zdnd11an1n64x5 FILLER_323_816 ();
 b15zdnd11an1n64x5 FILLER_323_880 ();
 b15zdnd11an1n64x5 FILLER_323_944 ();
 b15zdnd11an1n64x5 FILLER_323_1008 ();
 b15zdnd11an1n64x5 FILLER_323_1072 ();
 b15zdnd11an1n32x5 FILLER_323_1136 ();
 b15zdnd11an1n16x5 FILLER_323_1168 ();
 b15zdnd11an1n08x5 FILLER_323_1184 ();
 b15zdnd00an1n02x5 FILLER_323_1192 ();
 b15zdnd00an1n01x5 FILLER_323_1194 ();
 b15zdnd11an1n64x5 FILLER_323_1199 ();
 b15zdnd11an1n64x5 FILLER_323_1263 ();
 b15zdnd11an1n64x5 FILLER_323_1327 ();
 b15zdnd11an1n64x5 FILLER_323_1391 ();
 b15zdnd11an1n32x5 FILLER_323_1455 ();
 b15zdnd11an1n08x5 FILLER_323_1487 ();
 b15zdnd00an1n02x5 FILLER_323_1495 ();
 b15zdnd11an1n04x5 FILLER_323_1505 ();
 b15zdnd11an1n64x5 FILLER_323_1513 ();
 b15zdnd11an1n04x5 FILLER_323_1577 ();
 b15zdnd00an1n02x5 FILLER_323_1581 ();
 b15zdnd11an1n08x5 FILLER_323_1589 ();
 b15zdnd11an1n04x5 FILLER_323_1597 ();
 b15zdnd11an1n04x5 FILLER_323_1605 ();
 b15zdnd11an1n64x5 FILLER_323_1661 ();
 b15zdnd11an1n64x5 FILLER_323_1725 ();
 b15zdnd11an1n64x5 FILLER_323_1789 ();
 b15zdnd11an1n64x5 FILLER_323_1853 ();
 b15zdnd11an1n64x5 FILLER_323_1917 ();
 b15zdnd11an1n64x5 FILLER_323_1981 ();
 b15zdnd11an1n04x5 FILLER_323_2045 ();
 b15zdnd00an1n02x5 FILLER_323_2049 ();
 b15zdnd11an1n08x5 FILLER_323_2059 ();
 b15zdnd11an1n04x5 FILLER_323_2067 ();
 b15zdnd00an1n02x5 FILLER_323_2071 ();
 b15zdnd11an1n64x5 FILLER_323_2080 ();
 b15zdnd11an1n64x5 FILLER_323_2144 ();
 b15zdnd11an1n64x5 FILLER_323_2208 ();
 b15zdnd11an1n08x5 FILLER_323_2272 ();
 b15zdnd11an1n04x5 FILLER_323_2280 ();
 b15zdnd11an1n64x5 FILLER_324_8 ();
 b15zdnd11an1n64x5 FILLER_324_72 ();
 b15zdnd11an1n64x5 FILLER_324_136 ();
 b15zdnd11an1n64x5 FILLER_324_200 ();
 b15zdnd11an1n08x5 FILLER_324_264 ();
 b15zdnd00an1n02x5 FILLER_324_272 ();
 b15zdnd00an1n01x5 FILLER_324_274 ();
 b15zdnd11an1n04x5 FILLER_324_315 ();
 b15zdnd11an1n16x5 FILLER_324_322 ();
 b15zdnd11an1n08x5 FILLER_324_338 ();
 b15zdnd11an1n04x5 FILLER_324_346 ();
 b15zdnd00an1n01x5 FILLER_324_350 ();
 b15zdnd11an1n04x5 FILLER_324_367 ();
 b15zdnd11an1n16x5 FILLER_324_423 ();
 b15zdnd11an1n04x5 FILLER_324_439 ();
 b15zdnd11an1n08x5 FILLER_324_455 ();
 b15zdnd11an1n04x5 FILLER_324_463 ();
 b15zdnd00an1n01x5 FILLER_324_467 ();
 b15zdnd11an1n04x5 FILLER_324_484 ();
 b15zdnd00an1n02x5 FILLER_324_488 ();
 b15zdnd11an1n04x5 FILLER_324_505 ();
 b15zdnd11an1n04x5 FILLER_324_523 ();
 b15zdnd11an1n64x5 FILLER_324_531 ();
 b15zdnd11an1n64x5 FILLER_324_595 ();
 b15zdnd11an1n32x5 FILLER_324_659 ();
 b15zdnd11an1n16x5 FILLER_324_691 ();
 b15zdnd11an1n08x5 FILLER_324_707 ();
 b15zdnd00an1n02x5 FILLER_324_715 ();
 b15zdnd00an1n01x5 FILLER_324_717 ();
 b15zdnd11an1n32x5 FILLER_324_726 ();
 b15zdnd11an1n16x5 FILLER_324_758 ();
 b15zdnd11an1n08x5 FILLER_324_774 ();
 b15zdnd11an1n04x5 FILLER_324_782 ();
 b15zdnd00an1n01x5 FILLER_324_786 ();
 b15zdnd11an1n64x5 FILLER_324_829 ();
 b15zdnd11an1n64x5 FILLER_324_893 ();
 b15zdnd11an1n64x5 FILLER_324_957 ();
 b15zdnd11an1n64x5 FILLER_324_1021 ();
 b15zdnd11an1n64x5 FILLER_324_1085 ();
 b15zdnd11an1n32x5 FILLER_324_1149 ();
 b15zdnd11an1n08x5 FILLER_324_1181 ();
 b15zdnd00an1n02x5 FILLER_324_1189 ();
 b15zdnd11an1n04x5 FILLER_324_1200 ();
 b15zdnd11an1n64x5 FILLER_324_1216 ();
 b15zdnd11an1n64x5 FILLER_324_1280 ();
 b15zdnd11an1n64x5 FILLER_324_1344 ();
 b15zdnd11an1n64x5 FILLER_324_1408 ();
 b15zdnd11an1n32x5 FILLER_324_1472 ();
 b15zdnd00an1n02x5 FILLER_324_1504 ();
 b15zdnd11an1n64x5 FILLER_324_1511 ();
 b15zdnd11an1n32x5 FILLER_324_1575 ();
 b15zdnd11an1n16x5 FILLER_324_1607 ();
 b15zdnd11an1n08x5 FILLER_324_1623 ();
 b15zdnd11an1n04x5 FILLER_324_1631 ();
 b15zdnd11an1n64x5 FILLER_324_1638 ();
 b15zdnd11an1n64x5 FILLER_324_1702 ();
 b15zdnd11an1n64x5 FILLER_324_1766 ();
 b15zdnd11an1n64x5 FILLER_324_1830 ();
 b15zdnd11an1n64x5 FILLER_324_1894 ();
 b15zdnd11an1n64x5 FILLER_324_1958 ();
 b15zdnd11an1n16x5 FILLER_324_2022 ();
 b15zdnd11an1n08x5 FILLER_324_2038 ();
 b15zdnd11an1n04x5 FILLER_324_2046 ();
 b15zdnd11an1n64x5 FILLER_324_2075 ();
 b15zdnd11an1n08x5 FILLER_324_2139 ();
 b15zdnd11an1n04x5 FILLER_324_2147 ();
 b15zdnd00an1n02x5 FILLER_324_2151 ();
 b15zdnd00an1n01x5 FILLER_324_2153 ();
 b15zdnd11an1n64x5 FILLER_324_2162 ();
 b15zdnd11an1n32x5 FILLER_324_2226 ();
 b15zdnd11an1n16x5 FILLER_324_2258 ();
 b15zdnd00an1n02x5 FILLER_324_2274 ();
 b15zdnd11an1n64x5 FILLER_325_0 ();
 b15zdnd11an1n64x5 FILLER_325_64 ();
 b15zdnd11an1n64x5 FILLER_325_128 ();
 b15zdnd11an1n64x5 FILLER_325_192 ();
 b15zdnd11an1n16x5 FILLER_325_256 ();
 b15zdnd11an1n08x5 FILLER_325_272 ();
 b15zdnd00an1n01x5 FILLER_325_280 ();
 b15zdnd11an1n32x5 FILLER_325_323 ();
 b15zdnd11an1n08x5 FILLER_325_355 ();
 b15zdnd11an1n32x5 FILLER_325_405 ();
 b15zdnd11an1n08x5 FILLER_325_437 ();
 b15zdnd00an1n01x5 FILLER_325_445 ();
 b15zdnd11an1n32x5 FILLER_325_453 ();
 b15zdnd11an1n16x5 FILLER_325_485 ();
 b15zdnd11an1n08x5 FILLER_325_505 ();
 b15zdnd11an1n04x5 FILLER_325_513 ();
 b15zdnd11an1n04x5 FILLER_325_526 ();
 b15zdnd00an1n01x5 FILLER_325_530 ();
 b15zdnd11an1n64x5 FILLER_325_534 ();
 b15zdnd11an1n64x5 FILLER_325_598 ();
 b15zdnd11an1n32x5 FILLER_325_662 ();
 b15zdnd11an1n04x5 FILLER_325_694 ();
 b15zdnd00an1n02x5 FILLER_325_698 ();
 b15zdnd00an1n01x5 FILLER_325_700 ();
 b15zdnd11an1n04x5 FILLER_325_741 ();
 b15zdnd11an1n64x5 FILLER_325_748 ();
 b15zdnd11an1n64x5 FILLER_325_812 ();
 b15zdnd11an1n32x5 FILLER_325_876 ();
 b15zdnd11an1n04x5 FILLER_325_908 ();
 b15zdnd00an1n01x5 FILLER_325_912 ();
 b15zdnd11an1n64x5 FILLER_325_928 ();
 b15zdnd11an1n32x5 FILLER_325_992 ();
 b15zdnd00an1n02x5 FILLER_325_1024 ();
 b15zdnd00an1n01x5 FILLER_325_1026 ();
 b15zdnd11an1n16x5 FILLER_325_1041 ();
 b15zdnd11an1n04x5 FILLER_325_1057 ();
 b15zdnd00an1n02x5 FILLER_325_1061 ();
 b15zdnd11an1n04x5 FILLER_325_1078 ();
 b15zdnd11an1n64x5 FILLER_325_1090 ();
 b15zdnd11an1n64x5 FILLER_325_1154 ();
 b15zdnd11an1n16x5 FILLER_325_1218 ();
 b15zdnd11an1n04x5 FILLER_325_1234 ();
 b15zdnd00an1n02x5 FILLER_325_1238 ();
 b15zdnd11an1n16x5 FILLER_325_1251 ();
 b15zdnd11an1n04x5 FILLER_325_1267 ();
 b15zdnd00an1n01x5 FILLER_325_1271 ();
 b15zdnd11an1n64x5 FILLER_325_1282 ();
 b15zdnd11an1n64x5 FILLER_325_1346 ();
 b15zdnd11an1n64x5 FILLER_325_1410 ();
 b15zdnd11an1n16x5 FILLER_325_1474 ();
 b15zdnd00an1n02x5 FILLER_325_1490 ();
 b15zdnd11an1n64x5 FILLER_325_1497 ();
 b15zdnd11an1n64x5 FILLER_325_1561 ();
 b15zdnd11an1n64x5 FILLER_325_1625 ();
 b15zdnd11an1n64x5 FILLER_325_1689 ();
 b15zdnd11an1n64x5 FILLER_325_1753 ();
 b15zdnd11an1n64x5 FILLER_325_1817 ();
 b15zdnd11an1n32x5 FILLER_325_1881 ();
 b15zdnd11an1n08x5 FILLER_325_1913 ();
 b15zdnd00an1n02x5 FILLER_325_1921 ();
 b15zdnd00an1n01x5 FILLER_325_1923 ();
 b15zdnd11an1n04x5 FILLER_325_1927 ();
 b15zdnd11an1n64x5 FILLER_325_1934 ();
 b15zdnd11an1n32x5 FILLER_325_1998 ();
 b15zdnd11an1n08x5 FILLER_325_2030 ();
 b15zdnd11an1n04x5 FILLER_325_2038 ();
 b15zdnd00an1n02x5 FILLER_325_2042 ();
 b15zdnd11an1n04x5 FILLER_325_2054 ();
 b15zdnd11an1n08x5 FILLER_325_2064 ();
 b15zdnd00an1n01x5 FILLER_325_2072 ();
 b15zdnd11an1n64x5 FILLER_325_2085 ();
 b15zdnd11an1n64x5 FILLER_325_2149 ();
 b15zdnd11an1n64x5 FILLER_325_2213 ();
 b15zdnd11an1n04x5 FILLER_325_2277 ();
 b15zdnd00an1n02x5 FILLER_325_2281 ();
 b15zdnd00an1n01x5 FILLER_325_2283 ();
 b15zdnd11an1n64x5 FILLER_326_8 ();
 b15zdnd11an1n64x5 FILLER_326_72 ();
 b15zdnd11an1n64x5 FILLER_326_136 ();
 b15zdnd11an1n64x5 FILLER_326_200 ();
 b15zdnd11an1n16x5 FILLER_326_264 ();
 b15zdnd11an1n08x5 FILLER_326_280 ();
 b15zdnd00an1n01x5 FILLER_326_288 ();
 b15zdnd11an1n04x5 FILLER_326_307 ();
 b15zdnd11an1n64x5 FILLER_326_314 ();
 b15zdnd11an1n08x5 FILLER_326_378 ();
 b15zdnd00an1n02x5 FILLER_326_386 ();
 b15zdnd00an1n01x5 FILLER_326_388 ();
 b15zdnd11an1n04x5 FILLER_326_392 ();
 b15zdnd11an1n16x5 FILLER_326_399 ();
 b15zdnd11an1n04x5 FILLER_326_415 ();
 b15zdnd11an1n32x5 FILLER_326_461 ();
 b15zdnd11an1n04x5 FILLER_326_493 ();
 b15zdnd00an1n01x5 FILLER_326_497 ();
 b15zdnd11an1n64x5 FILLER_326_513 ();
 b15zdnd11an1n64x5 FILLER_326_577 ();
 b15zdnd11an1n64x5 FILLER_326_641 ();
 b15zdnd11an1n08x5 FILLER_326_705 ();
 b15zdnd11an1n04x5 FILLER_326_713 ();
 b15zdnd00an1n01x5 FILLER_326_717 ();
 b15zdnd11an1n04x5 FILLER_326_726 ();
 b15zdnd00an1n02x5 FILLER_326_730 ();
 b15zdnd00an1n01x5 FILLER_326_732 ();
 b15zdnd11an1n32x5 FILLER_326_736 ();
 b15zdnd11an1n16x5 FILLER_326_768 ();
 b15zdnd11an1n04x5 FILLER_326_784 ();
 b15zdnd11an1n64x5 FILLER_326_797 ();
 b15zdnd11an1n64x5 FILLER_326_861 ();
 b15zdnd11an1n64x5 FILLER_326_925 ();
 b15zdnd11an1n16x5 FILLER_326_989 ();
 b15zdnd11an1n08x5 FILLER_326_1005 ();
 b15zdnd11an1n04x5 FILLER_326_1013 ();
 b15zdnd00an1n01x5 FILLER_326_1017 ();
 b15zdnd11an1n64x5 FILLER_326_1022 ();
 b15zdnd11an1n64x5 FILLER_326_1086 ();
 b15zdnd11an1n64x5 FILLER_326_1150 ();
 b15zdnd11an1n64x5 FILLER_326_1214 ();
 b15zdnd11an1n04x5 FILLER_326_1287 ();
 b15zdnd11an1n32x5 FILLER_326_1298 ();
 b15zdnd11an1n04x5 FILLER_326_1330 ();
 b15zdnd00an1n01x5 FILLER_326_1334 ();
 b15zdnd11an1n16x5 FILLER_326_1345 ();
 b15zdnd00an1n02x5 FILLER_326_1361 ();
 b15zdnd11an1n64x5 FILLER_326_1371 ();
 b15zdnd11an1n32x5 FILLER_326_1435 ();
 b15zdnd11an1n16x5 FILLER_326_1467 ();
 b15zdnd11an1n08x5 FILLER_326_1483 ();
 b15zdnd11an1n04x5 FILLER_326_1491 ();
 b15zdnd00an1n01x5 FILLER_326_1495 ();
 b15zdnd11an1n64x5 FILLER_326_1510 ();
 b15zdnd11an1n64x5 FILLER_326_1574 ();
 b15zdnd11an1n16x5 FILLER_326_1638 ();
 b15zdnd11an1n04x5 FILLER_326_1654 ();
 b15zdnd00an1n01x5 FILLER_326_1658 ();
 b15zdnd11an1n08x5 FILLER_326_1701 ();
 b15zdnd00an1n02x5 FILLER_326_1709 ();
 b15zdnd11an1n64x5 FILLER_326_1714 ();
 b15zdnd11an1n16x5 FILLER_326_1778 ();
 b15zdnd11an1n08x5 FILLER_326_1794 ();
 b15zdnd11an1n04x5 FILLER_326_1805 ();
 b15zdnd11an1n64x5 FILLER_326_1812 ();
 b15zdnd11an1n16x5 FILLER_326_1876 ();
 b15zdnd11an1n08x5 FILLER_326_1892 ();
 b15zdnd11an1n04x5 FILLER_326_1900 ();
 b15zdnd00an1n02x5 FILLER_326_1904 ();
 b15zdnd11an1n64x5 FILLER_326_1958 ();
 b15zdnd11an1n32x5 FILLER_326_2022 ();
 b15zdnd00an1n02x5 FILLER_326_2054 ();
 b15zdnd00an1n01x5 FILLER_326_2056 ();
 b15zdnd11an1n64x5 FILLER_326_2068 ();
 b15zdnd11an1n16x5 FILLER_326_2132 ();
 b15zdnd11an1n04x5 FILLER_326_2148 ();
 b15zdnd00an1n02x5 FILLER_326_2152 ();
 b15zdnd11an1n64x5 FILLER_326_2162 ();
 b15zdnd11an1n32x5 FILLER_326_2226 ();
 b15zdnd11an1n16x5 FILLER_326_2258 ();
 b15zdnd00an1n02x5 FILLER_326_2274 ();
 b15zdnd11an1n64x5 FILLER_327_0 ();
 b15zdnd11an1n64x5 FILLER_327_64 ();
 b15zdnd11an1n64x5 FILLER_327_128 ();
 b15zdnd11an1n64x5 FILLER_327_192 ();
 b15zdnd11an1n64x5 FILLER_327_256 ();
 b15zdnd11an1n64x5 FILLER_327_320 ();
 b15zdnd11an1n64x5 FILLER_327_384 ();
 b15zdnd11an1n64x5 FILLER_327_448 ();
 b15zdnd11an1n64x5 FILLER_327_518 ();
 b15zdnd11an1n64x5 FILLER_327_582 ();
 b15zdnd11an1n64x5 FILLER_327_646 ();
 b15zdnd11an1n64x5 FILLER_327_710 ();
 b15zdnd11an1n64x5 FILLER_327_774 ();
 b15zdnd11an1n08x5 FILLER_327_838 ();
 b15zdnd11an1n04x5 FILLER_327_846 ();
 b15zdnd00an1n02x5 FILLER_327_850 ();
 b15zdnd00an1n01x5 FILLER_327_852 ();
 b15zdnd11an1n04x5 FILLER_327_859 ();
 b15zdnd11an1n16x5 FILLER_327_874 ();
 b15zdnd11an1n08x5 FILLER_327_890 ();
 b15zdnd11an1n04x5 FILLER_327_898 ();
 b15zdnd00an1n02x5 FILLER_327_902 ();
 b15zdnd00an1n01x5 FILLER_327_904 ();
 b15zdnd11an1n64x5 FILLER_327_928 ();
 b15zdnd11an1n64x5 FILLER_327_992 ();
 b15zdnd11an1n64x5 FILLER_327_1056 ();
 b15zdnd11an1n64x5 FILLER_327_1120 ();
 b15zdnd11an1n64x5 FILLER_327_1184 ();
 b15zdnd11an1n64x5 FILLER_327_1248 ();
 b15zdnd11an1n64x5 FILLER_327_1312 ();
 b15zdnd11an1n64x5 FILLER_327_1376 ();
 b15zdnd11an1n32x5 FILLER_327_1440 ();
 b15zdnd11an1n16x5 FILLER_327_1472 ();
 b15zdnd11an1n08x5 FILLER_327_1488 ();
 b15zdnd11an1n04x5 FILLER_327_1496 ();
 b15zdnd00an1n02x5 FILLER_327_1500 ();
 b15zdnd11an1n64x5 FILLER_327_1518 ();
 b15zdnd11an1n64x5 FILLER_327_1582 ();
 b15zdnd11an1n16x5 FILLER_327_1646 ();
 b15zdnd11an1n04x5 FILLER_327_1662 ();
 b15zdnd00an1n02x5 FILLER_327_1666 ();
 b15zdnd11an1n04x5 FILLER_327_1710 ();
 b15zdnd11an1n64x5 FILLER_327_1717 ();
 b15zdnd11an1n08x5 FILLER_327_1781 ();
 b15zdnd11an1n08x5 FILLER_327_1794 ();
 b15zdnd00an1n02x5 FILLER_327_1802 ();
 b15zdnd11an1n64x5 FILLER_327_1846 ();
 b15zdnd11an1n16x5 FILLER_327_1910 ();
 b15zdnd11an1n04x5 FILLER_327_1926 ();
 b15zdnd00an1n01x5 FILLER_327_1930 ();
 b15zdnd11an1n64x5 FILLER_327_1934 ();
 b15zdnd11an1n32x5 FILLER_327_1998 ();
 b15zdnd11an1n16x5 FILLER_327_2030 ();
 b15zdnd11an1n08x5 FILLER_327_2046 ();
 b15zdnd11an1n04x5 FILLER_327_2054 ();
 b15zdnd00an1n02x5 FILLER_327_2058 ();
 b15zdnd11an1n08x5 FILLER_327_2063 ();
 b15zdnd11an1n04x5 FILLER_327_2071 ();
 b15zdnd11an1n64x5 FILLER_327_2117 ();
 b15zdnd11an1n64x5 FILLER_327_2181 ();
 b15zdnd11an1n32x5 FILLER_327_2245 ();
 b15zdnd11an1n04x5 FILLER_327_2277 ();
 b15zdnd00an1n02x5 FILLER_327_2281 ();
 b15zdnd00an1n01x5 FILLER_327_2283 ();
 b15zdnd11an1n64x5 FILLER_328_8 ();
 b15zdnd11an1n64x5 FILLER_328_72 ();
 b15zdnd11an1n64x5 FILLER_328_136 ();
 b15zdnd11an1n64x5 FILLER_328_200 ();
 b15zdnd11an1n32x5 FILLER_328_264 ();
 b15zdnd11an1n08x5 FILLER_328_296 ();
 b15zdnd11an1n04x5 FILLER_328_304 ();
 b15zdnd00an1n02x5 FILLER_328_308 ();
 b15zdnd11an1n64x5 FILLER_328_316 ();
 b15zdnd11an1n64x5 FILLER_328_380 ();
 b15zdnd11an1n64x5 FILLER_328_444 ();
 b15zdnd11an1n64x5 FILLER_328_508 ();
 b15zdnd11an1n64x5 FILLER_328_572 ();
 b15zdnd11an1n64x5 FILLER_328_636 ();
 b15zdnd11an1n16x5 FILLER_328_700 ();
 b15zdnd00an1n02x5 FILLER_328_716 ();
 b15zdnd11an1n64x5 FILLER_328_726 ();
 b15zdnd11an1n64x5 FILLER_328_790 ();
 b15zdnd11an1n64x5 FILLER_328_854 ();
 b15zdnd11an1n64x5 FILLER_328_918 ();
 b15zdnd11an1n64x5 FILLER_328_982 ();
 b15zdnd11an1n16x5 FILLER_328_1046 ();
 b15zdnd11an1n08x5 FILLER_328_1062 ();
 b15zdnd11an1n04x5 FILLER_328_1070 ();
 b15zdnd00an1n02x5 FILLER_328_1074 ();
 b15zdnd00an1n01x5 FILLER_328_1076 ();
 b15zdnd11an1n64x5 FILLER_328_1102 ();
 b15zdnd11an1n16x5 FILLER_328_1166 ();
 b15zdnd00an1n01x5 FILLER_328_1182 ();
 b15zdnd11an1n32x5 FILLER_328_1195 ();
 b15zdnd11an1n08x5 FILLER_328_1227 ();
 b15zdnd11an1n04x5 FILLER_328_1235 ();
 b15zdnd00an1n01x5 FILLER_328_1239 ();
 b15zdnd11an1n64x5 FILLER_328_1252 ();
 b15zdnd11an1n64x5 FILLER_328_1316 ();
 b15zdnd11an1n64x5 FILLER_328_1380 ();
 b15zdnd11an1n32x5 FILLER_328_1444 ();
 b15zdnd11an1n16x5 FILLER_328_1476 ();
 b15zdnd11an1n04x5 FILLER_328_1492 ();
 b15zdnd11an1n64x5 FILLER_328_1507 ();
 b15zdnd11an1n64x5 FILLER_328_1571 ();
 b15zdnd11an1n32x5 FILLER_328_1635 ();
 b15zdnd11an1n16x5 FILLER_328_1667 ();
 b15zdnd00an1n02x5 FILLER_328_1683 ();
 b15zdnd00an1n01x5 FILLER_328_1685 ();
 b15zdnd11an1n32x5 FILLER_328_1738 ();
 b15zdnd11an1n08x5 FILLER_328_1770 ();
 b15zdnd00an1n01x5 FILLER_328_1778 ();
 b15zdnd11an1n64x5 FILLER_328_1831 ();
 b15zdnd11an1n64x5 FILLER_328_1895 ();
 b15zdnd11an1n64x5 FILLER_328_1959 ();
 b15zdnd11an1n32x5 FILLER_328_2023 ();
 b15zdnd00an1n02x5 FILLER_328_2055 ();
 b15zdnd00an1n01x5 FILLER_328_2057 ();
 b15zdnd11an1n32x5 FILLER_328_2100 ();
 b15zdnd11an1n16x5 FILLER_328_2132 ();
 b15zdnd11an1n04x5 FILLER_328_2148 ();
 b15zdnd00an1n02x5 FILLER_328_2152 ();
 b15zdnd11an1n64x5 FILLER_328_2162 ();
 b15zdnd11an1n32x5 FILLER_328_2226 ();
 b15zdnd11an1n16x5 FILLER_328_2258 ();
 b15zdnd00an1n02x5 FILLER_328_2274 ();
 b15zdnd11an1n64x5 FILLER_329_0 ();
 b15zdnd11an1n64x5 FILLER_329_64 ();
 b15zdnd11an1n64x5 FILLER_329_128 ();
 b15zdnd11an1n64x5 FILLER_329_192 ();
 b15zdnd11an1n64x5 FILLER_329_256 ();
 b15zdnd11an1n64x5 FILLER_329_320 ();
 b15zdnd11an1n64x5 FILLER_329_384 ();
 b15zdnd11an1n64x5 FILLER_329_448 ();
 b15zdnd11an1n64x5 FILLER_329_512 ();
 b15zdnd11an1n64x5 FILLER_329_576 ();
 b15zdnd11an1n64x5 FILLER_329_640 ();
 b15zdnd11an1n64x5 FILLER_329_704 ();
 b15zdnd11an1n08x5 FILLER_329_768 ();
 b15zdnd00an1n02x5 FILLER_329_776 ();
 b15zdnd00an1n01x5 FILLER_329_778 ();
 b15zdnd11an1n64x5 FILLER_329_831 ();
 b15zdnd11an1n08x5 FILLER_329_895 ();
 b15zdnd11an1n04x5 FILLER_329_903 ();
 b15zdnd00an1n02x5 FILLER_329_907 ();
 b15zdnd11an1n08x5 FILLER_329_922 ();
 b15zdnd11an1n04x5 FILLER_329_930 ();
 b15zdnd11an1n08x5 FILLER_329_940 ();
 b15zdnd11an1n04x5 FILLER_329_948 ();
 b15zdnd00an1n02x5 FILLER_329_952 ();
 b15zdnd00an1n01x5 FILLER_329_954 ();
 b15zdnd11an1n16x5 FILLER_329_959 ();
 b15zdnd11an1n08x5 FILLER_329_975 ();
 b15zdnd11an1n04x5 FILLER_329_983 ();
 b15zdnd00an1n02x5 FILLER_329_987 ();
 b15zdnd11an1n64x5 FILLER_329_1009 ();
 b15zdnd11an1n32x5 FILLER_329_1073 ();
 b15zdnd11an1n16x5 FILLER_329_1105 ();
 b15zdnd00an1n02x5 FILLER_329_1121 ();
 b15zdnd11an1n64x5 FILLER_329_1148 ();
 b15zdnd11an1n64x5 FILLER_329_1212 ();
 b15zdnd11an1n64x5 FILLER_329_1276 ();
 b15zdnd11an1n64x5 FILLER_329_1340 ();
 b15zdnd11an1n64x5 FILLER_329_1404 ();
 b15zdnd11an1n64x5 FILLER_329_1468 ();
 b15zdnd11an1n64x5 FILLER_329_1532 ();
 b15zdnd11an1n64x5 FILLER_329_1596 ();
 b15zdnd11an1n32x5 FILLER_329_1660 ();
 b15zdnd11an1n16x5 FILLER_329_1692 ();
 b15zdnd11an1n04x5 FILLER_329_1708 ();
 b15zdnd11an1n64x5 FILLER_329_1715 ();
 b15zdnd00an1n01x5 FILLER_329_1779 ();
 b15zdnd11an1n04x5 FILLER_329_1785 ();
 b15zdnd00an1n01x5 FILLER_329_1789 ();
 b15zdnd11an1n04x5 FILLER_329_1793 ();
 b15zdnd11an1n64x5 FILLER_329_1839 ();
 b15zdnd11an1n64x5 FILLER_329_1903 ();
 b15zdnd11an1n64x5 FILLER_329_1967 ();
 b15zdnd11an1n08x5 FILLER_329_2031 ();
 b15zdnd11an1n04x5 FILLER_329_2039 ();
 b15zdnd00an1n02x5 FILLER_329_2043 ();
 b15zdnd00an1n01x5 FILLER_329_2045 ();
 b15zdnd11an1n64x5 FILLER_329_2088 ();
 b15zdnd11an1n64x5 FILLER_329_2152 ();
 b15zdnd11an1n64x5 FILLER_329_2216 ();
 b15zdnd11an1n04x5 FILLER_329_2280 ();
 b15zdnd11an1n64x5 FILLER_330_8 ();
 b15zdnd11an1n64x5 FILLER_330_72 ();
 b15zdnd11an1n64x5 FILLER_330_136 ();
 b15zdnd11an1n16x5 FILLER_330_200 ();
 b15zdnd00an1n02x5 FILLER_330_216 ();
 b15zdnd00an1n01x5 FILLER_330_218 ();
 b15zdnd11an1n64x5 FILLER_330_223 ();
 b15zdnd11an1n64x5 FILLER_330_287 ();
 b15zdnd11an1n64x5 FILLER_330_351 ();
 b15zdnd11an1n64x5 FILLER_330_415 ();
 b15zdnd11an1n64x5 FILLER_330_479 ();
 b15zdnd11an1n64x5 FILLER_330_543 ();
 b15zdnd11an1n64x5 FILLER_330_607 ();
 b15zdnd11an1n32x5 FILLER_330_671 ();
 b15zdnd11an1n08x5 FILLER_330_703 ();
 b15zdnd11an1n04x5 FILLER_330_711 ();
 b15zdnd00an1n02x5 FILLER_330_715 ();
 b15zdnd00an1n01x5 FILLER_330_717 ();
 b15zdnd11an1n64x5 FILLER_330_726 ();
 b15zdnd11an1n08x5 FILLER_330_790 ();
 b15zdnd00an1n01x5 FILLER_330_798 ();
 b15zdnd11an1n04x5 FILLER_330_802 ();
 b15zdnd11an1n64x5 FILLER_330_809 ();
 b15zdnd11an1n16x5 FILLER_330_873 ();
 b15zdnd11an1n08x5 FILLER_330_889 ();
 b15zdnd00an1n01x5 FILLER_330_897 ();
 b15zdnd11an1n16x5 FILLER_330_917 ();
 b15zdnd11an1n16x5 FILLER_330_943 ();
 b15zdnd00an1n02x5 FILLER_330_959 ();
 b15zdnd11an1n16x5 FILLER_330_971 ();
 b15zdnd11an1n64x5 FILLER_330_991 ();
 b15zdnd11an1n64x5 FILLER_330_1055 ();
 b15zdnd11an1n64x5 FILLER_330_1119 ();
 b15zdnd11an1n64x5 FILLER_330_1183 ();
 b15zdnd11an1n64x5 FILLER_330_1247 ();
 b15zdnd11an1n64x5 FILLER_330_1311 ();
 b15zdnd11an1n64x5 FILLER_330_1375 ();
 b15zdnd11an1n32x5 FILLER_330_1439 ();
 b15zdnd11an1n16x5 FILLER_330_1471 ();
 b15zdnd11an1n08x5 FILLER_330_1487 ();
 b15zdnd00an1n02x5 FILLER_330_1495 ();
 b15zdnd00an1n01x5 FILLER_330_1497 ();
 b15zdnd11an1n04x5 FILLER_330_1504 ();
 b15zdnd11an1n64x5 FILLER_330_1515 ();
 b15zdnd11an1n64x5 FILLER_330_1579 ();
 b15zdnd11an1n32x5 FILLER_330_1643 ();
 b15zdnd00an1n01x5 FILLER_330_1675 ();
 b15zdnd11an1n64x5 FILLER_330_1694 ();
 b15zdnd11an1n08x5 FILLER_330_1758 ();
 b15zdnd11an1n04x5 FILLER_330_1766 ();
 b15zdnd11an1n04x5 FILLER_330_1774 ();
 b15zdnd11an1n04x5 FILLER_330_1789 ();
 b15zdnd11an1n64x5 FILLER_330_1835 ();
 b15zdnd11an1n08x5 FILLER_330_1899 ();
 b15zdnd11an1n04x5 FILLER_330_1907 ();
 b15zdnd00an1n01x5 FILLER_330_1911 ();
 b15zdnd11an1n16x5 FILLER_330_1915 ();
 b15zdnd00an1n01x5 FILLER_330_1931 ();
 b15zdnd11an1n64x5 FILLER_330_1974 ();
 b15zdnd11an1n64x5 FILLER_330_2038 ();
 b15zdnd11an1n32x5 FILLER_330_2102 ();
 b15zdnd11an1n16x5 FILLER_330_2134 ();
 b15zdnd11an1n04x5 FILLER_330_2150 ();
 b15zdnd11an1n64x5 FILLER_330_2162 ();
 b15zdnd11an1n32x5 FILLER_330_2226 ();
 b15zdnd11an1n16x5 FILLER_330_2258 ();
 b15zdnd00an1n02x5 FILLER_330_2274 ();
 b15zdnd11an1n64x5 FILLER_331_0 ();
 b15zdnd11an1n64x5 FILLER_331_64 ();
 b15zdnd11an1n64x5 FILLER_331_128 ();
 b15zdnd11an1n16x5 FILLER_331_192 ();
 b15zdnd00an1n02x5 FILLER_331_208 ();
 b15zdnd00an1n01x5 FILLER_331_210 ();
 b15zdnd11an1n04x5 FILLER_331_231 ();
 b15zdnd11an1n64x5 FILLER_331_266 ();
 b15zdnd11an1n64x5 FILLER_331_330 ();
 b15zdnd11an1n64x5 FILLER_331_394 ();
 b15zdnd11an1n64x5 FILLER_331_458 ();
 b15zdnd11an1n08x5 FILLER_331_522 ();
 b15zdnd00an1n01x5 FILLER_331_530 ();
 b15zdnd11an1n64x5 FILLER_331_573 ();
 b15zdnd11an1n64x5 FILLER_331_637 ();
 b15zdnd11an1n64x5 FILLER_331_701 ();
 b15zdnd11an1n32x5 FILLER_331_765 ();
 b15zdnd11an1n04x5 FILLER_331_797 ();
 b15zdnd11an1n64x5 FILLER_331_804 ();
 b15zdnd11an1n32x5 FILLER_331_868 ();
 b15zdnd11an1n08x5 FILLER_331_900 ();
 b15zdnd00an1n02x5 FILLER_331_908 ();
 b15zdnd00an1n01x5 FILLER_331_910 ();
 b15zdnd11an1n32x5 FILLER_331_921 ();
 b15zdnd11an1n08x5 FILLER_331_953 ();
 b15zdnd11an1n04x5 FILLER_331_961 ();
 b15zdnd00an1n02x5 FILLER_331_965 ();
 b15zdnd11an1n16x5 FILLER_331_976 ();
 b15zdnd00an1n02x5 FILLER_331_992 ();
 b15zdnd11an1n64x5 FILLER_331_1007 ();
 b15zdnd11an1n64x5 FILLER_331_1071 ();
 b15zdnd11an1n64x5 FILLER_331_1135 ();
 b15zdnd11an1n32x5 FILLER_331_1199 ();
 b15zdnd00an1n01x5 FILLER_331_1231 ();
 b15zdnd11an1n64x5 FILLER_331_1242 ();
 b15zdnd11an1n64x5 FILLER_331_1306 ();
 b15zdnd11an1n64x5 FILLER_331_1370 ();
 b15zdnd11an1n64x5 FILLER_331_1434 ();
 b15zdnd11an1n64x5 FILLER_331_1498 ();
 b15zdnd11an1n32x5 FILLER_331_1562 ();
 b15zdnd11an1n04x5 FILLER_331_1594 ();
 b15zdnd00an1n02x5 FILLER_331_1598 ();
 b15zdnd00an1n01x5 FILLER_331_1600 ();
 b15zdnd11an1n08x5 FILLER_331_1653 ();
 b15zdnd00an1n02x5 FILLER_331_1661 ();
 b15zdnd00an1n01x5 FILLER_331_1663 ();
 b15zdnd11an1n64x5 FILLER_331_1668 ();
 b15zdnd11an1n16x5 FILLER_331_1732 ();
 b15zdnd00an1n02x5 FILLER_331_1748 ();
 b15zdnd00an1n01x5 FILLER_331_1750 ();
 b15zdnd11an1n04x5 FILLER_331_1793 ();
 b15zdnd00an1n01x5 FILLER_331_1797 ();
 b15zdnd11an1n04x5 FILLER_331_1805 ();
 b15zdnd00an1n02x5 FILLER_331_1809 ();
 b15zdnd11an1n32x5 FILLER_331_1853 ();
 b15zdnd11an1n04x5 FILLER_331_1885 ();
 b15zdnd00an1n01x5 FILLER_331_1889 ();
 b15zdnd11an1n64x5 FILLER_331_1932 ();
 b15zdnd11an1n16x5 FILLER_331_1996 ();
 b15zdnd11an1n08x5 FILLER_331_2012 ();
 b15zdnd11an1n04x5 FILLER_331_2020 ();
 b15zdnd00an1n01x5 FILLER_331_2024 ();
 b15zdnd11an1n64x5 FILLER_331_2077 ();
 b15zdnd11an1n64x5 FILLER_331_2141 ();
 b15zdnd11an1n64x5 FILLER_331_2205 ();
 b15zdnd11an1n08x5 FILLER_331_2269 ();
 b15zdnd11an1n04x5 FILLER_331_2277 ();
 b15zdnd00an1n02x5 FILLER_331_2281 ();
 b15zdnd00an1n01x5 FILLER_331_2283 ();
 b15zdnd11an1n64x5 FILLER_332_8 ();
 b15zdnd11an1n64x5 FILLER_332_72 ();
 b15zdnd11an1n32x5 FILLER_332_136 ();
 b15zdnd11an1n16x5 FILLER_332_168 ();
 b15zdnd11an1n04x5 FILLER_332_184 ();
 b15zdnd11an1n64x5 FILLER_332_220 ();
 b15zdnd11an1n64x5 FILLER_332_284 ();
 b15zdnd11an1n64x5 FILLER_332_348 ();
 b15zdnd11an1n64x5 FILLER_332_412 ();
 b15zdnd11an1n32x5 FILLER_332_476 ();
 b15zdnd11an1n16x5 FILLER_332_508 ();
 b15zdnd11an1n08x5 FILLER_332_524 ();
 b15zdnd00an1n02x5 FILLER_332_532 ();
 b15zdnd00an1n01x5 FILLER_332_534 ();
 b15zdnd11an1n64x5 FILLER_332_577 ();
 b15zdnd11an1n64x5 FILLER_332_641 ();
 b15zdnd11an1n08x5 FILLER_332_705 ();
 b15zdnd11an1n04x5 FILLER_332_713 ();
 b15zdnd00an1n01x5 FILLER_332_717 ();
 b15zdnd11an1n64x5 FILLER_332_726 ();
 b15zdnd11an1n08x5 FILLER_332_790 ();
 b15zdnd11an1n04x5 FILLER_332_798 ();
 b15zdnd00an1n01x5 FILLER_332_802 ();
 b15zdnd11an1n64x5 FILLER_332_845 ();
 b15zdnd11an1n04x5 FILLER_332_909 ();
 b15zdnd00an1n02x5 FILLER_332_913 ();
 b15zdnd11an1n64x5 FILLER_332_919 ();
 b15zdnd11an1n64x5 FILLER_332_983 ();
 b15zdnd11an1n64x5 FILLER_332_1047 ();
 b15zdnd11an1n64x5 FILLER_332_1111 ();
 b15zdnd11an1n64x5 FILLER_332_1175 ();
 b15zdnd11an1n64x5 FILLER_332_1239 ();
 b15zdnd11an1n64x5 FILLER_332_1303 ();
 b15zdnd11an1n64x5 FILLER_332_1367 ();
 b15zdnd11an1n64x5 FILLER_332_1431 ();
 b15zdnd11an1n64x5 FILLER_332_1495 ();
 b15zdnd11an1n32x5 FILLER_332_1559 ();
 b15zdnd11an1n16x5 FILLER_332_1591 ();
 b15zdnd11an1n08x5 FILLER_332_1607 ();
 b15zdnd11an1n04x5 FILLER_332_1615 ();
 b15zdnd11an1n04x5 FILLER_332_1622 ();
 b15zdnd11an1n64x5 FILLER_332_1629 ();
 b15zdnd11an1n64x5 FILLER_332_1693 ();
 b15zdnd11an1n16x5 FILLER_332_1757 ();
 b15zdnd11an1n08x5 FILLER_332_1773 ();
 b15zdnd11an1n04x5 FILLER_332_1781 ();
 b15zdnd11an1n04x5 FILLER_332_1798 ();
 b15zdnd11an1n04x5 FILLER_332_1807 ();
 b15zdnd11an1n64x5 FILLER_332_1814 ();
 b15zdnd11an1n32x5 FILLER_332_1878 ();
 b15zdnd00an1n02x5 FILLER_332_1910 ();
 b15zdnd11an1n64x5 FILLER_332_1915 ();
 b15zdnd11an1n64x5 FILLER_332_1979 ();
 b15zdnd00an1n02x5 FILLER_332_2043 ();
 b15zdnd00an1n01x5 FILLER_332_2045 ();
 b15zdnd11an1n04x5 FILLER_332_2049 ();
 b15zdnd11an1n64x5 FILLER_332_2056 ();
 b15zdnd11an1n32x5 FILLER_332_2120 ();
 b15zdnd00an1n02x5 FILLER_332_2152 ();
 b15zdnd11an1n64x5 FILLER_332_2162 ();
 b15zdnd11an1n32x5 FILLER_332_2226 ();
 b15zdnd11an1n16x5 FILLER_332_2258 ();
 b15zdnd00an1n02x5 FILLER_332_2274 ();
 b15zdnd11an1n32x5 FILLER_333_0 ();
 b15zdnd11an1n04x5 FILLER_333_32 ();
 b15zdnd00an1n02x5 FILLER_333_36 ();
 b15zdnd11an1n64x5 FILLER_333_42 ();
 b15zdnd11an1n64x5 FILLER_333_106 ();
 b15zdnd11an1n32x5 FILLER_333_170 ();
 b15zdnd11an1n08x5 FILLER_333_202 ();
 b15zdnd11an1n04x5 FILLER_333_210 ();
 b15zdnd11an1n04x5 FILLER_333_217 ();
 b15zdnd11an1n64x5 FILLER_333_224 ();
 b15zdnd11an1n64x5 FILLER_333_288 ();
 b15zdnd11an1n64x5 FILLER_333_352 ();
 b15zdnd11an1n64x5 FILLER_333_416 ();
 b15zdnd11an1n64x5 FILLER_333_480 ();
 b15zdnd11an1n64x5 FILLER_333_544 ();
 b15zdnd11an1n64x5 FILLER_333_608 ();
 b15zdnd11an1n64x5 FILLER_333_672 ();
 b15zdnd11an1n64x5 FILLER_333_736 ();
 b15zdnd11an1n64x5 FILLER_333_800 ();
 b15zdnd11an1n32x5 FILLER_333_864 ();
 b15zdnd11an1n16x5 FILLER_333_896 ();
 b15zdnd11an1n04x5 FILLER_333_912 ();
 b15zdnd00an1n02x5 FILLER_333_916 ();
 b15zdnd00an1n01x5 FILLER_333_918 ();
 b15zdnd11an1n04x5 FILLER_333_923 ();
 b15zdnd11an1n64x5 FILLER_333_939 ();
 b15zdnd11an1n64x5 FILLER_333_1003 ();
 b15zdnd11an1n64x5 FILLER_333_1067 ();
 b15zdnd11an1n64x5 FILLER_333_1131 ();
 b15zdnd11an1n64x5 FILLER_333_1195 ();
 b15zdnd11an1n64x5 FILLER_333_1259 ();
 b15zdnd11an1n64x5 FILLER_333_1323 ();
 b15zdnd11an1n64x5 FILLER_333_1387 ();
 b15zdnd11an1n32x5 FILLER_333_1451 ();
 b15zdnd11an1n16x5 FILLER_333_1483 ();
 b15zdnd11an1n64x5 FILLER_333_1502 ();
 b15zdnd11an1n32x5 FILLER_333_1566 ();
 b15zdnd11an1n16x5 FILLER_333_1598 ();
 b15zdnd11an1n08x5 FILLER_333_1614 ();
 b15zdnd00an1n02x5 FILLER_333_1622 ();
 b15zdnd00an1n01x5 FILLER_333_1624 ();
 b15zdnd11an1n64x5 FILLER_333_1628 ();
 b15zdnd11an1n64x5 FILLER_333_1692 ();
 b15zdnd11an1n16x5 FILLER_333_1756 ();
 b15zdnd11an1n08x5 FILLER_333_1772 ();
 b15zdnd00an1n02x5 FILLER_333_1780 ();
 b15zdnd00an1n01x5 FILLER_333_1782 ();
 b15zdnd11an1n64x5 FILLER_333_1796 ();
 b15zdnd11an1n16x5 FILLER_333_1860 ();
 b15zdnd11an1n08x5 FILLER_333_1876 ();
 b15zdnd00an1n02x5 FILLER_333_1884 ();
 b15zdnd00an1n01x5 FILLER_333_1886 ();
 b15zdnd11an1n64x5 FILLER_333_1939 ();
 b15zdnd11an1n32x5 FILLER_333_2003 ();
 b15zdnd00an1n02x5 FILLER_333_2035 ();
 b15zdnd00an1n01x5 FILLER_333_2037 ();
 b15zdnd11an1n64x5 FILLER_333_2041 ();
 b15zdnd11an1n64x5 FILLER_333_2105 ();
 b15zdnd11an1n64x5 FILLER_333_2169 ();
 b15zdnd11an1n32x5 FILLER_333_2233 ();
 b15zdnd11an1n16x5 FILLER_333_2265 ();
 b15zdnd00an1n02x5 FILLER_333_2281 ();
 b15zdnd00an1n01x5 FILLER_333_2283 ();
 b15zdnd11an1n64x5 FILLER_334_8 ();
 b15zdnd11an1n64x5 FILLER_334_72 ();
 b15zdnd11an1n32x5 FILLER_334_136 ();
 b15zdnd11an1n04x5 FILLER_334_168 ();
 b15zdnd00an1n02x5 FILLER_334_172 ();
 b15zdnd11an1n04x5 FILLER_334_177 ();
 b15zdnd11an1n64x5 FILLER_334_184 ();
 b15zdnd11an1n64x5 FILLER_334_248 ();
 b15zdnd11an1n32x5 FILLER_334_312 ();
 b15zdnd11an1n16x5 FILLER_334_344 ();
 b15zdnd00an1n01x5 FILLER_334_360 ();
 b15zdnd11an1n64x5 FILLER_334_371 ();
 b15zdnd11an1n64x5 FILLER_334_435 ();
 b15zdnd11an1n64x5 FILLER_334_499 ();
 b15zdnd11an1n64x5 FILLER_334_563 ();
 b15zdnd11an1n64x5 FILLER_334_627 ();
 b15zdnd11an1n08x5 FILLER_334_691 ();
 b15zdnd00an1n02x5 FILLER_334_699 ();
 b15zdnd00an1n01x5 FILLER_334_701 ();
 b15zdnd00an1n02x5 FILLER_334_716 ();
 b15zdnd11an1n32x5 FILLER_334_726 ();
 b15zdnd11an1n16x5 FILLER_334_758 ();
 b15zdnd11an1n08x5 FILLER_334_774 ();
 b15zdnd00an1n01x5 FILLER_334_782 ();
 b15zdnd11an1n64x5 FILLER_334_786 ();
 b15zdnd11an1n64x5 FILLER_334_850 ();
 b15zdnd11an1n32x5 FILLER_334_914 ();
 b15zdnd00an1n01x5 FILLER_334_946 ();
 b15zdnd11an1n64x5 FILLER_334_963 ();
 b15zdnd11an1n08x5 FILLER_334_1027 ();
 b15zdnd00an1n01x5 FILLER_334_1035 ();
 b15zdnd11an1n64x5 FILLER_334_1078 ();
 b15zdnd11an1n64x5 FILLER_334_1142 ();
 b15zdnd11an1n64x5 FILLER_334_1206 ();
 b15zdnd11an1n64x5 FILLER_334_1270 ();
 b15zdnd11an1n64x5 FILLER_334_1334 ();
 b15zdnd11an1n64x5 FILLER_334_1398 ();
 b15zdnd11an1n16x5 FILLER_334_1462 ();
 b15zdnd11an1n08x5 FILLER_334_1478 ();
 b15zdnd11an1n04x5 FILLER_334_1486 ();
 b15zdnd00an1n01x5 FILLER_334_1490 ();
 b15zdnd11an1n16x5 FILLER_334_1494 ();
 b15zdnd11an1n04x5 FILLER_334_1510 ();
 b15zdnd00an1n01x5 FILLER_334_1514 ();
 b15zdnd11an1n64x5 FILLER_334_1519 ();
 b15zdnd11an1n64x5 FILLER_334_1583 ();
 b15zdnd11an1n64x5 FILLER_334_1647 ();
 b15zdnd11an1n64x5 FILLER_334_1711 ();
 b15zdnd11an1n64x5 FILLER_334_1775 ();
 b15zdnd11an1n64x5 FILLER_334_1839 ();
 b15zdnd11an1n08x5 FILLER_334_1903 ();
 b15zdnd00an1n01x5 FILLER_334_1911 ();
 b15zdnd11an1n64x5 FILLER_334_1915 ();
 b15zdnd11an1n64x5 FILLER_334_1979 ();
 b15zdnd11an1n64x5 FILLER_334_2043 ();
 b15zdnd11an1n32x5 FILLER_334_2107 ();
 b15zdnd11an1n08x5 FILLER_334_2139 ();
 b15zdnd11an1n04x5 FILLER_334_2147 ();
 b15zdnd00an1n02x5 FILLER_334_2151 ();
 b15zdnd00an1n01x5 FILLER_334_2153 ();
 b15zdnd11an1n64x5 FILLER_334_2162 ();
 b15zdnd11an1n32x5 FILLER_334_2226 ();
 b15zdnd11an1n16x5 FILLER_334_2258 ();
 b15zdnd00an1n02x5 FILLER_334_2274 ();
 b15zdnd11an1n64x5 FILLER_335_0 ();
 b15zdnd11an1n64x5 FILLER_335_64 ();
 b15zdnd11an1n32x5 FILLER_335_128 ();
 b15zdnd00an1n02x5 FILLER_335_160 ();
 b15zdnd00an1n01x5 FILLER_335_162 ();
 b15zdnd11an1n04x5 FILLER_335_166 ();
 b15zdnd11an1n64x5 FILLER_335_212 ();
 b15zdnd11an1n64x5 FILLER_335_276 ();
 b15zdnd11an1n64x5 FILLER_335_340 ();
 b15zdnd11an1n64x5 FILLER_335_404 ();
 b15zdnd11an1n64x5 FILLER_335_468 ();
 b15zdnd11an1n64x5 FILLER_335_532 ();
 b15zdnd11an1n64x5 FILLER_335_596 ();
 b15zdnd11an1n64x5 FILLER_335_660 ();
 b15zdnd11an1n32x5 FILLER_335_724 ();
 b15zdnd11an1n64x5 FILLER_335_808 ();
 b15zdnd11an1n32x5 FILLER_335_872 ();
 b15zdnd00an1n02x5 FILLER_335_904 ();
 b15zdnd11an1n64x5 FILLER_335_922 ();
 b15zdnd11an1n64x5 FILLER_335_986 ();
 b15zdnd11an1n08x5 FILLER_335_1050 ();
 b15zdnd11an1n04x5 FILLER_335_1058 ();
 b15zdnd11an1n16x5 FILLER_335_1107 ();
 b15zdnd11an1n08x5 FILLER_335_1123 ();
 b15zdnd11an1n04x5 FILLER_335_1131 ();
 b15zdnd11an1n64x5 FILLER_335_1160 ();
 b15zdnd11an1n64x5 FILLER_335_1224 ();
 b15zdnd11an1n64x5 FILLER_335_1288 ();
 b15zdnd11an1n64x5 FILLER_335_1352 ();
 b15zdnd11an1n32x5 FILLER_335_1416 ();
 b15zdnd11an1n16x5 FILLER_335_1448 ();
 b15zdnd00an1n02x5 FILLER_335_1464 ();
 b15zdnd11an1n04x5 FILLER_335_1518 ();
 b15zdnd11an1n64x5 FILLER_335_1564 ();
 b15zdnd11an1n64x5 FILLER_335_1628 ();
 b15zdnd11an1n64x5 FILLER_335_1692 ();
 b15zdnd11an1n32x5 FILLER_335_1756 ();
 b15zdnd11an1n08x5 FILLER_335_1788 ();
 b15zdnd11an1n64x5 FILLER_335_1806 ();
 b15zdnd11an1n64x5 FILLER_335_1870 ();
 b15zdnd11an1n64x5 FILLER_335_1934 ();
 b15zdnd11an1n64x5 FILLER_335_1998 ();
 b15zdnd11an1n64x5 FILLER_335_2062 ();
 b15zdnd11an1n64x5 FILLER_335_2126 ();
 b15zdnd11an1n64x5 FILLER_335_2190 ();
 b15zdnd11an1n16x5 FILLER_335_2254 ();
 b15zdnd11an1n08x5 FILLER_335_2270 ();
 b15zdnd11an1n04x5 FILLER_335_2278 ();
 b15zdnd00an1n02x5 FILLER_335_2282 ();
 b15zdnd11an1n64x5 FILLER_336_8 ();
 b15zdnd11an1n64x5 FILLER_336_72 ();
 b15zdnd11an1n16x5 FILLER_336_136 ();
 b15zdnd00an1n02x5 FILLER_336_152 ();
 b15zdnd11an1n64x5 FILLER_336_206 ();
 b15zdnd11an1n64x5 FILLER_336_270 ();
 b15zdnd11an1n64x5 FILLER_336_334 ();
 b15zdnd11an1n64x5 FILLER_336_398 ();
 b15zdnd11an1n64x5 FILLER_336_462 ();
 b15zdnd11an1n64x5 FILLER_336_526 ();
 b15zdnd11an1n64x5 FILLER_336_590 ();
 b15zdnd11an1n64x5 FILLER_336_654 ();
 b15zdnd11an1n04x5 FILLER_336_726 ();
 b15zdnd00an1n02x5 FILLER_336_730 ();
 b15zdnd00an1n01x5 FILLER_336_732 ();
 b15zdnd11an1n16x5 FILLER_336_758 ();
 b15zdnd11an1n04x5 FILLER_336_777 ();
 b15zdnd11an1n64x5 FILLER_336_784 ();
 b15zdnd11an1n32x5 FILLER_336_848 ();
 b15zdnd11an1n16x5 FILLER_336_880 ();
 b15zdnd11an1n08x5 FILLER_336_896 ();
 b15zdnd00an1n02x5 FILLER_336_904 ();
 b15zdnd11an1n64x5 FILLER_336_922 ();
 b15zdnd11an1n64x5 FILLER_336_986 ();
 b15zdnd11an1n64x5 FILLER_336_1050 ();
 b15zdnd11an1n64x5 FILLER_336_1114 ();
 b15zdnd11an1n64x5 FILLER_336_1178 ();
 b15zdnd11an1n64x5 FILLER_336_1242 ();
 b15zdnd11an1n32x5 FILLER_336_1306 ();
 b15zdnd11an1n08x5 FILLER_336_1338 ();
 b15zdnd00an1n02x5 FILLER_336_1346 ();
 b15zdnd11an1n64x5 FILLER_336_1390 ();
 b15zdnd11an1n16x5 FILLER_336_1454 ();
 b15zdnd11an1n08x5 FILLER_336_1470 ();
 b15zdnd11an1n04x5 FILLER_336_1478 ();
 b15zdnd00an1n02x5 FILLER_336_1482 ();
 b15zdnd11an1n04x5 FILLER_336_1487 ();
 b15zdnd11an1n08x5 FILLER_336_1494 ();
 b15zdnd00an1n02x5 FILLER_336_1502 ();
 b15zdnd00an1n01x5 FILLER_336_1504 ();
 b15zdnd11an1n64x5 FILLER_336_1510 ();
 b15zdnd11an1n64x5 FILLER_336_1574 ();
 b15zdnd11an1n64x5 FILLER_336_1638 ();
 b15zdnd11an1n64x5 FILLER_336_1702 ();
 b15zdnd11an1n64x5 FILLER_336_1766 ();
 b15zdnd11an1n64x5 FILLER_336_1830 ();
 b15zdnd11an1n64x5 FILLER_336_1894 ();
 b15zdnd11an1n64x5 FILLER_336_1958 ();
 b15zdnd11an1n64x5 FILLER_336_2022 ();
 b15zdnd11an1n64x5 FILLER_336_2086 ();
 b15zdnd11an1n04x5 FILLER_336_2150 ();
 b15zdnd11an1n64x5 FILLER_336_2162 ();
 b15zdnd11an1n32x5 FILLER_336_2226 ();
 b15zdnd11an1n16x5 FILLER_336_2258 ();
 b15zdnd00an1n02x5 FILLER_336_2274 ();
 b15zdnd11an1n64x5 FILLER_337_0 ();
 b15zdnd11an1n64x5 FILLER_337_64 ();
 b15zdnd11an1n64x5 FILLER_337_128 ();
 b15zdnd11an1n64x5 FILLER_337_192 ();
 b15zdnd11an1n64x5 FILLER_337_256 ();
 b15zdnd11an1n64x5 FILLER_337_320 ();
 b15zdnd11an1n64x5 FILLER_337_384 ();
 b15zdnd11an1n08x5 FILLER_337_448 ();
 b15zdnd11an1n04x5 FILLER_337_456 ();
 b15zdnd00an1n01x5 FILLER_337_460 ();
 b15zdnd11an1n04x5 FILLER_337_464 ();
 b15zdnd11an1n64x5 FILLER_337_473 ();
 b15zdnd11an1n64x5 FILLER_337_537 ();
 b15zdnd11an1n64x5 FILLER_337_601 ();
 b15zdnd11an1n64x5 FILLER_337_665 ();
 b15zdnd11an1n64x5 FILLER_337_729 ();
 b15zdnd11an1n64x5 FILLER_337_793 ();
 b15zdnd11an1n64x5 FILLER_337_857 ();
 b15zdnd11an1n64x5 FILLER_337_921 ();
 b15zdnd11an1n64x5 FILLER_337_985 ();
 b15zdnd11an1n32x5 FILLER_337_1049 ();
 b15zdnd11an1n16x5 FILLER_337_1081 ();
 b15zdnd11an1n04x5 FILLER_337_1097 ();
 b15zdnd00an1n02x5 FILLER_337_1101 ();
 b15zdnd11an1n32x5 FILLER_337_1128 ();
 b15zdnd00an1n01x5 FILLER_337_1160 ();
 b15zdnd11an1n64x5 FILLER_337_1192 ();
 b15zdnd11an1n32x5 FILLER_337_1256 ();
 b15zdnd11an1n08x5 FILLER_337_1288 ();
 b15zdnd00an1n02x5 FILLER_337_1296 ();
 b15zdnd00an1n01x5 FILLER_337_1298 ();
 b15zdnd11an1n64x5 FILLER_337_1341 ();
 b15zdnd11an1n64x5 FILLER_337_1405 ();
 b15zdnd11an1n32x5 FILLER_337_1469 ();
 b15zdnd11an1n64x5 FILLER_337_1514 ();
 b15zdnd11an1n64x5 FILLER_337_1578 ();
 b15zdnd11an1n64x5 FILLER_337_1642 ();
 b15zdnd11an1n64x5 FILLER_337_1706 ();
 b15zdnd11an1n64x5 FILLER_337_1770 ();
 b15zdnd11an1n32x5 FILLER_337_1834 ();
 b15zdnd11an1n08x5 FILLER_337_1866 ();
 b15zdnd11an1n04x5 FILLER_337_1874 ();
 b15zdnd00an1n01x5 FILLER_337_1878 ();
 b15zdnd11an1n64x5 FILLER_337_1921 ();
 b15zdnd11an1n64x5 FILLER_337_1985 ();
 b15zdnd11an1n64x5 FILLER_337_2049 ();
 b15zdnd11an1n64x5 FILLER_337_2113 ();
 b15zdnd11an1n64x5 FILLER_337_2177 ();
 b15zdnd11an1n32x5 FILLER_337_2241 ();
 b15zdnd11an1n08x5 FILLER_337_2273 ();
 b15zdnd00an1n02x5 FILLER_337_2281 ();
 b15zdnd00an1n01x5 FILLER_337_2283 ();
 b15zdnd11an1n64x5 FILLER_338_8 ();
 b15zdnd11an1n64x5 FILLER_338_72 ();
 b15zdnd11an1n32x5 FILLER_338_136 ();
 b15zdnd11an1n16x5 FILLER_338_168 ();
 b15zdnd11an1n08x5 FILLER_338_184 ();
 b15zdnd11an1n04x5 FILLER_338_192 ();
 b15zdnd00an1n02x5 FILLER_338_196 ();
 b15zdnd00an1n01x5 FILLER_338_198 ();
 b15zdnd11an1n64x5 FILLER_338_210 ();
 b15zdnd11an1n64x5 FILLER_338_274 ();
 b15zdnd11an1n64x5 FILLER_338_338 ();
 b15zdnd11an1n64x5 FILLER_338_402 ();
 b15zdnd11an1n32x5 FILLER_338_466 ();
 b15zdnd11an1n16x5 FILLER_338_498 ();
 b15zdnd11an1n04x5 FILLER_338_514 ();
 b15zdnd11an1n64x5 FILLER_338_521 ();
 b15zdnd11an1n64x5 FILLER_338_585 ();
 b15zdnd11an1n64x5 FILLER_338_649 ();
 b15zdnd11an1n04x5 FILLER_338_713 ();
 b15zdnd00an1n01x5 FILLER_338_717 ();
 b15zdnd11an1n64x5 FILLER_338_726 ();
 b15zdnd11an1n64x5 FILLER_338_790 ();
 b15zdnd11an1n64x5 FILLER_338_854 ();
 b15zdnd11an1n64x5 FILLER_338_918 ();
 b15zdnd11an1n64x5 FILLER_338_982 ();
 b15zdnd11an1n64x5 FILLER_338_1046 ();
 b15zdnd11an1n64x5 FILLER_338_1110 ();
 b15zdnd11an1n08x5 FILLER_338_1174 ();
 b15zdnd11an1n04x5 FILLER_338_1182 ();
 b15zdnd00an1n02x5 FILLER_338_1186 ();
 b15zdnd11an1n32x5 FILLER_338_1196 ();
 b15zdnd11an1n16x5 FILLER_338_1228 ();
 b15zdnd00an1n02x5 FILLER_338_1244 ();
 b15zdnd11an1n64x5 FILLER_338_1261 ();
 b15zdnd11an1n64x5 FILLER_338_1325 ();
 b15zdnd11an1n64x5 FILLER_338_1389 ();
 b15zdnd11an1n64x5 FILLER_338_1453 ();
 b15zdnd11an1n64x5 FILLER_338_1517 ();
 b15zdnd11an1n64x5 FILLER_338_1581 ();
 b15zdnd11an1n64x5 FILLER_338_1645 ();
 b15zdnd11an1n64x5 FILLER_338_1709 ();
 b15zdnd11an1n64x5 FILLER_338_1773 ();
 b15zdnd11an1n64x5 FILLER_338_1837 ();
 b15zdnd11an1n64x5 FILLER_338_1901 ();
 b15zdnd11an1n64x5 FILLER_338_1965 ();
 b15zdnd11an1n64x5 FILLER_338_2029 ();
 b15zdnd11an1n32x5 FILLER_338_2093 ();
 b15zdnd11an1n16x5 FILLER_338_2125 ();
 b15zdnd11an1n08x5 FILLER_338_2141 ();
 b15zdnd11an1n04x5 FILLER_338_2149 ();
 b15zdnd00an1n01x5 FILLER_338_2153 ();
 b15zdnd11an1n64x5 FILLER_338_2162 ();
 b15zdnd11an1n32x5 FILLER_338_2226 ();
 b15zdnd11an1n16x5 FILLER_338_2258 ();
 b15zdnd00an1n02x5 FILLER_338_2274 ();
 b15zdnd11an1n64x5 FILLER_339_0 ();
 b15zdnd11an1n64x5 FILLER_339_64 ();
 b15zdnd11an1n64x5 FILLER_339_128 ();
 b15zdnd11an1n64x5 FILLER_339_192 ();
 b15zdnd11an1n64x5 FILLER_339_256 ();
 b15zdnd11an1n64x5 FILLER_339_320 ();
 b15zdnd11an1n64x5 FILLER_339_384 ();
 b15zdnd11an1n32x5 FILLER_339_448 ();
 b15zdnd11an1n08x5 FILLER_339_480 ();
 b15zdnd00an1n02x5 FILLER_339_488 ();
 b15zdnd00an1n01x5 FILLER_339_490 ();
 b15zdnd11an1n64x5 FILLER_339_543 ();
 b15zdnd11an1n64x5 FILLER_339_607 ();
 b15zdnd11an1n64x5 FILLER_339_671 ();
 b15zdnd11an1n64x5 FILLER_339_735 ();
 b15zdnd11an1n64x5 FILLER_339_799 ();
 b15zdnd11an1n64x5 FILLER_339_863 ();
 b15zdnd11an1n64x5 FILLER_339_927 ();
 b15zdnd11an1n16x5 FILLER_339_991 ();
 b15zdnd11an1n64x5 FILLER_339_1011 ();
 b15zdnd11an1n64x5 FILLER_339_1075 ();
 b15zdnd11an1n32x5 FILLER_339_1139 ();
 b15zdnd11an1n04x5 FILLER_339_1171 ();
 b15zdnd11an1n32x5 FILLER_339_1191 ();
 b15zdnd11an1n16x5 FILLER_339_1223 ();
 b15zdnd11an1n08x5 FILLER_339_1239 ();
 b15zdnd11an1n04x5 FILLER_339_1247 ();
 b15zdnd11an1n32x5 FILLER_339_1257 ();
 b15zdnd11an1n08x5 FILLER_339_1289 ();
 b15zdnd00an1n01x5 FILLER_339_1297 ();
 b15zdnd11an1n64x5 FILLER_339_1310 ();
 b15zdnd11an1n16x5 FILLER_339_1374 ();
 b15zdnd11an1n64x5 FILLER_339_1405 ();
 b15zdnd11an1n64x5 FILLER_339_1469 ();
 b15zdnd11an1n64x5 FILLER_339_1533 ();
 b15zdnd11an1n64x5 FILLER_339_1597 ();
 b15zdnd11an1n64x5 FILLER_339_1661 ();
 b15zdnd11an1n64x5 FILLER_339_1725 ();
 b15zdnd11an1n64x5 FILLER_339_1789 ();
 b15zdnd11an1n32x5 FILLER_339_1853 ();
 b15zdnd11an1n08x5 FILLER_339_1885 ();
 b15zdnd00an1n02x5 FILLER_339_1893 ();
 b15zdnd00an1n01x5 FILLER_339_1895 ();
 b15zdnd11an1n64x5 FILLER_339_1938 ();
 b15zdnd11an1n64x5 FILLER_339_2002 ();
 b15zdnd11an1n64x5 FILLER_339_2066 ();
 b15zdnd11an1n64x5 FILLER_339_2130 ();
 b15zdnd11an1n64x5 FILLER_339_2194 ();
 b15zdnd11an1n16x5 FILLER_339_2258 ();
 b15zdnd11an1n08x5 FILLER_339_2274 ();
 b15zdnd00an1n02x5 FILLER_339_2282 ();
 b15zdnd11an1n64x5 FILLER_340_8 ();
 b15zdnd11an1n64x5 FILLER_340_72 ();
 b15zdnd11an1n64x5 FILLER_340_136 ();
 b15zdnd11an1n64x5 FILLER_340_200 ();
 b15zdnd11an1n64x5 FILLER_340_264 ();
 b15zdnd11an1n64x5 FILLER_340_328 ();
 b15zdnd11an1n64x5 FILLER_340_392 ();
 b15zdnd11an1n32x5 FILLER_340_456 ();
 b15zdnd11an1n16x5 FILLER_340_488 ();
 b15zdnd11an1n04x5 FILLER_340_504 ();
 b15zdnd00an1n01x5 FILLER_340_508 ();
 b15zdnd11an1n04x5 FILLER_340_512 ();
 b15zdnd11an1n64x5 FILLER_340_519 ();
 b15zdnd11an1n32x5 FILLER_340_583 ();
 b15zdnd11an1n08x5 FILLER_340_615 ();
 b15zdnd00an1n01x5 FILLER_340_623 ();
 b15zdnd11an1n04x5 FILLER_340_631 ();
 b15zdnd00an1n01x5 FILLER_340_635 ();
 b15zdnd11an1n64x5 FILLER_340_640 ();
 b15zdnd11an1n08x5 FILLER_340_704 ();
 b15zdnd11an1n04x5 FILLER_340_712 ();
 b15zdnd00an1n02x5 FILLER_340_716 ();
 b15zdnd11an1n64x5 FILLER_340_726 ();
 b15zdnd11an1n64x5 FILLER_340_790 ();
 b15zdnd11an1n64x5 FILLER_340_854 ();
 b15zdnd11an1n64x5 FILLER_340_918 ();
 b15zdnd11an1n64x5 FILLER_340_982 ();
 b15zdnd11an1n64x5 FILLER_340_1046 ();
 b15zdnd11an1n08x5 FILLER_340_1110 ();
 b15zdnd00an1n02x5 FILLER_340_1118 ();
 b15zdnd00an1n01x5 FILLER_340_1120 ();
 b15zdnd11an1n04x5 FILLER_340_1139 ();
 b15zdnd00an1n01x5 FILLER_340_1143 ();
 b15zdnd11an1n32x5 FILLER_340_1169 ();
 b15zdnd11an1n08x5 FILLER_340_1201 ();
 b15zdnd11an1n04x5 FILLER_340_1209 ();
 b15zdnd00an1n02x5 FILLER_340_1213 ();
 b15zdnd11an1n64x5 FILLER_340_1218 ();
 b15zdnd11an1n64x5 FILLER_340_1282 ();
 b15zdnd11an1n64x5 FILLER_340_1346 ();
 b15zdnd11an1n64x5 FILLER_340_1410 ();
 b15zdnd11an1n64x5 FILLER_340_1474 ();
 b15zdnd11an1n64x5 FILLER_340_1538 ();
 b15zdnd11an1n16x5 FILLER_340_1602 ();
 b15zdnd11an1n08x5 FILLER_340_1618 ();
 b15zdnd11an1n04x5 FILLER_340_1626 ();
 b15zdnd11an1n04x5 FILLER_340_1633 ();
 b15zdnd00an1n01x5 FILLER_340_1637 ();
 b15zdnd11an1n64x5 FILLER_340_1641 ();
 b15zdnd11an1n64x5 FILLER_340_1705 ();
 b15zdnd11an1n64x5 FILLER_340_1769 ();
 b15zdnd11an1n64x5 FILLER_340_1833 ();
 b15zdnd11an1n64x5 FILLER_340_1897 ();
 b15zdnd11an1n64x5 FILLER_340_1961 ();
 b15zdnd11an1n64x5 FILLER_340_2025 ();
 b15zdnd11an1n64x5 FILLER_340_2089 ();
 b15zdnd00an1n01x5 FILLER_340_2153 ();
 b15zdnd11an1n64x5 FILLER_340_2162 ();
 b15zdnd11an1n32x5 FILLER_340_2226 ();
 b15zdnd11an1n16x5 FILLER_340_2258 ();
 b15zdnd00an1n02x5 FILLER_340_2274 ();
 b15zdnd11an1n64x5 FILLER_341_0 ();
 b15zdnd11an1n64x5 FILLER_341_64 ();
 b15zdnd11an1n64x5 FILLER_341_128 ();
 b15zdnd11an1n64x5 FILLER_341_192 ();
 b15zdnd11an1n64x5 FILLER_341_256 ();
 b15zdnd11an1n64x5 FILLER_341_320 ();
 b15zdnd11an1n64x5 FILLER_341_384 ();
 b15zdnd11an1n64x5 FILLER_341_448 ();
 b15zdnd11an1n64x5 FILLER_341_512 ();
 b15zdnd11an1n32x5 FILLER_341_576 ();
 b15zdnd11an1n08x5 FILLER_341_608 ();
 b15zdnd11an1n04x5 FILLER_341_616 ();
 b15zdnd00an1n02x5 FILLER_341_620 ();
 b15zdnd11an1n08x5 FILLER_341_632 ();
 b15zdnd11an1n04x5 FILLER_341_645 ();
 b15zdnd11an1n64x5 FILLER_341_652 ();
 b15zdnd11an1n64x5 FILLER_341_716 ();
 b15zdnd11an1n64x5 FILLER_341_780 ();
 b15zdnd11an1n64x5 FILLER_341_844 ();
 b15zdnd11an1n64x5 FILLER_341_908 ();
 b15zdnd11an1n32x5 FILLER_341_972 ();
 b15zdnd00an1n02x5 FILLER_341_1004 ();
 b15zdnd11an1n16x5 FILLER_341_1030 ();
 b15zdnd11an1n08x5 FILLER_341_1046 ();
 b15zdnd11an1n04x5 FILLER_341_1054 ();
 b15zdnd00an1n02x5 FILLER_341_1058 ();
 b15zdnd00an1n01x5 FILLER_341_1060 ();
 b15zdnd11an1n64x5 FILLER_341_1068 ();
 b15zdnd11an1n64x5 FILLER_341_1132 ();
 b15zdnd11an1n64x5 FILLER_341_1196 ();
 b15zdnd11an1n32x5 FILLER_341_1260 ();
 b15zdnd11an1n08x5 FILLER_341_1292 ();
 b15zdnd11an1n04x5 FILLER_341_1300 ();
 b15zdnd00an1n02x5 FILLER_341_1304 ();
 b15zdnd00an1n01x5 FILLER_341_1306 ();
 b15zdnd11an1n64x5 FILLER_341_1325 ();
 b15zdnd11an1n64x5 FILLER_341_1389 ();
 b15zdnd11an1n64x5 FILLER_341_1453 ();
 b15zdnd11an1n64x5 FILLER_341_1517 ();
 b15zdnd11an1n16x5 FILLER_341_1581 ();
 b15zdnd00an1n02x5 FILLER_341_1597 ();
 b15zdnd11an1n08x5 FILLER_341_1639 ();
 b15zdnd00an1n02x5 FILLER_341_1647 ();
 b15zdnd11an1n64x5 FILLER_341_1658 ();
 b15zdnd11an1n64x5 FILLER_341_1722 ();
 b15zdnd11an1n64x5 FILLER_341_1786 ();
 b15zdnd11an1n64x5 FILLER_341_1850 ();
 b15zdnd11an1n64x5 FILLER_341_1914 ();
 b15zdnd11an1n64x5 FILLER_341_1978 ();
 b15zdnd11an1n64x5 FILLER_341_2042 ();
 b15zdnd11an1n64x5 FILLER_341_2106 ();
 b15zdnd11an1n64x5 FILLER_341_2170 ();
 b15zdnd11an1n32x5 FILLER_341_2234 ();
 b15zdnd11an1n16x5 FILLER_341_2266 ();
 b15zdnd00an1n02x5 FILLER_341_2282 ();
 b15zdnd11an1n64x5 FILLER_342_8 ();
 b15zdnd11an1n64x5 FILLER_342_72 ();
 b15zdnd11an1n64x5 FILLER_342_136 ();
 b15zdnd11an1n16x5 FILLER_342_200 ();
 b15zdnd11an1n64x5 FILLER_342_221 ();
 b15zdnd11an1n64x5 FILLER_342_285 ();
 b15zdnd11an1n64x5 FILLER_342_349 ();
 b15zdnd11an1n64x5 FILLER_342_413 ();
 b15zdnd11an1n64x5 FILLER_342_477 ();
 b15zdnd11an1n64x5 FILLER_342_541 ();
 b15zdnd11an1n16x5 FILLER_342_605 ();
 b15zdnd00an1n02x5 FILLER_342_621 ();
 b15zdnd11an1n04x5 FILLER_342_636 ();
 b15zdnd00an1n02x5 FILLER_342_640 ();
 b15zdnd00an1n01x5 FILLER_342_642 ();
 b15zdnd11an1n04x5 FILLER_342_652 ();
 b15zdnd11an1n32x5 FILLER_342_662 ();
 b15zdnd11an1n16x5 FILLER_342_694 ();
 b15zdnd11an1n08x5 FILLER_342_710 ();
 b15zdnd11an1n64x5 FILLER_342_726 ();
 b15zdnd11an1n64x5 FILLER_342_790 ();
 b15zdnd11an1n64x5 FILLER_342_854 ();
 b15zdnd11an1n64x5 FILLER_342_918 ();
 b15zdnd11an1n64x5 FILLER_342_982 ();
 b15zdnd11an1n32x5 FILLER_342_1046 ();
 b15zdnd11an1n08x5 FILLER_342_1078 ();
 b15zdnd00an1n01x5 FILLER_342_1086 ();
 b15zdnd11an1n04x5 FILLER_342_1090 ();
 b15zdnd11an1n64x5 FILLER_342_1101 ();
 b15zdnd11an1n64x5 FILLER_342_1165 ();
 b15zdnd11an1n64x5 FILLER_342_1229 ();
 b15zdnd11an1n08x5 FILLER_342_1293 ();
 b15zdnd11an1n32x5 FILLER_342_1325 ();
 b15zdnd11an1n16x5 FILLER_342_1357 ();
 b15zdnd11an1n08x5 FILLER_342_1373 ();
 b15zdnd00an1n02x5 FILLER_342_1381 ();
 b15zdnd00an1n01x5 FILLER_342_1383 ();
 b15zdnd11an1n64x5 FILLER_342_1394 ();
 b15zdnd11an1n64x5 FILLER_342_1458 ();
 b15zdnd11an1n64x5 FILLER_342_1522 ();
 b15zdnd11an1n64x5 FILLER_342_1586 ();
 b15zdnd11an1n64x5 FILLER_342_1650 ();
 b15zdnd11an1n64x5 FILLER_342_1714 ();
 b15zdnd11an1n64x5 FILLER_342_1778 ();
 b15zdnd11an1n64x5 FILLER_342_1842 ();
 b15zdnd11an1n64x5 FILLER_342_1906 ();
 b15zdnd11an1n64x5 FILLER_342_1970 ();
 b15zdnd11an1n64x5 FILLER_342_2034 ();
 b15zdnd11an1n32x5 FILLER_342_2098 ();
 b15zdnd11an1n16x5 FILLER_342_2130 ();
 b15zdnd11an1n08x5 FILLER_342_2146 ();
 b15zdnd11an1n64x5 FILLER_342_2162 ();
 b15zdnd11an1n32x5 FILLER_342_2226 ();
 b15zdnd11an1n16x5 FILLER_342_2258 ();
 b15zdnd00an1n02x5 FILLER_342_2274 ();
 b15zdnd11an1n64x5 FILLER_343_0 ();
 b15zdnd11an1n64x5 FILLER_343_64 ();
 b15zdnd11an1n64x5 FILLER_343_128 ();
 b15zdnd11an1n16x5 FILLER_343_192 ();
 b15zdnd11an1n08x5 FILLER_343_208 ();
 b15zdnd00an1n02x5 FILLER_343_216 ();
 b15zdnd00an1n01x5 FILLER_343_218 ();
 b15zdnd11an1n64x5 FILLER_343_261 ();
 b15zdnd11an1n64x5 FILLER_343_325 ();
 b15zdnd11an1n64x5 FILLER_343_389 ();
 b15zdnd11an1n64x5 FILLER_343_453 ();
 b15zdnd11an1n64x5 FILLER_343_517 ();
 b15zdnd11an1n16x5 FILLER_343_581 ();
 b15zdnd11an1n08x5 FILLER_343_597 ();
 b15zdnd11an1n04x5 FILLER_343_605 ();
 b15zdnd00an1n02x5 FILLER_343_609 ();
 b15zdnd11an1n04x5 FILLER_343_653 ();
 b15zdnd11an1n04x5 FILLER_343_665 ();
 b15zdnd11an1n64x5 FILLER_343_675 ();
 b15zdnd11an1n64x5 FILLER_343_739 ();
 b15zdnd11an1n64x5 FILLER_343_803 ();
 b15zdnd11an1n64x5 FILLER_343_867 ();
 b15zdnd11an1n64x5 FILLER_343_931 ();
 b15zdnd11an1n64x5 FILLER_343_995 ();
 b15zdnd00an1n01x5 FILLER_343_1059 ();
 b15zdnd11an1n64x5 FILLER_343_1112 ();
 b15zdnd11an1n64x5 FILLER_343_1176 ();
 b15zdnd11an1n32x5 FILLER_343_1240 ();
 b15zdnd11an1n04x5 FILLER_343_1272 ();
 b15zdnd00an1n02x5 FILLER_343_1276 ();
 b15zdnd00an1n01x5 FILLER_343_1278 ();
 b15zdnd11an1n04x5 FILLER_343_1297 ();
 b15zdnd11an1n64x5 FILLER_343_1311 ();
 b15zdnd11an1n64x5 FILLER_343_1375 ();
 b15zdnd11an1n64x5 FILLER_343_1439 ();
 b15zdnd11an1n64x5 FILLER_343_1503 ();
 b15zdnd11an1n64x5 FILLER_343_1567 ();
 b15zdnd11an1n64x5 FILLER_343_1631 ();
 b15zdnd11an1n64x5 FILLER_343_1695 ();
 b15zdnd11an1n32x5 FILLER_343_1759 ();
 b15zdnd11an1n04x5 FILLER_343_1791 ();
 b15zdnd00an1n01x5 FILLER_343_1795 ();
 b15zdnd11an1n08x5 FILLER_343_1800 ();
 b15zdnd11an1n04x5 FILLER_343_1808 ();
 b15zdnd00an1n01x5 FILLER_343_1812 ();
 b15zdnd11an1n64x5 FILLER_343_1816 ();
 b15zdnd11an1n16x5 FILLER_343_1880 ();
 b15zdnd11an1n04x5 FILLER_343_1896 ();
 b15zdnd00an1n02x5 FILLER_343_1900 ();
 b15zdnd11an1n64x5 FILLER_343_1907 ();
 b15zdnd11an1n64x5 FILLER_343_1971 ();
 b15zdnd11an1n64x5 FILLER_343_2035 ();
 b15zdnd11an1n64x5 FILLER_343_2099 ();
 b15zdnd11an1n64x5 FILLER_343_2163 ();
 b15zdnd11an1n32x5 FILLER_343_2227 ();
 b15zdnd11an1n16x5 FILLER_343_2259 ();
 b15zdnd11an1n08x5 FILLER_343_2275 ();
 b15zdnd00an1n01x5 FILLER_343_2283 ();
 b15zdnd11an1n64x5 FILLER_344_8 ();
 b15zdnd11an1n64x5 FILLER_344_72 ();
 b15zdnd11an1n64x5 FILLER_344_136 ();
 b15zdnd11an1n32x5 FILLER_344_200 ();
 b15zdnd11an1n08x5 FILLER_344_232 ();
 b15zdnd00an1n01x5 FILLER_344_240 ();
 b15zdnd11an1n32x5 FILLER_344_266 ();
 b15zdnd11an1n08x5 FILLER_344_298 ();
 b15zdnd00an1n02x5 FILLER_344_306 ();
 b15zdnd11an1n64x5 FILLER_344_348 ();
 b15zdnd11an1n64x5 FILLER_344_412 ();
 b15zdnd11an1n64x5 FILLER_344_476 ();
 b15zdnd11an1n64x5 FILLER_344_540 ();
 b15zdnd11an1n08x5 FILLER_344_604 ();
 b15zdnd11an1n04x5 FILLER_344_612 ();
 b15zdnd11an1n04x5 FILLER_344_658 ();
 b15zdnd11an1n08x5 FILLER_344_704 ();
 b15zdnd11an1n04x5 FILLER_344_712 ();
 b15zdnd00an1n02x5 FILLER_344_716 ();
 b15zdnd11an1n64x5 FILLER_344_726 ();
 b15zdnd11an1n64x5 FILLER_344_790 ();
 b15zdnd11an1n64x5 FILLER_344_854 ();
 b15zdnd11an1n64x5 FILLER_344_918 ();
 b15zdnd11an1n64x5 FILLER_344_982 ();
 b15zdnd11an1n32x5 FILLER_344_1046 ();
 b15zdnd11an1n04x5 FILLER_344_1078 ();
 b15zdnd00an1n02x5 FILLER_344_1082 ();
 b15zdnd00an1n01x5 FILLER_344_1084 ();
 b15zdnd11an1n64x5 FILLER_344_1088 ();
 b15zdnd11an1n64x5 FILLER_344_1152 ();
 b15zdnd11an1n64x5 FILLER_344_1216 ();
 b15zdnd11an1n16x5 FILLER_344_1280 ();
 b15zdnd11an1n08x5 FILLER_344_1296 ();
 b15zdnd00an1n02x5 FILLER_344_1304 ();
 b15zdnd00an1n01x5 FILLER_344_1306 ();
 b15zdnd11an1n64x5 FILLER_344_1326 ();
 b15zdnd11an1n64x5 FILLER_344_1390 ();
 b15zdnd11an1n64x5 FILLER_344_1454 ();
 b15zdnd11an1n64x5 FILLER_344_1518 ();
 b15zdnd11an1n64x5 FILLER_344_1582 ();
 b15zdnd11an1n64x5 FILLER_344_1646 ();
 b15zdnd11an1n64x5 FILLER_344_1710 ();
 b15zdnd11an1n04x5 FILLER_344_1774 ();
 b15zdnd11an1n64x5 FILLER_344_1818 ();
 b15zdnd11an1n64x5 FILLER_344_1882 ();
 b15zdnd11an1n64x5 FILLER_344_1946 ();
 b15zdnd11an1n08x5 FILLER_344_2010 ();
 b15zdnd11an1n04x5 FILLER_344_2018 ();
 b15zdnd00an1n02x5 FILLER_344_2022 ();
 b15zdnd11an1n04x5 FILLER_344_2027 ();
 b15zdnd11an1n04x5 FILLER_344_2034 ();
 b15zdnd11an1n64x5 FILLER_344_2041 ();
 b15zdnd11an1n32x5 FILLER_344_2105 ();
 b15zdnd11an1n16x5 FILLER_344_2137 ();
 b15zdnd00an1n01x5 FILLER_344_2153 ();
 b15zdnd11an1n64x5 FILLER_344_2162 ();
 b15zdnd11an1n32x5 FILLER_344_2226 ();
 b15zdnd11an1n16x5 FILLER_344_2258 ();
 b15zdnd00an1n02x5 FILLER_344_2274 ();
 b15zdnd11an1n64x5 FILLER_345_0 ();
 b15zdnd11an1n64x5 FILLER_345_64 ();
 b15zdnd11an1n64x5 FILLER_345_128 ();
 b15zdnd11an1n32x5 FILLER_345_192 ();
 b15zdnd11an1n16x5 FILLER_345_224 ();
 b15zdnd11an1n08x5 FILLER_345_240 ();
 b15zdnd11an1n04x5 FILLER_345_248 ();
 b15zdnd00an1n02x5 FILLER_345_252 ();
 b15zdnd00an1n01x5 FILLER_345_254 ();
 b15zdnd11an1n64x5 FILLER_345_259 ();
 b15zdnd11an1n08x5 FILLER_345_323 ();
 b15zdnd11an1n04x5 FILLER_345_331 ();
 b15zdnd00an1n02x5 FILLER_345_335 ();
 b15zdnd11an1n04x5 FILLER_345_340 ();
 b15zdnd00an1n02x5 FILLER_345_344 ();
 b15zdnd11an1n08x5 FILLER_345_349 ();
 b15zdnd11an1n08x5 FILLER_345_368 ();
 b15zdnd00an1n01x5 FILLER_345_376 ();
 b15zdnd11an1n08x5 FILLER_345_385 ();
 b15zdnd00an1n01x5 FILLER_345_393 ();
 b15zdnd11an1n64x5 FILLER_345_399 ();
 b15zdnd11an1n64x5 FILLER_345_463 ();
 b15zdnd11an1n64x5 FILLER_345_527 ();
 b15zdnd11an1n16x5 FILLER_345_591 ();
 b15zdnd11an1n08x5 FILLER_345_607 ();
 b15zdnd11an1n04x5 FILLER_345_624 ();
 b15zdnd11an1n04x5 FILLER_345_670 ();
 b15zdnd00an1n01x5 FILLER_345_674 ();
 b15zdnd11an1n04x5 FILLER_345_678 ();
 b15zdnd11an1n64x5 FILLER_345_724 ();
 b15zdnd11an1n32x5 FILLER_345_788 ();
 b15zdnd11an1n08x5 FILLER_345_820 ();
 b15zdnd00an1n02x5 FILLER_345_828 ();
 b15zdnd00an1n01x5 FILLER_345_830 ();
 b15zdnd11an1n16x5 FILLER_345_873 ();
 b15zdnd11an1n08x5 FILLER_345_889 ();
 b15zdnd11an1n04x5 FILLER_345_897 ();
 b15zdnd00an1n02x5 FILLER_345_901 ();
 b15zdnd11an1n16x5 FILLER_345_924 ();
 b15zdnd11an1n08x5 FILLER_345_940 ();
 b15zdnd00an1n02x5 FILLER_345_948 ();
 b15zdnd00an1n01x5 FILLER_345_950 ();
 b15zdnd11an1n16x5 FILLER_345_955 ();
 b15zdnd11an1n08x5 FILLER_345_971 ();
 b15zdnd00an1n01x5 FILLER_345_979 ();
 b15zdnd11an1n64x5 FILLER_345_994 ();
 b15zdnd11an1n16x5 FILLER_345_1058 ();
 b15zdnd11an1n08x5 FILLER_345_1074 ();
 b15zdnd11an1n04x5 FILLER_345_1082 ();
 b15zdnd11an1n64x5 FILLER_345_1089 ();
 b15zdnd11an1n64x5 FILLER_345_1153 ();
 b15zdnd11an1n64x5 FILLER_345_1217 ();
 b15zdnd11an1n64x5 FILLER_345_1281 ();
 b15zdnd11an1n16x5 FILLER_345_1345 ();
 b15zdnd11an1n08x5 FILLER_345_1361 ();
 b15zdnd11an1n04x5 FILLER_345_1369 ();
 b15zdnd00an1n01x5 FILLER_345_1373 ();
 b15zdnd11an1n64x5 FILLER_345_1386 ();
 b15zdnd11an1n64x5 FILLER_345_1450 ();
 b15zdnd11an1n64x5 FILLER_345_1514 ();
 b15zdnd11an1n64x5 FILLER_345_1578 ();
 b15zdnd11an1n64x5 FILLER_345_1642 ();
 b15zdnd11an1n64x5 FILLER_345_1706 ();
 b15zdnd11an1n32x5 FILLER_345_1770 ();
 b15zdnd11an1n08x5 FILLER_345_1802 ();
 b15zdnd11an1n04x5 FILLER_345_1810 ();
 b15zdnd00an1n02x5 FILLER_345_1814 ();
 b15zdnd11an1n64x5 FILLER_345_1819 ();
 b15zdnd11an1n64x5 FILLER_345_1883 ();
 b15zdnd11an1n32x5 FILLER_345_1947 ();
 b15zdnd11an1n16x5 FILLER_345_1979 ();
 b15zdnd11an1n08x5 FILLER_345_1995 ();
 b15zdnd00an1n02x5 FILLER_345_2003 ();
 b15zdnd00an1n01x5 FILLER_345_2005 ();
 b15zdnd11an1n04x5 FILLER_345_2058 ();
 b15zdnd11an1n64x5 FILLER_345_2065 ();
 b15zdnd11an1n64x5 FILLER_345_2129 ();
 b15zdnd11an1n64x5 FILLER_345_2193 ();
 b15zdnd11an1n16x5 FILLER_345_2257 ();
 b15zdnd11an1n08x5 FILLER_345_2273 ();
 b15zdnd00an1n02x5 FILLER_345_2281 ();
 b15zdnd00an1n01x5 FILLER_345_2283 ();
 b15zdnd11an1n64x5 FILLER_346_8 ();
 b15zdnd11an1n64x5 FILLER_346_72 ();
 b15zdnd11an1n64x5 FILLER_346_136 ();
 b15zdnd11an1n32x5 FILLER_346_200 ();
 b15zdnd11an1n04x5 FILLER_346_232 ();
 b15zdnd00an1n01x5 FILLER_346_236 ();
 b15zdnd11an1n04x5 FILLER_346_245 ();
 b15zdnd11an1n32x5 FILLER_346_276 ();
 b15zdnd11an1n08x5 FILLER_346_308 ();
 b15zdnd11an1n04x5 FILLER_346_316 ();
 b15zdnd00an1n02x5 FILLER_346_320 ();
 b15zdnd00an1n01x5 FILLER_346_322 ();
 b15zdnd11an1n32x5 FILLER_346_335 ();
 b15zdnd11an1n04x5 FILLER_346_367 ();
 b15zdnd00an1n02x5 FILLER_346_371 ();
 b15zdnd11an1n04x5 FILLER_346_382 ();
 b15zdnd11an1n64x5 FILLER_346_426 ();
 b15zdnd11an1n64x5 FILLER_346_490 ();
 b15zdnd11an1n64x5 FILLER_346_554 ();
 b15zdnd00an1n02x5 FILLER_346_618 ();
 b15zdnd11an1n04x5 FILLER_346_623 ();
 b15zdnd11an1n04x5 FILLER_346_669 ();
 b15zdnd00an1n02x5 FILLER_346_715 ();
 b15zdnd00an1n01x5 FILLER_346_717 ();
 b15zdnd11an1n64x5 FILLER_346_726 ();
 b15zdnd11an1n64x5 FILLER_346_790 ();
 b15zdnd11an1n08x5 FILLER_346_854 ();
 b15zdnd00an1n02x5 FILLER_346_862 ();
 b15zdnd11an1n32x5 FILLER_346_876 ();
 b15zdnd11an1n04x5 FILLER_346_908 ();
 b15zdnd00an1n02x5 FILLER_346_912 ();
 b15zdnd11an1n64x5 FILLER_346_945 ();
 b15zdnd11an1n64x5 FILLER_346_1009 ();
 b15zdnd11an1n64x5 FILLER_346_1073 ();
 b15zdnd11an1n64x5 FILLER_346_1137 ();
 b15zdnd11an1n64x5 FILLER_346_1201 ();
 b15zdnd11an1n64x5 FILLER_346_1265 ();
 b15zdnd11an1n64x5 FILLER_346_1329 ();
 b15zdnd11an1n64x5 FILLER_346_1393 ();
 b15zdnd11an1n64x5 FILLER_346_1457 ();
 b15zdnd11an1n64x5 FILLER_346_1521 ();
 b15zdnd11an1n16x5 FILLER_346_1585 ();
 b15zdnd00an1n01x5 FILLER_346_1601 ();
 b15zdnd11an1n04x5 FILLER_346_1644 ();
 b15zdnd00an1n02x5 FILLER_346_1648 ();
 b15zdnd00an1n01x5 FILLER_346_1650 ();
 b15zdnd11an1n64x5 FILLER_346_1693 ();
 b15zdnd11an1n64x5 FILLER_346_1757 ();
 b15zdnd11an1n64x5 FILLER_346_1821 ();
 b15zdnd11an1n64x5 FILLER_346_1885 ();
 b15zdnd11an1n64x5 FILLER_346_1949 ();
 b15zdnd11an1n16x5 FILLER_346_2013 ();
 b15zdnd11an1n64x5 FILLER_346_2081 ();
 b15zdnd11an1n08x5 FILLER_346_2145 ();
 b15zdnd00an1n01x5 FILLER_346_2153 ();
 b15zdnd11an1n64x5 FILLER_346_2162 ();
 b15zdnd11an1n32x5 FILLER_346_2226 ();
 b15zdnd11an1n16x5 FILLER_346_2258 ();
 b15zdnd00an1n02x5 FILLER_346_2274 ();
 b15zdnd11an1n64x5 FILLER_347_0 ();
 b15zdnd11an1n64x5 FILLER_347_64 ();
 b15zdnd11an1n64x5 FILLER_347_128 ();
 b15zdnd11an1n16x5 FILLER_347_192 ();
 b15zdnd11an1n08x5 FILLER_347_208 ();
 b15zdnd11an1n04x5 FILLER_347_216 ();
 b15zdnd00an1n02x5 FILLER_347_220 ();
 b15zdnd11an1n64x5 FILLER_347_264 ();
 b15zdnd11an1n32x5 FILLER_347_328 ();
 b15zdnd11an1n16x5 FILLER_347_360 ();
 b15zdnd11an1n08x5 FILLER_347_376 ();
 b15zdnd11an1n04x5 FILLER_347_426 ();
 b15zdnd11an1n64x5 FILLER_347_433 ();
 b15zdnd11an1n64x5 FILLER_347_497 ();
 b15zdnd11an1n32x5 FILLER_347_561 ();
 b15zdnd00an1n01x5 FILLER_347_593 ();
 b15zdnd11an1n04x5 FILLER_347_646 ();
 b15zdnd11an1n64x5 FILLER_347_702 ();
 b15zdnd11an1n64x5 FILLER_347_766 ();
 b15zdnd11an1n64x5 FILLER_347_830 ();
 b15zdnd11an1n08x5 FILLER_347_894 ();
 b15zdnd11an1n64x5 FILLER_347_916 ();
 b15zdnd11an1n64x5 FILLER_347_988 ();
 b15zdnd11an1n08x5 FILLER_347_1052 ();
 b15zdnd11an1n04x5 FILLER_347_1060 ();
 b15zdnd00an1n01x5 FILLER_347_1064 ();
 b15zdnd11an1n64x5 FILLER_347_1080 ();
 b15zdnd11an1n32x5 FILLER_347_1144 ();
 b15zdnd11an1n16x5 FILLER_347_1176 ();
 b15zdnd11an1n08x5 FILLER_347_1192 ();
 b15zdnd11an1n04x5 FILLER_347_1200 ();
 b15zdnd00an1n02x5 FILLER_347_1204 ();
 b15zdnd00an1n01x5 FILLER_347_1206 ();
 b15zdnd11an1n64x5 FILLER_347_1222 ();
 b15zdnd11an1n64x5 FILLER_347_1286 ();
 b15zdnd11an1n64x5 FILLER_347_1350 ();
 b15zdnd11an1n64x5 FILLER_347_1414 ();
 b15zdnd11an1n64x5 FILLER_347_1478 ();
 b15zdnd11an1n64x5 FILLER_347_1542 ();
 b15zdnd11an1n64x5 FILLER_347_1606 ();
 b15zdnd11an1n64x5 FILLER_347_1670 ();
 b15zdnd11an1n64x5 FILLER_347_1734 ();
 b15zdnd11an1n64x5 FILLER_347_1798 ();
 b15zdnd11an1n64x5 FILLER_347_1862 ();
 b15zdnd11an1n32x5 FILLER_347_1926 ();
 b15zdnd11an1n08x5 FILLER_347_1958 ();
 b15zdnd11an1n04x5 FILLER_347_1966 ();
 b15zdnd00an1n01x5 FILLER_347_1970 ();
 b15zdnd11an1n64x5 FILLER_347_1977 ();
 b15zdnd11an1n04x5 FILLER_347_2041 ();
 b15zdnd00an1n01x5 FILLER_347_2045 ();
 b15zdnd11an1n04x5 FILLER_347_2049 ();
 b15zdnd11an1n64x5 FILLER_347_2095 ();
 b15zdnd11an1n64x5 FILLER_347_2159 ();
 b15zdnd11an1n32x5 FILLER_347_2223 ();
 b15zdnd11an1n16x5 FILLER_347_2255 ();
 b15zdnd11an1n08x5 FILLER_347_2271 ();
 b15zdnd11an1n04x5 FILLER_347_2279 ();
 b15zdnd00an1n01x5 FILLER_347_2283 ();
 b15zdnd11an1n64x5 FILLER_348_8 ();
 b15zdnd11an1n64x5 FILLER_348_72 ();
 b15zdnd11an1n64x5 FILLER_348_136 ();
 b15zdnd11an1n16x5 FILLER_348_200 ();
 b15zdnd11an1n08x5 FILLER_348_216 ();
 b15zdnd11an1n04x5 FILLER_348_224 ();
 b15zdnd00an1n02x5 FILLER_348_228 ();
 b15zdnd11an1n08x5 FILLER_348_233 ();
 b15zdnd11an1n04x5 FILLER_348_241 ();
 b15zdnd00an1n01x5 FILLER_348_245 ();
 b15zdnd11an1n64x5 FILLER_348_288 ();
 b15zdnd11an1n32x5 FILLER_348_352 ();
 b15zdnd11an1n08x5 FILLER_348_384 ();
 b15zdnd11an1n04x5 FILLER_348_392 ();
 b15zdnd00an1n02x5 FILLER_348_396 ();
 b15zdnd00an1n01x5 FILLER_348_398 ();
 b15zdnd11an1n04x5 FILLER_348_411 ();
 b15zdnd00an1n02x5 FILLER_348_415 ();
 b15zdnd00an1n01x5 FILLER_348_417 ();
 b15zdnd11an1n64x5 FILLER_348_421 ();
 b15zdnd11an1n64x5 FILLER_348_485 ();
 b15zdnd11an1n64x5 FILLER_348_549 ();
 b15zdnd11an1n04x5 FILLER_348_616 ();
 b15zdnd11an1n08x5 FILLER_348_623 ();
 b15zdnd00an1n02x5 FILLER_348_631 ();
 b15zdnd00an1n01x5 FILLER_348_633 ();
 b15zdnd11an1n04x5 FILLER_348_640 ();
 b15zdnd00an1n01x5 FILLER_348_644 ();
 b15zdnd11an1n16x5 FILLER_348_687 ();
 b15zdnd11an1n08x5 FILLER_348_703 ();
 b15zdnd11an1n04x5 FILLER_348_711 ();
 b15zdnd00an1n02x5 FILLER_348_715 ();
 b15zdnd00an1n01x5 FILLER_348_717 ();
 b15zdnd11an1n64x5 FILLER_348_726 ();
 b15zdnd11an1n64x5 FILLER_348_790 ();
 b15zdnd11an1n32x5 FILLER_348_854 ();
 b15zdnd11an1n16x5 FILLER_348_886 ();
 b15zdnd11an1n04x5 FILLER_348_902 ();
 b15zdnd00an1n02x5 FILLER_348_906 ();
 b15zdnd00an1n01x5 FILLER_348_908 ();
 b15zdnd11an1n04x5 FILLER_348_913 ();
 b15zdnd11an1n64x5 FILLER_348_931 ();
 b15zdnd11an1n64x5 FILLER_348_995 ();
 b15zdnd11an1n64x5 FILLER_348_1059 ();
 b15zdnd11an1n64x5 FILLER_348_1123 ();
 b15zdnd11an1n32x5 FILLER_348_1187 ();
 b15zdnd11an1n04x5 FILLER_348_1219 ();
 b15zdnd11an1n64x5 FILLER_348_1226 ();
 b15zdnd11an1n08x5 FILLER_348_1290 ();
 b15zdnd11an1n64x5 FILLER_348_1316 ();
 b15zdnd11an1n64x5 FILLER_348_1380 ();
 b15zdnd11an1n64x5 FILLER_348_1444 ();
 b15zdnd11an1n64x5 FILLER_348_1508 ();
 b15zdnd11an1n64x5 FILLER_348_1572 ();
 b15zdnd11an1n64x5 FILLER_348_1636 ();
 b15zdnd11an1n32x5 FILLER_348_1700 ();
 b15zdnd00an1n01x5 FILLER_348_1732 ();
 b15zdnd11an1n04x5 FILLER_348_1736 ();
 b15zdnd11an1n32x5 FILLER_348_1743 ();
 b15zdnd11an1n16x5 FILLER_348_1775 ();
 b15zdnd11an1n04x5 FILLER_348_1791 ();
 b15zdnd00an1n02x5 FILLER_348_1795 ();
 b15zdnd00an1n01x5 FILLER_348_1797 ();
 b15zdnd11an1n64x5 FILLER_348_1802 ();
 b15zdnd11an1n16x5 FILLER_348_1866 ();
 b15zdnd11an1n08x5 FILLER_348_1882 ();
 b15zdnd11an1n04x5 FILLER_348_1890 ();
 b15zdnd00an1n01x5 FILLER_348_1894 ();
 b15zdnd11an1n64x5 FILLER_348_1898 ();
 b15zdnd11an1n64x5 FILLER_348_1962 ();
 b15zdnd11an1n16x5 FILLER_348_2026 ();
 b15zdnd11an1n08x5 FILLER_348_2042 ();
 b15zdnd11an1n04x5 FILLER_348_2050 ();
 b15zdnd11an1n64x5 FILLER_348_2057 ();
 b15zdnd11an1n32x5 FILLER_348_2121 ();
 b15zdnd00an1n01x5 FILLER_348_2153 ();
 b15zdnd11an1n64x5 FILLER_348_2162 ();
 b15zdnd11an1n32x5 FILLER_348_2226 ();
 b15zdnd11an1n16x5 FILLER_348_2258 ();
 b15zdnd00an1n02x5 FILLER_348_2274 ();
 b15zdnd11an1n64x5 FILLER_349_0 ();
 b15zdnd11an1n64x5 FILLER_349_64 ();
 b15zdnd11an1n64x5 FILLER_349_128 ();
 b15zdnd11an1n08x5 FILLER_349_192 ();
 b15zdnd00an1n02x5 FILLER_349_200 ();
 b15zdnd00an1n01x5 FILLER_349_202 ();
 b15zdnd11an1n64x5 FILLER_349_255 ();
 b15zdnd11an1n64x5 FILLER_349_319 ();
 b15zdnd11an1n16x5 FILLER_349_383 ();
 b15zdnd00an1n01x5 FILLER_349_399 ();
 b15zdnd11an1n04x5 FILLER_349_404 ();
 b15zdnd11an1n64x5 FILLER_349_411 ();
 b15zdnd11an1n64x5 FILLER_349_475 ();
 b15zdnd11an1n64x5 FILLER_349_539 ();
 b15zdnd11an1n64x5 FILLER_349_603 ();
 b15zdnd00an1n01x5 FILLER_349_667 ();
 b15zdnd11an1n04x5 FILLER_349_671 ();
 b15zdnd11an1n64x5 FILLER_349_678 ();
 b15zdnd11an1n64x5 FILLER_349_742 ();
 b15zdnd11an1n64x5 FILLER_349_806 ();
 b15zdnd11an1n64x5 FILLER_349_870 ();
 b15zdnd11an1n64x5 FILLER_349_934 ();
 b15zdnd11an1n64x5 FILLER_349_998 ();
 b15zdnd11an1n64x5 FILLER_349_1062 ();
 b15zdnd11an1n64x5 FILLER_349_1126 ();
 b15zdnd11an1n32x5 FILLER_349_1190 ();
 b15zdnd11an1n64x5 FILLER_349_1246 ();
 b15zdnd11an1n64x5 FILLER_349_1310 ();
 b15zdnd11an1n64x5 FILLER_349_1374 ();
 b15zdnd11an1n64x5 FILLER_349_1438 ();
 b15zdnd11an1n64x5 FILLER_349_1502 ();
 b15zdnd11an1n64x5 FILLER_349_1566 ();
 b15zdnd11an1n64x5 FILLER_349_1630 ();
 b15zdnd11an1n16x5 FILLER_349_1694 ();
 b15zdnd11an1n04x5 FILLER_349_1710 ();
 b15zdnd00an1n01x5 FILLER_349_1714 ();
 b15zdnd11an1n64x5 FILLER_349_1767 ();
 b15zdnd11an1n64x5 FILLER_349_1831 ();
 b15zdnd11an1n16x5 FILLER_349_1898 ();
 b15zdnd11an1n08x5 FILLER_349_1914 ();
 b15zdnd11an1n04x5 FILLER_349_1922 ();
 b15zdnd00an1n02x5 FILLER_349_1926 ();
 b15zdnd11an1n64x5 FILLER_349_1959 ();
 b15zdnd11an1n64x5 FILLER_349_2023 ();
 b15zdnd11an1n64x5 FILLER_349_2087 ();
 b15zdnd11an1n64x5 FILLER_349_2151 ();
 b15zdnd11an1n64x5 FILLER_349_2215 ();
 b15zdnd11an1n04x5 FILLER_349_2279 ();
 b15zdnd00an1n01x5 FILLER_349_2283 ();
 b15zdnd11an1n64x5 FILLER_350_8 ();
 b15zdnd11an1n64x5 FILLER_350_72 ();
 b15zdnd11an1n64x5 FILLER_350_136 ();
 b15zdnd11an1n16x5 FILLER_350_200 ();
 b15zdnd11an1n04x5 FILLER_350_216 ();
 b15zdnd00an1n01x5 FILLER_350_220 ();
 b15zdnd11an1n04x5 FILLER_350_224 ();
 b15zdnd11an1n64x5 FILLER_350_231 ();
 b15zdnd11an1n64x5 FILLER_350_295 ();
 b15zdnd11an1n64x5 FILLER_350_359 ();
 b15zdnd11an1n64x5 FILLER_350_423 ();
 b15zdnd11an1n16x5 FILLER_350_487 ();
 b15zdnd11an1n08x5 FILLER_350_503 ();
 b15zdnd11an1n04x5 FILLER_350_511 ();
 b15zdnd00an1n02x5 FILLER_350_515 ();
 b15zdnd00an1n01x5 FILLER_350_517 ();
 b15zdnd11an1n64x5 FILLER_350_521 ();
 b15zdnd11an1n64x5 FILLER_350_585 ();
 b15zdnd11an1n64x5 FILLER_350_649 ();
 b15zdnd11an1n04x5 FILLER_350_713 ();
 b15zdnd00an1n01x5 FILLER_350_717 ();
 b15zdnd11an1n64x5 FILLER_350_726 ();
 b15zdnd11an1n64x5 FILLER_350_790 ();
 b15zdnd11an1n64x5 FILLER_350_854 ();
 b15zdnd11an1n04x5 FILLER_350_918 ();
 b15zdnd11an1n64x5 FILLER_350_926 ();
 b15zdnd11an1n64x5 FILLER_350_990 ();
 b15zdnd11an1n64x5 FILLER_350_1054 ();
 b15zdnd11an1n64x5 FILLER_350_1118 ();
 b15zdnd11an1n64x5 FILLER_350_1182 ();
 b15zdnd11an1n64x5 FILLER_350_1246 ();
 b15zdnd11an1n32x5 FILLER_350_1310 ();
 b15zdnd11an1n16x5 FILLER_350_1342 ();
 b15zdnd11an1n08x5 FILLER_350_1358 ();
 b15zdnd11an1n04x5 FILLER_350_1366 ();
 b15zdnd11an1n64x5 FILLER_350_1385 ();
 b15zdnd11an1n64x5 FILLER_350_1449 ();
 b15zdnd11an1n64x5 FILLER_350_1513 ();
 b15zdnd11an1n64x5 FILLER_350_1577 ();
 b15zdnd11an1n64x5 FILLER_350_1641 ();
 b15zdnd11an1n32x5 FILLER_350_1705 ();
 b15zdnd00an1n02x5 FILLER_350_1737 ();
 b15zdnd00an1n01x5 FILLER_350_1739 ();
 b15zdnd11an1n64x5 FILLER_350_1743 ();
 b15zdnd11an1n32x5 FILLER_350_1807 ();
 b15zdnd11an1n16x5 FILLER_350_1839 ();
 b15zdnd11an1n08x5 FILLER_350_1855 ();
 b15zdnd11an1n04x5 FILLER_350_1863 ();
 b15zdnd00an1n02x5 FILLER_350_1867 ();
 b15zdnd00an1n01x5 FILLER_350_1869 ();
 b15zdnd11an1n04x5 FILLER_350_1922 ();
 b15zdnd11an1n64x5 FILLER_350_1968 ();
 b15zdnd11an1n64x5 FILLER_350_2032 ();
 b15zdnd11an1n32x5 FILLER_350_2096 ();
 b15zdnd11an1n16x5 FILLER_350_2128 ();
 b15zdnd11an1n08x5 FILLER_350_2144 ();
 b15zdnd00an1n02x5 FILLER_350_2152 ();
 b15zdnd11an1n64x5 FILLER_350_2162 ();
 b15zdnd11an1n32x5 FILLER_350_2226 ();
 b15zdnd11an1n16x5 FILLER_350_2258 ();
 b15zdnd00an1n02x5 FILLER_350_2274 ();
 b15zdnd11an1n64x5 FILLER_351_0 ();
 b15zdnd11an1n64x5 FILLER_351_64 ();
 b15zdnd11an1n64x5 FILLER_351_128 ();
 b15zdnd11an1n64x5 FILLER_351_192 ();
 b15zdnd11an1n64x5 FILLER_351_256 ();
 b15zdnd11an1n64x5 FILLER_351_320 ();
 b15zdnd11an1n64x5 FILLER_351_384 ();
 b15zdnd11an1n32x5 FILLER_351_448 ();
 b15zdnd11an1n08x5 FILLER_351_480 ();
 b15zdnd00an1n02x5 FILLER_351_488 ();
 b15zdnd00an1n01x5 FILLER_351_490 ();
 b15zdnd11an1n64x5 FILLER_351_543 ();
 b15zdnd11an1n64x5 FILLER_351_607 ();
 b15zdnd11an1n64x5 FILLER_351_671 ();
 b15zdnd11an1n64x5 FILLER_351_735 ();
 b15zdnd11an1n64x5 FILLER_351_799 ();
 b15zdnd11an1n64x5 FILLER_351_863 ();
 b15zdnd11an1n64x5 FILLER_351_927 ();
 b15zdnd11an1n64x5 FILLER_351_991 ();
 b15zdnd11an1n64x5 FILLER_351_1055 ();
 b15zdnd11an1n64x5 FILLER_351_1119 ();
 b15zdnd11an1n32x5 FILLER_351_1183 ();
 b15zdnd11an1n04x5 FILLER_351_1215 ();
 b15zdnd00an1n02x5 FILLER_351_1219 ();
 b15zdnd00an1n01x5 FILLER_351_1221 ();
 b15zdnd11an1n64x5 FILLER_351_1237 ();
 b15zdnd11an1n64x5 FILLER_351_1301 ();
 b15zdnd11an1n64x5 FILLER_351_1365 ();
 b15zdnd11an1n64x5 FILLER_351_1429 ();
 b15zdnd11an1n64x5 FILLER_351_1493 ();
 b15zdnd11an1n64x5 FILLER_351_1557 ();
 b15zdnd11an1n16x5 FILLER_351_1621 ();
 b15zdnd11an1n04x5 FILLER_351_1637 ();
 b15zdnd11an1n64x5 FILLER_351_1693 ();
 b15zdnd11an1n64x5 FILLER_351_1757 ();
 b15zdnd11an1n64x5 FILLER_351_1821 ();
 b15zdnd11an1n08x5 FILLER_351_1885 ();
 b15zdnd00an1n02x5 FILLER_351_1893 ();
 b15zdnd00an1n01x5 FILLER_351_1895 ();
 b15zdnd11an1n32x5 FILLER_351_1899 ();
 b15zdnd11an1n16x5 FILLER_351_1931 ();
 b15zdnd00an1n02x5 FILLER_351_1947 ();
 b15zdnd00an1n01x5 FILLER_351_1949 ();
 b15zdnd11an1n04x5 FILLER_351_1959 ();
 b15zdnd11an1n64x5 FILLER_351_1979 ();
 b15zdnd11an1n64x5 FILLER_351_2043 ();
 b15zdnd11an1n64x5 FILLER_351_2107 ();
 b15zdnd11an1n64x5 FILLER_351_2171 ();
 b15zdnd11an1n32x5 FILLER_351_2235 ();
 b15zdnd11an1n16x5 FILLER_351_2267 ();
 b15zdnd00an1n01x5 FILLER_351_2283 ();
 b15zdnd11an1n64x5 FILLER_352_8 ();
 b15zdnd11an1n64x5 FILLER_352_72 ();
 b15zdnd11an1n64x5 FILLER_352_136 ();
 b15zdnd11an1n64x5 FILLER_352_200 ();
 b15zdnd11an1n64x5 FILLER_352_264 ();
 b15zdnd11an1n64x5 FILLER_352_328 ();
 b15zdnd11an1n08x5 FILLER_352_392 ();
 b15zdnd00an1n02x5 FILLER_352_400 ();
 b15zdnd11an1n64x5 FILLER_352_414 ();
 b15zdnd11an1n16x5 FILLER_352_478 ();
 b15zdnd11an1n08x5 FILLER_352_494 ();
 b15zdnd11an1n04x5 FILLER_352_502 ();
 b15zdnd00an1n02x5 FILLER_352_506 ();
 b15zdnd00an1n01x5 FILLER_352_508 ();
 b15zdnd11an1n04x5 FILLER_352_512 ();
 b15zdnd11an1n64x5 FILLER_352_519 ();
 b15zdnd11an1n64x5 FILLER_352_583 ();
 b15zdnd11an1n64x5 FILLER_352_647 ();
 b15zdnd11an1n04x5 FILLER_352_711 ();
 b15zdnd00an1n02x5 FILLER_352_715 ();
 b15zdnd00an1n01x5 FILLER_352_717 ();
 b15zdnd11an1n32x5 FILLER_352_726 ();
 b15zdnd11an1n16x5 FILLER_352_758 ();
 b15zdnd11an1n08x5 FILLER_352_774 ();
 b15zdnd11an1n04x5 FILLER_352_782 ();
 b15zdnd00an1n02x5 FILLER_352_786 ();
 b15zdnd11an1n64x5 FILLER_352_791 ();
 b15zdnd11an1n64x5 FILLER_352_855 ();
 b15zdnd11an1n64x5 FILLER_352_919 ();
 b15zdnd11an1n32x5 FILLER_352_983 ();
 b15zdnd11an1n16x5 FILLER_352_1015 ();
 b15zdnd11an1n08x5 FILLER_352_1031 ();
 b15zdnd11an1n04x5 FILLER_352_1039 ();
 b15zdnd00an1n01x5 FILLER_352_1043 ();
 b15zdnd11an1n32x5 FILLER_352_1075 ();
 b15zdnd11an1n16x5 FILLER_352_1107 ();
 b15zdnd11an1n08x5 FILLER_352_1123 ();
 b15zdnd00an1n02x5 FILLER_352_1131 ();
 b15zdnd11an1n64x5 FILLER_352_1147 ();
 b15zdnd11an1n64x5 FILLER_352_1211 ();
 b15zdnd11an1n64x5 FILLER_352_1275 ();
 b15zdnd11an1n64x5 FILLER_352_1339 ();
 b15zdnd11an1n64x5 FILLER_352_1403 ();
 b15zdnd11an1n64x5 FILLER_352_1467 ();
 b15zdnd11an1n64x5 FILLER_352_1531 ();
 b15zdnd11an1n32x5 FILLER_352_1595 ();
 b15zdnd11an1n16x5 FILLER_352_1627 ();
 b15zdnd11an1n08x5 FILLER_352_1643 ();
 b15zdnd11an1n04x5 FILLER_352_1651 ();
 b15zdnd00an1n02x5 FILLER_352_1655 ();
 b15zdnd11an1n04x5 FILLER_352_1699 ();
 b15zdnd11an1n64x5 FILLER_352_1717 ();
 b15zdnd11an1n64x5 FILLER_352_1781 ();
 b15zdnd11an1n64x5 FILLER_352_1845 ();
 b15zdnd11an1n64x5 FILLER_352_1909 ();
 b15zdnd11an1n64x5 FILLER_352_1973 ();
 b15zdnd11an1n64x5 FILLER_352_2037 ();
 b15zdnd11an1n32x5 FILLER_352_2101 ();
 b15zdnd11an1n16x5 FILLER_352_2133 ();
 b15zdnd11an1n04x5 FILLER_352_2149 ();
 b15zdnd00an1n01x5 FILLER_352_2153 ();
 b15zdnd11an1n64x5 FILLER_352_2162 ();
 b15zdnd11an1n32x5 FILLER_352_2226 ();
 b15zdnd11an1n16x5 FILLER_352_2258 ();
 b15zdnd00an1n02x5 FILLER_352_2274 ();
 b15zdnd11an1n64x5 FILLER_353_0 ();
 b15zdnd11an1n64x5 FILLER_353_64 ();
 b15zdnd11an1n64x5 FILLER_353_128 ();
 b15zdnd11an1n64x5 FILLER_353_192 ();
 b15zdnd11an1n64x5 FILLER_353_256 ();
 b15zdnd11an1n64x5 FILLER_353_320 ();
 b15zdnd11an1n16x5 FILLER_353_384 ();
 b15zdnd11an1n04x5 FILLER_353_400 ();
 b15zdnd00an1n02x5 FILLER_353_404 ();
 b15zdnd00an1n01x5 FILLER_353_406 ();
 b15zdnd11an1n64x5 FILLER_353_412 ();
 b15zdnd11an1n64x5 FILLER_353_476 ();
 b15zdnd11an1n64x5 FILLER_353_540 ();
 b15zdnd11an1n64x5 FILLER_353_604 ();
 b15zdnd11an1n64x5 FILLER_353_668 ();
 b15zdnd11an1n16x5 FILLER_353_732 ();
 b15zdnd11an1n04x5 FILLER_353_748 ();
 b15zdnd11an1n64x5 FILLER_353_792 ();
 b15zdnd11an1n16x5 FILLER_353_856 ();
 b15zdnd11an1n04x5 FILLER_353_872 ();
 b15zdnd00an1n02x5 FILLER_353_876 ();
 b15zdnd11an1n04x5 FILLER_353_882 ();
 b15zdnd11an1n08x5 FILLER_353_895 ();
 b15zdnd11an1n04x5 FILLER_353_903 ();
 b15zdnd00an1n02x5 FILLER_353_907 ();
 b15zdnd11an1n32x5 FILLER_353_913 ();
 b15zdnd11an1n08x5 FILLER_353_945 ();
 b15zdnd00an1n02x5 FILLER_353_953 ();
 b15zdnd00an1n01x5 FILLER_353_955 ();
 b15zdnd11an1n64x5 FILLER_353_981 ();
 b15zdnd11an1n16x5 FILLER_353_1045 ();
 b15zdnd11an1n08x5 FILLER_353_1061 ();
 b15zdnd11an1n64x5 FILLER_353_1100 ();
 b15zdnd00an1n02x5 FILLER_353_1164 ();
 b15zdnd11an1n16x5 FILLER_353_1192 ();
 b15zdnd00an1n02x5 FILLER_353_1208 ();
 b15zdnd00an1n01x5 FILLER_353_1210 ();
 b15zdnd11an1n04x5 FILLER_353_1222 ();
 b15zdnd11an1n64x5 FILLER_353_1235 ();
 b15zdnd11an1n08x5 FILLER_353_1299 ();
 b15zdnd11an1n04x5 FILLER_353_1307 ();
 b15zdnd00an1n01x5 FILLER_353_1311 ();
 b15zdnd11an1n64x5 FILLER_353_1354 ();
 b15zdnd11an1n64x5 FILLER_353_1418 ();
 b15zdnd11an1n64x5 FILLER_353_1482 ();
 b15zdnd11an1n64x5 FILLER_353_1546 ();
 b15zdnd11an1n32x5 FILLER_353_1610 ();
 b15zdnd11an1n16x5 FILLER_353_1642 ();
 b15zdnd00an1n02x5 FILLER_353_1658 ();
 b15zdnd11an1n04x5 FILLER_353_1663 ();
 b15zdnd11an1n04x5 FILLER_353_1670 ();
 b15zdnd11an1n64x5 FILLER_353_1677 ();
 b15zdnd11an1n32x5 FILLER_353_1741 ();
 b15zdnd11an1n16x5 FILLER_353_1773 ();
 b15zdnd11an1n08x5 FILLER_353_1789 ();
 b15zdnd00an1n02x5 FILLER_353_1797 ();
 b15zdnd11an1n64x5 FILLER_353_1841 ();
 b15zdnd11an1n64x5 FILLER_353_1905 ();
 b15zdnd11an1n64x5 FILLER_353_1979 ();
 b15zdnd11an1n64x5 FILLER_353_2043 ();
 b15zdnd11an1n64x5 FILLER_353_2107 ();
 b15zdnd11an1n64x5 FILLER_353_2171 ();
 b15zdnd11an1n32x5 FILLER_353_2235 ();
 b15zdnd11an1n16x5 FILLER_353_2267 ();
 b15zdnd00an1n01x5 FILLER_353_2283 ();
 b15zdnd00an1n02x5 FILLER_354_8 ();
 b15zdnd11an1n64x5 FILLER_354_15 ();
 b15zdnd11an1n64x5 FILLER_354_79 ();
 b15zdnd11an1n64x5 FILLER_354_143 ();
 b15zdnd11an1n64x5 FILLER_354_207 ();
 b15zdnd11an1n64x5 FILLER_354_271 ();
 b15zdnd11an1n64x5 FILLER_354_335 ();
 b15zdnd11an1n64x5 FILLER_354_399 ();
 b15zdnd11an1n64x5 FILLER_354_463 ();
 b15zdnd11an1n64x5 FILLER_354_527 ();
 b15zdnd11an1n64x5 FILLER_354_591 ();
 b15zdnd11an1n32x5 FILLER_354_655 ();
 b15zdnd11an1n16x5 FILLER_354_687 ();
 b15zdnd11an1n08x5 FILLER_354_703 ();
 b15zdnd11an1n04x5 FILLER_354_711 ();
 b15zdnd00an1n02x5 FILLER_354_715 ();
 b15zdnd00an1n01x5 FILLER_354_717 ();
 b15zdnd11an1n32x5 FILLER_354_726 ();
 b15zdnd11an1n16x5 FILLER_354_758 ();
 b15zdnd11an1n08x5 FILLER_354_774 ();
 b15zdnd11an1n04x5 FILLER_354_782 ();
 b15zdnd00an1n02x5 FILLER_354_786 ();
 b15zdnd11an1n64x5 FILLER_354_791 ();
 b15zdnd11an1n32x5 FILLER_354_855 ();
 b15zdnd11an1n16x5 FILLER_354_887 ();
 b15zdnd11an1n64x5 FILLER_354_922 ();
 b15zdnd11an1n64x5 FILLER_354_986 ();
 b15zdnd11an1n32x5 FILLER_354_1050 ();
 b15zdnd11an1n04x5 FILLER_354_1082 ();
 b15zdnd00an1n02x5 FILLER_354_1086 ();
 b15zdnd00an1n01x5 FILLER_354_1088 ();
 b15zdnd11an1n64x5 FILLER_354_1114 ();
 b15zdnd11an1n32x5 FILLER_354_1178 ();
 b15zdnd11an1n16x5 FILLER_354_1210 ();
 b15zdnd00an1n02x5 FILLER_354_1226 ();
 b15zdnd11an1n08x5 FILLER_354_1252 ();
 b15zdnd00an1n02x5 FILLER_354_1260 ();
 b15zdnd00an1n01x5 FILLER_354_1262 ();
 b15zdnd11an1n64x5 FILLER_354_1305 ();
 b15zdnd11an1n32x5 FILLER_354_1369 ();
 b15zdnd11an1n08x5 FILLER_354_1401 ();
 b15zdnd11an1n04x5 FILLER_354_1409 ();
 b15zdnd11an1n04x5 FILLER_354_1416 ();
 b15zdnd11an1n64x5 FILLER_354_1423 ();
 b15zdnd11an1n32x5 FILLER_354_1487 ();
 b15zdnd11an1n16x5 FILLER_354_1519 ();
 b15zdnd11an1n08x5 FILLER_354_1535 ();
 b15zdnd00an1n01x5 FILLER_354_1543 ();
 b15zdnd11an1n64x5 FILLER_354_1553 ();
 b15zdnd11an1n64x5 FILLER_354_1617 ();
 b15zdnd11an1n64x5 FILLER_354_1681 ();
 b15zdnd11an1n64x5 FILLER_354_1745 ();
 b15zdnd11an1n64x5 FILLER_354_1809 ();
 b15zdnd11an1n64x5 FILLER_354_1873 ();
 b15zdnd11an1n08x5 FILLER_354_1937 ();
 b15zdnd00an1n02x5 FILLER_354_1945 ();
 b15zdnd11an1n04x5 FILLER_354_1950 ();
 b15zdnd00an1n02x5 FILLER_354_1954 ();
 b15zdnd00an1n01x5 FILLER_354_1956 ();
 b15zdnd11an1n64x5 FILLER_354_1972 ();
 b15zdnd11an1n64x5 FILLER_354_2036 ();
 b15zdnd11an1n32x5 FILLER_354_2100 ();
 b15zdnd11an1n16x5 FILLER_354_2132 ();
 b15zdnd11an1n04x5 FILLER_354_2148 ();
 b15zdnd00an1n02x5 FILLER_354_2152 ();
 b15zdnd11an1n64x5 FILLER_354_2162 ();
 b15zdnd11an1n32x5 FILLER_354_2226 ();
 b15zdnd11an1n16x5 FILLER_354_2258 ();
 b15zdnd00an1n02x5 FILLER_354_2274 ();
 b15zdnd11an1n64x5 FILLER_355_0 ();
 b15zdnd11an1n64x5 FILLER_355_64 ();
 b15zdnd11an1n64x5 FILLER_355_128 ();
 b15zdnd11an1n64x5 FILLER_355_192 ();
 b15zdnd11an1n64x5 FILLER_355_256 ();
 b15zdnd11an1n64x5 FILLER_355_320 ();
 b15zdnd11an1n08x5 FILLER_355_384 ();
 b15zdnd11an1n04x5 FILLER_355_392 ();
 b15zdnd00an1n02x5 FILLER_355_396 ();
 b15zdnd11an1n64x5 FILLER_355_440 ();
 b15zdnd11an1n64x5 FILLER_355_504 ();
 b15zdnd11an1n64x5 FILLER_355_568 ();
 b15zdnd11an1n64x5 FILLER_355_632 ();
 b15zdnd11an1n64x5 FILLER_355_696 ();
 b15zdnd11an1n64x5 FILLER_355_760 ();
 b15zdnd11an1n32x5 FILLER_355_824 ();
 b15zdnd11an1n16x5 FILLER_355_856 ();
 b15zdnd11an1n08x5 FILLER_355_872 ();
 b15zdnd00an1n02x5 FILLER_355_880 ();
 b15zdnd00an1n01x5 FILLER_355_882 ();
 b15zdnd11an1n04x5 FILLER_355_914 ();
 b15zdnd11an1n04x5 FILLER_355_935 ();
 b15zdnd11an1n64x5 FILLER_355_954 ();
 b15zdnd11an1n64x5 FILLER_355_1018 ();
 b15zdnd11an1n16x5 FILLER_355_1082 ();
 b15zdnd11an1n04x5 FILLER_355_1098 ();
 b15zdnd00an1n01x5 FILLER_355_1102 ();
 b15zdnd11an1n64x5 FILLER_355_1128 ();
 b15zdnd11an1n64x5 FILLER_355_1192 ();
 b15zdnd11an1n64x5 FILLER_355_1256 ();
 b15zdnd11an1n32x5 FILLER_355_1320 ();
 b15zdnd11an1n08x5 FILLER_355_1352 ();
 b15zdnd11an1n04x5 FILLER_355_1360 ();
 b15zdnd00an1n02x5 FILLER_355_1364 ();
 b15zdnd00an1n01x5 FILLER_355_1366 ();
 b15zdnd11an1n08x5 FILLER_355_1392 ();
 b15zdnd11an1n04x5 FILLER_355_1400 ();
 b15zdnd11an1n64x5 FILLER_355_1446 ();
 b15zdnd11an1n64x5 FILLER_355_1510 ();
 b15zdnd11an1n64x5 FILLER_355_1574 ();
 b15zdnd11an1n64x5 FILLER_355_1638 ();
 b15zdnd11an1n64x5 FILLER_355_1702 ();
 b15zdnd11an1n32x5 FILLER_355_1766 ();
 b15zdnd11an1n16x5 FILLER_355_1798 ();
 b15zdnd11an1n08x5 FILLER_355_1814 ();
 b15zdnd11an1n04x5 FILLER_355_1825 ();
 b15zdnd11an1n64x5 FILLER_355_1832 ();
 b15zdnd11an1n64x5 FILLER_355_1896 ();
 b15zdnd00an1n02x5 FILLER_355_1960 ();
 b15zdnd11an1n64x5 FILLER_355_1975 ();
 b15zdnd11an1n64x5 FILLER_355_2039 ();
 b15zdnd11an1n64x5 FILLER_355_2103 ();
 b15zdnd11an1n64x5 FILLER_355_2167 ();
 b15zdnd11an1n32x5 FILLER_355_2231 ();
 b15zdnd11an1n16x5 FILLER_355_2263 ();
 b15zdnd11an1n04x5 FILLER_355_2279 ();
 b15zdnd00an1n01x5 FILLER_355_2283 ();
 b15zdnd11an1n64x5 FILLER_356_8 ();
 b15zdnd11an1n64x5 FILLER_356_72 ();
 b15zdnd11an1n64x5 FILLER_356_136 ();
 b15zdnd11an1n64x5 FILLER_356_200 ();
 b15zdnd11an1n64x5 FILLER_356_264 ();
 b15zdnd11an1n64x5 FILLER_356_328 ();
 b15zdnd11an1n64x5 FILLER_356_392 ();
 b15zdnd11an1n64x5 FILLER_356_456 ();
 b15zdnd11an1n64x5 FILLER_356_520 ();
 b15zdnd11an1n64x5 FILLER_356_584 ();
 b15zdnd11an1n64x5 FILLER_356_648 ();
 b15zdnd11an1n04x5 FILLER_356_712 ();
 b15zdnd00an1n02x5 FILLER_356_716 ();
 b15zdnd11an1n32x5 FILLER_356_726 ();
 b15zdnd11an1n16x5 FILLER_356_758 ();
 b15zdnd11an1n08x5 FILLER_356_774 ();
 b15zdnd11an1n04x5 FILLER_356_782 ();
 b15zdnd00an1n02x5 FILLER_356_786 ();
 b15zdnd00an1n01x5 FILLER_356_788 ();
 b15zdnd11an1n64x5 FILLER_356_792 ();
 b15zdnd11an1n32x5 FILLER_356_856 ();
 b15zdnd11an1n08x5 FILLER_356_888 ();
 b15zdnd11an1n04x5 FILLER_356_896 ();
 b15zdnd00an1n02x5 FILLER_356_900 ();
 b15zdnd11an1n64x5 FILLER_356_917 ();
 b15zdnd11an1n64x5 FILLER_356_981 ();
 b15zdnd11an1n64x5 FILLER_356_1045 ();
 b15zdnd11an1n64x5 FILLER_356_1109 ();
 b15zdnd11an1n32x5 FILLER_356_1173 ();
 b15zdnd11an1n64x5 FILLER_356_1215 ();
 b15zdnd11an1n04x5 FILLER_356_1279 ();
 b15zdnd00an1n01x5 FILLER_356_1283 ();
 b15zdnd11an1n32x5 FILLER_356_1302 ();
 b15zdnd11an1n16x5 FILLER_356_1334 ();
 b15zdnd11an1n04x5 FILLER_356_1350 ();
 b15zdnd00an1n02x5 FILLER_356_1354 ();
 b15zdnd11an1n08x5 FILLER_356_1374 ();
 b15zdnd11an1n04x5 FILLER_356_1382 ();
 b15zdnd00an1n02x5 FILLER_356_1386 ();
 b15zdnd11an1n64x5 FILLER_356_1440 ();
 b15zdnd11an1n64x5 FILLER_356_1504 ();
 b15zdnd11an1n64x5 FILLER_356_1568 ();
 b15zdnd11an1n64x5 FILLER_356_1632 ();
 b15zdnd11an1n64x5 FILLER_356_1696 ();
 b15zdnd11an1n32x5 FILLER_356_1760 ();
 b15zdnd11an1n04x5 FILLER_356_1792 ();
 b15zdnd00an1n01x5 FILLER_356_1796 ();
 b15zdnd11an1n64x5 FILLER_356_1849 ();
 b15zdnd11an1n32x5 FILLER_356_1913 ();
 b15zdnd11an1n16x5 FILLER_356_1945 ();
 b15zdnd00an1n02x5 FILLER_356_1961 ();
 b15zdnd11an1n64x5 FILLER_356_1968 ();
 b15zdnd11an1n64x5 FILLER_356_2032 ();
 b15zdnd11an1n32x5 FILLER_356_2096 ();
 b15zdnd11an1n16x5 FILLER_356_2128 ();
 b15zdnd11an1n08x5 FILLER_356_2144 ();
 b15zdnd00an1n02x5 FILLER_356_2152 ();
 b15zdnd11an1n64x5 FILLER_356_2162 ();
 b15zdnd11an1n32x5 FILLER_356_2226 ();
 b15zdnd11an1n16x5 FILLER_356_2258 ();
 b15zdnd00an1n02x5 FILLER_356_2274 ();
 b15zdnd11an1n64x5 FILLER_357_0 ();
 b15zdnd11an1n64x5 FILLER_357_64 ();
 b15zdnd11an1n64x5 FILLER_357_128 ();
 b15zdnd11an1n64x5 FILLER_357_192 ();
 b15zdnd11an1n64x5 FILLER_357_256 ();
 b15zdnd11an1n64x5 FILLER_357_320 ();
 b15zdnd11an1n64x5 FILLER_357_384 ();
 b15zdnd11an1n64x5 FILLER_357_448 ();
 b15zdnd11an1n64x5 FILLER_357_512 ();
 b15zdnd11an1n64x5 FILLER_357_576 ();
 b15zdnd11an1n64x5 FILLER_357_640 ();
 b15zdnd11an1n32x5 FILLER_357_704 ();
 b15zdnd11an1n16x5 FILLER_357_736 ();
 b15zdnd00an1n02x5 FILLER_357_752 ();
 b15zdnd00an1n01x5 FILLER_357_754 ();
 b15zdnd11an1n04x5 FILLER_357_795 ();
 b15zdnd11an1n64x5 FILLER_357_802 ();
 b15zdnd11an1n64x5 FILLER_357_866 ();
 b15zdnd11an1n32x5 FILLER_357_930 ();
 b15zdnd11an1n16x5 FILLER_357_962 ();
 b15zdnd11an1n64x5 FILLER_357_993 ();
 b15zdnd11an1n64x5 FILLER_357_1057 ();
 b15zdnd11an1n64x5 FILLER_357_1121 ();
 b15zdnd11an1n32x5 FILLER_357_1185 ();
 b15zdnd11an1n04x5 FILLER_357_1217 ();
 b15zdnd00an1n02x5 FILLER_357_1221 ();
 b15zdnd11an1n64x5 FILLER_357_1238 ();
 b15zdnd11an1n64x5 FILLER_357_1302 ();
 b15zdnd11an1n32x5 FILLER_357_1366 ();
 b15zdnd11an1n16x5 FILLER_357_1398 ();
 b15zdnd11an1n64x5 FILLER_357_1417 ();
 b15zdnd11an1n64x5 FILLER_357_1481 ();
 b15zdnd11an1n64x5 FILLER_357_1545 ();
 b15zdnd11an1n64x5 FILLER_357_1609 ();
 b15zdnd11an1n64x5 FILLER_357_1673 ();
 b15zdnd11an1n64x5 FILLER_357_1737 ();
 b15zdnd11an1n16x5 FILLER_357_1801 ();
 b15zdnd11an1n04x5 FILLER_357_1817 ();
 b15zdnd00an1n02x5 FILLER_357_1821 ();
 b15zdnd11an1n64x5 FILLER_357_1826 ();
 b15zdnd11an1n64x5 FILLER_357_1890 ();
 b15zdnd11an1n08x5 FILLER_357_1954 ();
 b15zdnd11an1n04x5 FILLER_357_1962 ();
 b15zdnd11an1n16x5 FILLER_357_1977 ();
 b15zdnd11an1n04x5 FILLER_357_2003 ();
 b15zdnd11an1n64x5 FILLER_357_2011 ();
 b15zdnd11an1n64x5 FILLER_357_2075 ();
 b15zdnd11an1n64x5 FILLER_357_2139 ();
 b15zdnd11an1n64x5 FILLER_357_2203 ();
 b15zdnd11an1n16x5 FILLER_357_2267 ();
 b15zdnd00an1n01x5 FILLER_357_2283 ();
 b15zdnd11an1n64x5 FILLER_358_8 ();
 b15zdnd11an1n64x5 FILLER_358_72 ();
 b15zdnd11an1n64x5 FILLER_358_136 ();
 b15zdnd11an1n64x5 FILLER_358_200 ();
 b15zdnd11an1n64x5 FILLER_358_264 ();
 b15zdnd11an1n64x5 FILLER_358_328 ();
 b15zdnd11an1n64x5 FILLER_358_392 ();
 b15zdnd11an1n64x5 FILLER_358_456 ();
 b15zdnd11an1n64x5 FILLER_358_520 ();
 b15zdnd11an1n64x5 FILLER_358_584 ();
 b15zdnd11an1n64x5 FILLER_358_648 ();
 b15zdnd11an1n04x5 FILLER_358_712 ();
 b15zdnd00an1n02x5 FILLER_358_716 ();
 b15zdnd11an1n64x5 FILLER_358_726 ();
 b15zdnd11an1n64x5 FILLER_358_790 ();
 b15zdnd11an1n64x5 FILLER_358_854 ();
 b15zdnd11an1n64x5 FILLER_358_918 ();
 b15zdnd11an1n64x5 FILLER_358_982 ();
 b15zdnd11an1n64x5 FILLER_358_1046 ();
 b15zdnd11an1n16x5 FILLER_358_1110 ();
 b15zdnd11an1n08x5 FILLER_358_1126 ();
 b15zdnd00an1n02x5 FILLER_358_1134 ();
 b15zdnd11an1n04x5 FILLER_358_1151 ();
 b15zdnd00an1n02x5 FILLER_358_1155 ();
 b15zdnd00an1n01x5 FILLER_358_1157 ();
 b15zdnd11an1n64x5 FILLER_358_1176 ();
 b15zdnd11an1n32x5 FILLER_358_1240 ();
 b15zdnd11an1n16x5 FILLER_358_1272 ();
 b15zdnd11an1n04x5 FILLER_358_1288 ();
 b15zdnd00an1n02x5 FILLER_358_1292 ();
 b15zdnd11an1n04x5 FILLER_358_1312 ();
 b15zdnd11an1n64x5 FILLER_358_1336 ();
 b15zdnd11an1n64x5 FILLER_358_1400 ();
 b15zdnd11an1n32x5 FILLER_358_1464 ();
 b15zdnd11an1n16x5 FILLER_358_1496 ();
 b15zdnd11an1n04x5 FILLER_358_1512 ();
 b15zdnd11an1n04x5 FILLER_358_1543 ();
 b15zdnd11an1n64x5 FILLER_358_1550 ();
 b15zdnd11an1n64x5 FILLER_358_1614 ();
 b15zdnd11an1n64x5 FILLER_358_1678 ();
 b15zdnd11an1n64x5 FILLER_358_1742 ();
 b15zdnd11an1n64x5 FILLER_358_1806 ();
 b15zdnd11an1n64x5 FILLER_358_1870 ();
 b15zdnd11an1n64x5 FILLER_358_1934 ();
 b15zdnd11an1n64x5 FILLER_358_1998 ();
 b15zdnd11an1n64x5 FILLER_358_2062 ();
 b15zdnd11an1n16x5 FILLER_358_2126 ();
 b15zdnd11an1n08x5 FILLER_358_2142 ();
 b15zdnd11an1n04x5 FILLER_358_2150 ();
 b15zdnd11an1n64x5 FILLER_358_2162 ();
 b15zdnd11an1n32x5 FILLER_358_2226 ();
 b15zdnd11an1n16x5 FILLER_358_2258 ();
 b15zdnd00an1n02x5 FILLER_358_2274 ();
 b15zdnd11an1n64x5 FILLER_359_0 ();
 b15zdnd11an1n64x5 FILLER_359_64 ();
 b15zdnd11an1n64x5 FILLER_359_128 ();
 b15zdnd11an1n16x5 FILLER_359_192 ();
 b15zdnd11an1n08x5 FILLER_359_208 ();
 b15zdnd11an1n04x5 FILLER_359_216 ();
 b15zdnd00an1n02x5 FILLER_359_220 ();
 b15zdnd00an1n01x5 FILLER_359_222 ();
 b15zdnd11an1n64x5 FILLER_359_265 ();
 b15zdnd11an1n64x5 FILLER_359_329 ();
 b15zdnd11an1n16x5 FILLER_359_393 ();
 b15zdnd11an1n04x5 FILLER_359_409 ();
 b15zdnd11an1n04x5 FILLER_359_416 ();
 b15zdnd00an1n01x5 FILLER_359_420 ();
 b15zdnd11an1n64x5 FILLER_359_424 ();
 b15zdnd11an1n64x5 FILLER_359_488 ();
 b15zdnd11an1n64x5 FILLER_359_552 ();
 b15zdnd11an1n64x5 FILLER_359_616 ();
 b15zdnd11an1n64x5 FILLER_359_680 ();
 b15zdnd11an1n64x5 FILLER_359_744 ();
 b15zdnd11an1n16x5 FILLER_359_808 ();
 b15zdnd11an1n04x5 FILLER_359_824 ();
 b15zdnd00an1n02x5 FILLER_359_828 ();
 b15zdnd00an1n01x5 FILLER_359_830 ();
 b15zdnd11an1n08x5 FILLER_359_873 ();
 b15zdnd11an1n64x5 FILLER_359_899 ();
 b15zdnd11an1n64x5 FILLER_359_963 ();
 b15zdnd11an1n64x5 FILLER_359_1027 ();
 b15zdnd11an1n64x5 FILLER_359_1091 ();
 b15zdnd11an1n32x5 FILLER_359_1155 ();
 b15zdnd11an1n16x5 FILLER_359_1187 ();
 b15zdnd11an1n08x5 FILLER_359_1203 ();
 b15zdnd11an1n04x5 FILLER_359_1211 ();
 b15zdnd00an1n01x5 FILLER_359_1215 ();
 b15zdnd11an1n04x5 FILLER_359_1240 ();
 b15zdnd11an1n64x5 FILLER_359_1259 ();
 b15zdnd11an1n16x5 FILLER_359_1323 ();
 b15zdnd11an1n04x5 FILLER_359_1339 ();
 b15zdnd00an1n02x5 FILLER_359_1343 ();
 b15zdnd11an1n64x5 FILLER_359_1360 ();
 b15zdnd11an1n64x5 FILLER_359_1424 ();
 b15zdnd11an1n16x5 FILLER_359_1488 ();
 b15zdnd11an1n08x5 FILLER_359_1504 ();
 b15zdnd00an1n02x5 FILLER_359_1512 ();
 b15zdnd00an1n01x5 FILLER_359_1514 ();
 b15zdnd11an1n64x5 FILLER_359_1567 ();
 b15zdnd11an1n64x5 FILLER_359_1631 ();
 b15zdnd11an1n64x5 FILLER_359_1695 ();
 b15zdnd11an1n64x5 FILLER_359_1759 ();
 b15zdnd11an1n64x5 FILLER_359_1823 ();
 b15zdnd11an1n64x5 FILLER_359_1887 ();
 b15zdnd11an1n64x5 FILLER_359_1951 ();
 b15zdnd11an1n64x5 FILLER_359_2015 ();
 b15zdnd11an1n64x5 FILLER_359_2079 ();
 b15zdnd11an1n64x5 FILLER_359_2143 ();
 b15zdnd11an1n64x5 FILLER_359_2207 ();
 b15zdnd11an1n08x5 FILLER_359_2271 ();
 b15zdnd11an1n04x5 FILLER_359_2279 ();
 b15zdnd00an1n01x5 FILLER_359_2283 ();
 b15zdnd11an1n64x5 FILLER_360_8 ();
 b15zdnd11an1n64x5 FILLER_360_72 ();
 b15zdnd11an1n64x5 FILLER_360_136 ();
 b15zdnd11an1n04x5 FILLER_360_200 ();
 b15zdnd00an1n02x5 FILLER_360_204 ();
 b15zdnd00an1n01x5 FILLER_360_206 ();
 b15zdnd11an1n64x5 FILLER_360_259 ();
 b15zdnd11an1n64x5 FILLER_360_323 ();
 b15zdnd11an1n04x5 FILLER_360_387 ();
 b15zdnd00an1n02x5 FILLER_360_391 ();
 b15zdnd11an1n64x5 FILLER_360_425 ();
 b15zdnd11an1n64x5 FILLER_360_489 ();
 b15zdnd11an1n64x5 FILLER_360_553 ();
 b15zdnd11an1n64x5 FILLER_360_617 ();
 b15zdnd11an1n32x5 FILLER_360_681 ();
 b15zdnd11an1n04x5 FILLER_360_713 ();
 b15zdnd00an1n01x5 FILLER_360_717 ();
 b15zdnd11an1n64x5 FILLER_360_726 ();
 b15zdnd11an1n64x5 FILLER_360_790 ();
 b15zdnd11an1n32x5 FILLER_360_854 ();
 b15zdnd11an1n08x5 FILLER_360_886 ();
 b15zdnd00an1n02x5 FILLER_360_894 ();
 b15zdnd00an1n01x5 FILLER_360_896 ();
 b15zdnd11an1n64x5 FILLER_360_928 ();
 b15zdnd11an1n64x5 FILLER_360_992 ();
 b15zdnd11an1n64x5 FILLER_360_1056 ();
 b15zdnd11an1n16x5 FILLER_360_1120 ();
 b15zdnd11an1n04x5 FILLER_360_1136 ();
 b15zdnd00an1n01x5 FILLER_360_1140 ();
 b15zdnd11an1n64x5 FILLER_360_1181 ();
 b15zdnd11an1n64x5 FILLER_360_1245 ();
 b15zdnd11an1n64x5 FILLER_360_1309 ();
 b15zdnd11an1n64x5 FILLER_360_1373 ();
 b15zdnd11an1n64x5 FILLER_360_1437 ();
 b15zdnd11an1n04x5 FILLER_360_1501 ();
 b15zdnd00an1n02x5 FILLER_360_1505 ();
 b15zdnd11an1n04x5 FILLER_360_1559 ();
 b15zdnd11an1n04x5 FILLER_360_1566 ();
 b15zdnd11an1n16x5 FILLER_360_1573 ();
 b15zdnd11an1n08x5 FILLER_360_1589 ();
 b15zdnd00an1n02x5 FILLER_360_1597 ();
 b15zdnd11an1n04x5 FILLER_360_1641 ();
 b15zdnd00an1n02x5 FILLER_360_1645 ();
 b15zdnd00an1n01x5 FILLER_360_1647 ();
 b15zdnd11an1n64x5 FILLER_360_1690 ();
 b15zdnd11an1n64x5 FILLER_360_1754 ();
 b15zdnd11an1n64x5 FILLER_360_1818 ();
 b15zdnd11an1n64x5 FILLER_360_1882 ();
 b15zdnd11an1n64x5 FILLER_360_1946 ();
 b15zdnd11an1n64x5 FILLER_360_2010 ();
 b15zdnd11an1n64x5 FILLER_360_2074 ();
 b15zdnd11an1n16x5 FILLER_360_2138 ();
 b15zdnd11an1n64x5 FILLER_360_2162 ();
 b15zdnd11an1n32x5 FILLER_360_2226 ();
 b15zdnd11an1n16x5 FILLER_360_2258 ();
 b15zdnd00an1n02x5 FILLER_360_2274 ();
 b15zdnd11an1n64x5 FILLER_361_0 ();
 b15zdnd11an1n64x5 FILLER_361_64 ();
 b15zdnd11an1n64x5 FILLER_361_128 ();
 b15zdnd11an1n32x5 FILLER_361_192 ();
 b15zdnd00an1n02x5 FILLER_361_224 ();
 b15zdnd00an1n01x5 FILLER_361_226 ();
 b15zdnd11an1n04x5 FILLER_361_230 ();
 b15zdnd11an1n64x5 FILLER_361_237 ();
 b15zdnd11an1n64x5 FILLER_361_301 ();
 b15zdnd11an1n64x5 FILLER_361_365 ();
 b15zdnd11an1n64x5 FILLER_361_429 ();
 b15zdnd11an1n64x5 FILLER_361_493 ();
 b15zdnd11an1n64x5 FILLER_361_557 ();
 b15zdnd11an1n64x5 FILLER_361_621 ();
 b15zdnd11an1n64x5 FILLER_361_685 ();
 b15zdnd11an1n64x5 FILLER_361_749 ();
 b15zdnd11an1n64x5 FILLER_361_813 ();
 b15zdnd11an1n64x5 FILLER_361_877 ();
 b15zdnd11an1n64x5 FILLER_361_941 ();
 b15zdnd11an1n64x5 FILLER_361_1005 ();
 b15zdnd11an1n32x5 FILLER_361_1069 ();
 b15zdnd11an1n08x5 FILLER_361_1101 ();
 b15zdnd00an1n02x5 FILLER_361_1109 ();
 b15zdnd00an1n01x5 FILLER_361_1111 ();
 b15zdnd11an1n64x5 FILLER_361_1143 ();
 b15zdnd11an1n64x5 FILLER_361_1207 ();
 b15zdnd11an1n64x5 FILLER_361_1271 ();
 b15zdnd11an1n64x5 FILLER_361_1335 ();
 b15zdnd11an1n64x5 FILLER_361_1399 ();
 b15zdnd11an1n32x5 FILLER_361_1463 ();
 b15zdnd11an1n08x5 FILLER_361_1495 ();
 b15zdnd00an1n02x5 FILLER_361_1503 ();
 b15zdnd00an1n01x5 FILLER_361_1505 ();
 b15zdnd11an1n04x5 FILLER_361_1558 ();
 b15zdnd11an1n64x5 FILLER_361_1571 ();
 b15zdnd11an1n64x5 FILLER_361_1635 ();
 b15zdnd11an1n64x5 FILLER_361_1699 ();
 b15zdnd11an1n64x5 FILLER_361_1763 ();
 b15zdnd11an1n64x5 FILLER_361_1827 ();
 b15zdnd11an1n64x5 FILLER_361_1891 ();
 b15zdnd11an1n08x5 FILLER_361_1955 ();
 b15zdnd00an1n02x5 FILLER_361_1963 ();
 b15zdnd11an1n64x5 FILLER_361_2007 ();
 b15zdnd11an1n64x5 FILLER_361_2071 ();
 b15zdnd11an1n64x5 FILLER_361_2135 ();
 b15zdnd11an1n64x5 FILLER_361_2199 ();
 b15zdnd11an1n16x5 FILLER_361_2263 ();
 b15zdnd11an1n04x5 FILLER_361_2279 ();
 b15zdnd00an1n01x5 FILLER_361_2283 ();
 b15zdnd11an1n64x5 FILLER_362_8 ();
 b15zdnd11an1n64x5 FILLER_362_72 ();
 b15zdnd11an1n64x5 FILLER_362_136 ();
 b15zdnd11an1n32x5 FILLER_362_200 ();
 b15zdnd11an1n64x5 FILLER_362_235 ();
 b15zdnd11an1n64x5 FILLER_362_299 ();
 b15zdnd11an1n64x5 FILLER_362_363 ();
 b15zdnd11an1n64x5 FILLER_362_427 ();
 b15zdnd11an1n64x5 FILLER_362_491 ();
 b15zdnd11an1n64x5 FILLER_362_555 ();
 b15zdnd11an1n64x5 FILLER_362_619 ();
 b15zdnd11an1n32x5 FILLER_362_683 ();
 b15zdnd00an1n02x5 FILLER_362_715 ();
 b15zdnd00an1n01x5 FILLER_362_717 ();
 b15zdnd11an1n64x5 FILLER_362_726 ();
 b15zdnd11an1n64x5 FILLER_362_790 ();
 b15zdnd11an1n64x5 FILLER_362_854 ();
 b15zdnd11an1n64x5 FILLER_362_918 ();
 b15zdnd11an1n08x5 FILLER_362_982 ();
 b15zdnd11an1n04x5 FILLER_362_990 ();
 b15zdnd00an1n02x5 FILLER_362_994 ();
 b15zdnd11an1n64x5 FILLER_362_1014 ();
 b15zdnd11an1n64x5 FILLER_362_1078 ();
 b15zdnd11an1n64x5 FILLER_362_1142 ();
 b15zdnd11an1n64x5 FILLER_362_1206 ();
 b15zdnd11an1n64x5 FILLER_362_1270 ();
 b15zdnd11an1n64x5 FILLER_362_1334 ();
 b15zdnd11an1n64x5 FILLER_362_1398 ();
 b15zdnd11an1n32x5 FILLER_362_1462 ();
 b15zdnd11an1n08x5 FILLER_362_1494 ();
 b15zdnd00an1n02x5 FILLER_362_1502 ();
 b15zdnd11an1n04x5 FILLER_362_1507 ();
 b15zdnd11an1n04x5 FILLER_362_1563 ();
 b15zdnd11an1n64x5 FILLER_362_1570 ();
 b15zdnd11an1n64x5 FILLER_362_1634 ();
 b15zdnd11an1n64x5 FILLER_362_1698 ();
 b15zdnd11an1n64x5 FILLER_362_1762 ();
 b15zdnd11an1n64x5 FILLER_362_1826 ();
 b15zdnd11an1n64x5 FILLER_362_1890 ();
 b15zdnd00an1n02x5 FILLER_362_1954 ();
 b15zdnd00an1n01x5 FILLER_362_1956 ();
 b15zdnd11an1n64x5 FILLER_362_1999 ();
 b15zdnd11an1n64x5 FILLER_362_2063 ();
 b15zdnd11an1n16x5 FILLER_362_2127 ();
 b15zdnd11an1n08x5 FILLER_362_2143 ();
 b15zdnd00an1n02x5 FILLER_362_2151 ();
 b15zdnd00an1n01x5 FILLER_362_2153 ();
 b15zdnd11an1n64x5 FILLER_362_2162 ();
 b15zdnd11an1n32x5 FILLER_362_2226 ();
 b15zdnd11an1n16x5 FILLER_362_2258 ();
 b15zdnd00an1n02x5 FILLER_362_2274 ();
 b15zdnd11an1n64x5 FILLER_363_0 ();
 b15zdnd11an1n64x5 FILLER_363_64 ();
 b15zdnd11an1n64x5 FILLER_363_128 ();
 b15zdnd11an1n64x5 FILLER_363_192 ();
 b15zdnd11an1n64x5 FILLER_363_256 ();
 b15zdnd11an1n64x5 FILLER_363_320 ();
 b15zdnd11an1n64x5 FILLER_363_384 ();
 b15zdnd11an1n64x5 FILLER_363_448 ();
 b15zdnd11an1n64x5 FILLER_363_512 ();
 b15zdnd11an1n64x5 FILLER_363_576 ();
 b15zdnd11an1n64x5 FILLER_363_640 ();
 b15zdnd11an1n32x5 FILLER_363_704 ();
 b15zdnd11an1n16x5 FILLER_363_736 ();
 b15zdnd00an1n02x5 FILLER_363_752 ();
 b15zdnd00an1n01x5 FILLER_363_754 ();
 b15zdnd11an1n64x5 FILLER_363_797 ();
 b15zdnd11an1n32x5 FILLER_363_861 ();
 b15zdnd11an1n16x5 FILLER_363_893 ();
 b15zdnd00an1n02x5 FILLER_363_909 ();
 b15zdnd00an1n01x5 FILLER_363_911 ();
 b15zdnd11an1n64x5 FILLER_363_921 ();
 b15zdnd11an1n32x5 FILLER_363_985 ();
 b15zdnd11an1n08x5 FILLER_363_1017 ();
 b15zdnd11an1n04x5 FILLER_363_1025 ();
 b15zdnd00an1n02x5 FILLER_363_1029 ();
 b15zdnd00an1n01x5 FILLER_363_1031 ();
 b15zdnd11an1n64x5 FILLER_363_1044 ();
 b15zdnd11an1n32x5 FILLER_363_1108 ();
 b15zdnd11an1n08x5 FILLER_363_1140 ();
 b15zdnd00an1n01x5 FILLER_363_1148 ();
 b15zdnd11an1n04x5 FILLER_363_1189 ();
 b15zdnd11an1n16x5 FILLER_363_1224 ();
 b15zdnd11an1n64x5 FILLER_363_1250 ();
 b15zdnd11an1n64x5 FILLER_363_1314 ();
 b15zdnd11an1n64x5 FILLER_363_1378 ();
 b15zdnd11an1n64x5 FILLER_363_1442 ();
 b15zdnd11an1n08x5 FILLER_363_1506 ();
 b15zdnd11an1n04x5 FILLER_363_1514 ();
 b15zdnd11an1n04x5 FILLER_363_1521 ();
 b15zdnd00an1n01x5 FILLER_363_1525 ();
 b15zdnd11an1n04x5 FILLER_363_1529 ();
 b15zdnd11an1n04x5 FILLER_363_1536 ();
 b15zdnd11an1n04x5 FILLER_363_1543 ();
 b15zdnd00an1n02x5 FILLER_363_1547 ();
 b15zdnd00an1n01x5 FILLER_363_1549 ();
 b15zdnd11an1n64x5 FILLER_363_1553 ();
 b15zdnd11an1n64x5 FILLER_363_1617 ();
 b15zdnd11an1n64x5 FILLER_363_1681 ();
 b15zdnd11an1n64x5 FILLER_363_1745 ();
 b15zdnd11an1n64x5 FILLER_363_1809 ();
 b15zdnd11an1n64x5 FILLER_363_1873 ();
 b15zdnd11an1n32x5 FILLER_363_1937 ();
 b15zdnd11an1n16x5 FILLER_363_1969 ();
 b15zdnd11an1n64x5 FILLER_363_2027 ();
 b15zdnd11an1n64x5 FILLER_363_2091 ();
 b15zdnd11an1n64x5 FILLER_363_2155 ();
 b15zdnd11an1n64x5 FILLER_363_2219 ();
 b15zdnd00an1n01x5 FILLER_363_2283 ();
 b15zdnd11an1n64x5 FILLER_364_8 ();
 b15zdnd11an1n64x5 FILLER_364_72 ();
 b15zdnd11an1n64x5 FILLER_364_136 ();
 b15zdnd11an1n64x5 FILLER_364_200 ();
 b15zdnd11an1n64x5 FILLER_364_264 ();
 b15zdnd11an1n32x5 FILLER_364_328 ();
 b15zdnd11an1n16x5 FILLER_364_360 ();
 b15zdnd00an1n02x5 FILLER_364_376 ();
 b15zdnd00an1n01x5 FILLER_364_378 ();
 b15zdnd11an1n64x5 FILLER_364_421 ();
 b15zdnd11an1n64x5 FILLER_364_485 ();
 b15zdnd11an1n64x5 FILLER_364_549 ();
 b15zdnd11an1n64x5 FILLER_364_613 ();
 b15zdnd11an1n32x5 FILLER_364_677 ();
 b15zdnd11an1n08x5 FILLER_364_709 ();
 b15zdnd00an1n01x5 FILLER_364_717 ();
 b15zdnd11an1n64x5 FILLER_364_726 ();
 b15zdnd11an1n64x5 FILLER_364_790 ();
 b15zdnd11an1n64x5 FILLER_364_854 ();
 b15zdnd11an1n64x5 FILLER_364_918 ();
 b15zdnd11an1n64x5 FILLER_364_982 ();
 b15zdnd11an1n16x5 FILLER_364_1046 ();
 b15zdnd11an1n04x5 FILLER_364_1072 ();
 b15zdnd11an1n64x5 FILLER_364_1107 ();
 b15zdnd11an1n64x5 FILLER_364_1171 ();
 b15zdnd11an1n08x5 FILLER_364_1235 ();
 b15zdnd00an1n01x5 FILLER_364_1243 ();
 b15zdnd11an1n64x5 FILLER_364_1262 ();
 b15zdnd11an1n64x5 FILLER_364_1326 ();
 b15zdnd11an1n64x5 FILLER_364_1390 ();
 b15zdnd11an1n32x5 FILLER_364_1454 ();
 b15zdnd11an1n16x5 FILLER_364_1486 ();
 b15zdnd11an1n08x5 FILLER_364_1502 ();
 b15zdnd11an1n04x5 FILLER_364_1510 ();
 b15zdnd00an1n02x5 FILLER_364_1514 ();
 b15zdnd11an1n04x5 FILLER_364_1525 ();
 b15zdnd11an1n04x5 FILLER_364_1532 ();
 b15zdnd11an1n04x5 FILLER_364_1539 ();
 b15zdnd11an1n64x5 FILLER_364_1546 ();
 b15zdnd11an1n64x5 FILLER_364_1610 ();
 b15zdnd11an1n64x5 FILLER_364_1674 ();
 b15zdnd11an1n32x5 FILLER_364_1738 ();
 b15zdnd11an1n16x5 FILLER_364_1770 ();
 b15zdnd11an1n08x5 FILLER_364_1786 ();
 b15zdnd11an1n04x5 FILLER_364_1794 ();
 b15zdnd00an1n02x5 FILLER_364_1798 ();
 b15zdnd11an1n64x5 FILLER_364_1805 ();
 b15zdnd11an1n64x5 FILLER_364_1869 ();
 b15zdnd11an1n64x5 FILLER_364_1933 ();
 b15zdnd11an1n64x5 FILLER_364_1997 ();
 b15zdnd11an1n64x5 FILLER_364_2061 ();
 b15zdnd11an1n16x5 FILLER_364_2125 ();
 b15zdnd11an1n08x5 FILLER_364_2141 ();
 b15zdnd11an1n04x5 FILLER_364_2149 ();
 b15zdnd00an1n01x5 FILLER_364_2153 ();
 b15zdnd11an1n64x5 FILLER_364_2162 ();
 b15zdnd11an1n32x5 FILLER_364_2226 ();
 b15zdnd11an1n16x5 FILLER_364_2258 ();
 b15zdnd00an1n02x5 FILLER_364_2274 ();
 b15zdnd11an1n64x5 FILLER_365_0 ();
 b15zdnd11an1n64x5 FILLER_365_64 ();
 b15zdnd11an1n64x5 FILLER_365_128 ();
 b15zdnd11an1n64x5 FILLER_365_192 ();
 b15zdnd11an1n64x5 FILLER_365_256 ();
 b15zdnd11an1n64x5 FILLER_365_320 ();
 b15zdnd11an1n64x5 FILLER_365_384 ();
 b15zdnd11an1n32x5 FILLER_365_448 ();
 b15zdnd00an1n02x5 FILLER_365_480 ();
 b15zdnd11an1n64x5 FILLER_365_524 ();
 b15zdnd11an1n64x5 FILLER_365_588 ();
 b15zdnd11an1n64x5 FILLER_365_652 ();
 b15zdnd11an1n64x5 FILLER_365_716 ();
 b15zdnd11an1n64x5 FILLER_365_780 ();
 b15zdnd11an1n64x5 FILLER_365_844 ();
 b15zdnd11an1n64x5 FILLER_365_908 ();
 b15zdnd11an1n08x5 FILLER_365_972 ();
 b15zdnd11an1n04x5 FILLER_365_980 ();
 b15zdnd11an1n32x5 FILLER_365_988 ();
 b15zdnd11an1n08x5 FILLER_365_1020 ();
 b15zdnd11an1n04x5 FILLER_365_1028 ();
 b15zdnd00an1n02x5 FILLER_365_1032 ();
 b15zdnd00an1n01x5 FILLER_365_1034 ();
 b15zdnd11an1n64x5 FILLER_365_1042 ();
 b15zdnd11an1n32x5 FILLER_365_1106 ();
 b15zdnd11an1n04x5 FILLER_365_1138 ();
 b15zdnd00an1n02x5 FILLER_365_1142 ();
 b15zdnd11an1n64x5 FILLER_365_1169 ();
 b15zdnd11an1n32x5 FILLER_365_1233 ();
 b15zdnd11an1n08x5 FILLER_365_1265 ();
 b15zdnd11an1n04x5 FILLER_365_1273 ();
 b15zdnd11an1n64x5 FILLER_365_1308 ();
 b15zdnd11an1n64x5 FILLER_365_1372 ();
 b15zdnd11an1n64x5 FILLER_365_1436 ();
 b15zdnd11an1n64x5 FILLER_365_1500 ();
 b15zdnd11an1n64x5 FILLER_365_1564 ();
 b15zdnd11an1n64x5 FILLER_365_1628 ();
 b15zdnd11an1n64x5 FILLER_365_1692 ();
 b15zdnd11an1n08x5 FILLER_365_1756 ();
 b15zdnd11an1n04x5 FILLER_365_1764 ();
 b15zdnd00an1n02x5 FILLER_365_1768 ();
 b15zdnd11an1n64x5 FILLER_365_1778 ();
 b15zdnd11an1n64x5 FILLER_365_1842 ();
 b15zdnd11an1n64x5 FILLER_365_1906 ();
 b15zdnd11an1n64x5 FILLER_365_1970 ();
 b15zdnd11an1n64x5 FILLER_365_2034 ();
 b15zdnd11an1n64x5 FILLER_365_2098 ();
 b15zdnd11an1n64x5 FILLER_365_2162 ();
 b15zdnd11an1n32x5 FILLER_365_2226 ();
 b15zdnd11an1n16x5 FILLER_365_2258 ();
 b15zdnd11an1n08x5 FILLER_365_2274 ();
 b15zdnd00an1n02x5 FILLER_365_2282 ();
 b15zdnd11an1n64x5 FILLER_366_8 ();
 b15zdnd11an1n64x5 FILLER_366_72 ();
 b15zdnd11an1n64x5 FILLER_366_136 ();
 b15zdnd11an1n64x5 FILLER_366_200 ();
 b15zdnd11an1n64x5 FILLER_366_264 ();
 b15zdnd11an1n08x5 FILLER_366_328 ();
 b15zdnd00an1n01x5 FILLER_366_336 ();
 b15zdnd11an1n64x5 FILLER_366_369 ();
 b15zdnd11an1n64x5 FILLER_366_433 ();
 b15zdnd11an1n64x5 FILLER_366_497 ();
 b15zdnd11an1n64x5 FILLER_366_561 ();
 b15zdnd11an1n64x5 FILLER_366_625 ();
 b15zdnd11an1n16x5 FILLER_366_689 ();
 b15zdnd11an1n08x5 FILLER_366_705 ();
 b15zdnd11an1n04x5 FILLER_366_713 ();
 b15zdnd00an1n01x5 FILLER_366_717 ();
 b15zdnd11an1n32x5 FILLER_366_726 ();
 b15zdnd00an1n02x5 FILLER_366_758 ();
 b15zdnd11an1n64x5 FILLER_366_802 ();
 b15zdnd11an1n64x5 FILLER_366_866 ();
 b15zdnd11an1n64x5 FILLER_366_930 ();
 b15zdnd11an1n32x5 FILLER_366_994 ();
 b15zdnd11an1n16x5 FILLER_366_1026 ();
 b15zdnd00an1n01x5 FILLER_366_1042 ();
 b15zdnd11an1n32x5 FILLER_366_1063 ();
 b15zdnd11an1n04x5 FILLER_366_1095 ();
 b15zdnd00an1n02x5 FILLER_366_1099 ();
 b15zdnd00an1n01x5 FILLER_366_1101 ();
 b15zdnd11an1n64x5 FILLER_366_1127 ();
 b15zdnd11an1n64x5 FILLER_366_1191 ();
 b15zdnd11an1n64x5 FILLER_366_1255 ();
 b15zdnd11an1n64x5 FILLER_366_1319 ();
 b15zdnd11an1n64x5 FILLER_366_1383 ();
 b15zdnd11an1n64x5 FILLER_366_1447 ();
 b15zdnd11an1n64x5 FILLER_366_1511 ();
 b15zdnd11an1n64x5 FILLER_366_1575 ();
 b15zdnd11an1n64x5 FILLER_366_1639 ();
 b15zdnd00an1n02x5 FILLER_366_1703 ();
 b15zdnd11an1n16x5 FILLER_366_1757 ();
 b15zdnd00an1n02x5 FILLER_366_1773 ();
 b15zdnd00an1n01x5 FILLER_366_1775 ();
 b15zdnd11an1n64x5 FILLER_366_1781 ();
 b15zdnd11an1n64x5 FILLER_366_1845 ();
 b15zdnd11an1n64x5 FILLER_366_1909 ();
 b15zdnd11an1n64x5 FILLER_366_1973 ();
 b15zdnd11an1n64x5 FILLER_366_2037 ();
 b15zdnd11an1n32x5 FILLER_366_2101 ();
 b15zdnd11an1n16x5 FILLER_366_2133 ();
 b15zdnd11an1n04x5 FILLER_366_2149 ();
 b15zdnd00an1n01x5 FILLER_366_2153 ();
 b15zdnd11an1n64x5 FILLER_366_2162 ();
 b15zdnd11an1n32x5 FILLER_366_2226 ();
 b15zdnd11an1n16x5 FILLER_366_2258 ();
 b15zdnd00an1n02x5 FILLER_366_2274 ();
 b15zdnd11an1n64x5 FILLER_367_0 ();
 b15zdnd11an1n64x5 FILLER_367_64 ();
 b15zdnd11an1n64x5 FILLER_367_128 ();
 b15zdnd11an1n64x5 FILLER_367_192 ();
 b15zdnd11an1n64x5 FILLER_367_256 ();
 b15zdnd11an1n32x5 FILLER_367_320 ();
 b15zdnd11an1n04x5 FILLER_367_352 ();
 b15zdnd00an1n02x5 FILLER_367_356 ();
 b15zdnd11an1n04x5 FILLER_367_361 ();
 b15zdnd11an1n64x5 FILLER_367_368 ();
 b15zdnd11an1n64x5 FILLER_367_432 ();
 b15zdnd11an1n64x5 FILLER_367_496 ();
 b15zdnd11an1n64x5 FILLER_367_560 ();
 b15zdnd11an1n64x5 FILLER_367_624 ();
 b15zdnd11an1n08x5 FILLER_367_688 ();
 b15zdnd11an1n04x5 FILLER_367_696 ();
 b15zdnd00an1n02x5 FILLER_367_700 ();
 b15zdnd11an1n64x5 FILLER_367_706 ();
 b15zdnd11an1n64x5 FILLER_367_770 ();
 b15zdnd11an1n64x5 FILLER_367_834 ();
 b15zdnd11an1n08x5 FILLER_367_898 ();
 b15zdnd11an1n04x5 FILLER_367_906 ();
 b15zdnd00an1n02x5 FILLER_367_910 ();
 b15zdnd11an1n64x5 FILLER_367_925 ();
 b15zdnd11an1n64x5 FILLER_367_989 ();
 b15zdnd11an1n32x5 FILLER_367_1053 ();
 b15zdnd11an1n08x5 FILLER_367_1085 ();
 b15zdnd11an1n04x5 FILLER_367_1093 ();
 b15zdnd11an1n64x5 FILLER_367_1137 ();
 b15zdnd11an1n64x5 FILLER_367_1201 ();
 b15zdnd11an1n32x5 FILLER_367_1265 ();
 b15zdnd11an1n16x5 FILLER_367_1297 ();
 b15zdnd11an1n08x5 FILLER_367_1313 ();
 b15zdnd11an1n04x5 FILLER_367_1321 ();
 b15zdnd00an1n02x5 FILLER_367_1325 ();
 b15zdnd00an1n01x5 FILLER_367_1327 ();
 b15zdnd11an1n08x5 FILLER_367_1338 ();
 b15zdnd11an1n04x5 FILLER_367_1346 ();
 b15zdnd11an1n08x5 FILLER_367_1365 ();
 b15zdnd11an1n04x5 FILLER_367_1373 ();
 b15zdnd00an1n02x5 FILLER_367_1377 ();
 b15zdnd11an1n64x5 FILLER_367_1388 ();
 b15zdnd11an1n64x5 FILLER_367_1452 ();
 b15zdnd11an1n04x5 FILLER_367_1516 ();
 b15zdnd00an1n02x5 FILLER_367_1520 ();
 b15zdnd11an1n04x5 FILLER_367_1564 ();
 b15zdnd00an1n01x5 FILLER_367_1568 ();
 b15zdnd11an1n64x5 FILLER_367_1611 ();
 b15zdnd11an1n32x5 FILLER_367_1675 ();
 b15zdnd11an1n16x5 FILLER_367_1707 ();
 b15zdnd11an1n04x5 FILLER_367_1726 ();
 b15zdnd11an1n32x5 FILLER_367_1733 ();
 b15zdnd11an1n04x5 FILLER_367_1765 ();
 b15zdnd00an1n02x5 FILLER_367_1769 ();
 b15zdnd11an1n08x5 FILLER_367_1778 ();
 b15zdnd11an1n04x5 FILLER_367_1786 ();
 b15zdnd00an1n01x5 FILLER_367_1790 ();
 b15zdnd11an1n64x5 FILLER_367_1797 ();
 b15zdnd11an1n64x5 FILLER_367_1861 ();
 b15zdnd11an1n32x5 FILLER_367_1925 ();
 b15zdnd11an1n04x5 FILLER_367_1957 ();
 b15zdnd00an1n02x5 FILLER_367_1961 ();
 b15zdnd00an1n01x5 FILLER_367_1963 ();
 b15zdnd11an1n04x5 FILLER_367_1967 ();
 b15zdnd11an1n64x5 FILLER_367_1974 ();
 b15zdnd11an1n64x5 FILLER_367_2038 ();
 b15zdnd11an1n64x5 FILLER_367_2102 ();
 b15zdnd11an1n64x5 FILLER_367_2166 ();
 b15zdnd11an1n32x5 FILLER_367_2230 ();
 b15zdnd11an1n16x5 FILLER_367_2262 ();
 b15zdnd11an1n04x5 FILLER_367_2278 ();
 b15zdnd00an1n02x5 FILLER_367_2282 ();
 b15zdnd11an1n64x5 FILLER_368_8 ();
 b15zdnd11an1n64x5 FILLER_368_72 ();
 b15zdnd11an1n64x5 FILLER_368_136 ();
 b15zdnd11an1n64x5 FILLER_368_200 ();
 b15zdnd11an1n64x5 FILLER_368_264 ();
 b15zdnd11an1n64x5 FILLER_368_328 ();
 b15zdnd11an1n64x5 FILLER_368_392 ();
 b15zdnd11an1n64x5 FILLER_368_456 ();
 b15zdnd11an1n64x5 FILLER_368_520 ();
 b15zdnd11an1n64x5 FILLER_368_584 ();
 b15zdnd11an1n16x5 FILLER_368_648 ();
 b15zdnd11an1n04x5 FILLER_368_664 ();
 b15zdnd00an1n02x5 FILLER_368_668 ();
 b15zdnd00an1n01x5 FILLER_368_670 ();
 b15zdnd11an1n16x5 FILLER_368_699 ();
 b15zdnd00an1n02x5 FILLER_368_715 ();
 b15zdnd00an1n01x5 FILLER_368_717 ();
 b15zdnd11an1n64x5 FILLER_368_726 ();
 b15zdnd11an1n64x5 FILLER_368_790 ();
 b15zdnd11an1n64x5 FILLER_368_854 ();
 b15zdnd11an1n64x5 FILLER_368_918 ();
 b15zdnd11an1n64x5 FILLER_368_982 ();
 b15zdnd11an1n64x5 FILLER_368_1046 ();
 b15zdnd11an1n64x5 FILLER_368_1110 ();
 b15zdnd11an1n64x5 FILLER_368_1174 ();
 b15zdnd11an1n64x5 FILLER_368_1238 ();
 b15zdnd11an1n64x5 FILLER_368_1302 ();
 b15zdnd11an1n64x5 FILLER_368_1366 ();
 b15zdnd11an1n32x5 FILLER_368_1430 ();
 b15zdnd11an1n16x5 FILLER_368_1462 ();
 b15zdnd11an1n08x5 FILLER_368_1478 ();
 b15zdnd11an1n04x5 FILLER_368_1486 ();
 b15zdnd00an1n02x5 FILLER_368_1490 ();
 b15zdnd00an1n01x5 FILLER_368_1492 ();
 b15zdnd11an1n04x5 FILLER_368_1535 ();
 b15zdnd00an1n01x5 FILLER_368_1539 ();
 b15zdnd11an1n64x5 FILLER_368_1582 ();
 b15zdnd11an1n64x5 FILLER_368_1646 ();
 b15zdnd11an1n16x5 FILLER_368_1710 ();
 b15zdnd11an1n04x5 FILLER_368_1726 ();
 b15zdnd00an1n01x5 FILLER_368_1730 ();
 b15zdnd11an1n32x5 FILLER_368_1734 ();
 b15zdnd11an1n08x5 FILLER_368_1766 ();
 b15zdnd00an1n01x5 FILLER_368_1774 ();
 b15zdnd11an1n64x5 FILLER_368_1796 ();
 b15zdnd11an1n64x5 FILLER_368_1860 ();
 b15zdnd11an1n16x5 FILLER_368_1924 ();
 b15zdnd11an1n04x5 FILLER_368_1940 ();
 b15zdnd00an1n02x5 FILLER_368_1944 ();
 b15zdnd11an1n64x5 FILLER_368_1998 ();
 b15zdnd11an1n64x5 FILLER_368_2062 ();
 b15zdnd11an1n16x5 FILLER_368_2126 ();
 b15zdnd11an1n08x5 FILLER_368_2142 ();
 b15zdnd11an1n04x5 FILLER_368_2150 ();
 b15zdnd11an1n64x5 FILLER_368_2162 ();
 b15zdnd11an1n32x5 FILLER_368_2226 ();
 b15zdnd11an1n16x5 FILLER_368_2258 ();
 b15zdnd00an1n02x5 FILLER_368_2274 ();
 b15zdnd11an1n64x5 FILLER_369_0 ();
 b15zdnd11an1n64x5 FILLER_369_64 ();
 b15zdnd11an1n64x5 FILLER_369_128 ();
 b15zdnd11an1n64x5 FILLER_369_192 ();
 b15zdnd11an1n64x5 FILLER_369_256 ();
 b15zdnd11an1n64x5 FILLER_369_320 ();
 b15zdnd11an1n64x5 FILLER_369_384 ();
 b15zdnd11an1n64x5 FILLER_369_448 ();
 b15zdnd11an1n16x5 FILLER_369_512 ();
 b15zdnd11an1n08x5 FILLER_369_528 ();
 b15zdnd11an1n04x5 FILLER_369_536 ();
 b15zdnd00an1n02x5 FILLER_369_540 ();
 b15zdnd00an1n01x5 FILLER_369_542 ();
 b15zdnd11an1n04x5 FILLER_369_575 ();
 b15zdnd11an1n64x5 FILLER_369_582 ();
 b15zdnd11an1n32x5 FILLER_369_646 ();
 b15zdnd11an1n08x5 FILLER_369_678 ();
 b15zdnd00an1n01x5 FILLER_369_686 ();
 b15zdnd11an1n04x5 FILLER_369_690 ();
 b15zdnd00an1n02x5 FILLER_369_694 ();
 b15zdnd11an1n64x5 FILLER_369_699 ();
 b15zdnd11an1n32x5 FILLER_369_763 ();
 b15zdnd11an1n16x5 FILLER_369_795 ();
 b15zdnd00an1n02x5 FILLER_369_811 ();
 b15zdnd00an1n01x5 FILLER_369_813 ();
 b15zdnd11an1n64x5 FILLER_369_817 ();
 b15zdnd11an1n64x5 FILLER_369_881 ();
 b15zdnd11an1n64x5 FILLER_369_945 ();
 b15zdnd11an1n64x5 FILLER_369_1009 ();
 b15zdnd11an1n64x5 FILLER_369_1073 ();
 b15zdnd11an1n64x5 FILLER_369_1137 ();
 b15zdnd11an1n64x5 FILLER_369_1201 ();
 b15zdnd11an1n64x5 FILLER_369_1265 ();
 b15zdnd11an1n64x5 FILLER_369_1329 ();
 b15zdnd11an1n64x5 FILLER_369_1393 ();
 b15zdnd11an1n32x5 FILLER_369_1457 ();
 b15zdnd11an1n16x5 FILLER_369_1489 ();
 b15zdnd00an1n01x5 FILLER_369_1505 ();
 b15zdnd11an1n04x5 FILLER_369_1548 ();
 b15zdnd11an1n64x5 FILLER_369_1594 ();
 b15zdnd11an1n64x5 FILLER_369_1658 ();
 b15zdnd11an1n32x5 FILLER_369_1722 ();
 b15zdnd11an1n16x5 FILLER_369_1754 ();
 b15zdnd11an1n08x5 FILLER_369_1770 ();
 b15zdnd11an1n04x5 FILLER_369_1781 ();
 b15zdnd11an1n64x5 FILLER_369_1789 ();
 b15zdnd11an1n64x5 FILLER_369_1853 ();
 b15zdnd11an1n32x5 FILLER_369_1917 ();
 b15zdnd11an1n16x5 FILLER_369_1949 ();
 b15zdnd11an1n04x5 FILLER_369_1965 ();
 b15zdnd00an1n02x5 FILLER_369_1969 ();
 b15zdnd11an1n64x5 FILLER_369_1974 ();
 b15zdnd11an1n64x5 FILLER_369_2038 ();
 b15zdnd11an1n64x5 FILLER_369_2102 ();
 b15zdnd11an1n64x5 FILLER_369_2166 ();
 b15zdnd11an1n32x5 FILLER_369_2230 ();
 b15zdnd11an1n16x5 FILLER_369_2262 ();
 b15zdnd11an1n04x5 FILLER_369_2278 ();
 b15zdnd00an1n02x5 FILLER_369_2282 ();
 b15zdnd11an1n64x5 FILLER_370_8 ();
 b15zdnd11an1n64x5 FILLER_370_72 ();
 b15zdnd11an1n64x5 FILLER_370_136 ();
 b15zdnd11an1n64x5 FILLER_370_200 ();
 b15zdnd11an1n64x5 FILLER_370_264 ();
 b15zdnd11an1n64x5 FILLER_370_328 ();
 b15zdnd11an1n64x5 FILLER_370_392 ();
 b15zdnd11an1n64x5 FILLER_370_456 ();
 b15zdnd11an1n32x5 FILLER_370_520 ();
 b15zdnd11an1n08x5 FILLER_370_552 ();
 b15zdnd11an1n04x5 FILLER_370_560 ();
 b15zdnd00an1n02x5 FILLER_370_564 ();
 b15zdnd00an1n01x5 FILLER_370_566 ();
 b15zdnd11an1n64x5 FILLER_370_570 ();
 b15zdnd11an1n64x5 FILLER_370_634 ();
 b15zdnd11an1n16x5 FILLER_370_698 ();
 b15zdnd11an1n04x5 FILLER_370_714 ();
 b15zdnd11an1n32x5 FILLER_370_726 ();
 b15zdnd11an1n16x5 FILLER_370_758 ();
 b15zdnd11an1n04x5 FILLER_370_774 ();
 b15zdnd00an1n02x5 FILLER_370_778 ();
 b15zdnd11an1n64x5 FILLER_370_820 ();
 b15zdnd11an1n64x5 FILLER_370_884 ();
 b15zdnd11an1n64x5 FILLER_370_948 ();
 b15zdnd11an1n64x5 FILLER_370_1012 ();
 b15zdnd11an1n64x5 FILLER_370_1076 ();
 b15zdnd11an1n64x5 FILLER_370_1140 ();
 b15zdnd11an1n64x5 FILLER_370_1204 ();
 b15zdnd11an1n16x5 FILLER_370_1268 ();
 b15zdnd11an1n08x5 FILLER_370_1284 ();
 b15zdnd00an1n02x5 FILLER_370_1292 ();
 b15zdnd11an1n64x5 FILLER_370_1336 ();
 b15zdnd11an1n64x5 FILLER_370_1400 ();
 b15zdnd11an1n32x5 FILLER_370_1464 ();
 b15zdnd11an1n16x5 FILLER_370_1496 ();
 b15zdnd00an1n01x5 FILLER_370_1512 ();
 b15zdnd11an1n04x5 FILLER_370_1555 ();
 b15zdnd00an1n02x5 FILLER_370_1559 ();
 b15zdnd00an1n01x5 FILLER_370_1561 ();
 b15zdnd11an1n64x5 FILLER_370_1604 ();
 b15zdnd11an1n64x5 FILLER_370_1668 ();
 b15zdnd11an1n32x5 FILLER_370_1732 ();
 b15zdnd00an1n02x5 FILLER_370_1764 ();
 b15zdnd00an1n01x5 FILLER_370_1766 ();
 b15zdnd11an1n64x5 FILLER_370_1809 ();
 b15zdnd11an1n64x5 FILLER_370_1873 ();
 b15zdnd11an1n64x5 FILLER_370_1937 ();
 b15zdnd11an1n64x5 FILLER_370_2001 ();
 b15zdnd11an1n64x5 FILLER_370_2065 ();
 b15zdnd11an1n16x5 FILLER_370_2129 ();
 b15zdnd11an1n08x5 FILLER_370_2145 ();
 b15zdnd00an1n01x5 FILLER_370_2153 ();
 b15zdnd11an1n64x5 FILLER_370_2162 ();
 b15zdnd11an1n32x5 FILLER_370_2226 ();
 b15zdnd11an1n16x5 FILLER_370_2258 ();
 b15zdnd00an1n02x5 FILLER_370_2274 ();
 b15zdnd11an1n64x5 FILLER_371_0 ();
 b15zdnd11an1n64x5 FILLER_371_64 ();
 b15zdnd11an1n64x5 FILLER_371_128 ();
 b15zdnd11an1n64x5 FILLER_371_192 ();
 b15zdnd11an1n64x5 FILLER_371_256 ();
 b15zdnd11an1n64x5 FILLER_371_320 ();
 b15zdnd11an1n64x5 FILLER_371_384 ();
 b15zdnd11an1n64x5 FILLER_371_448 ();
 b15zdnd11an1n64x5 FILLER_371_512 ();
 b15zdnd11an1n64x5 FILLER_371_576 ();
 b15zdnd11an1n32x5 FILLER_371_640 ();
 b15zdnd11an1n16x5 FILLER_371_672 ();
 b15zdnd00an1n02x5 FILLER_371_688 ();
 b15zdnd00an1n01x5 FILLER_371_690 ();
 b15zdnd11an1n32x5 FILLER_371_695 ();
 b15zdnd11an1n16x5 FILLER_371_727 ();
 b15zdnd11an1n08x5 FILLER_371_743 ();
 b15zdnd00an1n02x5 FILLER_371_751 ();
 b15zdnd00an1n01x5 FILLER_371_753 ();
 b15zdnd11an1n16x5 FILLER_371_796 ();
 b15zdnd00an1n02x5 FILLER_371_812 ();
 b15zdnd11an1n64x5 FILLER_371_817 ();
 b15zdnd11an1n64x5 FILLER_371_881 ();
 b15zdnd11an1n64x5 FILLER_371_945 ();
 b15zdnd11an1n64x5 FILLER_371_1009 ();
 b15zdnd11an1n64x5 FILLER_371_1073 ();
 b15zdnd11an1n64x5 FILLER_371_1137 ();
 b15zdnd11an1n64x5 FILLER_371_1201 ();
 b15zdnd11an1n64x5 FILLER_371_1265 ();
 b15zdnd11an1n64x5 FILLER_371_1329 ();
 b15zdnd11an1n64x5 FILLER_371_1393 ();
 b15zdnd11an1n64x5 FILLER_371_1457 ();
 b15zdnd11an1n64x5 FILLER_371_1521 ();
 b15zdnd11an1n64x5 FILLER_371_1585 ();
 b15zdnd11an1n64x5 FILLER_371_1649 ();
 b15zdnd11an1n64x5 FILLER_371_1713 ();
 b15zdnd11an1n64x5 FILLER_371_1777 ();
 b15zdnd11an1n64x5 FILLER_371_1841 ();
 b15zdnd11an1n64x5 FILLER_371_1905 ();
 b15zdnd11an1n64x5 FILLER_371_1969 ();
 b15zdnd11an1n64x5 FILLER_371_2033 ();
 b15zdnd11an1n64x5 FILLER_371_2097 ();
 b15zdnd11an1n64x5 FILLER_371_2161 ();
 b15zdnd11an1n32x5 FILLER_371_2225 ();
 b15zdnd11an1n16x5 FILLER_371_2257 ();
 b15zdnd11an1n08x5 FILLER_371_2273 ();
 b15zdnd00an1n02x5 FILLER_371_2281 ();
 b15zdnd00an1n01x5 FILLER_371_2283 ();
 b15zdnd11an1n64x5 FILLER_372_8 ();
 b15zdnd11an1n64x5 FILLER_372_72 ();
 b15zdnd11an1n64x5 FILLER_372_136 ();
 b15zdnd11an1n64x5 FILLER_372_200 ();
 b15zdnd11an1n64x5 FILLER_372_264 ();
 b15zdnd11an1n64x5 FILLER_372_328 ();
 b15zdnd11an1n64x5 FILLER_372_392 ();
 b15zdnd11an1n64x5 FILLER_372_456 ();
 b15zdnd11an1n64x5 FILLER_372_520 ();
 b15zdnd11an1n64x5 FILLER_372_584 ();
 b15zdnd11an1n64x5 FILLER_372_648 ();
 b15zdnd11an1n04x5 FILLER_372_712 ();
 b15zdnd00an1n02x5 FILLER_372_716 ();
 b15zdnd11an1n64x5 FILLER_372_726 ();
 b15zdnd11an1n64x5 FILLER_372_790 ();
 b15zdnd11an1n32x5 FILLER_372_854 ();
 b15zdnd11an1n16x5 FILLER_372_886 ();
 b15zdnd11an1n08x5 FILLER_372_902 ();
 b15zdnd11an1n04x5 FILLER_372_910 ();
 b15zdnd00an1n02x5 FILLER_372_914 ();
 b15zdnd00an1n01x5 FILLER_372_916 ();
 b15zdnd11an1n64x5 FILLER_372_927 ();
 b15zdnd11an1n64x5 FILLER_372_991 ();
 b15zdnd11an1n64x5 FILLER_372_1055 ();
 b15zdnd11an1n64x5 FILLER_372_1119 ();
 b15zdnd11an1n32x5 FILLER_372_1183 ();
 b15zdnd11an1n16x5 FILLER_372_1215 ();
 b15zdnd11an1n08x5 FILLER_372_1231 ();
 b15zdnd11an1n04x5 FILLER_372_1239 ();
 b15zdnd00an1n02x5 FILLER_372_1243 ();
 b15zdnd11an1n64x5 FILLER_372_1287 ();
 b15zdnd11an1n64x5 FILLER_372_1351 ();
 b15zdnd11an1n64x5 FILLER_372_1415 ();
 b15zdnd11an1n64x5 FILLER_372_1479 ();
 b15zdnd11an1n64x5 FILLER_372_1543 ();
 b15zdnd11an1n64x5 FILLER_372_1607 ();
 b15zdnd11an1n64x5 FILLER_372_1671 ();
 b15zdnd11an1n64x5 FILLER_372_1735 ();
 b15zdnd11an1n64x5 FILLER_372_1799 ();
 b15zdnd11an1n64x5 FILLER_372_1863 ();
 b15zdnd11an1n64x5 FILLER_372_1927 ();
 b15zdnd11an1n64x5 FILLER_372_1991 ();
 b15zdnd11an1n64x5 FILLER_372_2055 ();
 b15zdnd11an1n32x5 FILLER_372_2119 ();
 b15zdnd00an1n02x5 FILLER_372_2151 ();
 b15zdnd00an1n01x5 FILLER_372_2153 ();
 b15zdnd11an1n64x5 FILLER_372_2162 ();
 b15zdnd11an1n32x5 FILLER_372_2226 ();
 b15zdnd11an1n16x5 FILLER_372_2258 ();
 b15zdnd00an1n02x5 FILLER_372_2274 ();
 b15zdnd11an1n64x5 FILLER_373_0 ();
 b15zdnd11an1n64x5 FILLER_373_64 ();
 b15zdnd11an1n64x5 FILLER_373_128 ();
 b15zdnd11an1n64x5 FILLER_373_192 ();
 b15zdnd11an1n64x5 FILLER_373_256 ();
 b15zdnd11an1n64x5 FILLER_373_320 ();
 b15zdnd11an1n64x5 FILLER_373_384 ();
 b15zdnd11an1n64x5 FILLER_373_448 ();
 b15zdnd11an1n64x5 FILLER_373_512 ();
 b15zdnd11an1n64x5 FILLER_373_576 ();
 b15zdnd11an1n32x5 FILLER_373_640 ();
 b15zdnd11an1n08x5 FILLER_373_672 ();
 b15zdnd11an1n32x5 FILLER_373_722 ();
 b15zdnd11an1n04x5 FILLER_373_754 ();
 b15zdnd00an1n02x5 FILLER_373_758 ();
 b15zdnd00an1n01x5 FILLER_373_760 ();
 b15zdnd11an1n64x5 FILLER_373_803 ();
 b15zdnd11an1n32x5 FILLER_373_867 ();
 b15zdnd11an1n08x5 FILLER_373_899 ();
 b15zdnd00an1n02x5 FILLER_373_907 ();
 b15zdnd00an1n01x5 FILLER_373_909 ();
 b15zdnd11an1n64x5 FILLER_373_916 ();
 b15zdnd11an1n64x5 FILLER_373_980 ();
 b15zdnd11an1n64x5 FILLER_373_1044 ();
 b15zdnd11an1n64x5 FILLER_373_1108 ();
 b15zdnd11an1n64x5 FILLER_373_1172 ();
 b15zdnd11an1n64x5 FILLER_373_1236 ();
 b15zdnd11an1n64x5 FILLER_373_1300 ();
 b15zdnd11an1n64x5 FILLER_373_1364 ();
 b15zdnd11an1n64x5 FILLER_373_1428 ();
 b15zdnd11an1n32x5 FILLER_373_1492 ();
 b15zdnd00an1n01x5 FILLER_373_1524 ();
 b15zdnd11an1n64x5 FILLER_373_1567 ();
 b15zdnd11an1n64x5 FILLER_373_1631 ();
 b15zdnd11an1n64x5 FILLER_373_1695 ();
 b15zdnd11an1n16x5 FILLER_373_1759 ();
 b15zdnd11an1n08x5 FILLER_373_1775 ();
 b15zdnd11an1n04x5 FILLER_373_1783 ();
 b15zdnd00an1n02x5 FILLER_373_1787 ();
 b15zdnd00an1n01x5 FILLER_373_1789 ();
 b15zdnd11an1n64x5 FILLER_373_1799 ();
 b15zdnd11an1n64x5 FILLER_373_1863 ();
 b15zdnd11an1n64x5 FILLER_373_1927 ();
 b15zdnd11an1n64x5 FILLER_373_1991 ();
 b15zdnd11an1n64x5 FILLER_373_2055 ();
 b15zdnd11an1n64x5 FILLER_373_2119 ();
 b15zdnd11an1n64x5 FILLER_373_2183 ();
 b15zdnd11an1n32x5 FILLER_373_2247 ();
 b15zdnd11an1n04x5 FILLER_373_2279 ();
 b15zdnd00an1n01x5 FILLER_373_2283 ();
 b15zdnd11an1n64x5 FILLER_374_8 ();
 b15zdnd11an1n64x5 FILLER_374_72 ();
 b15zdnd11an1n64x5 FILLER_374_136 ();
 b15zdnd11an1n64x5 FILLER_374_200 ();
 b15zdnd11an1n64x5 FILLER_374_264 ();
 b15zdnd11an1n64x5 FILLER_374_328 ();
 b15zdnd11an1n64x5 FILLER_374_392 ();
 b15zdnd11an1n64x5 FILLER_374_456 ();
 b15zdnd11an1n64x5 FILLER_374_520 ();
 b15zdnd11an1n64x5 FILLER_374_584 ();
 b15zdnd11an1n64x5 FILLER_374_648 ();
 b15zdnd11an1n04x5 FILLER_374_712 ();
 b15zdnd00an1n02x5 FILLER_374_716 ();
 b15zdnd11an1n64x5 FILLER_374_726 ();
 b15zdnd11an1n64x5 FILLER_374_790 ();
 b15zdnd11an1n32x5 FILLER_374_854 ();
 b15zdnd11an1n16x5 FILLER_374_886 ();
 b15zdnd11an1n08x5 FILLER_374_902 ();
 b15zdnd00an1n02x5 FILLER_374_910 ();
 b15zdnd00an1n01x5 FILLER_374_912 ();
 b15zdnd11an1n64x5 FILLER_374_944 ();
 b15zdnd11an1n64x5 FILLER_374_1008 ();
 b15zdnd11an1n08x5 FILLER_374_1072 ();
 b15zdnd00an1n02x5 FILLER_374_1080 ();
 b15zdnd11an1n64x5 FILLER_374_1124 ();
 b15zdnd11an1n64x5 FILLER_374_1188 ();
 b15zdnd11an1n64x5 FILLER_374_1252 ();
 b15zdnd11an1n64x5 FILLER_374_1316 ();
 b15zdnd11an1n64x5 FILLER_374_1380 ();
 b15zdnd11an1n32x5 FILLER_374_1444 ();
 b15zdnd11an1n16x5 FILLER_374_1476 ();
 b15zdnd11an1n08x5 FILLER_374_1492 ();
 b15zdnd00an1n02x5 FILLER_374_1500 ();
 b15zdnd11an1n16x5 FILLER_374_1544 ();
 b15zdnd11an1n08x5 FILLER_374_1560 ();
 b15zdnd00an1n02x5 FILLER_374_1568 ();
 b15zdnd00an1n01x5 FILLER_374_1570 ();
 b15zdnd11an1n64x5 FILLER_374_1613 ();
 b15zdnd11an1n64x5 FILLER_374_1677 ();
 b15zdnd11an1n16x5 FILLER_374_1741 ();
 b15zdnd11an1n08x5 FILLER_374_1757 ();
 b15zdnd11an1n04x5 FILLER_374_1765 ();
 b15zdnd00an1n01x5 FILLER_374_1769 ();
 b15zdnd11an1n64x5 FILLER_374_1784 ();
 b15zdnd11an1n64x5 FILLER_374_1848 ();
 b15zdnd11an1n64x5 FILLER_374_1912 ();
 b15zdnd11an1n64x5 FILLER_374_1976 ();
 b15zdnd11an1n64x5 FILLER_374_2040 ();
 b15zdnd11an1n32x5 FILLER_374_2104 ();
 b15zdnd11an1n16x5 FILLER_374_2136 ();
 b15zdnd00an1n02x5 FILLER_374_2152 ();
 b15zdnd11an1n64x5 FILLER_374_2162 ();
 b15zdnd11an1n32x5 FILLER_374_2226 ();
 b15zdnd11an1n16x5 FILLER_374_2258 ();
 b15zdnd00an1n02x5 FILLER_374_2274 ();
 b15zdnd11an1n64x5 FILLER_375_0 ();
 b15zdnd11an1n64x5 FILLER_375_64 ();
 b15zdnd11an1n64x5 FILLER_375_128 ();
 b15zdnd11an1n64x5 FILLER_375_192 ();
 b15zdnd11an1n64x5 FILLER_375_256 ();
 b15zdnd11an1n64x5 FILLER_375_320 ();
 b15zdnd11an1n64x5 FILLER_375_384 ();
 b15zdnd11an1n64x5 FILLER_375_448 ();
 b15zdnd11an1n64x5 FILLER_375_512 ();
 b15zdnd11an1n64x5 FILLER_375_576 ();
 b15zdnd11an1n64x5 FILLER_375_640 ();
 b15zdnd11an1n64x5 FILLER_375_704 ();
 b15zdnd11an1n64x5 FILLER_375_768 ();
 b15zdnd11an1n16x5 FILLER_375_832 ();
 b15zdnd11an1n08x5 FILLER_375_890 ();
 b15zdnd11an1n04x5 FILLER_375_898 ();
 b15zdnd00an1n02x5 FILLER_375_902 ();
 b15zdnd11an1n64x5 FILLER_375_920 ();
 b15zdnd11an1n64x5 FILLER_375_984 ();
 b15zdnd11an1n64x5 FILLER_375_1048 ();
 b15zdnd11an1n64x5 FILLER_375_1112 ();
 b15zdnd11an1n16x5 FILLER_375_1176 ();
 b15zdnd11an1n04x5 FILLER_375_1192 ();
 b15zdnd00an1n02x5 FILLER_375_1196 ();
 b15zdnd00an1n01x5 FILLER_375_1198 ();
 b15zdnd11an1n64x5 FILLER_375_1202 ();
 b15zdnd11an1n64x5 FILLER_375_1266 ();
 b15zdnd11an1n64x5 FILLER_375_1330 ();
 b15zdnd11an1n64x5 FILLER_375_1394 ();
 b15zdnd11an1n16x5 FILLER_375_1458 ();
 b15zdnd00an1n01x5 FILLER_375_1474 ();
 b15zdnd11an1n04x5 FILLER_375_1517 ();
 b15zdnd00an1n01x5 FILLER_375_1521 ();
 b15zdnd11an1n64x5 FILLER_375_1564 ();
 b15zdnd11an1n64x5 FILLER_375_1628 ();
 b15zdnd11an1n32x5 FILLER_375_1692 ();
 b15zdnd11an1n08x5 FILLER_375_1724 ();
 b15zdnd11an1n04x5 FILLER_375_1732 ();
 b15zdnd00an1n01x5 FILLER_375_1736 ();
 b15zdnd11an1n64x5 FILLER_375_1755 ();
 b15zdnd11an1n64x5 FILLER_375_1819 ();
 b15zdnd11an1n64x5 FILLER_375_1883 ();
 b15zdnd11an1n64x5 FILLER_375_1947 ();
 b15zdnd11an1n64x5 FILLER_375_2011 ();
 b15zdnd11an1n64x5 FILLER_375_2075 ();
 b15zdnd11an1n64x5 FILLER_375_2139 ();
 b15zdnd11an1n64x5 FILLER_375_2203 ();
 b15zdnd11an1n16x5 FILLER_375_2267 ();
 b15zdnd00an1n01x5 FILLER_375_2283 ();
 b15zdnd11an1n64x5 FILLER_376_8 ();
 b15zdnd11an1n64x5 FILLER_376_72 ();
 b15zdnd11an1n64x5 FILLER_376_136 ();
 b15zdnd11an1n64x5 FILLER_376_200 ();
 b15zdnd11an1n64x5 FILLER_376_264 ();
 b15zdnd11an1n64x5 FILLER_376_328 ();
 b15zdnd11an1n64x5 FILLER_376_392 ();
 b15zdnd11an1n64x5 FILLER_376_456 ();
 b15zdnd11an1n64x5 FILLER_376_520 ();
 b15zdnd11an1n64x5 FILLER_376_584 ();
 b15zdnd11an1n64x5 FILLER_376_648 ();
 b15zdnd11an1n04x5 FILLER_376_712 ();
 b15zdnd00an1n02x5 FILLER_376_716 ();
 b15zdnd11an1n16x5 FILLER_376_726 ();
 b15zdnd11an1n08x5 FILLER_376_742 ();
 b15zdnd00an1n01x5 FILLER_376_750 ();
 b15zdnd11an1n04x5 FILLER_376_793 ();
 b15zdnd11an1n04x5 FILLER_376_800 ();
 b15zdnd00an1n01x5 FILLER_376_804 ();
 b15zdnd11an1n32x5 FILLER_376_847 ();
 b15zdnd11an1n16x5 FILLER_376_879 ();
 b15zdnd11an1n08x5 FILLER_376_895 ();
 b15zdnd11an1n04x5 FILLER_376_903 ();
 b15zdnd00an1n02x5 FILLER_376_907 ();
 b15zdnd11an1n04x5 FILLER_376_921 ();
 b15zdnd11an1n04x5 FILLER_376_931 ();
 b15zdnd11an1n64x5 FILLER_376_946 ();
 b15zdnd11an1n64x5 FILLER_376_1010 ();
 b15zdnd11an1n64x5 FILLER_376_1074 ();
 b15zdnd11an1n16x5 FILLER_376_1138 ();
 b15zdnd11an1n08x5 FILLER_376_1154 ();
 b15zdnd00an1n02x5 FILLER_376_1162 ();
 b15zdnd11an1n04x5 FILLER_376_1204 ();
 b15zdnd11an1n64x5 FILLER_376_1211 ();
 b15zdnd11an1n64x5 FILLER_376_1275 ();
 b15zdnd11an1n32x5 FILLER_376_1339 ();
 b15zdnd11an1n08x5 FILLER_376_1371 ();
 b15zdnd11an1n04x5 FILLER_376_1379 ();
 b15zdnd00an1n01x5 FILLER_376_1383 ();
 b15zdnd11an1n64x5 FILLER_376_1399 ();
 b15zdnd11an1n32x5 FILLER_376_1463 ();
 b15zdnd11an1n16x5 FILLER_376_1495 ();
 b15zdnd00an1n01x5 FILLER_376_1511 ();
 b15zdnd11an1n04x5 FILLER_376_1554 ();
 b15zdnd00an1n02x5 FILLER_376_1558 ();
 b15zdnd00an1n01x5 FILLER_376_1560 ();
 b15zdnd11an1n64x5 FILLER_376_1603 ();
 b15zdnd11an1n64x5 FILLER_376_1667 ();
 b15zdnd11an1n32x5 FILLER_376_1731 ();
 b15zdnd11an1n16x5 FILLER_376_1763 ();
 b15zdnd11an1n04x5 FILLER_376_1779 ();
 b15zdnd11an1n04x5 FILLER_376_1787 ();
 b15zdnd11an1n64x5 FILLER_376_1796 ();
 b15zdnd11an1n64x5 FILLER_376_1860 ();
 b15zdnd11an1n64x5 FILLER_376_1924 ();
 b15zdnd11an1n64x5 FILLER_376_1988 ();
 b15zdnd11an1n64x5 FILLER_376_2052 ();
 b15zdnd11an1n32x5 FILLER_376_2116 ();
 b15zdnd11an1n04x5 FILLER_376_2148 ();
 b15zdnd00an1n02x5 FILLER_376_2152 ();
 b15zdnd11an1n64x5 FILLER_376_2162 ();
 b15zdnd11an1n32x5 FILLER_376_2226 ();
 b15zdnd11an1n16x5 FILLER_376_2258 ();
 b15zdnd00an1n02x5 FILLER_376_2274 ();
 b15zdnd11an1n64x5 FILLER_377_0 ();
 b15zdnd11an1n64x5 FILLER_377_64 ();
 b15zdnd11an1n64x5 FILLER_377_128 ();
 b15zdnd11an1n64x5 FILLER_377_192 ();
 b15zdnd11an1n64x5 FILLER_377_256 ();
 b15zdnd11an1n64x5 FILLER_377_320 ();
 b15zdnd11an1n64x5 FILLER_377_384 ();
 b15zdnd11an1n64x5 FILLER_377_448 ();
 b15zdnd11an1n64x5 FILLER_377_512 ();
 b15zdnd11an1n64x5 FILLER_377_576 ();
 b15zdnd11an1n64x5 FILLER_377_640 ();
 b15zdnd11an1n32x5 FILLER_377_704 ();
 b15zdnd11an1n16x5 FILLER_377_736 ();
 b15zdnd11an1n08x5 FILLER_377_752 ();
 b15zdnd11an1n04x5 FILLER_377_760 ();
 b15zdnd00an1n02x5 FILLER_377_764 ();
 b15zdnd00an1n01x5 FILLER_377_766 ();
 b15zdnd11an1n64x5 FILLER_377_809 ();
 b15zdnd11an1n32x5 FILLER_377_873 ();
 b15zdnd11an1n08x5 FILLER_377_905 ();
 b15zdnd11an1n04x5 FILLER_377_913 ();
 b15zdnd00an1n02x5 FILLER_377_917 ();
 b15zdnd00an1n01x5 FILLER_377_919 ();
 b15zdnd11an1n16x5 FILLER_377_933 ();
 b15zdnd11an1n08x5 FILLER_377_949 ();
 b15zdnd11an1n04x5 FILLER_377_957 ();
 b15zdnd11an1n64x5 FILLER_377_986 ();
 b15zdnd11an1n64x5 FILLER_377_1050 ();
 b15zdnd11an1n64x5 FILLER_377_1114 ();
 b15zdnd11an1n08x5 FILLER_377_1178 ();
 b15zdnd00an1n02x5 FILLER_377_1186 ();
 b15zdnd00an1n01x5 FILLER_377_1188 ();
 b15zdnd11an1n64x5 FILLER_377_1192 ();
 b15zdnd11an1n64x5 FILLER_377_1256 ();
 b15zdnd11an1n08x5 FILLER_377_1320 ();
 b15zdnd00an1n01x5 FILLER_377_1328 ();
 b15zdnd11an1n04x5 FILLER_377_1332 ();
 b15zdnd11an1n64x5 FILLER_377_1339 ();
 b15zdnd11an1n16x5 FILLER_377_1403 ();
 b15zdnd11an1n04x5 FILLER_377_1422 ();
 b15zdnd11an1n64x5 FILLER_377_1466 ();
 b15zdnd11an1n04x5 FILLER_377_1530 ();
 b15zdnd00an1n02x5 FILLER_377_1534 ();
 b15zdnd00an1n01x5 FILLER_377_1536 ();
 b15zdnd11an1n64x5 FILLER_377_1579 ();
 b15zdnd11an1n64x5 FILLER_377_1643 ();
 b15zdnd11an1n64x5 FILLER_377_1707 ();
 b15zdnd11an1n64x5 FILLER_377_1771 ();
 b15zdnd11an1n64x5 FILLER_377_1835 ();
 b15zdnd11an1n64x5 FILLER_377_1899 ();
 b15zdnd11an1n64x5 FILLER_377_1963 ();
 b15zdnd11an1n64x5 FILLER_377_2027 ();
 b15zdnd11an1n64x5 FILLER_377_2091 ();
 b15zdnd11an1n64x5 FILLER_377_2155 ();
 b15zdnd11an1n64x5 FILLER_377_2219 ();
 b15zdnd00an1n01x5 FILLER_377_2283 ();
 b15zdnd11an1n64x5 FILLER_378_8 ();
 b15zdnd11an1n64x5 FILLER_378_72 ();
 b15zdnd11an1n64x5 FILLER_378_136 ();
 b15zdnd11an1n64x5 FILLER_378_200 ();
 b15zdnd11an1n64x5 FILLER_378_264 ();
 b15zdnd11an1n64x5 FILLER_378_328 ();
 b15zdnd11an1n64x5 FILLER_378_392 ();
 b15zdnd11an1n64x5 FILLER_378_456 ();
 b15zdnd11an1n64x5 FILLER_378_520 ();
 b15zdnd11an1n64x5 FILLER_378_584 ();
 b15zdnd11an1n64x5 FILLER_378_648 ();
 b15zdnd11an1n04x5 FILLER_378_712 ();
 b15zdnd00an1n02x5 FILLER_378_716 ();
 b15zdnd11an1n08x5 FILLER_378_726 ();
 b15zdnd00an1n02x5 FILLER_378_734 ();
 b15zdnd11an1n08x5 FILLER_378_746 ();
 b15zdnd00an1n02x5 FILLER_378_754 ();
 b15zdnd00an1n01x5 FILLER_378_756 ();
 b15zdnd11an1n04x5 FILLER_378_797 ();
 b15zdnd11an1n64x5 FILLER_378_804 ();
 b15zdnd00an1n02x5 FILLER_378_868 ();
 b15zdnd11an1n64x5 FILLER_378_884 ();
 b15zdnd00an1n02x5 FILLER_378_948 ();
 b15zdnd00an1n01x5 FILLER_378_950 ();
 b15zdnd11an1n64x5 FILLER_378_971 ();
 b15zdnd11an1n32x5 FILLER_378_1035 ();
 b15zdnd00an1n02x5 FILLER_378_1067 ();
 b15zdnd00an1n01x5 FILLER_378_1069 ();
 b15zdnd11an1n64x5 FILLER_378_1073 ();
 b15zdnd11an1n04x5 FILLER_378_1137 ();
 b15zdnd00an1n01x5 FILLER_378_1141 ();
 b15zdnd11an1n04x5 FILLER_378_1168 ();
 b15zdnd11an1n04x5 FILLER_378_1196 ();
 b15zdnd11an1n64x5 FILLER_378_1203 ();
 b15zdnd11an1n32x5 FILLER_378_1267 ();
 b15zdnd11an1n08x5 FILLER_378_1299 ();
 b15zdnd11an1n04x5 FILLER_378_1307 ();
 b15zdnd11an1n32x5 FILLER_378_1363 ();
 b15zdnd00an1n01x5 FILLER_378_1395 ();
 b15zdnd11an1n16x5 FILLER_378_1448 ();
 b15zdnd11an1n04x5 FILLER_378_1464 ();
 b15zdnd00an1n01x5 FILLER_378_1468 ();
 b15zdnd11an1n64x5 FILLER_378_1475 ();
 b15zdnd11an1n64x5 FILLER_378_1539 ();
 b15zdnd11an1n64x5 FILLER_378_1603 ();
 b15zdnd11an1n64x5 FILLER_378_1667 ();
 b15zdnd11an1n64x5 FILLER_378_1731 ();
 b15zdnd11an1n64x5 FILLER_378_1795 ();
 b15zdnd11an1n64x5 FILLER_378_1859 ();
 b15zdnd11an1n64x5 FILLER_378_1923 ();
 b15zdnd11an1n64x5 FILLER_378_1987 ();
 b15zdnd11an1n64x5 FILLER_378_2051 ();
 b15zdnd11an1n32x5 FILLER_378_2115 ();
 b15zdnd11an1n04x5 FILLER_378_2147 ();
 b15zdnd00an1n02x5 FILLER_378_2151 ();
 b15zdnd00an1n01x5 FILLER_378_2153 ();
 b15zdnd11an1n64x5 FILLER_378_2162 ();
 b15zdnd11an1n32x5 FILLER_378_2226 ();
 b15zdnd11an1n16x5 FILLER_378_2258 ();
 b15zdnd00an1n02x5 FILLER_378_2274 ();
 b15zdnd11an1n64x5 FILLER_379_0 ();
 b15zdnd11an1n64x5 FILLER_379_64 ();
 b15zdnd11an1n64x5 FILLER_379_128 ();
 b15zdnd11an1n64x5 FILLER_379_192 ();
 b15zdnd11an1n64x5 FILLER_379_256 ();
 b15zdnd11an1n64x5 FILLER_379_320 ();
 b15zdnd11an1n64x5 FILLER_379_384 ();
 b15zdnd11an1n64x5 FILLER_379_448 ();
 b15zdnd11an1n64x5 FILLER_379_512 ();
 b15zdnd11an1n64x5 FILLER_379_576 ();
 b15zdnd11an1n32x5 FILLER_379_640 ();
 b15zdnd11an1n08x5 FILLER_379_672 ();
 b15zdnd11an1n04x5 FILLER_379_680 ();
 b15zdnd00an1n01x5 FILLER_379_684 ();
 b15zdnd11an1n04x5 FILLER_379_727 ();
 b15zdnd11an1n04x5 FILLER_379_751 ();
 b15zdnd11an1n64x5 FILLER_379_759 ();
 b15zdnd11an1n64x5 FILLER_379_823 ();
 b15zdnd00an1n02x5 FILLER_379_887 ();
 b15zdnd11an1n04x5 FILLER_379_920 ();
 b15zdnd11an1n04x5 FILLER_379_930 ();
 b15zdnd00an1n01x5 FILLER_379_934 ();
 b15zdnd11an1n16x5 FILLER_379_959 ();
 b15zdnd11an1n08x5 FILLER_379_975 ();
 b15zdnd11an1n04x5 FILLER_379_983 ();
 b15zdnd00an1n01x5 FILLER_379_987 ();
 b15zdnd11an1n16x5 FILLER_379_1019 ();
 b15zdnd11an1n08x5 FILLER_379_1035 ();
 b15zdnd11an1n32x5 FILLER_379_1095 ();
 b15zdnd11an1n16x5 FILLER_379_1127 ();
 b15zdnd11an1n08x5 FILLER_379_1143 ();
 b15zdnd00an1n01x5 FILLER_379_1151 ();
 b15zdnd11an1n04x5 FILLER_379_1159 ();
 b15zdnd00an1n01x5 FILLER_379_1163 ();
 b15zdnd11an1n04x5 FILLER_379_1216 ();
 b15zdnd11an1n16x5 FILLER_379_1223 ();
 b15zdnd11an1n08x5 FILLER_379_1239 ();
 b15zdnd00an1n01x5 FILLER_379_1247 ();
 b15zdnd11an1n64x5 FILLER_379_1262 ();
 b15zdnd11an1n08x5 FILLER_379_1326 ();
 b15zdnd00an1n02x5 FILLER_379_1334 ();
 b15zdnd00an1n01x5 FILLER_379_1336 ();
 b15zdnd11an1n04x5 FILLER_379_1340 ();
 b15zdnd11an1n04x5 FILLER_379_1352 ();
 b15zdnd11an1n16x5 FILLER_379_1398 ();
 b15zdnd11an1n04x5 FILLER_379_1417 ();
 b15zdnd11an1n08x5 FILLER_379_1424 ();
 b15zdnd00an1n01x5 FILLER_379_1432 ();
 b15zdnd11an1n64x5 FILLER_379_1450 ();
 b15zdnd11an1n64x5 FILLER_379_1514 ();
 b15zdnd11an1n64x5 FILLER_379_1578 ();
 b15zdnd11an1n64x5 FILLER_379_1642 ();
 b15zdnd11an1n64x5 FILLER_379_1706 ();
 b15zdnd11an1n04x5 FILLER_379_1770 ();
 b15zdnd11an1n64x5 FILLER_379_1778 ();
 b15zdnd11an1n64x5 FILLER_379_1842 ();
 b15zdnd11an1n64x5 FILLER_379_1906 ();
 b15zdnd11an1n64x5 FILLER_379_1970 ();
 b15zdnd11an1n64x5 FILLER_379_2034 ();
 b15zdnd11an1n64x5 FILLER_379_2098 ();
 b15zdnd11an1n64x5 FILLER_379_2162 ();
 b15zdnd11an1n32x5 FILLER_379_2226 ();
 b15zdnd11an1n16x5 FILLER_379_2258 ();
 b15zdnd11an1n08x5 FILLER_379_2274 ();
 b15zdnd00an1n02x5 FILLER_379_2282 ();
 b15zdnd11an1n64x5 FILLER_380_8 ();
 b15zdnd11an1n64x5 FILLER_380_72 ();
 b15zdnd11an1n64x5 FILLER_380_136 ();
 b15zdnd11an1n64x5 FILLER_380_200 ();
 b15zdnd11an1n64x5 FILLER_380_264 ();
 b15zdnd11an1n64x5 FILLER_380_328 ();
 b15zdnd11an1n64x5 FILLER_380_392 ();
 b15zdnd11an1n64x5 FILLER_380_456 ();
 b15zdnd11an1n64x5 FILLER_380_520 ();
 b15zdnd11an1n64x5 FILLER_380_584 ();
 b15zdnd11an1n32x5 FILLER_380_648 ();
 b15zdnd11an1n16x5 FILLER_380_680 ();
 b15zdnd11an1n08x5 FILLER_380_696 ();
 b15zdnd00an1n02x5 FILLER_380_704 ();
 b15zdnd00an1n02x5 FILLER_380_716 ();
 b15zdnd00an1n02x5 FILLER_380_726 ();
 b15zdnd11an1n32x5 FILLER_380_770 ();
 b15zdnd11an1n16x5 FILLER_380_802 ();
 b15zdnd11an1n08x5 FILLER_380_818 ();
 b15zdnd11an1n64x5 FILLER_380_868 ();
 b15zdnd11an1n16x5 FILLER_380_932 ();
 b15zdnd11an1n04x5 FILLER_380_948 ();
 b15zdnd00an1n02x5 FILLER_380_952 ();
 b15zdnd11an1n16x5 FILLER_380_958 ();
 b15zdnd11an1n04x5 FILLER_380_974 ();
 b15zdnd00an1n02x5 FILLER_380_978 ();
 b15zdnd11an1n16x5 FILLER_380_994 ();
 b15zdnd11an1n08x5 FILLER_380_1010 ();
 b15zdnd11an1n04x5 FILLER_380_1018 ();
 b15zdnd00an1n02x5 FILLER_380_1022 ();
 b15zdnd11an1n16x5 FILLER_380_1037 ();
 b15zdnd11an1n08x5 FILLER_380_1053 ();
 b15zdnd11an1n04x5 FILLER_380_1064 ();
 b15zdnd11an1n32x5 FILLER_380_1071 ();
 b15zdnd11an1n04x5 FILLER_380_1148 ();
 b15zdnd00an1n01x5 FILLER_380_1152 ();
 b15zdnd11an1n08x5 FILLER_380_1195 ();
 b15zdnd00an1n02x5 FILLER_380_1203 ();
 b15zdnd00an1n01x5 FILLER_380_1205 ();
 b15zdnd11an1n04x5 FILLER_380_1213 ();
 b15zdnd00an1n01x5 FILLER_380_1217 ();
 b15zdnd11an1n32x5 FILLER_380_1249 ();
 b15zdnd11an1n16x5 FILLER_380_1281 ();
 b15zdnd11an1n08x5 FILLER_380_1297 ();
 b15zdnd11an1n04x5 FILLER_380_1305 ();
 b15zdnd00an1n02x5 FILLER_380_1309 ();
 b15zdnd00an1n01x5 FILLER_380_1311 ();
 b15zdnd11an1n32x5 FILLER_380_1357 ();
 b15zdnd11an1n04x5 FILLER_380_1389 ();
 b15zdnd11an1n16x5 FILLER_380_1407 ();
 b15zdnd11an1n04x5 FILLER_380_1423 ();
 b15zdnd00an1n02x5 FILLER_380_1427 ();
 b15zdnd11an1n16x5 FILLER_380_1444 ();
 b15zdnd11an1n04x5 FILLER_380_1460 ();
 b15zdnd00an1n02x5 FILLER_380_1464 ();
 b15zdnd00an1n01x5 FILLER_380_1466 ();
 b15zdnd11an1n64x5 FILLER_380_1492 ();
 b15zdnd11an1n64x5 FILLER_380_1556 ();
 b15zdnd11an1n64x5 FILLER_380_1620 ();
 b15zdnd11an1n64x5 FILLER_380_1684 ();
 b15zdnd11an1n64x5 FILLER_380_1748 ();
 b15zdnd11an1n32x5 FILLER_380_1812 ();
 b15zdnd11an1n08x5 FILLER_380_1844 ();
 b15zdnd00an1n02x5 FILLER_380_1852 ();
 b15zdnd11an1n64x5 FILLER_380_1880 ();
 b15zdnd11an1n64x5 FILLER_380_1944 ();
 b15zdnd11an1n64x5 FILLER_380_2008 ();
 b15zdnd11an1n64x5 FILLER_380_2072 ();
 b15zdnd11an1n16x5 FILLER_380_2136 ();
 b15zdnd00an1n02x5 FILLER_380_2152 ();
 b15zdnd11an1n64x5 FILLER_380_2162 ();
 b15zdnd11an1n32x5 FILLER_380_2226 ();
 b15zdnd11an1n16x5 FILLER_380_2258 ();
 b15zdnd00an1n02x5 FILLER_380_2274 ();
 b15zdnd11an1n64x5 FILLER_381_0 ();
 b15zdnd11an1n64x5 FILLER_381_64 ();
 b15zdnd11an1n64x5 FILLER_381_128 ();
 b15zdnd11an1n64x5 FILLER_381_192 ();
 b15zdnd11an1n64x5 FILLER_381_256 ();
 b15zdnd11an1n64x5 FILLER_381_320 ();
 b15zdnd11an1n64x5 FILLER_381_384 ();
 b15zdnd11an1n64x5 FILLER_381_448 ();
 b15zdnd11an1n64x5 FILLER_381_512 ();
 b15zdnd11an1n64x5 FILLER_381_576 ();
 b15zdnd11an1n64x5 FILLER_381_640 ();
 b15zdnd11an1n04x5 FILLER_381_746 ();
 b15zdnd00an1n02x5 FILLER_381_750 ();
 b15zdnd00an1n01x5 FILLER_381_752 ();
 b15zdnd11an1n04x5 FILLER_381_795 ();
 b15zdnd00an1n02x5 FILLER_381_799 ();
 b15zdnd11an1n32x5 FILLER_381_804 ();
 b15zdnd11an1n16x5 FILLER_381_836 ();
 b15zdnd11an1n04x5 FILLER_381_852 ();
 b15zdnd11an1n64x5 FILLER_381_898 ();
 b15zdnd11an1n64x5 FILLER_381_962 ();
 b15zdnd11an1n32x5 FILLER_381_1026 ();
 b15zdnd11an1n16x5 FILLER_381_1058 ();
 b15zdnd11an1n08x5 FILLER_381_1074 ();
 b15zdnd00an1n02x5 FILLER_381_1082 ();
 b15zdnd11an1n08x5 FILLER_381_1129 ();
 b15zdnd00an1n01x5 FILLER_381_1137 ();
 b15zdnd11an1n04x5 FILLER_381_1180 ();
 b15zdnd11an1n08x5 FILLER_381_1210 ();
 b15zdnd00an1n02x5 FILLER_381_1218 ();
 b15zdnd11an1n04x5 FILLER_381_1265 ();
 b15zdnd11an1n16x5 FILLER_381_1289 ();
 b15zdnd11an1n04x5 FILLER_381_1305 ();
 b15zdnd11an1n32x5 FILLER_381_1327 ();
 b15zdnd11an1n08x5 FILLER_381_1359 ();
 b15zdnd11an1n04x5 FILLER_381_1367 ();
 b15zdnd00an1n02x5 FILLER_381_1371 ();
 b15zdnd11an1n04x5 FILLER_381_1418 ();
 b15zdnd00an1n01x5 FILLER_381_1422 ();
 b15zdnd11an1n64x5 FILLER_381_1433 ();
 b15zdnd11an1n08x5 FILLER_381_1497 ();
 b15zdnd00an1n01x5 FILLER_381_1505 ();
 b15zdnd11an1n64x5 FILLER_381_1537 ();
 b15zdnd11an1n64x5 FILLER_381_1601 ();
 b15zdnd11an1n64x5 FILLER_381_1665 ();
 b15zdnd11an1n64x5 FILLER_381_1729 ();
 b15zdnd11an1n64x5 FILLER_381_1793 ();
 b15zdnd11an1n08x5 FILLER_381_1857 ();
 b15zdnd11an1n64x5 FILLER_381_1872 ();
 b15zdnd11an1n64x5 FILLER_381_1936 ();
 b15zdnd11an1n64x5 FILLER_381_2000 ();
 b15zdnd11an1n64x5 FILLER_381_2064 ();
 b15zdnd11an1n64x5 FILLER_381_2128 ();
 b15zdnd11an1n64x5 FILLER_381_2192 ();
 b15zdnd11an1n16x5 FILLER_381_2256 ();
 b15zdnd11an1n08x5 FILLER_381_2272 ();
 b15zdnd11an1n04x5 FILLER_381_2280 ();
 b15zdnd11an1n64x5 FILLER_382_8 ();
 b15zdnd11an1n64x5 FILLER_382_72 ();
 b15zdnd11an1n64x5 FILLER_382_136 ();
 b15zdnd11an1n64x5 FILLER_382_200 ();
 b15zdnd11an1n64x5 FILLER_382_264 ();
 b15zdnd11an1n64x5 FILLER_382_328 ();
 b15zdnd11an1n64x5 FILLER_382_392 ();
 b15zdnd11an1n64x5 FILLER_382_456 ();
 b15zdnd11an1n64x5 FILLER_382_520 ();
 b15zdnd11an1n64x5 FILLER_382_584 ();
 b15zdnd11an1n32x5 FILLER_382_648 ();
 b15zdnd11an1n08x5 FILLER_382_680 ();
 b15zdnd11an1n08x5 FILLER_382_698 ();
 b15zdnd00an1n02x5 FILLER_382_716 ();
 b15zdnd00an1n02x5 FILLER_382_726 ();
 b15zdnd11an1n04x5 FILLER_382_740 ();
 b15zdnd00an1n01x5 FILLER_382_744 ();
 b15zdnd11an1n16x5 FILLER_382_787 ();
 b15zdnd11an1n08x5 FILLER_382_803 ();
 b15zdnd00an1n02x5 FILLER_382_811 ();
 b15zdnd00an1n01x5 FILLER_382_813 ();
 b15zdnd11an1n16x5 FILLER_382_820 ();
 b15zdnd00an1n01x5 FILLER_382_836 ();
 b15zdnd11an1n04x5 FILLER_382_848 ();
 b15zdnd11an1n64x5 FILLER_382_856 ();
 b15zdnd11an1n64x5 FILLER_382_920 ();
 b15zdnd11an1n32x5 FILLER_382_984 ();
 b15zdnd11an1n16x5 FILLER_382_1016 ();
 b15zdnd11an1n08x5 FILLER_382_1032 ();
 b15zdnd11an1n04x5 FILLER_382_1040 ();
 b15zdnd00an1n02x5 FILLER_382_1044 ();
 b15zdnd00an1n01x5 FILLER_382_1046 ();
 b15zdnd11an1n16x5 FILLER_382_1092 ();
 b15zdnd11an1n04x5 FILLER_382_1108 ();
 b15zdnd00an1n01x5 FILLER_382_1112 ();
 b15zdnd11an1n16x5 FILLER_382_1127 ();
 b15zdnd00an1n01x5 FILLER_382_1143 ();
 b15zdnd11an1n04x5 FILLER_382_1189 ();
 b15zdnd11an1n32x5 FILLER_382_1197 ();
 b15zdnd11an1n16x5 FILLER_382_1229 ();
 b15zdnd11an1n08x5 FILLER_382_1245 ();
 b15zdnd11an1n04x5 FILLER_382_1253 ();
 b15zdnd00an1n02x5 FILLER_382_1257 ();
 b15zdnd11an1n64x5 FILLER_382_1266 ();
 b15zdnd11an1n64x5 FILLER_382_1330 ();
 b15zdnd11an1n16x5 FILLER_382_1394 ();
 b15zdnd11an1n08x5 FILLER_382_1410 ();
 b15zdnd11an1n04x5 FILLER_382_1418 ();
 b15zdnd00an1n02x5 FILLER_382_1422 ();
 b15zdnd11an1n04x5 FILLER_382_1469 ();
 b15zdnd11an1n64x5 FILLER_382_1491 ();
 b15zdnd11an1n64x5 FILLER_382_1555 ();
 b15zdnd11an1n64x5 FILLER_382_1619 ();
 b15zdnd11an1n64x5 FILLER_382_1683 ();
 b15zdnd11an1n64x5 FILLER_382_1747 ();
 b15zdnd11an1n64x5 FILLER_382_1811 ();
 b15zdnd11an1n64x5 FILLER_382_1875 ();
 b15zdnd11an1n64x5 FILLER_382_1939 ();
 b15zdnd11an1n64x5 FILLER_382_2003 ();
 b15zdnd11an1n64x5 FILLER_382_2067 ();
 b15zdnd11an1n16x5 FILLER_382_2131 ();
 b15zdnd11an1n04x5 FILLER_382_2147 ();
 b15zdnd00an1n02x5 FILLER_382_2151 ();
 b15zdnd00an1n01x5 FILLER_382_2153 ();
 b15zdnd11an1n64x5 FILLER_382_2162 ();
 b15zdnd11an1n32x5 FILLER_382_2226 ();
 b15zdnd11an1n16x5 FILLER_382_2258 ();
 b15zdnd00an1n02x5 FILLER_382_2274 ();
 b15zdnd11an1n64x5 FILLER_383_0 ();
 b15zdnd11an1n64x5 FILLER_383_64 ();
 b15zdnd11an1n64x5 FILLER_383_128 ();
 b15zdnd11an1n64x5 FILLER_383_192 ();
 b15zdnd11an1n64x5 FILLER_383_256 ();
 b15zdnd11an1n64x5 FILLER_383_320 ();
 b15zdnd11an1n64x5 FILLER_383_384 ();
 b15zdnd11an1n64x5 FILLER_383_448 ();
 b15zdnd11an1n64x5 FILLER_383_512 ();
 b15zdnd11an1n64x5 FILLER_383_576 ();
 b15zdnd11an1n64x5 FILLER_383_640 ();
 b15zdnd00an1n02x5 FILLER_383_704 ();
 b15zdnd00an1n01x5 FILLER_383_706 ();
 b15zdnd11an1n04x5 FILLER_383_749 ();
 b15zdnd11an1n64x5 FILLER_383_795 ();
 b15zdnd11an1n32x5 FILLER_383_859 ();
 b15zdnd11an1n16x5 FILLER_383_891 ();
 b15zdnd11an1n08x5 FILLER_383_907 ();
 b15zdnd00an1n02x5 FILLER_383_915 ();
 b15zdnd11an1n64x5 FILLER_383_959 ();
 b15zdnd11an1n64x5 FILLER_383_1023 ();
 b15zdnd11an1n16x5 FILLER_383_1087 ();
 b15zdnd11an1n08x5 FILLER_383_1103 ();
 b15zdnd11an1n04x5 FILLER_383_1114 ();
 b15zdnd11an1n04x5 FILLER_383_1138 ();
 b15zdnd11an1n16x5 FILLER_383_1184 ();
 b15zdnd11an1n08x5 FILLER_383_1200 ();
 b15zdnd00an1n02x5 FILLER_383_1208 ();
 b15zdnd11an1n32x5 FILLER_383_1252 ();
 b15zdnd11an1n16x5 FILLER_383_1284 ();
 b15zdnd11an1n04x5 FILLER_383_1300 ();
 b15zdnd00an1n01x5 FILLER_383_1304 ();
 b15zdnd11an1n64x5 FILLER_383_1347 ();
 b15zdnd11an1n64x5 FILLER_383_1411 ();
 b15zdnd11an1n64x5 FILLER_383_1475 ();
 b15zdnd11an1n64x5 FILLER_383_1539 ();
 b15zdnd11an1n64x5 FILLER_383_1603 ();
 b15zdnd11an1n64x5 FILLER_383_1667 ();
 b15zdnd11an1n64x5 FILLER_383_1731 ();
 b15zdnd11an1n64x5 FILLER_383_1795 ();
 b15zdnd11an1n64x5 FILLER_383_1859 ();
 b15zdnd11an1n64x5 FILLER_383_1923 ();
 b15zdnd11an1n64x5 FILLER_383_1987 ();
 b15zdnd11an1n64x5 FILLER_383_2051 ();
 b15zdnd11an1n64x5 FILLER_383_2115 ();
 b15zdnd11an1n64x5 FILLER_383_2179 ();
 b15zdnd11an1n32x5 FILLER_383_2243 ();
 b15zdnd11an1n08x5 FILLER_383_2275 ();
 b15zdnd00an1n01x5 FILLER_383_2283 ();
 b15zdnd11an1n64x5 FILLER_384_8 ();
 b15zdnd11an1n64x5 FILLER_384_72 ();
 b15zdnd11an1n64x5 FILLER_384_136 ();
 b15zdnd11an1n64x5 FILLER_384_200 ();
 b15zdnd11an1n64x5 FILLER_384_264 ();
 b15zdnd11an1n64x5 FILLER_384_328 ();
 b15zdnd11an1n64x5 FILLER_384_392 ();
 b15zdnd11an1n64x5 FILLER_384_456 ();
 b15zdnd11an1n64x5 FILLER_384_520 ();
 b15zdnd11an1n64x5 FILLER_384_584 ();
 b15zdnd11an1n64x5 FILLER_384_648 ();
 b15zdnd11an1n04x5 FILLER_384_712 ();
 b15zdnd00an1n02x5 FILLER_384_716 ();
 b15zdnd00an1n02x5 FILLER_384_726 ();
 b15zdnd11an1n64x5 FILLER_384_770 ();
 b15zdnd11an1n64x5 FILLER_384_834 ();
 b15zdnd11an1n64x5 FILLER_384_898 ();
 b15zdnd11an1n64x5 FILLER_384_962 ();
 b15zdnd11an1n64x5 FILLER_384_1026 ();
 b15zdnd11an1n64x5 FILLER_384_1090 ();
 b15zdnd11an1n04x5 FILLER_384_1154 ();
 b15zdnd00an1n02x5 FILLER_384_1158 ();
 b15zdnd11an1n32x5 FILLER_384_1202 ();
 b15zdnd11an1n04x5 FILLER_384_1234 ();
 b15zdnd00an1n02x5 FILLER_384_1238 ();
 b15zdnd00an1n01x5 FILLER_384_1240 ();
 b15zdnd11an1n64x5 FILLER_384_1245 ();
 b15zdnd11an1n64x5 FILLER_384_1309 ();
 b15zdnd11an1n64x5 FILLER_384_1373 ();
 b15zdnd11an1n16x5 FILLER_384_1437 ();
 b15zdnd11an1n04x5 FILLER_384_1453 ();
 b15zdnd00an1n01x5 FILLER_384_1457 ();
 b15zdnd11an1n64x5 FILLER_384_1500 ();
 b15zdnd11an1n64x5 FILLER_384_1564 ();
 b15zdnd11an1n64x5 FILLER_384_1628 ();
 b15zdnd11an1n64x5 FILLER_384_1692 ();
 b15zdnd11an1n64x5 FILLER_384_1756 ();
 b15zdnd11an1n64x5 FILLER_384_1820 ();
 b15zdnd11an1n64x5 FILLER_384_1884 ();
 b15zdnd11an1n64x5 FILLER_384_1948 ();
 b15zdnd11an1n64x5 FILLER_384_2012 ();
 b15zdnd11an1n64x5 FILLER_384_2076 ();
 b15zdnd11an1n08x5 FILLER_384_2140 ();
 b15zdnd11an1n04x5 FILLER_384_2148 ();
 b15zdnd00an1n02x5 FILLER_384_2152 ();
 b15zdnd11an1n64x5 FILLER_384_2162 ();
 b15zdnd11an1n32x5 FILLER_384_2226 ();
 b15zdnd11an1n16x5 FILLER_384_2258 ();
 b15zdnd00an1n02x5 FILLER_384_2274 ();
 b15zdnd11an1n64x5 FILLER_385_0 ();
 b15zdnd11an1n64x5 FILLER_385_64 ();
 b15zdnd11an1n64x5 FILLER_385_128 ();
 b15zdnd11an1n64x5 FILLER_385_192 ();
 b15zdnd11an1n64x5 FILLER_385_256 ();
 b15zdnd11an1n64x5 FILLER_385_320 ();
 b15zdnd11an1n64x5 FILLER_385_384 ();
 b15zdnd11an1n64x5 FILLER_385_448 ();
 b15zdnd11an1n64x5 FILLER_385_512 ();
 b15zdnd11an1n64x5 FILLER_385_576 ();
 b15zdnd11an1n32x5 FILLER_385_640 ();
 b15zdnd11an1n16x5 FILLER_385_672 ();
 b15zdnd11an1n04x5 FILLER_385_688 ();
 b15zdnd00an1n02x5 FILLER_385_692 ();
 b15zdnd11an1n04x5 FILLER_385_736 ();
 b15zdnd00an1n01x5 FILLER_385_740 ();
 b15zdnd11an1n64x5 FILLER_385_783 ();
 b15zdnd11an1n64x5 FILLER_385_847 ();
 b15zdnd11an1n64x5 FILLER_385_911 ();
 b15zdnd11an1n64x5 FILLER_385_975 ();
 b15zdnd11an1n64x5 FILLER_385_1039 ();
 b15zdnd11an1n64x5 FILLER_385_1103 ();
 b15zdnd11an1n32x5 FILLER_385_1167 ();
 b15zdnd11an1n08x5 FILLER_385_1199 ();
 b15zdnd00an1n02x5 FILLER_385_1207 ();
 b15zdnd11an1n16x5 FILLER_385_1213 ();
 b15zdnd11an1n08x5 FILLER_385_1229 ();
 b15zdnd11an1n04x5 FILLER_385_1242 ();
 b15zdnd11an1n04x5 FILLER_385_1251 ();
 b15zdnd00an1n02x5 FILLER_385_1255 ();
 b15zdnd11an1n16x5 FILLER_385_1262 ();
 b15zdnd11an1n08x5 FILLER_385_1278 ();
 b15zdnd11an1n04x5 FILLER_385_1286 ();
 b15zdnd11an1n04x5 FILLER_385_1296 ();
 b15zdnd00an1n01x5 FILLER_385_1300 ();
 b15zdnd11an1n64x5 FILLER_385_1305 ();
 b15zdnd11an1n64x5 FILLER_385_1369 ();
 b15zdnd11an1n64x5 FILLER_385_1433 ();
 b15zdnd11an1n64x5 FILLER_385_1497 ();
 b15zdnd11an1n64x5 FILLER_385_1561 ();
 b15zdnd11an1n64x5 FILLER_385_1625 ();
 b15zdnd11an1n64x5 FILLER_385_1689 ();
 b15zdnd11an1n64x5 FILLER_385_1753 ();
 b15zdnd11an1n64x5 FILLER_385_1817 ();
 b15zdnd11an1n64x5 FILLER_385_1881 ();
 b15zdnd11an1n64x5 FILLER_385_1945 ();
 b15zdnd11an1n64x5 FILLER_385_2009 ();
 b15zdnd11an1n64x5 FILLER_385_2073 ();
 b15zdnd11an1n64x5 FILLER_385_2137 ();
 b15zdnd11an1n64x5 FILLER_385_2201 ();
 b15zdnd11an1n16x5 FILLER_385_2265 ();
 b15zdnd00an1n02x5 FILLER_385_2281 ();
 b15zdnd00an1n01x5 FILLER_385_2283 ();
 b15zdnd11an1n64x5 FILLER_386_8 ();
 b15zdnd11an1n64x5 FILLER_386_72 ();
 b15zdnd11an1n64x5 FILLER_386_136 ();
 b15zdnd11an1n64x5 FILLER_386_200 ();
 b15zdnd11an1n64x5 FILLER_386_264 ();
 b15zdnd11an1n64x5 FILLER_386_328 ();
 b15zdnd11an1n64x5 FILLER_386_392 ();
 b15zdnd11an1n64x5 FILLER_386_456 ();
 b15zdnd11an1n64x5 FILLER_386_520 ();
 b15zdnd11an1n64x5 FILLER_386_584 ();
 b15zdnd11an1n16x5 FILLER_386_648 ();
 b15zdnd11an1n08x5 FILLER_386_664 ();
 b15zdnd00an1n02x5 FILLER_386_672 ();
 b15zdnd00an1n02x5 FILLER_386_716 ();
 b15zdnd00an1n02x5 FILLER_386_726 ();
 b15zdnd00an1n01x5 FILLER_386_728 ();
 b15zdnd11an1n16x5 FILLER_386_733 ();
 b15zdnd11an1n08x5 FILLER_386_749 ();
 b15zdnd11an1n04x5 FILLER_386_757 ();
 b15zdnd00an1n01x5 FILLER_386_761 ();
 b15zdnd11an1n08x5 FILLER_386_766 ();
 b15zdnd11an1n04x5 FILLER_386_774 ();
 b15zdnd00an1n02x5 FILLER_386_778 ();
 b15zdnd00an1n01x5 FILLER_386_780 ();
 b15zdnd11an1n32x5 FILLER_386_786 ();
 b15zdnd11an1n16x5 FILLER_386_818 ();
 b15zdnd11an1n08x5 FILLER_386_834 ();
 b15zdnd00an1n02x5 FILLER_386_842 ();
 b15zdnd00an1n01x5 FILLER_386_844 ();
 b15zdnd11an1n08x5 FILLER_386_887 ();
 b15zdnd00an1n01x5 FILLER_386_895 ();
 b15zdnd11an1n64x5 FILLER_386_902 ();
 b15zdnd11an1n32x5 FILLER_386_966 ();
 b15zdnd11an1n16x5 FILLER_386_998 ();
 b15zdnd11an1n08x5 FILLER_386_1014 ();
 b15zdnd11an1n04x5 FILLER_386_1022 ();
 b15zdnd00an1n01x5 FILLER_386_1026 ();
 b15zdnd11an1n64x5 FILLER_386_1031 ();
 b15zdnd11an1n64x5 FILLER_386_1095 ();
 b15zdnd11an1n32x5 FILLER_386_1159 ();
 b15zdnd11an1n08x5 FILLER_386_1191 ();
 b15zdnd11an1n04x5 FILLER_386_1199 ();
 b15zdnd00an1n02x5 FILLER_386_1203 ();
 b15zdnd11an1n04x5 FILLER_386_1209 ();
 b15zdnd11an1n08x5 FILLER_386_1219 ();
 b15zdnd11an1n04x5 FILLER_386_1227 ();
 b15zdnd00an1n02x5 FILLER_386_1231 ();
 b15zdnd00an1n01x5 FILLER_386_1233 ();
 b15zdnd11an1n04x5 FILLER_386_1241 ();
 b15zdnd00an1n02x5 FILLER_386_1245 ();
 b15zdnd11an1n04x5 FILLER_386_1253 ();
 b15zdnd00an1n02x5 FILLER_386_1257 ();
 b15zdnd00an1n01x5 FILLER_386_1259 ();
 b15zdnd11an1n04x5 FILLER_386_1267 ();
 b15zdnd11an1n04x5 FILLER_386_1278 ();
 b15zdnd11an1n04x5 FILLER_386_1289 ();
 b15zdnd00an1n02x5 FILLER_386_1293 ();
 b15zdnd11an1n04x5 FILLER_386_1299 ();
 b15zdnd11an1n08x5 FILLER_386_1307 ();
 b15zdnd00an1n01x5 FILLER_386_1315 ();
 b15zdnd11an1n64x5 FILLER_386_1321 ();
 b15zdnd11an1n64x5 FILLER_386_1385 ();
 b15zdnd11an1n32x5 FILLER_386_1449 ();
 b15zdnd00an1n02x5 FILLER_386_1481 ();
 b15zdnd00an1n01x5 FILLER_386_1483 ();
 b15zdnd11an1n16x5 FILLER_386_1488 ();
 b15zdnd11an1n08x5 FILLER_386_1504 ();
 b15zdnd11an1n04x5 FILLER_386_1512 ();
 b15zdnd11an1n04x5 FILLER_386_1520 ();
 b15zdnd00an1n02x5 FILLER_386_1524 ();
 b15zdnd00an1n01x5 FILLER_386_1526 ();
 b15zdnd11an1n04x5 FILLER_386_1531 ();
 b15zdnd11an1n04x5 FILLER_386_1539 ();
 b15zdnd11an1n04x5 FILLER_386_1547 ();
 b15zdnd11an1n64x5 FILLER_386_1555 ();
 b15zdnd11an1n64x5 FILLER_386_1619 ();
 b15zdnd11an1n64x5 FILLER_386_1683 ();
 b15zdnd11an1n64x5 FILLER_386_1747 ();
 b15zdnd11an1n64x5 FILLER_386_1811 ();
 b15zdnd11an1n64x5 FILLER_386_1875 ();
 b15zdnd11an1n64x5 FILLER_386_1939 ();
 b15zdnd11an1n64x5 FILLER_386_2003 ();
 b15zdnd11an1n64x5 FILLER_386_2067 ();
 b15zdnd11an1n16x5 FILLER_386_2131 ();
 b15zdnd11an1n04x5 FILLER_386_2147 ();
 b15zdnd00an1n02x5 FILLER_386_2151 ();
 b15zdnd00an1n01x5 FILLER_386_2153 ();
 b15zdnd11an1n64x5 FILLER_386_2162 ();
 b15zdnd11an1n32x5 FILLER_386_2226 ();
 b15zdnd11an1n16x5 FILLER_386_2258 ();
 b15zdnd00an1n02x5 FILLER_386_2274 ();
 b15zdnd11an1n64x5 FILLER_387_0 ();
 b15zdnd11an1n64x5 FILLER_387_64 ();
 b15zdnd11an1n64x5 FILLER_387_128 ();
 b15zdnd11an1n64x5 FILLER_387_192 ();
 b15zdnd11an1n64x5 FILLER_387_256 ();
 b15zdnd11an1n64x5 FILLER_387_320 ();
 b15zdnd11an1n64x5 FILLER_387_384 ();
 b15zdnd11an1n64x5 FILLER_387_448 ();
 b15zdnd11an1n64x5 FILLER_387_512 ();
 b15zdnd11an1n64x5 FILLER_387_576 ();
 b15zdnd11an1n32x5 FILLER_387_640 ();
 b15zdnd11an1n04x5 FILLER_387_672 ();
 b15zdnd00an1n01x5 FILLER_387_676 ();
 b15zdnd11an1n04x5 FILLER_387_681 ();
 b15zdnd11an1n04x5 FILLER_387_689 ();
 b15zdnd11an1n04x5 FILLER_387_697 ();
 b15zdnd11an1n04x5 FILLER_387_705 ();
 b15zdnd11an1n04x5 FILLER_387_751 ();
 b15zdnd00an1n02x5 FILLER_387_755 ();
 b15zdnd11an1n64x5 FILLER_387_799 ();
 b15zdnd11an1n04x5 FILLER_387_863 ();
 b15zdnd11an1n16x5 FILLER_387_871 ();
 b15zdnd11an1n08x5 FILLER_387_887 ();
 b15zdnd11an1n04x5 FILLER_387_895 ();
 b15zdnd00an1n01x5 FILLER_387_899 ();
 b15zdnd11an1n32x5 FILLER_387_906 ();
 b15zdnd11an1n16x5 FILLER_387_938 ();
 b15zdnd00an1n02x5 FILLER_387_954 ();
 b15zdnd11an1n32x5 FILLER_387_963 ();
 b15zdnd11an1n16x5 FILLER_387_995 ();
 b15zdnd11an1n08x5 FILLER_387_1011 ();
 b15zdnd11an1n04x5 FILLER_387_1019 ();
 b15zdnd00an1n02x5 FILLER_387_1023 ();
 b15zdnd00an1n01x5 FILLER_387_1025 ();
 b15zdnd11an1n32x5 FILLER_387_1034 ();
 b15zdnd00an1n02x5 FILLER_387_1066 ();
 b15zdnd11an1n16x5 FILLER_387_1075 ();
 b15zdnd11an1n08x5 FILLER_387_1091 ();
 b15zdnd11an1n04x5 FILLER_387_1103 ();
 b15zdnd11an1n04x5 FILLER_387_1111 ();
 b15zdnd11an1n08x5 FILLER_387_1119 ();
 b15zdnd00an1n01x5 FILLER_387_1127 ();
 b15zdnd11an1n16x5 FILLER_387_1134 ();
 b15zdnd11an1n08x5 FILLER_387_1150 ();
 b15zdnd11an1n04x5 FILLER_387_1158 ();
 b15zdnd00an1n02x5 FILLER_387_1162 ();
 b15zdnd11an1n16x5 FILLER_387_1168 ();
 b15zdnd11an1n04x5 FILLER_387_1184 ();
 b15zdnd00an1n02x5 FILLER_387_1188 ();
 b15zdnd00an1n01x5 FILLER_387_1190 ();
 b15zdnd11an1n04x5 FILLER_387_1195 ();
 b15zdnd11an1n04x5 FILLER_387_1205 ();
 b15zdnd11an1n04x5 FILLER_387_1213 ();
 b15zdnd11an1n08x5 FILLER_387_1224 ();
 b15zdnd11an1n04x5 FILLER_387_1243 ();
 b15zdnd00an1n02x5 FILLER_387_1247 ();
 b15zdnd11an1n04x5 FILLER_387_1255 ();
 b15zdnd00an1n02x5 FILLER_387_1259 ();
 b15zdnd00an1n01x5 FILLER_387_1261 ();
 b15zdnd11an1n04x5 FILLER_387_1282 ();
 b15zdnd11an1n04x5 FILLER_387_1292 ();
 b15zdnd11an1n04x5 FILLER_387_1302 ();
 b15zdnd11an1n04x5 FILLER_387_1311 ();
 b15zdnd11an1n64x5 FILLER_387_1321 ();
 b15zdnd11an1n32x5 FILLER_387_1385 ();
 b15zdnd00an1n02x5 FILLER_387_1417 ();
 b15zdnd11an1n04x5 FILLER_387_1423 ();
 b15zdnd00an1n02x5 FILLER_387_1427 ();
 b15zdnd00an1n01x5 FILLER_387_1429 ();
 b15zdnd11an1n04x5 FILLER_387_1435 ();
 b15zdnd11an1n08x5 FILLER_387_1443 ();
 b15zdnd11an1n16x5 FILLER_387_1456 ();
 b15zdnd11an1n04x5 FILLER_387_1472 ();
 b15zdnd11an1n04x5 FILLER_387_1480 ();
 b15zdnd00an1n02x5 FILLER_387_1484 ();
 b15zdnd00an1n01x5 FILLER_387_1486 ();
 b15zdnd11an1n04x5 FILLER_387_1491 ();
 b15zdnd11an1n08x5 FILLER_387_1499 ();
 b15zdnd11an1n04x5 FILLER_387_1507 ();
 b15zdnd00an1n01x5 FILLER_387_1511 ();
 b15zdnd11an1n04x5 FILLER_387_1554 ();
 b15zdnd11an1n04x5 FILLER_387_1562 ();
 b15zdnd11an1n04x5 FILLER_387_1570 ();
 b15zdnd11an1n08x5 FILLER_387_1578 ();
 b15zdnd00an1n02x5 FILLER_387_1586 ();
 b15zdnd00an1n01x5 FILLER_387_1588 ();
 b15zdnd11an1n64x5 FILLER_387_1631 ();
 b15zdnd11an1n64x5 FILLER_387_1695 ();
 b15zdnd11an1n64x5 FILLER_387_1759 ();
 b15zdnd11an1n64x5 FILLER_387_1823 ();
 b15zdnd11an1n64x5 FILLER_387_1887 ();
 b15zdnd11an1n64x5 FILLER_387_1951 ();
 b15zdnd11an1n64x5 FILLER_387_2015 ();
 b15zdnd11an1n64x5 FILLER_387_2079 ();
 b15zdnd11an1n64x5 FILLER_387_2143 ();
 b15zdnd11an1n64x5 FILLER_387_2207 ();
 b15zdnd11an1n08x5 FILLER_387_2271 ();
 b15zdnd11an1n04x5 FILLER_387_2279 ();
 b15zdnd00an1n01x5 FILLER_387_2283 ();
 b15zdnd11an1n64x5 FILLER_388_8 ();
 b15zdnd11an1n64x5 FILLER_388_72 ();
 b15zdnd11an1n64x5 FILLER_388_136 ();
 b15zdnd11an1n64x5 FILLER_388_200 ();
 b15zdnd11an1n64x5 FILLER_388_264 ();
 b15zdnd11an1n64x5 FILLER_388_328 ();
 b15zdnd11an1n64x5 FILLER_388_392 ();
 b15zdnd11an1n64x5 FILLER_388_456 ();
 b15zdnd11an1n64x5 FILLER_388_520 ();
 b15zdnd11an1n64x5 FILLER_388_584 ();
 b15zdnd11an1n16x5 FILLER_388_648 ();
 b15zdnd00an1n02x5 FILLER_388_664 ();
 b15zdnd11an1n04x5 FILLER_388_670 ();
 b15zdnd00an1n02x5 FILLER_388_716 ();
 b15zdnd11an1n08x5 FILLER_388_726 ();
 b15zdnd11an1n04x5 FILLER_388_738 ();
 b15zdnd11an1n04x5 FILLER_388_746 ();
 b15zdnd11an1n04x5 FILLER_388_754 ();
 b15zdnd11an1n32x5 FILLER_388_800 ();
 b15zdnd00an1n01x5 FILLER_388_832 ();
 b15zdnd11an1n08x5 FILLER_388_837 ();
 b15zdnd11an1n08x5 FILLER_388_887 ();
 b15zdnd00an1n02x5 FILLER_388_895 ();
 b15zdnd11an1n04x5 FILLER_388_905 ();
 b15zdnd11an1n16x5 FILLER_388_917 ();
 b15zdnd11an1n08x5 FILLER_388_933 ();
 b15zdnd00an1n02x5 FILLER_388_941 ();
 b15zdnd00an1n01x5 FILLER_388_943 ();
 b15zdnd11an1n04x5 FILLER_388_950 ();
 b15zdnd00an1n01x5 FILLER_388_954 ();
 b15zdnd11an1n04x5 FILLER_388_961 ();
 b15zdnd00an1n02x5 FILLER_388_965 ();
 b15zdnd11an1n16x5 FILLER_388_972 ();
 b15zdnd11an1n04x5 FILLER_388_988 ();
 b15zdnd11an1n08x5 FILLER_388_1006 ();
 b15zdnd00an1n02x5 FILLER_388_1014 ();
 b15zdnd11an1n16x5 FILLER_388_1024 ();
 b15zdnd11an1n04x5 FILLER_388_1040 ();
 b15zdnd11an1n04x5 FILLER_388_1048 ();
 b15zdnd11an1n04x5 FILLER_388_1056 ();
 b15zdnd11an1n04x5 FILLER_388_1071 ();
 b15zdnd00an1n01x5 FILLER_388_1075 ();
 b15zdnd11an1n04x5 FILLER_388_1084 ();
 b15zdnd11an1n08x5 FILLER_388_1095 ();
 b15zdnd11an1n04x5 FILLER_388_1103 ();
 b15zdnd11an1n08x5 FILLER_388_1127 ();
 b15zdnd00an1n02x5 FILLER_388_1135 ();
 b15zdnd00an1n01x5 FILLER_388_1137 ();
 b15zdnd11an1n04x5 FILLER_388_1146 ();
 b15zdnd11an1n04x5 FILLER_388_1155 ();
 b15zdnd11an1n16x5 FILLER_388_1163 ();
 b15zdnd11an1n04x5 FILLER_388_1179 ();
 b15zdnd00an1n02x5 FILLER_388_1183 ();
 b15zdnd11an1n08x5 FILLER_388_1192 ();
 b15zdnd00an1n02x5 FILLER_388_1200 ();
 b15zdnd00an1n01x5 FILLER_388_1202 ();
 b15zdnd11an1n04x5 FILLER_388_1245 ();
 b15zdnd11an1n04x5 FILLER_388_1260 ();
 b15zdnd00an1n02x5 FILLER_388_1264 ();
 b15zdnd00an1n01x5 FILLER_388_1266 ();
 b15zdnd11an1n04x5 FILLER_388_1287 ();
 b15zdnd11an1n04x5 FILLER_388_1317 ();
 b15zdnd11an1n64x5 FILLER_388_1328 ();
 b15zdnd11an1n04x5 FILLER_388_1392 ();
 b15zdnd00an1n01x5 FILLER_388_1396 ();
 b15zdnd11an1n04x5 FILLER_388_1423 ();
 b15zdnd11an1n04x5 FILLER_388_1447 ();
 b15zdnd11an1n04x5 FILLER_388_1465 ();
 b15zdnd11an1n04x5 FILLER_388_1473 ();
 b15zdnd00an1n01x5 FILLER_388_1477 ();
 b15zdnd11an1n04x5 FILLER_388_1520 ();
 b15zdnd11an1n08x5 FILLER_388_1528 ();
 b15zdnd11an1n04x5 FILLER_388_1578 ();
 b15zdnd11an1n16x5 FILLER_388_1624 ();
 b15zdnd00an1n02x5 FILLER_388_1640 ();
 b15zdnd00an1n01x5 FILLER_388_1642 ();
 b15zdnd11an1n16x5 FILLER_388_1647 ();
 b15zdnd11an1n64x5 FILLER_388_1667 ();
 b15zdnd11an1n64x5 FILLER_388_1731 ();
 b15zdnd11an1n64x5 FILLER_388_1795 ();
 b15zdnd11an1n64x5 FILLER_388_1859 ();
 b15zdnd11an1n64x5 FILLER_388_1923 ();
 b15zdnd11an1n64x5 FILLER_388_1987 ();
 b15zdnd11an1n64x5 FILLER_388_2051 ();
 b15zdnd11an1n32x5 FILLER_388_2115 ();
 b15zdnd11an1n04x5 FILLER_388_2147 ();
 b15zdnd00an1n02x5 FILLER_388_2151 ();
 b15zdnd00an1n01x5 FILLER_388_2153 ();
 b15zdnd11an1n64x5 FILLER_388_2162 ();
 b15zdnd11an1n32x5 FILLER_388_2226 ();
 b15zdnd11an1n16x5 FILLER_388_2258 ();
 b15zdnd00an1n02x5 FILLER_388_2274 ();
 b15zdnd11an1n64x5 FILLER_389_0 ();
 b15zdnd11an1n64x5 FILLER_389_64 ();
 b15zdnd11an1n64x5 FILLER_389_128 ();
 b15zdnd11an1n64x5 FILLER_389_192 ();
 b15zdnd11an1n64x5 FILLER_389_256 ();
 b15zdnd11an1n64x5 FILLER_389_320 ();
 b15zdnd11an1n64x5 FILLER_389_384 ();
 b15zdnd11an1n64x5 FILLER_389_448 ();
 b15zdnd11an1n64x5 FILLER_389_512 ();
 b15zdnd11an1n04x5 FILLER_389_576 ();
 b15zdnd00an1n01x5 FILLER_389_580 ();
 b15zdnd11an1n64x5 FILLER_389_585 ();
 b15zdnd11an1n08x5 FILLER_389_649 ();
 b15zdnd00an1n02x5 FILLER_389_657 ();
 b15zdnd00an1n01x5 FILLER_389_659 ();
 b15zdnd11an1n08x5 FILLER_389_665 ();
 b15zdnd00an1n01x5 FILLER_389_673 ();
 b15zdnd11an1n04x5 FILLER_389_716 ();
 b15zdnd11an1n04x5 FILLER_389_762 ();
 b15zdnd11an1n04x5 FILLER_389_808 ();
 b15zdnd00an1n02x5 FILLER_389_812 ();
 b15zdnd11an1n08x5 FILLER_389_818 ();
 b15zdnd11an1n04x5 FILLER_389_826 ();
 b15zdnd11an1n16x5 FILLER_389_834 ();
 b15zdnd11an1n08x5 FILLER_389_850 ();
 b15zdnd11an1n04x5 FILLER_389_865 ();
 b15zdnd11an1n04x5 FILLER_389_911 ();
 b15zdnd11an1n04x5 FILLER_389_921 ();
 b15zdnd11an1n04x5 FILLER_389_933 ();
 b15zdnd11an1n04x5 FILLER_389_945 ();
 b15zdnd11an1n08x5 FILLER_389_954 ();
 b15zdnd11an1n08x5 FILLER_389_967 ();
 b15zdnd00an1n01x5 FILLER_389_975 ();
 b15zdnd11an1n08x5 FILLER_389_982 ();
 b15zdnd00an1n02x5 FILLER_389_990 ();
 b15zdnd00an1n01x5 FILLER_389_992 ();
 b15zdnd11an1n16x5 FILLER_389_1004 ();
 b15zdnd11an1n04x5 FILLER_389_1031 ();
 b15zdnd11an1n08x5 FILLER_389_1039 ();
 b15zdnd00an1n02x5 FILLER_389_1047 ();
 b15zdnd11an1n04x5 FILLER_389_1055 ();
 b15zdnd11an1n04x5 FILLER_389_1067 ();
 b15zdnd11an1n08x5 FILLER_389_1082 ();
 b15zdnd00an1n02x5 FILLER_389_1090 ();
 b15zdnd11an1n04x5 FILLER_389_1100 ();
 b15zdnd11an1n16x5 FILLER_389_1146 ();
 b15zdnd00an1n02x5 FILLER_389_1162 ();
 b15zdnd11an1n04x5 FILLER_389_1168 ();
 b15zdnd11an1n04x5 FILLER_389_1176 ();
 b15zdnd00an1n01x5 FILLER_389_1180 ();
 b15zdnd11an1n04x5 FILLER_389_1186 ();
 b15zdnd00an1n02x5 FILLER_389_1190 ();
 b15zdnd00an1n01x5 FILLER_389_1192 ();
 b15zdnd11an1n04x5 FILLER_389_1235 ();
 b15zdnd00an1n02x5 FILLER_389_1239 ();
 b15zdnd00an1n01x5 FILLER_389_1241 ();
 b15zdnd11an1n08x5 FILLER_389_1284 ();
 b15zdnd00an1n02x5 FILLER_389_1292 ();
 b15zdnd11an1n08x5 FILLER_389_1336 ();
 b15zdnd11an1n04x5 FILLER_389_1348 ();
 b15zdnd11an1n04x5 FILLER_389_1363 ();
 b15zdnd11an1n32x5 FILLER_389_1375 ();
 b15zdnd11an1n16x5 FILLER_389_1407 ();
 b15zdnd00an1n02x5 FILLER_389_1423 ();
 b15zdnd00an1n01x5 FILLER_389_1425 ();
 b15zdnd11an1n04x5 FILLER_389_1468 ();
 b15zdnd11an1n04x5 FILLER_389_1514 ();
 b15zdnd11an1n04x5 FILLER_389_1560 ();
 b15zdnd11an1n04x5 FILLER_389_1606 ();
 b15zdnd11an1n16x5 FILLER_389_1614 ();
 b15zdnd11an1n04x5 FILLER_389_1630 ();
 b15zdnd00an1n02x5 FILLER_389_1634 ();
 b15zdnd00an1n01x5 FILLER_389_1636 ();
 b15zdnd11an1n32x5 FILLER_389_1679 ();
 b15zdnd11an1n16x5 FILLER_389_1711 ();
 b15zdnd00an1n02x5 FILLER_389_1727 ();
 b15zdnd11an1n64x5 FILLER_389_1734 ();
 b15zdnd11an1n64x5 FILLER_389_1798 ();
 b15zdnd11an1n64x5 FILLER_389_1862 ();
 b15zdnd11an1n64x5 FILLER_389_1926 ();
 b15zdnd11an1n64x5 FILLER_389_1990 ();
 b15zdnd11an1n64x5 FILLER_389_2054 ();
 b15zdnd11an1n64x5 FILLER_389_2118 ();
 b15zdnd11an1n64x5 FILLER_389_2182 ();
 b15zdnd11an1n32x5 FILLER_389_2246 ();
 b15zdnd11an1n04x5 FILLER_389_2278 ();
 b15zdnd00an1n02x5 FILLER_389_2282 ();
endmodule
