module trng_mapcore (
    input       valid,
    input       clk,
    input       rst_n,
    input  pllMap_pkg::pllmap2pll pllmap_i,
    output pllMap_pkg::pllmap2pll pllcontrol



);


endmodule