///////////////////////////////////////////////////////////////////////////////
// Intel Confidential                                                        
///////////////////////////////////////////////////////////////////////////////
// Copyright 2021 Intel Corporation.                                         
// The information contained herein is the proprietary and confidential      
// information of Intel or its licensors, and is supplied subject to, and    
// may be used only in accordance with, previously executed agreements       
// with Intel ,                                                                                                   
// EXCEPT AS MAY OTHERWISE BE AGREED IN WRITING:                            
// (1) ALL MATERIALS FURNISHED BY INTEL HEREUNDER ARE PROVIDED "AS IS"      
//      WITHOUT WARRANTY OF ANY KIND;                            
// (2) INTEL SPECIFICALLY DISCLAIMS ANY WARRANTY OF NONINFRINGEMENT, FITNESS 
//      FOR A PARTICULAR PURPOSE OR MERCHANTABILITY; AND                     
// (3) INTEL WILL NOT BE LIABLE FOR ANY COSTS OF PROCUREMENT OF SUBSTITUTES, 
//      LOSS OF PROFITS, INTERRUPTION OF BUSINESS, OR                       
//      FOR ANY OTHER SPECIAL, CONSEQUENTIAL OR INCIDENTAL DAMAGES,        
//      HOWEVER CAUSED, WHETHER FOR BREACH OF WARRANTY, CONTRACT,            
//      TORT, NEGLIGENCE, STRICT LIABILITY OR OTHERWISE.

//##module names of all CBBs are changed 
//
// Model built by create_model on Thu Oct  5 15:55:22 CDT 2017
//
// collage-pragma translate_off
`timescale 1ps / 1ps
//=============================================================================
//
// Description:
//   <Enter Description Here>
//
//=============================================================================
`ifndef ip2211ringpll_SOC_MACROS_VH
`define ip2211ringpll_SOC_MACROS_VH

////`include "vlv_macro_tech_map.vh"
`ifndef ip2211ringpll_SVA_OFF
// //`include "intel_checkers.sv"
`endif

`define ip2211ringpll_RST_LATCH_P(q,i,clock,rst)                           \
`ifdef INTC_SIM                                                   \
   `ifdef  ip2211ringpll_MACRO_ATTRIBUTE                                   \
      `undef ip2211ringpll_MACRO_ATTRIBUTE                                 \
      `ip2211ringpll_RST_LATCH(q,i,(~(clock)),rst)                         \
      `define ip2211ringpll_MACRO_ATTRIBUTE                                \
   `else                                                     \
      `ip2211ringpll_RST_LATCH(q,i,(~(clock)),rst)                         \
   `endif                                                    \
`else                                                        \
  logic \clkb_``q;                                           \
  `ip2211ringpll_CLKINV(\clkb_``q,(clock))                                 \
  `ip2211ringpll_RST_LATCH(q,i,\clkb_``q,rst)                              \
`endif


//THIS macro is causing problems during synthesis, use ip2211ringpll_LATCH_P instead

//`define ASYNC_RST_LATCH_P(q,i,clock,rst)                      \
//   always_latch                                             \
//      begin                                                 \
//         if      (~rst) q <= '0; /* lintra s-30529 */        \
//         else if (clock) q <= i;                            \
//      end /* lintra s-30500 */






//// New inverter for top level tie-offs
//// Usage is only for top level tie-offs so inverter won't be optimized away by synthesis
//`define INV_PRSRV(outb,in)                                          \
//`ifdef INTC_DC                                                           \
//     `LIB_INV_PRSRV(outb,in)                                        \
//`else                                                               \
//  assign outb = ~in ;     /* lintra s-35000, s-35006 */             \
//`endif          

//New macros for top level tie-offs
`define ip2211ringpll_TIEOFF_0_PRSRV(out)                                        \
`ifdef INTC_DC                                                          \
   `LIB_TIEOFF_0_PRSRV(out)  /* lintra s-30516 */                  \
`else                                                              \
   assign out = {$bits(out){1'b0}};                                \
`endif                                                             

`define ip2211ringpll_TIEOFF_1_PRSRV(out)                                        \
`ifdef INTC_DC                                                          \
   `LIB_TIEOFF_1_PRSRV(out) /* lintra s-30516 */                   \
`else                                                              \
   assign out = {$bits(out){1'b1}};                                \
`endif 








///============================================================================================
///
/// Flops and Drivers
///
///============================================================================================

// ip2211ringpll_MSFF macros:
//
// The standard ip2211ringpll_MSFF takes as its input both the gridclk and its counterpart clock enable. In real circuit
// implementation, these two signals ANDed together will give you your gated clock.
//
// If you create your own clock, (you are not using the MAKE_CLK_ENABLE() macro) then tie the clken off with 1'b1 as its
// input. Otherwise use the MAKE_CLK_ENABLE() macro and use gridclock as your clk input.
//
// If you are flopping an L phase signal, be sure to pass in ~gridclk as your clk and an L phase clken. The L phase
// clken should be created with the MAKE_CLK_ENABLE() macro, with all inputs of L phase.
//
`define ip2211ringpll_MSFF(q,i,clock)                                     \
   always_ff @(posedge clock)                               \
      begin                                                 \
         q <= i;                                            \
      end                                                   \
/* lintra s-30500 */

`define ip2211ringpll_MSFF_BLK(q,i,clock)                                 \
   logic [$bits(i)-1:0] \``dlyin_``q ;                      \
   assign  \``dlyin_``q = i;                                \
   always_ff @(posedge clock)                               \
      begin                                                 \
         q = \``dlyin_``q ;                                 \
      end                                                   \
/* lintra s-30500, s-31501, s-30531 */                      \

`define ip2211ringpll_MSFF_P(q,i,clock)                                   \
   always_ff @(negedge clock)                               \
      begin                                                 \
         q <= i;                                            \
      end                                                   \
/* lintra s-30500 */

`define ip2211ringpll_EN_MSFF(q,i,clock,enable)                           \
   always_ff @(posedge clock)                               \
      begin                                                 \
         if (enable) q <= i;                                \
       end                                                  \
/* lintra s-30500 */

`define ip2211ringpll_RST_MSFF(q,i,clock,rst)                             \
   always_ff @(posedge clock)                               \
      begin                                                 \
         if (rst) q <= '0;                                  \
         else     q <=  i;                                  \
      end                                                   \
/* lintra s-30500 */


`define ip2211ringpll_SET_MSFF(q,i,clock,set)                             \
   always_ff @(posedge clock)                               \
      begin                                                 \
         if (set) q <= {$bits(q){1'b1}};                    \
         else     q <=  i;                                  \
      end                                                   \
/* lintra s-30500 */                                        \


`define ip2211ringpll_RST_MSFF_P(q,i,clock,rst)                           \
   always_ff @(negedge clock)                               \
      begin                                                 \
         if (rst) q <= '0;                                  \
         else     q <=  i;                                  \
      end

`define ip2211ringpll_EN_RST_MSFF(q,i,clock,enable,rst)                   \
   always_ff @(posedge clock )                              \
      begin                                                 \
         if ( rst )         q <= '0 ;                       \
         else if ( enable ) q <= i ;                        \
      end                                                   \

/* lintra s-30500 */

`define ip2211ringpll_EN_RST_MSFF_P(q,i,clock,enable,rst)                 \
   always_ff @(negedge clock )                              \
      begin                                                 \
         if ( rst )         q <= '0 ;                       \
         else if ( enable ) q <= i ;                        \
      end


`define ip2211ringpll_EN_SET_MSFF(q,i,clock,enable,set)                   \
   always_ff @(posedge clock)                               \
      begin                                                 \
         if (set)         q <=  {$bits(q){1'b1}};           \
         else if (enable) q <=  i;                          \
      end                                                   \
/* lintra s-30500 */

`define ip2211ringpll_ASYNC_RST_MSFF(q,i,clock,rst)                       \
logic \``q``_rst ;                                           \
assign \``q``_rst = rst ;                                   \
   always_ff @(posedge clock or posedge \``q``_rst )        \
      begin                                                 \
         if ( \``q``_rst )  q <= '0;                        \
         else      q <= i;                                  \
      end                                                   \
/* lintra s-30500 */

`define ip2211ringpll_ASYNC_SET_MSFF(q,i,clock,set)                       \
   logic \``q``_set ;                                       \
   assign \``q``_set = set ;                                \
   always_ff @(posedge clock or posedge \``q``_set )        \
      begin                                                 \
         if (\``q``_set ) q <= {$bits(q){1'b1}};            \
         else                 q <= i;                       \
      end                                                   \
/* lintra s-30500, s-30531 */

`define ip2211ringpll_ASYNC_RST_MSFF_P(q,i,clock,rst)                     \
   always_ff @(negedge clock or posedge rst)                \
      begin                                                 \
         if (rst)  q <=  '0;                                \
         else      q <=  i;                                 \
   end

/* lintra s-30500, s-30531 */

`define ip2211ringpll_ASYNC_RSTD_MSFF(q,i,clock,rst,rstd)                 \
   always_ff @(posedge clock or posedge rst)                \
      begin                                                 \
         if (rst)  q <=  rstd;                              \
         else      q <=  i;                                 \
      end                                                   \
/* lintra s-30500 */

`define ip2211ringpll_EN_ASYNC_RSTD_MSFF(q,i,clock,enable,rst,rstd)       \
   always_ff @(posedge clock or posedge rst)                \
      begin                                                 \
         if (rst)  q <= rstd;                               \
         else if (enable) q <= i;                           \
      end                                                   \

/* lintra s-30500, s-30531 */

`define ip2211ringpll_ASYNC_SET_RST_MSFF(q,i,clock,set,rst)                \
   logic \``rst_``q ;                                        \
   logic \``set_``q ;                                        \
   assign \``rst_``q = rst ;                                 \
   assign \``set_``q = set ;                                 \
   always_ff @(posedge clock or posedge set or posedge rst ) \
      begin                                                  \
         if (rst)      q <=  {$bits(q){1'b0}};               \
         else if (set) q <=  {$bits(q){1'b1}};               \
         else                 q <= i;                        \
      end                                                   


/* lintra s-30500 */
`define ip2211ringpll_EN_ASYNC_RST_MSFF(q,i,clock,enable,rst)               \
   logic [$bits(i)-1:0] \``dlyin_``q ;                        \
   logic \``dlyen_``q ;                                       \
   assign  \``dlyin_``q = i;                                  \
   assign  \``dlyen_``q = enable;                             \
   always_ff @(posedge clock or posedge rst)                  \
      begin                                                   \
         if (rst)     q <=  '0;                                \
         else if (\``dlyen_``q ) q <=  \``dlyin_``q ;          \
      end                                                     \



///============================================================================================
///           META STABLE 2 ip2211ringpll_FLOP MACROS 
///============================================================================================
//`LIB_ASYNC_RST_2MSFF_META(q,i,clk,rstb) 

`define ip2211ringpll_ASYNC_RST_2MSFF_META(q,i,clkin,rst_b)                     \
//`ifdef INTC_DC                                                      \
//  ctech_lib_msff_async_rst_meta ctech_lib_msff_async_rst_meta_``q``(.o(q),.d(i),.clk(clkin),.rst(!rstb));  \
//`else                                                          \
`ifdef INTC_DC                                                      \
 ctech_lib_doublesync_rstb ctech_lib_doublesync_rstb``q``(.o(q),.d(i),.clk(clkin),.rstb(rst_b));  \
  //ctech_lib_doublesync_setb ctech_lib_doublesync_setb``q``(.o(q),.d(i),.clk(clkin),.setb(rstb));  \
`else                                                          \
 logic [$bits(i)-1:0] \``staged_``q ;                         \
  always_ff @(posedge clkin or negedge rst_b ) begin              \
    if ( ~rst_b )       \``staged_``q <= '0;                    \
    else               \``staged_``q <=  i;                    \
  end                                                          \
  always_ff @(posedge clkin or negedge rst_b) begin               \
    if ( ~rst_b )       q <= '0;                                \
    else               q <=  \``staged_``q ;                   \
  end                                                          \
`endif                                                         \

/* lintra s-30500 */

//`define ip2211ringpll_ASYNC_RST_2MSFF_META(q,i,clkin,rst_b)                     \
//ctech_lib_doublesync_rstb ctech_lib_doublesync_rstb``q``(.o(q),.d(i),.clk(clkin),.rstb(rst_b));

`define ip2211ringpll_CLKGATE_TE(q,cp,enab,tenab) \
`ifdef INTC_DC \
b15cilb81al1n02x5 ``q``clk_gate_tdr_data_out_reg_latch (.clkout(q), .clk(cp), .en(enab), .te(tenab));  \
`else \
logic ``q``_clko; \
always_latch  \
    begin \
      if (cp) ``q``_clko <= ~(enab|tenab); \
    end   \
assign q = ``q``_clko  | cp;       \
`endif

//`LIB_ASYNC_SET_2MSFF_META(q,i,clk,psb)
`define ip2211ringpll_ASYNC_SET_2MSFF_META(q,i,clkin,psb)                      \
//`ifdef INTC_DC                                                      \
//   ctech_lib_msff_async_set_meta ctech_lib_msff_async_set_meta_``q``(.o(q),.d(i),.clk(clkin),.set(!psb));\
//`else                                                          \
  logic [$bits(i)-1:0] \``staged_``q ;                         \
  always_ff @(posedge clkin or negedge psb ) begin               \
    if ( ~psb )        \``staged_``q <= '1;                    \
    else               \``staged_``q <=  i;                    \
  end                                                          \
  always_ff @(posedge clkin or negedge psb) begin                \
    if ( ~psb )        q <= '1;                                \
    else               q <=  \``staged_``q ;                   \
  end                                                          \
//`endif                                                         \
/* lintra s-30500 */



///============================================================================================
///          ADDING CLK BUFFER FOR TESTING
///============================================================================================
`define ip2211ringpll_CLK_BUF(clkout,clk)                     \
`ifdef INTC_DC                                                      \
  ctech_lib_clk_buf ctech_lib_clk_buf``clkout``(.clkout(clkout),.clk(clk));  \
`endif                                                         \
/* lintra s-30500 */



///============================================================================================
///           META STABLE ip2211ringpll_FLOP MACRO 
///============================================================================================
//***** NEEDS TO BE UPDATED BASED ON OUTCOME OF LIBRARY REQUEST *****
//`LIB_SOC_MSFF_META(q,i,clock)
`define ip2211ringpll_MSFF_META(q,i,clock)                                   \
//`ifdef INTC_DC                                                      \
//    ctech_lib_msff_meta_hard ctech_lib_msff_meta_hard_``q``(.o(q),.d(i),.clk(clock));   \
//`else                                                          \
 `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                        \
                                                               \
   `endif                                                      \
   always_ff @(posedge clock)                                  \
      begin                                                    \
         q <= i;                                               \
      end                                                      \
/* lintra s-30500 */                                           \
//`endif

//***** NEEDS TO BE UPDATED BASED ON OUTCOME OF LIBRARY REQUEST *****
/* lintra s-30500 */


`define ip2211ringpll_LATCH(q,i,clock)                                    \
   always_latch                                             \
      begin                                                 \
         if (clock) q <= i;                                 \
      end                                                   \
/* lintra s-30500 */

`define ip2211ringpll_LATCH_P(q,i,clock)                                  \
   always_latch                                             \
      begin                                                 \
         if (~clock) q <=  i;                               \
      end                                                   

`define ip2211ringpll_RST_LATCH(q,i,clock,rst)                            \
   always_latch                                             \
      begin                                                 \
         if (clock)                                         \
            if (rst) q <= '0;                               \
            else     q <=  i;                               \
      end                                                   \
/* lintra s-30500 */


`define ip2211ringpll_ASYNC_SET_LATCH(q,i,clock,set)                      \
   always_latch                                             \
     begin                                                  \
         if (set)          q <= '1; /* lintra s-30529 */    \
           else if (clock) q <=  i;                         \
             end                                            \
/* lintra s-30500 */

`define ip2211ringpll_ASYNC_RST_LATCH(q,i,clock,rst)                      \
   always_latch                                             \
      begin                                                 \
         if      (rst) q <= '0; /* lintra s-30529 */        \
         else if (clock) q <= i;                            \
      end /* lintra s-30500 */

`define ip2211ringpll_ASYNC_RST_LATCH_BLK(q,i,clock,rst)                  \
   always_latch                                             \
      begin                                                 \
         if      (rst) q = '0; /* lintra s-30529 */        \
         else if (clock) q = i;                             \
      end /* lintra s-30500 */

`define ip2211ringpll_EN_ASYNC_RST_LATCH(q,i,clock,enable,rst)            \
   always_latch                                             \
      begin                                                 \
         if      (rst)      q <= '0; /* lintra s-30529 */   \
         else if (clock & enable) q <=   i;                 \
      end /* lintra s-30500 */

/* lintra s-30500 */

`define ip2211ringpll_ASYNC_RSTD_LATCH_P(q,i,clock,rst,rstd) `ip2211ringpll_ASYNC_RSTD_LATCH(q,i,(~(clock)),rst,rstd)

`define ip2211ringpll_ASYNC_RSTD_LATCH(q,i,clock,rst,rstd)                \
   always_latch                                             \
      begin                                                 \
         if      (rst) q <= rstd;                           \
         else if (clock) q <=  i;                           \
      end                                                   \



/* lintra s-30500 */

`define ip2211ringpll_ASYNC_RST_SET(q,rst,set)                            \
  `ip2211ringpll_RST_LATCH(q,set,(set|rst),rst)

/* lintra s-30500 */

`define ip2211ringpll_LATCH_P_DESKEW(q,i,clock)                           \
   always_latch                                             \
      begin                                                 \
         if (~clock) q <=  i;                               \
      end                                                   \
/* lintra s-50500 */

`define ip2211ringpll_ASYNC_RST_MSFF_META(q,i,clk,rstb)                      \
`ifdef INTC_DC                                                      \
  `LIB_ASYNC_RST_MSFF_META(q,i,clk,rstb)                       \
`else                                                          \
                                                               \
  always_ff @(posedge clk or negedge rstb) begin               \
    if ( ~rstb )  q <= '0;                                     \
    else          q <=  i;                                     \
  end                                                          \
`endif                                                         \

// ----------------------------------
//  RESET DISTRIBUTION MACROS
// ----------------------------------
`define ip2211ringpll_MAKE_RST_DIST(irstoutb, iusyncout, iclk, irstinb, iusyncin) \
    ip2211ringpll_sync_rst_gen \``sync_rst_``irstoutb (                           \
         .rstoutb(irstoutb),                                        \
         .usyncout(iusyncout),                                      \
         .clk(iclk),                                                \
         .rstinb(irstinb),                                          \
         .usyncin(iusyncin)                                         \
   );                                                                  
/* lintra s-31500, s-33048, s-33049 */

///============================================================================================
///
/// IO Driver Macros
///
///============================================================================================
///
///
///   BUS TYPE MACRO                DESCRIPTION        UNDRIVEN VALUE* CONTENTION*
///  
///   TRI                         - Tri-State          'Z              Multiple Drivers

///   WAND                        - Wired-And          Weakpull 1      None 

///   WOR                         - Wired-Or           Weakpull 0      None 

///   *Semantics achieved only in conjunction with applicable, explict SUSTAIN, WEAKPULL, PRECHARGE, DRIVE macros
///    and relevant assertions
///
///   BUS DRIVER MACRO              DESCRIPTION
///
///   TRI_DRIVE     (Bus,En,Data) - Driver for busses of all Tri-State types
///   WAND_DRIVE    (Bus,En,Data) - WAND bus driver
///   WAND_WEAKPULL (Bus, En)     - WAND bus weak pull up
///   WOR_DRIVE     (Bus,En,Data) - WOR bus driver
///   WOR_WEAKPULL  (Bus, En)     - WOR bus weak pull down


`define ip2211ringpll_NO_SYNTH_WAND_WEAKPULL(Bus,En)                                                                   \
  `ifdef INTC_EMULATION                                                                                       \
        assign (weak1, highz0)   Bus = {$bits(Bus){1'b1}};                                               \
  `else                                                                                                  \
        assign (weak1, highz0)   Bus = En ? {$bits(Bus){1'b1}} : {$bits(Bus){1'bz}};                     \
  `endif

`define ip2211ringpll_NO_SYNTH_WAND_DRIVE(Bus,En,Data)                                                                 \
  `ifdef INTC_EMULATION                                                                                       \
        assign (strong0, highz1) Bus = En ? Data : {$bits(Bus){1'b1}};                                   \
  `else                                                                                                  \
        assign (strong0, highz1) Bus = En ? Data : {$bits(Bus){1'bz}};                                   \
  `endif

`define ip2211ringpll_NO_SYNTH_WOR_WEAKPULL(Bus,En)                                                                    \
  `ifdef INTC_EMULATION                                                                                       \
        assign (weak0, highz1)   Bus = {$bits(Bus){1'b0}};                                               \
  `else                                                                                                  \
        assign (weak0, highz1)   Bus = En ? {$bits(Bus){1'b0}} : {$bits(Bus){1'bz}};                     \
  `endif

`define ip2211ringpll_NO_SYNTH_WOR_DRIVE(Bus,En,Data)                                                                  \
  `ifdef INTC_EMULATION                                                                                       \
        assign (strong1, highz0) Bus = En ? Data : {$bits(Bus){1'b0}};                                   \
  `else                                                                                                  \
        assign (strong1, highz0) Bus = En ? Data : {$bits(Bus){1'bz}};                                   \
  `endif

`define ip2211ringpll_NO_SYNTH_WOR_TRI_DRIVE(Bus,En,Data) /* lintra s-50505 */                                         \
  `ifdef INTC_EMULATION                                                                                       \
        assign Bus = En ? Data : {$bits(Bus){1'b0}}; /* lintra s-23083 */                                \
  `else                                                                                                  \
        assign Bus = En ? Data : {$bits(Bus){1'bz}}; /* lintra s-23083 */                                \
  `endif



///============================================================================================

`define ip2211ringpll_SET_MSFF_BLK(q,i,clock,set)                                                                      \
   `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                                \
                                                                                                         \
   `endif                                                                                                \
   logic [$bits(i)-1:0] \``dlyin_``q ;                                                                   \
   logic \``dlyset_``q ;                                                                                 \
   assign  \``dlyin_``q = i;                                                                             \
   assign  \``dlyset_``q = set;                                                                          \
   always_ff @(posedge clock)                                                                            \
      begin                                                                                              \
         if ( \``dlyset_``q ) q = {$bits(q){1'b1}};                                                      \
         else     q =  \``dlyin_``q ;                                                                    \
      end    /* lintra s-30500, s-31501, s-30531 */
                                                      
`define ip2211ringpll_EN_RSTD_MSFF(q,i,clock,enable,rst,rstd)             \
   `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                   \
                                                            \
     `endif                                                 \
   always_ff @(posedge clock)                               \
      begin                                                 \
         if (rst)          q <=  rstd;                      \
         else if (enable)  q <=  i;                         \
      end /* lintra s-30500 */   
                                                     
//`define TRI_DRIVE(Bus,En,Data) /* lintra s-30505 */         \
//  `ifdef FALCON                                             \
//        assign Bus = {$bits(Bus){1'b1}};                    \
//      `else                                                 \
//        assign Bus = En ? Data : {$bits(Bus){1'bz}};        \
//  `endif

`define ip2211ringpll_MSFF_P_BLK(q,i,clock)                               \
   `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                   \
                                                            \
   `endif                                                   \
   logic [$bits(i)-1:0] \``dlyin_``q ;                      \
   assign  \``dlyin_``q = i;                                \
   always_ff @(negedge clock )                              \
      begin                                                 \
         q = \``dlyin_``q ;                                 \
      end /* lintra s-30500, s-30531 */

`define ip2211ringpll_ASYNC_RST_MSFF_BLK(q,i,clock,rst)                   \
   `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                   \
                                                            \
   `endif                                                   \
   logic [$bits(i)-1:0] \``dlyin_``q ;                      \
   assign  \``dlyin_``q = i;                                \
   wire \``q``_rst ;                                        \
   assign \``q``_rst = rst ;                                \
   always_ff @(posedge clock or posedge \``q``_rst )        \
      begin                                                 \
         if ( \``q``_rst )  q = '0;                         \
         else      q =  \``dlyin_``q ;                      \
      end /* lintra s-30500, s-31501, s-30531 */

///=====================================================================
/// sVID Macros - Should be Review , Aviel
///======================================================================  

`define ip2211ringpll_RSTD_MSFF(q,i,clock,rst,rstd)                 \
   always_ff @(posedge clock)                         \
      begin                                           \
         if (rst)  q <=  rstd;                        \
         else      q <= i;                            \
      end                                             \
/* lintra s-30500 */

`define ip2211ringpll_RSTD_MSFF_P(q,i,clock,rst,rstd)               \
   always_ff @(negedge clock)                         \
      begin                                           \
         if (rst)  q <=  rstd;                        \
         else      q <=  i;                           \
      end                                             \
/* lintra s-30500 */

// `define ip2211ringpll_RSTD_MSFF(q,i,clock,rst,rstd)                       \
// `ifdef SYNPLIFY_WA_COMPLEX_EVENT                            \
//    node \clock_``q ;                                        \
//    assign \clock_``q = clock ;                              \
//    always_ff @(posedge \clock_``q )                         \
//          if (rst) q <= rstd;                                \
//          else     q <=  i;                                  \
// `else                                                       \
// `ifdef INTC_SIM                                                  \
//    `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                   \
//                                                             \
//    `endif                                                   \
//    always_ff @(posedge clock)                               \
//       begin                                                 \
//          if (rst)                                           \
//             q <= rstd;                                      \
//          else                                               \
//             q <= i;                                         \
//       end                                                   \
// /* lintra s-30500 */                                        \
// `else                                                       \
//    node \``rst_``q ;                                        \
//    assign \``rst_``q = rst ;                                \
//    /* synopsys sync_set_reset `" \``rst_``q `" */           \
//    always_ff @(posedge  clock )                             \
//       begin                                                 \
//          if ( \``rst_``q )                                  \
//             q <= rstd;                                      \
//          else                                               \
//             q <= i;                                         \
//       end                                                   \
// `endif                                                      \
// `endif


`define ip2211ringpll_SET_RST_MSFF(q,i,clock,set,rst)                       \
   logic \``rst_``q ;                                         \
   logic \``set_``q ;                                         \
   assign \``rst_``q = rst ;                                  \
   assign \``set_``q = set ;                                  \
   always_ff @(posedge clock )                                \
      begin                                                   \
         if (rst)      q <=  {$bits(q){1'b0}};                \
         else if (set) q <=  {$bits(q){1'b1}};                \
         else          q <=  i;                               \
      end                                                   


// We currently don't have such library cells.
//
// `define ip2211ringpll_SET_RST_MSFF(q,i,clock,set,rst)                    \
// `ifdef INTC_SIM                                                 \
//    `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                  \
//                                                            \
//    `endif                                                  \
//    always_ff @(posedge clock)                              \
//       begin                                                \
//          if (rst)      q <= '0;                            \
//          else if (set) q <= '1;                            \
//          else          q <=  i;                            \
//       end                                                  \
// /* lintra s-30500 */                                       \
// `else                                                      \
//    node \``rst_``q ;                                       \
//    node \``set_``q ;                                       \
//    assign \``rst_``q = rst ;                               \
//    assign \``set_``q = set ;                               \
//    /* synopsys sync_set_reset `" \``rst_``q  , \``set_``q `" */ \
//    always_ff @(posedge clock )                             \
//       begin                                                \
//          if ( \``rst_``q )      q <= '0;                   \
//          else if ( \``set_``q ) q <= '1;                   \
//          else                 q <=  i;                     \
//       end                                                  \
// `endif



`define ip2211ringpll_RST_SET_MSFF(q,i,clock,rst,set)                       \
   logic \``rst_``q ;                                         \
   logic \``set_``q ;                                         \
   assign \``rst_``q = rst ;                                  \
   assign \``set_``q = set ;                                  \
   always_ff @(posedge clock )                                \
      begin                                                   \
         if (set)        q <=  {$bits(q){1'b1}};              \
         else if (rst)   q <=  {$bits(q){1'b0}};              \
         else            q <=  i;                             \
      end                                                   




// `define ip2211ringpll_RST_SET_MSFF(q,i,clock,rst,set)                      \
// `ifdef INTC_SIM                                                   \
//    `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                    \
//                                                              \
//    `endif                                                    \
//    always_ff @(posedge clock)                                \
//       begin                                                  \
//    `ifdef VAL4_OPTIMIZED                                     \
//        q <= (clock) ? ((set) ? '1 : ((rst) ? '0 : i)) : q;   \
//    `else                                                     \
//            if (set)      q <= '1;                            \
//            else if (rst) q <= '0;                            \
//            else          q <=  i;                            \
//    `endif                                                    \
//       end                                                    \
// `else                                                        \
// `ifdef INF                                                   \
//    node \rst_``q ;                                           \
//    node \set_``q ;                                           \
//    assign \rst_``q = (rst) ;                                 \
//    assign \set_``q = (set) ;                                 \
//    /* synopsys sync_set_reset `" \rst_``q  , \set_``q `" */  \
//    always_ff @(posedge clock )                               \
//       begin                                                  \
//          if ( \set_``q )      q <= {$bits(q){1'b1}};         \
//          else if ( \rst_``q ) q <= {$bits(q){1'b0}};         \
//          else                 q <=  i;                       \
//       end                                                    \
// `else                                                        \
//    localparam \w_``q = $bits(q);                             \
//    node [\w_``q -1:0] \qual_i_``q ;                          \
//    node [\w_``q -1:0] \ibit_``q ;                            \
//    yg0bfn00nn1d0 \ibbuf_``q <$typeof(q)> (.o(<(\ibit_``q )>),.a(<(i)>)); \
//    always_comb                                               \
//       if (set)   \qual_i_``q = {\w_``q  {1'b1}};             \
//       else                                                   \
//  if (rst) \qual_i_``q = {\w_``q  {1'b0}};                    \
//         else     \qual_i_``q = \ibit_``q ;                   \
//   /* synopsys keep_signal_name \``q  */                      \
//    `BASIC_FF \_reg``q <$typeof(q)> (.o(<(q)>),.clk(clock),.d(<(\qual_i_``q )>)); \
// `endif                                                       \
// `endif

///============================================================================================

/////////////////////////////////////////////////////////////////
// BEGIN - Multi-cycle path macros section
/////////////////////////////////////////////////////////////////


`define ip2211ringpll_MCP(MCP_source_sig, MCP_rx_enable, MCP_count_clk, MCP_rx_clk, phase_delay, macro_inst_name, clock_edges_aligned_at_destination, sampling_edge_or_phase) \
                                                                                                                                                                \
 `ifdef INTC_MCP_ON                                                                                                                                                  \
  logic signal_``macro_inst_name;                                                                                                                               \
  `ifndef ip2211ringpll_SVA_OFF                                                                                                                                               \
  SVA_``macro_inst_name : `ip2211ringpll_ASSERT_FORBIDDEN (signal_``macro_inst_name , 1'b0) `ip2211ringpll_ERR_MSG (`"MCP stability condition violated for assertion SVA_``macro_inst_name as MCP_source_sig was not stable for phase_delay phases before it was sampled`") ; \
  `endif                                                                                                                                                        \
                                                                                                                                                                \
  generate                                                                                                                                                      \
    if ((`"clock_edges_aligned_at_destination`" == "ALIGNED") && ((`"sampling_edge_or_phase`" == "RISING") || (`"sampling_edge_or_phase`" == "LOW")))           \
      soc_multi_cycle #(.N($bits(MCP_source_sig)), .PHASE(phase_delay), .CLOCKS_ALIGNED(1), .RX_SAMPLED_AT_POSEDGE(1)) mcpinst_``macro_inst_name (.out(signal_``macro_inst_name), .source_sig({>>{MCP_source_sig}}), .rx_clk(MCP_rx_clk), .rx_enable(MCP_rx_enable), .count_clk(MCP_count_clk)); \
    else if ((`"clock_edges_aligned_at_destination`" == "ALIGNED") && ((`"sampling_edge_or_phase`" == "FALLING") || (`"sampling_edge_or_phase`" == "HIGH")))    \
      soc_multi_cycle #(.N($bits(MCP_source_sig)), .PHASE(phase_delay), .CLOCKS_ALIGNED(1), .RX_SAMPLED_AT_POSEDGE(0)) mcpinst_``macro_inst_name (.out(signal_``macro_inst_name), .source_sig({>>{MCP_source_sig}}), .rx_clk(MCP_rx_clk), .rx_enable(MCP_rx_enable), .count_clk(MCP_count_clk)); \
    else if ((`"clock_edges_aligned_at_destination`" == "NOT_ALIGNED") && ((`"sampling_edge_or_phase`" == "RISING") || (`"sampling_edge_or_phase`" == "LOW")))  \
      soc_multi_cycle #(.N($bits(MCP_source_sig)), .PHASE(phase_delay), .CLOCKS_ALIGNED(0), .RX_SAMPLED_AT_POSEDGE(1)) mcpinst_``macro_inst_name (.out(signal_``macro_inst_name), .source_sig({>>{MCP_source_sig}}), .rx_clk(MCP_rx_clk), .rx_enable(MCP_rx_enable), .count_clk(MCP_count_clk)); \
    else if ((`"clock_edges_aligned_at_destination`" == "NOT_ALIGNED") && ((`"sampling_edge_or_phase`" == "FALLING") || (`"sampling_edge_or_phase`" == "HIGH"))) \
      soc_multi_cycle #(.N($bits(MCP_source_sig)), .PHASE(phase_delay), .CLOCKS_ALIGNED(0), .RX_SAMPLED_AT_POSEDGE(0)) mcpinst_``macro_inst_name (.out(signal_``macro_inst_name), .source_sig({>>{MCP_source_sig}}), .rx_clk(MCP_rx_clk), .rx_enable(MCP_rx_enable), .count_clk(MCP_count_clk)); \
    else                                                                                                                                                        \
      non_existent_mcp_module ip2211ringpll_bogus_mcp_instance();                                                                                                             \
  endgenerate                                                                                                                                                   \
`endif







/////////////////////////////////////////////////////////////////
// END - Multi-cycle path macros
/////////////////////////////////////////////////////////////////


// New Sequential definations... Lint friendly

`define ip2211ringpll_FLOP(_clk_,_rstB_,_in_,_out_) `ip2211ringpll_RST_MSFF(_out_,_in_,_clk_,(~_rstB_))
`define ip2211ringpll_FLOP_NORESET(_clk_,_in_,_out_) `ip2211ringpll_MSFF(_out_,_in_,_clk_)

`define ip2211ringpll_FLOP_ENABLED(_clk_,_rstB_,_en_,_in_,_out_) `ip2211ringpll_EN_RST_MSFF(_out_,_in_,_clk_,_en_,(~_rstB_))
`define ip2211ringpll_FLOP_SET(_clk_,_rstB_,_in_,_out_) `ip2211ringpll_SET_MSFF(_out_,_in_,_clk_,(~_rstB_))
`define ip2211ringpll_FLOP_ENABLED_SET(_clk_,_rstB_,_en_,_in_,_out_) `ip2211ringpll_EN_SET_MSFF(_out_,_in_,_clk_,_en_,(~_rstB_))
   
// `define MUX41(_sel_,_ina_,_inb_,_inc_,_ind_,_out_) assign _out_ = _sel_[1] ?  (_sel_[0] ? _ind_ : _inc_) : (_sel_[0] ? _inb_ : _ina_)
// `define MUX81(_sel_,_ina_,_inb_,_inc_,_ind_,_ine_,_inf_,_ing_,_inh_,_out_) assign _out_ = _sel_[2] ? (_sel_[1] ?  (_sel_[0] ? _inh_ : _ing_) : (_sel_[0] ? _inf_ : _ine_)) : (_sel_[1] ?  (_sel_[0] ? _ind_ : _inc_) : (_sel_[0] ? _inb_ : _ina_))   
// `define MUX161(_sel_,_ina_,_inb_,_inc_,_ind_,_ine_,_inf_,_ing_,_inh_,_ini_,_inj_,_ink_,_inl_,_inm_,_inn_,_ino_,_inp_,_out_) assign _out_ = _sel_[3] ? (_sel_[2] ? (_sel_[1] ?  (_sel_[0] ? _inp_ : _ino_) : (_sel_[0] ? _inn_ : _inm_)) : (_sel_[1] ?  (_sel_[0] ? _inl_ : _ink_) : (_sel_[0] ? _inj_ : _ini_))) : (_sel_[2] ? (_sel_[1] ?  (_sel_[0] ? _inh_ : _ing_) : (_sel_[0] ? _inf_ : _ine_)) : (_sel_[1] ?  (_sel_[0] ? _ind_ : _inc_) : (_sel_[0] ? _inb_ : _ina_)))  


  //                                84 2152 1
  //                                     15 2
  //                                     26 8
  //                                GG GGGG G
  //                                BB BBBB B  


 `define ip2211ringpll_DATA_2_TO_1_MUX(dataout, datin1, datain2, muxselect)                                    \
   `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                        \
   `endif                                                                                        \
   assign dataout = ((datin1&({$bits(dataout){muxselect}})) | (datain2&{$bits(dataout){~muxselect}})); \

  
`endif //  `ifndef ip2211ringpll_SOC_MACROS_VH



/*************************************************************************************************************************
*
*    MACROS NOT BEING USED BY ANYONE - COMMENTED OUT -  FOR ANY ISSUES
*
**************************************************************************************************************************/     

//
//
///* lintra s-30500 */
//
//`define NO_SYNTH_ASYNC_RST_MSFF_BLK(q,i,clock,rst)                   \
//   logic [$bits(i)-1:0] \``dlyin_``q ;                        \
//   assign  \``dlyin_``q = i;                                \
//   always_ff @(posedge clock or posedge rst)                \
//      begin                                                 \
//         if (rst)  q =  '0;                                  \
//         else      q =  \``dlyin_``q ;                        \
//      end                                                   \
//
//
//
//`define NO_SYNTH_ASYNC_RST_MSFF_P_BLK(q,i,clock,rst)                 \
//   logic [$bits(i)-1:0] \``dlyin_``q ;                        \
//   assign  \``dlyin_``q = i;                                \
//   always_ff @(negedge clock or posedge rst)                \
//      begin                                                 \
//         if (rst)  q =  '0;                                  \
//         else      q =  \``dlyin_``q ;                        \
//      end                                                   \
//
//
///* lintra s-30500 */
//
//`define NO_SYNTH_EN_ASYNC_RST_MSFF_BLK(q,i,clock,enable,rst)         \
//   logic [$bits(i)-1:0] \``dlyin_``q ;                        \
//   logic \``dlyen_``q ;                                       \
//   assign  \``dlyin_``q = i;                                \
//   assign  \``dlyen_``q = enable;                           \
//   always_ff @(posedge clock or posedge rst)                \
//      begin                                                 \
//         if (rst)     q =  '0;                               \
//         else if (\``dlyen_``q ) q =  \``dlyin_``q ;             \
//      end                                                   \
//
//
//`define ASYNC_RST_SET_B(q_b,rst,set)                          \
//   always_latch                                               \
//      begin                                                   \
//         if (set | rst)                                       \
//            if (rst) q_b =  '1; /* lintra s-30529, s-30531  */  \
//            else     q_b = '0;                                \
//      end                                                     \
//
//
//`define NO_SYNTH_TRI_DRIVE(Bus,En,Data) /* lintra s-30505 */              \
//  `ifdef INTC_EMULATION                                                          \
//        assign Bus = {$bits(Bus){1'b1}}; \
//  `else                                                                  \
//        assign Bus = En ? Data : {$bits(Bus){1'bz}}; \
//  `endif
//
//
//
//`define NO_SYNTH_WAND_TRI_DRIVE(Bus,En,Data) /* lintra s-30505 */          \
//  `ifdef INTC_EMULATION                                                          \
//        assign Bus = En ? Data : {$bits(Bus){1'b1}}; \
//  `else                                                                  \
//        assign Bus = En ? Data : {$bits(Bus){1'bz}}; \
//  `endif
//
//
//
//
//
//`define MCP_BNL     `BNL
//`define MCP_PUNIT   `PUNIT
//`define MCP_CCK     `CCK
//`define MCP_DUNIT   `DUNIT
//`define MCP_NORTHC  `NORTHC
//`define MCP_MUNIT   `MUNIT
//`define MCP_HUNIT   `HUNIT
//`define MCP_AUNIT   `AUNIT
//`define MCP_BUNIT   `BUNIT
//`define MCP_CUNIT   `CUNIT
//`define MCP_BLAUNCH_PATH  `BLAUNCH_PATH
//`define MCP_BRAM_PATH     `BRAM_PATH
//`define MCP_DISP_2D `DISP_2D
//`define MCP_GVD     `GVD
//`define MCP_GFX     `GFX
//`define MCP_VED     `VED
//`define MCP_VEC     `VEC
//`define MCP_FUS     `FUS
//`define MCP_DMIC    `DMIC
//
//
//
//
//`define MCP_LNCGFX(MCP_source_sig, MCP_rx_enable, MCP_count_clk, MCP_rx_clk, phase_delay, macro_inst_name, clock_edges_aligned_at_destination, sampling_edge_or_phase) \
//\
//`ifdef LNCGFX \
//`ip2211ringpll_MCP(MCP_source_sig, MCP_rx_enable, MCP_count_clk, MCP_rx_clk, phase_delay, macro_inst_name, clock_edges_aligned_at_destination, sampling_edge_or_phase) \
//`else \
//`MCP_LNCFC(MCP_source_sig, MCP_rx_enable, MCP_count_clk, MCP_rx_clk, phase_delay, macro_inst_name, clock_edges_aligned_at_destination, sampling_edge_or_phase) \
//`endif 
//
//
//`define MCP_LNCBFM(MCP_source_sig, MCP_rx_enable, MCP_count_clk, MCP_rx_clk, phase_delay, macro_inst_name, clock_edges_aligned_at_destination, sampling_edge_or_phase) \
//\
//`ifdef LNCBFM \
//`ip2211ringpll_MCP(MCP_source_sig, MCP_rx_enable, MCP_count_clk, MCP_rx_clk, phase_delay, macro_inst_name, clock_edges_aligned_at_destination, sampling_edge_or_phase) \
//`else \
//`MCP_LNCGFX(MCP_source_sig, MCP_rx_enable, MCP_count_clk, MCP_rx_clk, phase_delay, macro_inst_name, clock_edges_aligned_at_destination, sampling_edge_or_phase) \
//`endif
//
// `define MUX21(_sel_,_ina_,_inb_,_out_) assign _out_ = (_sel_ ? _inb_ : _ina_)
//
//`define FLOP_NORESET_NODELAY(_clk_,_in_,_out_) `ip2211ringpll_MSFF(_out_,_in_,_clk_)
//
//`define FLOP_NEGEDGE(_clk_,_rstB_,_in_,_out_) `ip2211ringpll_RST_MSFF_P(_out_,_in_,_clk_,(~_rstB_))
//`define FLOP_NEGEDGE_ENABLED(_clk_,_rstB_,_en_,_in_,_out_) `ip2211ringpll_EN_RST_MSFF_P(_out_,_in_,_clk_,_en_,(~_rstB_))
//
//`define FLOP_NEGEDGE_SET(_clk_,_rstB_,_in_,_out_) `SET_MSFF_P(_out_,_in_,_clk_,(~_rstB_))
//`define FLOP_NEGEDGE_ENABLED_SET(_clk_,_rstB_,_en_,_in_,_out_) `EN_SET_MSFF_P(_out_,_in_,_clk_,_en_,(~_rstB_))

/*************************************************************************************************************************
*
*    MACROS NOT BEING USED BY ANYONE - COMMENTED OUT -
*
**************************************************************************************************************************/     

//`define ASYNC_FLOP(_clk_,_rstB_,_in_,_out_) `ip2211ringpll_ASYNC_RST_MSFF(_out_,_in_,_clk_,(~_rstB_))
//`define ASYNC_FLOP_SET(_clk_,_rstB_,_in_,_out_) `ip2211ringpll_ASYNC_SET_MSFF(_out_,_in_,_clk_,(~_rstB_))               \
//
//`define ip2211ringpll_ASYNC_RST_MSFF_META(q,i,clk,rstb)                      \
//`ifdef INTC_DC                                                      \
//  `LIB_ASYNC_RST_MSFF_META(q,i,clk,rstb)                       \
//`else                                                          \
//                                                               \
//  always_ff @(posedge clk or negedge rstb) begin               \
//    if ( ~rstb )  q <= '0;                                     \
//    else          q <=  i;                                     \
//  end                                                          \
//`endif                                                         \
//
//// New BUFFER for 1ns of delay ***** ONLY FOR USE ON UNGATED SUPPLIES (VNN OR VNNAON)
//`define BUF_1NS_DELAY_UNGATED(out,in,vcc_in)                      \
//`ifdef INTC_DC                                                         \
//     `LIB_BUF_1NS_DELAY_UNGATED(out,in,vcc_in)                    \
//`else                                                             \
//  assign out = in ;     /* lintra s-35000, s-35006 */              \
//`endif         
//
//
//  //                              3333 3322 2222 2222 1111 1111
//  //                              5432 1098 7654 3210 9876 5432
// `define BUNIT_REAL_BANK_MASK 24'b0000_0001_0000_0000_0100_1111
// `define BUNIT_REAL_ROW_MASK  24'b0000_1111_1111_1111_1111_1110
// `define BUNIT_REAL_RANK_MASK 24'b0001_1110_0000_0000_0000_0000  
//
//

//  
// `define FUNCTIONL_ADDRESS    24'b0011_1110_0000_0000_0000_0000
//
///* lintra s-30500 */
//
////Same functionality as regular latch, but adding DE-SKEW to the name
////so that it is clear whenever this latch is instantiated it is intended to be 
////redundant to reduce mindelay problems between high-skew sequentials
//`define LATCH_DESKEW(q,i,clock)                             \
//   always_latch                                             \
//      begin                                                 \
//         if (clock) q <=  i;                                 \
//      end                                                   \
//
//
//`define ASYNC_RST_MSFFD(q,i,clock,rst)                       \
//wire \``q``_rst ;                                             \
//assign \``q``_rst = rst ;                                      \
//   always_ff @(posedge clock or posedge \``q``_rst )           \
//      begin                                                 \
//         if ( \``q``_rst )  q <=  '0;                      \
//         else      q <=  i;                                 \
//      end                                                   \
//
//`define ASYNC_RSTB_MSFF_HF_NONSCAN(q,i,clock,rstb)                      \
//  logic [$bits(q)-1:0] \``q``_nonscan ;                                 \
//  assign q = \``q``_nonscan ;                                           \
//`ifdef INTC_DC                                                               \
//   `LIB_ASYNC_RSTB_MSFF_HF_NONSCAN(q,i,clock,rstb)                      \
//`else                                                                   \
//   wire \``q``_rstb ;                                                   \
//   assign \``q``_rstb = rstb ;                                          \
//   always_ff @(posedge clock or negedge \``q``_rstb )                   \
//      begin                                                             \
//         if (~(\``q``_rstb ))  \``q``_nonscan <= '0;                    \
//         else      \``q``_nonscan <=  i;                                \
//      end                                                               \
//`endif
//
////============================================================================================
////
////  6 Bit Comparator
////
////============================================================================================
//`define COMPARATOR_6_BIT(out, in1, in2)                       \
//compare_6_bit \``compare_6_bit_``out (                        \
//                                  .iout(out),                 \
//                                  .iin1(in1),                 \
//                                  .iin2(in2)                  \
//                                 ); 
//
//module compare_6_bit(iout, iin1, iin2);
//output logic iout;
//input logic [5:0] iin1;
//input logic [5:0] iin2;
//`ifdef INTC_DC
//   `LIB_compare_6_bit(iout, iin1, iin2)
//`else 
//   assign iout = (iin1 == iin2);
//`endif        
//endmodule
//    
//`define LATCH_NEGEDGE(_le_,_in_,_out_) `LATCH_PD(_out_,_in_,_le_)
//
//`define LATCH_P_HF_NONSCAN(q,i,clock)                       \
//  logic [$bits(q)-1:0] \``q``_nonscan ;                     \
//  assign q = \``q``_nonscan ;                               \
//`ifdef INTC_DC                                                   \
//   `LIB_LATCH_P_HF_NONSCAN(q,i,clock)                       \
//`else                                                       \
//   always_latch                                             \
//      begin                                                 \
//         if (~clock) \``q``_nonscan <= i;                   \
//      end                                                   \
//`endif
//
///* lintra s-50500 */
//
//
//`define LATCH_PD(q,i,clock)                                  \
//   always_latch                                             \
//      begin                                                 \
//         if (~clock) q <= i;                                \
//      end                                                   \
//
///* lintra s-50500 */
//
////Creating a MSFF_NONSCAN to allow users to instantiate a flop which won't be added to the scan chain
////Note that in INTC_DC mode the library module creates an instance name integration can key off
////of as well as appending _nonscan to the output signal name. Both of which should ensure the
////cell is kept and not swapped out for a scan version.
//`define MSFF_NONSCAN(q,i,clock)                              \
//  logic [$bits(q)-1:0] \``q``_nonscan ;                      \
//  assign q = \``q``_nonscan ;                                \
//                                                             \
//  `ifdef INTC_DC                                                  \
//    `LIB_MSFF_NONSCAN(q,i,clock)                \
//  `else                                                      \
//    always_ff @(posedge clock)                               \
//      begin                                                  \
//         \``q``_nonscan <= i;                                \
//      end                                                    \
//  `endif
//
//// Data Mux for timing critical signals
//
//`define MUX_2TO1_HF(out,in1,in2,sel)                       \
//`ifdef INTC_DC                                                  \
//   `LIB_MUX_2TO1_HF(out,in1,in2,sel)                       \
//`else                                                      \
//   assign out = (in1 & sel) | (in2 & ~sel);                \
//`endif  
//
//`define MUX_2TO1_INV_HF(out,in1,in2,sel)                       \
//`ifdef INTC_DC                                                  \
//   `LIB_MUX_2TO1_INV_HF(out,in1,in2,sel)                       \
//`else                                                      \
//   assign out = ~((in1 & sel) | (in2 & ~sel));                \
//`endif        
//
//
//// Data Mux using NAND-NAND gates for timing critical signals
//`define NAND_3TO1MUX(iout,iin1,iin2,iin3,isel1,isel2,isel3)    \
//nand_3to1_mux \``nand_mux_``iout (                             \
//                                  .out(iout),                  \
//                                  .in1(iin1),                  \
//                                  .in2(iin2),                  \
//                                  .in3(iin3),                  \
//                                  .sel1(isel1),                \
//                                  .sel2(isel2),                \
//                                  .sel3(isel3)                 \
//                                 ); 
//
//module nand_3to1_mux(out,in1,in2,in3,sel1,sel2,sel3);
//output logic out;
//input logic in1;
//input logic in2;
//input logic in3;
//input logic sel1;
//input logic sel2;
//input logic sel3;
//`ifdef INTC_DC
//   `LIB_NAND_3TO1MUX(out,in1,in2,in3,sel1,sel2,sel3) 
//`else 
//  always_comb begin
//    casex({ sel1, 
//            sel2,
//            sel3 })
//      3'b100  : out = in1;
//      3'b010  : out = in2;
//      3'b001  : out = in3;
//      default : out = 1'b0;
//    endcase
//  end
//`endif        
//endmodule
//
//  `define OUTREG logic
//
//`define MCP_LNCFC(MCP_source_sig, MCP_rx_enable, MCP_count_clk, MCP_rx_clk, phase_delay, macro_inst_name, clock_edges_aligned_at_destination, sampling_edge_or_phase) \
//\
//`ifdef LNCFC \
//`ip2211ringpll_MCP(MCP_source_sig, MCP_rx_enable, MCP_count_clk, MCP_rx_clk, phase_delay, macro_inst_name, clock_edges_aligned_at_destination, sampling_edge_or_phase) \
//`endif

`ifndef ip2211ringpll_SOC_CLOCK_MACROS_VH
`define ip2211ringpll_SOC_CLOCK_MACROS_VH

////`include "vlv_macro_tech_map.vh"
//`include "soc_macros.sv"

//`define ip2211ringpll_MAKE_CLK_DIV2_RESET(ckdiv2rout,ckdiv2rin,ckdiv2clkin,ckdiv2resetin)       \
`define ip2211ringpll_CLK_FF(ckdiv2rout,ckdiv2rin,ckdiv2clkin,ckdiv2resetin)                      \
ip2211ringpll_clockdivffreset \``clockdivffreset_``ckdiv2rout (                                   \
                                               .ffoutreset(ckdiv2rout),             \
                                               .ffinreset(ckdiv2rin),               \
                                               .clockinreset(ckdiv2clkin),          \
                                               .resetckdivff(ckdiv2resetin)         \
                                              );



`define ip2211ringpll_CLK_FF_RESETB(ckdiv2rout,ckdiv2rin,ckdiv2clkin,ckdiv2resetinb)                      \
ip2211ringpll_clockdivffresetb \``clockdivffresetb_``ckdiv2rout (                                   \
                                               .ffoutreset(ckdiv2rout),             \
                                               .ffinreset(ckdiv2rin),               \
                                               .clockinreset(ckdiv2clkin),          \
                                               .resetckdivffb(ckdiv2resetinb)         \
                                              );





`define ip2211ringpll_MAKE_CLK_DIV2_RESET(ckdiv2rout,ckdiv2rin,ckdiv2clkin,ckdiv2resetin)                      \
ip2211ringpll_clockdivffreset \``clockdivffreset_``ckdiv2rout (                                   \
                                               .ffoutreset(ckdiv2rout),             \
                                               .ffinreset(ckdiv2rin),               \
                                               .clockinreset(ckdiv2clkin),          \
                                               .resetckdivff(ckdiv2resetin)         \
                                              );


                                              
//module ip2211ringpll_clockdivffreset (ffoutreset, ffinreset, clockinreset,resetckdivff);    
//output ffoutreset;
//input ffinreset;
//input clockinreset;
//input resetckdivff;
//reg ffoutreset;
//wire ffinreset, clockinreset, resetckdivff;   
//reg  ffin_inv;
//wire set; 
//`ifdef INTC_DC 
//     `LIB_clockdivffreset(ffoutreset, ffinreset, clockinreset,resetckdivff) --- fixed INTC_FEV issue
//     `LIB_clockdivffreset(ffoutreset, ~ffinreset, clockinreset,resetckdivff) 
//`else 
//always @(posedge (set) or posedge clockinreset)
//begin
//  if (set)
//    ffin_inv = 1'b1; /* lintra s-60028 */
//  else
//    ffin_inv = (~ffinreset); /* lintra s-60028 */
//end
//assign set = ~resetckdivff;
//assign ffoutreset = ~ffin_inv;
//`endif
//endmodule

// This was the previous behavioural model - changed on request
module ip2211ringpll_clockdivffreset (ffoutreset, ffinreset, clockinreset,resetckdivff);    
output ffoutreset;
input ffinreset;
input clockinreset;
input resetckdivff;
reg ffoutreset;
wire ffinreset, ffinresetb, clockinreset, resetckdivff;   
wire ffin_inv;
//`ifdef INTC_DC 
       //     assign ffinresetb = ~ffinreset;
       //     `LIB_clockdivffreset(ffoutreset, ffinresetb, clockinreset,resetckdivff)
      //	 d04cdc03wd0d0 ckdiv2ff1 (.clkout(ffoutreset), .d(ffinresetb), .clk(clockinreset), .rb(resetckdivff));
//     ctech_lib_clk_inv ctech_lib_clk_inv(.clk(ffinreset),.clkout(ffinresetb));
//     ctech_lib_clk_div2_reset ctech_lib_clk_div2_reset(.clkout(ffoutreset),.in(ffinresetb),.clk(clockinreset),.rst(!resetckdivff));
//`else 
always @(negedge (resetckdivff) or posedge clockinreset)
begin
  if (~(resetckdivff))
    ffoutreset = 1'b0; /* lintra s-60028 */
  else
    ffoutreset = (ffinreset); /* lintra s-60028 */
end
//`endif
endmodule

module ip2211ringpll_clockdivffresetb (ffoutreset, ffinreset, clockinreset,resetckdivffb);
output ffoutreset;
input ffinreset;
input clockinreset;
input resetckdivffb;
reg ffoutreset;
wire ffinreset, ffinresetb, clockinreset, resetckdivffb, resetckdivff;
wire ffin_inv;
//`ifdef INTC_DC
     //     assign ffinresetb = ~ffinreset;
     //     assign resetckdivff = ~resetckdivffb;
     //     `LIB_clockdivffreset(ffoutreset, ffinresetb, clockinreset,resetckdivff)
     //	d04cdc03wd0d0 ckdiv2ff1 (.clkout(ffoutreset), .d(ffinresetb), .clk(clockinreset), .rb(resetckdivff));
//    ctech_lib_clk_inv ctech_lib_clk_inv(.clk(ffinreset),.clkout(ffinresetb));
//    ctech_lib_clk_div2_reset ctech_lib_clk_div2_reset(.clkout(ffoutreset),.in(ffinresetb),.clk(clockinreset),.rst(resetckdivffb));
//`else 
always @(posedge (resetckdivffb) or posedge clockinreset)
begin
  if (resetckdivffb)
    ffoutreset = 1'b0; /* lintra s-60028 */
  else
    ffoutreset = (ffinreset); /* lintra s-60028 */
end
//`endif
endmodule


module ip2211ringpll_CLK_NAND_3TO1_MUX(out,in1,in2,in3,sel1,sel2,sel3);
output logic out;
input logic in1;
input logic in2;
input logic in3;
input logic sel1;
input logic sel2;
input logic sel3;
//`ifdef INTC_DC
             //   `LIB_CLK_NAND_3TO1MUX(out,in1,in2,in3,sel1,sel2,sel3)
//   wire sel3b;                                                                     
//   wire sel2b;                                                                     
//   wire sel1b;                                                                     
//   wire nor1;                                                                      
//   wire nor2;                                                                      
//   wire nor3;                                                                      
//   wire x1;                                                                        
//   wire x2;                                                                        
//   wire x3;                                                                        
//   wire x4;                                                                        
//   wire x4x;                                                                       
          //    d04inn00wd0f7 i1_out (.o1(sel3b),.a(sel3));                            
          //    d04inn00wd0f7 i2_out (.o1(sel2b),.a(sel2));                            
          //    d04inn00wd0f7 i3_out (.o1(sel1b),.a(sel1));                            
          //    d04non03wd0d7 i4_out (.o1(nor1),.a(sel3b),.b(sel2),.c(sel1));          
          //    d04non03wd0d7 i5_out (.o1(nor2),.a(sel3),.b(sel2b),.c(sel1));          
          //    d04non03wd0d7 i6_out (.o1(nor3),.a(sel3),.b(sel2),.c(sel1b));          
          //    d04gna00wd0d0 i7_out (.clk(in3),.en(nor1),.clkout(x1));                      
          //    d04gna00wd0d0 i8_out (.clk(in2),.en(nor2),.clkout(x2));                      
          //    d04gna00wd0d0 i9_out (.clk(in1),.en(nor3),.clkout(x3));                      
          //    d04gna02wd0e0 i10_out (.clkout(x4x),.clk1(x1),.clk2(x2));                     
          //    d04inn00wd0f7 i11_out (.o1(x4),.a(x4x));                               
          //    d04gna02wd0e0 i12_out (.clkout(out),.clk1(x4),.clk2(x3));     
//   assign sel3b = ~sel3;
//   assign sel2b = ~sel2;
//   assign sel1b = ~sel1;
//   assign nor1 = ~(sel3b|sel2|sel1);
//   assign nor2 = ~(sel3|sel2b|sel1); 
//   assign nor3 = ~(sel3|sel2|sel1b);                         
//   ctech_lib_clk_nand_en ctech_lib_clk_nand_en_1(.clk(in3),.en(nor1),.clkout(x1));
//   ctech_lib_clk_nand_en ctech_lib_clk_nand_en_2(.clk(in2),.en(nor2),.clkout(x2));
//   ctech_lib_clk_nand_en ctech_lib_clk_nand_en_3(.clk(in1),.en(nor3),.clkout(x3));           
//   ctech_lib_clk_nand ctech_lib_clk_nand_1(.clkout(x4x),.clk1(x1),.clk2(x2));                      
//   ctech_lib_clk_inv ctech_lib_clk_inv (.clk(x4x),.clkout(x4));
//   ctech_lib_clk_nand ctech_lib_clk_nand_2(.clkout(out),.clk1(x4),.clk2(x3)); 
//`else 
  always_comb begin
    casex({ sel1, 
            sel2,
            sel3 })
      3'b100  : out = in1;
      3'b010  : out = in2;
      3'b001  : out = in3;
      default : out = 1'b0;
    endcase
  end
//`endif        
endmodule

// gclatchen clock gate macro with disable
`define ip2211ringpll_MAKE_CLK_GCLATCHEN(gcenclkout,gcenin,gctein,gcclrbin,gcckin)    \
ip2211ringpll_clklocgclatchen \``clklocgclatchen_``gcenclkout  (                                   \
                                               .gcenclkoutx(gcenclkout),               \
                                               .gceninx(gcenin),                       \
                                               .gcteinx(gctein),                       \
                                               .gcclrbinx(gcclrbin),                   \
                                               .gcckinx(gcckin)                        \
                                             );

module ip2211ringpll_clklocgclatchen (gcenclkoutx, gceninx, gcteinx, gcclrbinx, gcckinx);
input gceninx;
input gcteinx;
input gcclrbinx;
input gcckinx;
output gcenclkoutx;

//`ifdef INTC_DC
         //   LIB_GCLATCHEN(gcenclkoutx,gceninx,gcteinx,gcclrbinx,gcckinx) 
         //     d04cgc02wd0d0 \ckgclatchen_dcszo (.clkout(gcenclkoutx),.clk(gcckinx),.en(gceninx),.te(gcteinx));  
//   ctech_lib_clk_gate_te_rst_ss ctech_lib_clk_gate_te_rst_ss(.clkout(gcenclkoutx),.clk(gcckinx),.en(gceninx),.te(gcteinx),.rst(!gcclrbinx),.ss(1'b0));                
//`else                                                                        
reg lq;                                                                      
                                                                             
always_latch                                                                 
begin : gclatchen0_internal_latches                                          
                                                                             
  if (( ~gcckinx) == 1'b1) lq <= gceninx;                                      
                                                                             
end // begin: gclatchen0_internal_latches                                    
                                                                             
assign gcenclkoutx = gcclrbinx & gcckinx & (gcteinx | lq);                       
//`endif                                                                       
endmodule


//Including clk_gate_te macro
`define ip2211ringpll_MAKE_CLK_GEN(gcenclkout,gcenin,gctein,gcckin)    \
ip2211ringpll_clkgateen \``ip2211ringpll_clkgateen``gcenclkout  (                                   \
                                               .gcenclkoutx(gcenclkout),               \
                                               .gceninx(gcenin),                       \
                                               .gcteinx(gctein),                       \
                                               .gcckinx(gcckin)                        \
                                             );

module ip2211ringpll_clkgateen (gcenclkoutx, gceninx, gcteinx, gcckinx);
input logic gceninx;
input logic gcteinx;
input logic gcckinx;
output logic gcenclkoutx;

`ifdef INTC_DC
   ctech_lib_clk_gate_te ctech_lib_clk_gate_te(.clkout(gcenclkoutx),.clk(gcckinx),.en(gceninx),.te(gcteinx));
`else
reg lq;

always_latch
begin : gclatchen0_internal_latches

  if (( ~gcckinx) == 1'b1) lq <= gceninx | gcteinx ;

end // begin: gclatchen0_internal_latches

assign gcenclkoutx = gcckinx & lq;
`endif
endmodule



`define ip2211ringpll_MAKE_CLK_INV(ckinvout,ckinvin)             \
ip2211ringpll_clkinv \``clkinv_``ckinvout (                        \
                           .clkout (ckinvout),     \
                           .clkin (ckinvin)        \
                          );

// clock inverter module
module ip2211ringpll_clkinv (clkout,clkin);
output clkout;
input clkin;
wire clkout,clkin;
//`ifdef INTC_DC
          //     `LIB_clkinv(clkout,clkin)
//	ctech_lib_clk_inv ctech_lib_clk_inv(.clkout(clkout),.clk(clkin));
//`else
assign clkout = ~clkin ;
//`endif
endmodule

//equal rise and flal time for two input clks


`define ip2211ringpll_MAKE_CLKNOR(clkout,clkin1,clkin2)                    \
ip2211ringpll_clknor \``clknor_``clkout  (                                     \
                          .ckoout (clkout),                     \
                          .ckoin1 (clkin1),                     \
                          .ckoin2 (clkin2)                      \
                         );

module ip2211ringpll_clknor (ckoout, ckoin1,ckoin2);
output ckoout;
input ckoin1;
input ckoin2;
wire ckoout,ckoin1,ckoin2;

//`ifdef INTC_DC
         //     `LIB_clknor(ckoout, ckoin1,ckoin2)
//      ctech_lib_clk_nor ctech_lib_clk_nor(.clkout(ckoout),.clk1(ckoin1),.clk2(ckoin2));
//`else
assign ckoout = (~(ckoin1|ckoin2));
//`endif
endmodule




`define ip2211ringpll_MAKE_CLK_DIV4_RESET(ckdiv4rout,ckdiv4rin,ckdiv4resetin)                 \
ip2211ringpll_clockdiv4ffreset \``clockdiv4ffreset_``ckdiv4rout (                             \
                                               .clk_out(ckdiv4rout),         	\
                                               .clk_in(ckdiv4rin),              \
                                               .reset_in(ckdiv4resetin)         \
                                              );




`define ip2211ringpll_CLK_GATE(o, clk, a)                                                                 \
 ip2211ringpll_soc_rbe_clk \``soc_rbe_clk_``o (                                                           \
                                  .ckrcbxpn  (o),                                           \
                                  .ckgridxpn (clk),                                         \
                                  .latrcben  (a)                                            \
                                );

`define ip2211ringpll_CLK_GATE_W_OVERRIDE(o, clk, pwrgate, override)                                      \
 clk_gate_kin \``clk_gate_kin_``o (                                                         \
                                  .ckrcbxpn1  (o),                                          \
                                  .ckgridxpn1 (clk),                                        \
                                  .latrcben1  (pwrgate),                                    \
                                  .testen1    (override)                                    \
                                );

//`LIB_SOC_CLKAND(outclk,inclk,enable) 
`define ip2211ringpll_CLKAND(outclk,inclk,enable)                                                         \
//`ifdef INTC_DC                                                                                   \
//    ctech_lib_clk_and_en \ctech_lib_clk_and_en_``outclk``_a (.clkout(outclk),.clk(inclk),.en(enable));\
//`else                                                                                       \
   `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                   \
                                                                                            \
   `endif                                                                                   \
   assign outclk = inclk & enable; /* lintra s-30004, s-31500 */                            \
//`endif 

module ip2211ringpll_clk_and(input logic a,b, output logic o);
//`ifdef INTC_DC
       //  `LIB_SOC_CLKAND(o,a,b)
//ctech_lib_clk_and ctech_lib_clk_and (.clk1(a), .clk2(b), .clkout(o));
//`else
  assign o = a & b;
//`endif
endmodule

//// Macro for MODQ simulation queue for clock tree in bus cluster
//`define CLKANDMODQ(outclk, inclk1, inclk0)                                                  \
//   soc_clkandmodq \``clkandmodq_``outclk ( /* lintra s-32002 */                             \
//      .outclkm (outclk),                                                                    \
//      .inclk1m (inclk1),                                                                    \
//      .inclk0m (inclk0)                                                                     \
//   );
//
//
//
//module soc_clkandmodq (outclkm,
//                   inclk1m,
//                   inclk0m);
//
//output outclkm;
//input inclk1m;
//input inclk0m;
//
//wire outclkm, inclk1m, inclk0m;
//
//assign outclkm = inclk1m & inclk0m;
//
//
//endmodule // soc_clkandmodq

// Clock buffer for "clocks in the datapath".  Usage of this macro requires a waiver.
`define ip2211ringpll_CLKAND_DP(outclk,inclk, enable)                                                     \
`ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                      \
                                                                                            \
`endif                                                                                      \
   always_comb outclk <= inclk & enable; /* lintra s-30003, s-31500, s-31503 */             \

//wire outclk``_tmp;  mnigri, removed from inside the macro, cause problem when outclk is of the form blabla[4] then adding _tmp is problematic, fails in INTC_DC
// its a MF macro technology !!!!  


// New clock buffer macro

//     `LIB_CLKBF_SOC(clkbufout,clkbufin)
`define ip2211ringpll_CLKBF(clkbufout,clkbufin)                                                           \
//`ifdef INTC_DC                                                                                   \
//     ctech_lib_clk_buf \ctech_lib_clk_buf_``clkbufout``c (.clkout(clkbufout),.clk(clkbufin));  \
// `else                                                                                      \
  `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                    \
                                                                                            \
   `endif                                                                                   \
     assign clkbufout =  (~(~(clkbufin)));                                                  \
// `endif

`define ip2211ringpll_CLKINV(clkinvout,clkinvin)                                                          \
//`ifdef INTC_DC                                                                                   \
//	ctech_lib_clk_inv iclk_lib_clk_inv_``clkinvout``(.clkout(clkinvout), .clk(clkinvin));  \
// `else                                                                                      \
  `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                    \
                                                                                            \
   `endif                                                                                   \
     assign clkinvout =  (~(clkinvin));                                                     \
// `endif

//     `LIB_clknan(o,ck1,ck2)
`define ip2211ringpll_CLK_NAND(o,ck1,ck2)                                                                 \
//`ifdef INTC_DC                                                                                   \
//     ctech_lib_clk_nand ctech_lib_clk_nand_``o``(.clkout(o),.clk1(ck1),.clk2(ck2));               \
//`else                                                                                       \
  assign o = ~(ck1 & ck2);                                                                  \
//`endif                                                                                      \


`define ip2211ringpll_CLK_NAND_EN(o,ck,en)                                                                \
//`ifdef INTC_DC                                                                                   \
//     `LIB_clknanen(o,ck,en)                                                                 \
//`else                                                                                       \
  assign o = ~(ck & en);                                                                    \
//`endif                                                                                      \

//`LIB_clknor(o,ck1,ck2)
`define ip2211ringpll_CLK_NOR(o,ck1,ck2)                                                                  \
//`ifdef INTC_DC                                                                                   \
//     ctech_lib_clk_nor ctech_lib_clk_nor_``o``(.clkout(o),.clk1(ck1),.clk2(ck2));           \
//`else                                                                                       \
  assign o = ~(ck1 | ck2);                                                                  \
//`endif                                                                                      \

`define ip2211ringpll_CLK_AND_EN(o,ck,en)                                                                 \
//`ifdef INTC_DC                                                                                   \
//    ctech_lib_clk_and_en ctech_lib_clk_and_en_``o``(.clkout(o),.clk(ck),.en(en));\
//`else                                                                                       \
  assign o = (ck & en);                                                                     \
//`endif                                                                                      \

//needed for BSCAN that requires to map a ctech macro  AND gate for non-clock signals, they are currently using a clk AND that is giving us timing problems because they are data signals

`define ip2211ringpll_DATAAND(outd,ind1,ind2)                                                             \
//`ifdef INTC_DC                                                                                   \
//      ctech_lib_and2 ctech_lib_and2_``outd``(.o(outd),.a(ind1),.b(ind2));                   \
//`else                                                                                       \
   `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                   \
   `endif                                                                                   \
   assign outd = ind1 & ind2; /* lintra s-30004, s-31500 */                                 \
//`endif


 `define ip2211ringpll_MAKE_CLK_2TO1MUX(clkmuxout,clkmuxin1,clkmuxin2,clkmuxselect)                       \
 ip2211ringpll_clk2to1mux \``clk2to1mux_``clkmuxout (                                                     \
                                     .ckmuxout (clkmuxout),                                 \
                                     .ckin1    (clkmuxin1),                                 \
                                     .ckin2    (clkmuxin2),                                 \
                                     .muxselect(clkmuxselect)                               \
                                    );

 
module ip2211ringpll_clk2to1mux (ckmuxout,ckin1,ckin2,muxselect);
output ckmuxout;
input ckin1;
input ckin2;
input muxselect;
wire ckmuxout,ckin1,ckin2,muxselect;
//`ifdef INTC_DC  
        //     `LIB_clk2to1mux(ckmuxout,ckin2,ckin1,muxselect)
//      ctech_lib_clk_mux_2to1 ctech_lib_clk_mux_2to1 (.clk1(ckin2), .clk2(ckin1), .s(muxselect), .clkout(ckmuxout));
//`else    
 assign ckmuxout = ((ckin1&~(muxselect)) | (ckin2&muxselect));
//`endif
endmodule

 `define ip2211ringpll_MAKE_DATA_2TO1MUX(clkmuxout,clkmuxin1,clkmuxin2,clkmuxselect)                 \
 ip2211ringpll_data2to1mux \``data2to1mux_``clkmuxout (                                              \
                                     .out (clkmuxout),                                 \
                                     .in1 (clkmuxin1),                                 \
                                     .in2 (clkmuxin2),                                 \
                                     .sel (clkmuxselect)                               \
                                    );

module ip2211ringpll_data2to1mux (out,in1,in2,sel);
output out;
input in1;
input in2;
input sel;
wire out,in1,in2,sel;
//`ifdef INTC_DC
       //     `LIB_MUX_2TO1_HF(out,in1,in2,sel)
//     ctech_lib_mux_2to1_hf ctech_lib_mux_2to1_hf(.out(out),.in1(in1),.in2(in2),.sel(sel));
//`else
  assign out = ((in1 & sel) | (in2 & ~sel));
//`endif
endmodule


/* -----\/----- EXCLUDED -----\/-----
`define MAKE_CLK_DELAY16(clkd16out,clkd16clkin,clkd16in0,clkd16in1,clkd16in2,clkd16in3,clkd16in4,clkd16in5,clkd16in6,clkd16in7,clkd16in8,clkd16in9,clkd16in10,clkd16in11,clkd16in12,clkd16in13,clkd16in14)                                   \
clk16delay \``clk16delay_``clkd16out (                                                      \
                                    .clk16delayout (clkd16out),                             \
                                    .clk16delayin (clkd16clkin),                            \
                                    .clk16in0 (clkd16in0),                                  \
                                    .clk16in1 (clkd16in1),                                  \
                                    .clk16in2 (clkd16in2),                                  \
                                    .clk16in3 (clkd16in3),                                  \
                                    .clk16in4 (clkd16in4),                                  \
                                    .clk16in5 (clkd16in5),                                  \
                                    .clk16in6 (clkd16in6),                                  \
                                    .clk16in7 (clkd16in7),                                  \
                                    .clk16in8 (clkd16in8),                                  \
                                    .clk16in9 (clkd16in9),                                  \
                                    .clk16in10 (clkd16in10),                                \
                                    .clk16in11 (clkd16in11),                                \
                                    .clk16in12 (clkd16in12),                                \
                                    .clk16in13 (clkd16in13),                                \
                                    .clk16in14 (clkd16in14)                                 \
                                  );

// Adjustable delay elements macros
module clk16delay (clk16delayout,clk16delayin,clk16in0,clk16in1,clk16in2,clk16in3,clk16in4,clk16in5,clk16in6,clk16in7,clk16in8,clk16in9,clk16in10,clk16in11,clk16in12,clk16in13,clk16in14);
output clk16delayout;
input clk16delayin;
input clk16in0;
input clk16in1;
input clk16in2;
input clk16in3;
input clk16in4;
input clk16in5;
input clk16in6;
input clk16in7;
input clk16in8;
input clk16in9;
input clk16in10;
input clk16in11;
input clk16in12;
input clk16in13;
input clk16in14;
wire clk16delayout,clk16delayin,clk16in0,clk16in1,clk16in2,clk16in3,clk16in4,clk16in5,clk16in6,clk16in7,clk16in8,clk16in9,clk16in10,clk16in11,clk16in12,clk16in13,clk16in14;
//`ifdef INTC_DC
             //     `LIB_clk16delay(clk16delayout,clk16delayin,clk16in0,clk16in1,clk16in2,clk16in3,clk16in4,clk16in5,clk16in6,clk16in7,clk16in8,clk16in9,clk16in10,clk16in11,clk16in12,clk16in13,clk16in14) 
//     ctech_lib_clk_16delay ctech_lib_clk_16delay(.clk16delayout(clk16delayout),.clk16delayin(clk16delayin),.clk16in0(clk16in0),.clk16in1(clk16in1),.clk16in2(clk16in2),.clk16in3(clk16in3),.clk16in4(clk16in4),.clk16in5(clk16in5),.clk16in6(clk16in6),.clk16in7(clk16in7),.clk16in8(clk16in8),.clk16in9(clk16in9),.clk16in10(clk16in10),.clk16in11(clk16in11),.clk16in12(clk16in12),.clk16in13(clk16in13),.clk16in14(clk16in14)); 
// `else
assign  clk16delayout = clk16delayin;
//`endif
endmodule                                  
 -----/\----- EXCLUDED -----/\----- */

/* -----\/----- EXCLUDED -----\/-----
//`define MAKE_CLK_
// clkdiv2 \``clk_div2_``cknameout (                                   \
//                                .div2cknameout (cknameout),          \
//                                .div2ipinckin (ipinckin),            \
//                                .div2usync (usync)                   \
//                               );

// creating FF module to be used by clock macros below
module clockdivff (ffout, ffin, clockin);    
output ffout;
input ffin;
input clockin;
reg ffout;
wire ffin, clockin;
//`ifdef INTC_DC 
        //     assign ffin_b = ~ffin;
        //     `LIB_clockdivff(ffout, ffin_b, clockin)
//       ctech_lib_clk_div2 ctech_lib_clk_div2(.clkout(ffout),.in(~ffin),.clk(clockin));
//`else                                                                         
 always @(posedge clockin)                                                
      begin                                                                  
         ffout = ffin; /-* lintra s-60028 *-/
      end  
//`endif
endmodule



module clkdiv2 (div2cknameout,div2ipinckin,div2usync);
output div2cknameout;
input div2ipinckin;
input div2usync;
reg div2cknameout;
wire div2ipinckin,div2usync;
 reg cknameout_ffout ;                                             
 wire cknameout_ffinvout ;                                         
 wire cknameout_andout ;                                           
always_latch                                                         
      begin                                                          
         if (~div2ipinckin) cknameout_ffout  = div2usync; /-* lintra s-60028 *-/
      end                                                            
assign cknameout_ffinvout  = (~(cknameout_ffout));              
//assign  cknameout_andout = (cknameout_ffinvout  & ~div2cknameout); 
assign  cknameout_andout = (cknameout_ffinvout  & div2cknameout);  // bug fix - the FF cell already make the invertion
clockdivff clockdivff_cknameout (                                 
                                  .ffout(div2cknameout),                 
                                  .ffin(cknameout_andout),         
                                  .clockin(div2ipinckin)                 
                                 );
endmodule
 -----/\----- EXCLUDED -----/\----- */
                               

`define ip2211ringpll_MAKE_CLK_OREN(ckorenout,ckorenckin,ckorenenin)              \
ip2211ringpll_clkoren \``clkoren_``ckorenout (                                    \
                              .clkorenout (ckorenout),              \
                              .clkorenckin (ckorenckin),            \
                              .clkorenenin (ckorenenin)             \
                             );

module ip2211ringpll_clkoren(clkorenout,clkorenckin,clkorenenin);
output clkorenout;
input clkorenckin;
input clkorenenin;
wire clkorenout,clkorenckin,clkorenenin;
wire clkorent1;
//`ifdef INTC_DC
        //     `LIB_clkoren(clkorenout,clkorenckin,clkorenenin)
//	ctech_lib_clk_or_en ctech_lib_clk_or_en(.clkout(clkorenout),.clk(clkorenckin),.en(clkorenenin));
 
//`else
assign clkorent1 = ~(clkorenckin|clkorenenin);
assign clkorenout = ~clkorent1;
//`endif
endmodule


`define ip2211ringpll_MAKE_CLKOR(clkorout,clkorin1,clkorin2)                    \
ip2211ringpll_clkor \``clkor_``clkorout  (                                      \
                          .ckoout (clkorout),                     \
                          .ckoin1 (clkorin1),                     \
                          .ckoin2 (clkorin2)                      \
                         );
module ip2211ringpll_clkor (ckoout, ckoin1,ckoin2);
output ckoout;
input ckoin1;
input ckoin2;
wire ckoout,ckoin1,ckoin2;
//`ifdef INTC_DC
       //     `LIB_clkor(ckoout, ckoin1,ckoin2)
// 	ctech_lib_clk_or ctech_lib_clk_or(.clkout(ckoout),.clk1(ckoin1),.clk2(ckoin2));
//`else   
assign ckoout = (~(~(ckoin1|ckoin2)));
//`endif
endmodule

// RBE clock ANDing logic.
//
module ip2211ringpll_soc_rbe_clk (output logic ckrcbxpn, input logic ckgridxpn, latrcben);  //lintra s-31506
logic latrcbenl; // rce state element
//`ifdef INTC_DC
         //     `LIB_soc_rbe_clk(ckrcbxpn,ckgridxpn,latrcben)
//	ctech_lib_latch_p ctech_lib_latch_p(.o(latrcbenl),.d(latrcben),.clkb(ckgridxpn));
//	ctech_lib_clk_and_en ctech_lib_clk_and_en(.clkout(ckrcbxpn),.clk(ckgridxpn),.en(latrcbenl));
	 
//`else
`ifndef INTC_VLV_FPGA_CLK_GATE
//   logic latrcbenl; // rce state element
  
  `ip2211ringpll_LATCH_P(latrcbenl, latrcben, ckgridxpn)
  `ip2211ringpll_CLKAND(ckrcbxpn, ckgridxpn, latrcbenl)
`else
assign ckrcbxpn = ckgridxpn;
`endif
//`endif
endmodule // ip2211ringpll_soc_rbe_clk                         

// RBE clock macro instantiating ip2211ringpll_soc_rbe_clk module above

`define ip2211ringpll_MAKE_SOC_RBE_CLK(ckrcbxpnout,ckgridxpnin,latrcbenin)                               \
 `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                    \
                                                                                           \
  `endif                                                                                   \
  ip2211ringpll_soc_rbe_clk \``soc_rbe_clk_``ckrcbxpnout (                                               \
                                          .ckrcbxpn (ckrcbxpnout),                         \
                                          .ckgridxpn (ckgridxpnin),                        \
                                          .latrcben (latrcbenin)                           \
                                         );

/* -----\/----- EXCLUDED -----\/-----
module qual_gen (
    input      clka,
    input      clkb,
    input      clka_usync,
    input      clkb_usync,
    input [5:0] clka_ratio,
    input [5:0] clkb_ratio,
    input       test_override,
    output reg  clka_qual,
    output reg  clkb_qual,
    output wire freq_match
                 
                  );

   reg[6:0]   clka_error;
   reg[6:0]   clkb_error;
   wire[6:0]  clka_ratio_adjusted;
   wire[6:0]  clkb_ratio_adjusted;
   wire[6:0]  clka_error_tmp;
   wire[6:0]  clkb_error_tmp;
   wire[6:0]  clka_ratio_adjusted_a;
   wire[6:0]  clka_ratio_adjusted_b;
   wire[6:0]  clkb_ratio_adjusted_a;
   wire[6:0]  clkb_ratio_adjusted_b;
   reg[5:0]   clka_ratio_fa;
   reg[5:0]   clkb_ratio_fa;
   reg[5:0]   clka_ratio_fb;
   reg[5:0]   clkb_ratio_fb;
   wire[6:0]  clka_ratio_twos;
   wire[6:0]  clkb_ratio_twos;

   assign     freq_match = clka_ratio == clkb_ratio;
   assign clka_ratio_adjusted[6:0] = {1'b0, clka_ratio[5:0]} + 7'b0000001;
   assign clkb_ratio_adjusted[6:0] = {1'b0, clkb_ratio[5:0]} + 7'b0000001;
   assign clka_ratio_adjusted_a[6:0] = {1'b0, clka_ratio_fa[5:0]} + 7'b0000001;
   assign clka_ratio_adjusted_b[6:0] = {1'b0, clka_ratio_fb[5:0]} + 7'b0000001;
   assign clkb_ratio_adjusted_a[6:0] = {1'b0, clkb_ratio_fa[5:0]} + 7'b0000001;
   assign clkb_ratio_adjusted_b[6:0] = {1'b0, clkb_ratio_fb[5:0]} + 7'b0000001;
   assign clka_ratio_twos[6:0]       = ~clka_ratio_adjusted[6:0] + 7'b0000001;
   assign clkb_ratio_twos[6:0]       = ~clkb_ratio_adjusted[6:0] + 7'b0000001;
   assign clka_error_tmp[6:0]      = {clkb_ratio_twos[6], clkb_ratio_twos[6:1]};
   assign clkb_error_tmp[6:0]      = {clka_ratio_twos[6], clka_ratio_twos[6:1]};

   always@(posedge clka)
     if(clka_usync)
       begin
	  clka_ratio_fa <= clka_ratio;
       end
     else
       begin
	  clka_ratio_fa <= clka_ratio_fa;
       end
   always@(posedge clka)
     if(clka_usync)
       begin
	  clkb_ratio_fa <= clkb_ratio;
       end
     else
       begin
	  clkb_ratio_fa <= clkb_ratio_fa;
       end
   always@(posedge clkb)
     if(clkb_usync)
       begin
	  clka_ratio_fb <= clka_ratio;
       end
     else
       begin
	  clka_ratio_fb <= clka_ratio_fb;
       end
   always@(posedge clkb)
     if(clkb_usync)
       begin
	  clkb_ratio_fb <= clkb_ratio;
       end
     else
       begin
	  clkb_ratio_fb <= clkb_ratio_fb;
       end
     
   always@(posedge clka)
     if(clka_usync)
       begin
          clka_error[6:0] <= clka_error_tmp[6:0];
       end
     else
       begin
         clka_error[6:0] <= clka_error[6] ?
                      (clka_error[6:0] + clka_ratio_adjusted_a[6:0] - clkb_ratio_adjusted_a[6:0]) :
                      (clka_error[6:0] - clkb_ratio_adjusted_a[6:0]);
       end
       
   always@(posedge clkb)
     if(clkb_usync)
       begin
          clkb_error[6:0] <= clkb_error_tmp[6:0];
       end
     else
       begin
         clkb_error[6:0] <= clkb_error[6] ?
                      (clkb_error[6:0] + clkb_ratio_adjusted_b[6:0] - clka_ratio_adjusted_b[6:0]) :
                      (clkb_error[6:0] - clka_ratio_adjusted_b[6:0]);
       end

   always_comb
     begin
        if (clka_ratio_fa[5:0] == clkb_ratio_fa[5:0] | test_override)
            begin
               clka_qual = 1'b1;
            end
        else if (clka_ratio_fa[5:0] > clkb_ratio_fa[5:0])
            begin
               clka_qual = clka_error[6];
            end
        else
            begin
               clka_qual = 1'b1;
            end   
     end // always_comb
   
   always_comb
     begin
        if (clka_ratio_fb[5:0] == clkb_ratio_fb[5:0] | test_override)
            begin
               clkb_qual = 1'b1;
            end
        else if (clka_ratio_fb[5:0] > clkb_ratio_fb[5:0])
            begin
               clkb_qual = 1'b1;
            end
        else
            begin
               clkb_qual = clkb_error[6];
            end   
     end
endmodule // qual_gen
 -----/\----- EXCLUDED -----/\----- */



// `define MAKE_CLK_SAMPLE_GEN(squash_clk, clk_sample, local_rstb, base_clk,reset_n, clk_enable, squash_div, test_override_en, test_override_div, test_over_div )                   \
// clk_sample_gen \``clk_sample_gen_``squash_clk (                                                                                                                                                                          \
//                                                             .squash_clk(squash_clk),                                                                                           \
//                                                             .clk_sample(clk_sample),                                                                                                                 \
//                                                             .local_rstb(local_rstb),                                                                                                                       \
//                                                             .base_clk(base_clk),                                                                                                           \
//                                                             .reset_n(reset_n),                                                                                                                                              \
//                                                             .clk_enable(clk_enable)                                                                                                                   \
//                                                             .squash_div(squash_div)                                                                                                                 \
//                                                             .test_override_en(test_override_en)                                                                                                       \
//                                                             .test_override_div(test_override_div)                                                                                                      \
//                                                             .test_over_div(test_over_div)                                                                                                      \
//                                                           );
// 
// module clk_sample_gen
//   #(parameter dWidth = 4) 
//     (
//    input logic                  base_clk,
//    input logic                  reset_n,      
//    input logic                  clk_enable,
//    input logic [(dWidth - 1):0] squash_div,
//    input logic                  test_override_en,
//    input logic                  test_override_div,
//    input logic [(dWidth - 1):0] test_over_div,
//    output logic                 local_rstb,
//    output logic                 clk_sample,
//    output logic                 squash_clk
// );
// 
//    logic  [(dWidth - 1):0] count, up_down_count;
//    logic                   clk_sample_i;
//    logic                   byp_div_atspeed;
//    logic                   test_mode_atspeed;
//    logic                   int_rstb, int_clk_enable, sync_clk_enable, int_squash_clk, temp_clk_en;
//    logic                       rst;
//    logic                   fall_edge_count;
//    logic                   fall_edge_clk;
//    
//        
// // synchronizing the reset and the enable to the output squash clock     
// `ip2211ringpll_ASYNC_RST_2MSFF_META(local_rstb, 1'b1, squash_clk , reset_n)
// 
// // synchronizing the internal reset and the enable to the base clock     
// `ip2211ringpll_ASYNC_RST_2MSFF_META(int_rstb, 1'b1, base_clk , reset_n)
// //`ip2211ringpll_ASYNC_RST_2MSFF_META(sync_clk_enable, int_clk_enable, base_clk , int_rstb)
// 
// // test mode will override the externa clock enable
// assign int_clk_enable = clk_enable | test_override_en;    
// 
//      // Using this to generate the clock adding the enable signal to the clock gate 
// `ip2211ringpll_CLK_GATE(squash_clk, base_clk, temp_clk_en)
// 
// //assign   temp_clk_en = (clk_sample_i & sync_clk_enable) | ~int_rstb;  
// assign   temp_clk_en = (clk_sample_i & int_clk_enable) | ~int_rstb; 
// 
//      // Standard up-down counter : squash_div must be stinkronized
//      // to base_clk which is not a end of CTS tree
// //   always @(posedge base_clk or negedge  int_rstb)
// //     if (~int_rstb)
// //    count <= 'b0;     // Divider initial 1 or 0
// //     else if (squash_div == 0)
// //    count <= 'b0;
// //     else if (((count < squash_div) & !test_override) || (test_override & (count < test_over_div)))
// //    count <= count + 1;
// //     else
// //    count <= 'b0;
// 
// 
// assign rst = ~int_rstb;
// assign up_down_count = ((squash_div != 0) & (((count < squash_div) & !test_override_div) || (test_override_div & (count < test_over_div)))) ? (count + 1) : 'b0;
// `ip2211ringpll_ASYNC_RST_MSFF(count,up_down_count,base_clk,rst)  
// 
//      // Falling edge used to clock forward the sample signal
// //   always @(negedge base_clk or negedge int_rstb)
// //     if (~int_rstb)
// //         clk_sample_i <= 'b1;     
// //     else if (~sync_clk_enable)    // I1 control
// //     clk_sample_i <= 'b0;
// //     else if ( count == 0 )
// //     clk_sample_i <= 'b1;
// //     else
// //     clk_sample_i <= 'b0;
// //
// //   assign clk_sample = clk_sample_i;
// 
// //assign fall_edge_count = (sync_clk_enable & ( count == 0 )) ? 1'b1: 1'b0;
// assign fall_edge_count = ( count == 0 ) ? 1'b1: 1'b0;
// //assign fall_edge_clk = ~base_clk;
// `ip2211ringpll_MAKE_CLK_INV (fall_edge_clk,base_clk)
// // CLOCK Sample needs to be 1 during reset
// `ip2211ringpll_ASYNC_SET_MSFF(clk_sample_i,fall_edge_count,fall_edge_clk,rst)  
// assign clk_sample = clk_sample_i;
// 
//    
// endmodule // clk_sample_gen


///============================================================================================
///
/// Clocks
///
///============================================================================================

// changing all the clock macros to add an extra module level of hierarchy



/* -----\/----- EXCLUDED -----\/-----
module det_clkdomainX #(parameter dWidth = 32, parameter fifo_depth = 10, parameter separation = 2) 
//  for synchronization that's done between two clocks that are derived from the same reference clock and use separation 1,
// this synchronizer must initiate it's rd/wr pointers at usync and not at reset!
// otherwise separation is not ensured.
// module det_clkdomainX must be abandoned and only this module det_clkdomainX_with_usync must be used.
(
                      input reset_ckRd,
                      input reset_ckWr,
                      input ckWr,
                      input ckRd,
                      input qualWr,
                      input qualRd,
                      input [dWidth-1:0] data_in,
                      output [dWidth-1:0] data_out
                      );

   logic [dWidth-1:0] det_clkdomainX_write_data_array[fifo_depth - 1:0];
   logic [dWidth-1:0] det_clkdomainX_read_data_mux;
   logic [fifo_depth - 1:0] wrptr;
   logic [fifo_depth - 1:0] rdptr;
   logic [fifo_depth - 1:0] start_ptr;
   logic write_clk;
   logic read_clk;

   `ip2211ringpll_CLK_GATE(write_clk, ckWr, qualWr)
   `ip2211ringpll_CLK_GATE(read_clk, ckRd, qualRd)
  
   // data path generation
   always @(posedge write_clk or negedge reset_ckWr)
     begin: write_clk_scope
        integer i;
        if (~reset_ckWr)
          begin
             for (i=0;i<fifo_depth;i=i+1)
               begin
                  det_clkdomainX_write_data_array[i] <= 0;
               end
          end
        else
          begin
             for (i=0;i<fifo_depth;i=i+1)
               begin
                  if (wrptr[i])
                    det_clkdomainX_write_data_array[i] <= data_in;
               end
          end
     end

   always @(posedge read_clk or negedge reset_ckRd)
     begin: read_clk_scope
        integer i;
        if (~reset_ckRd)
          begin
             det_clkdomainX_read_data_mux <= 0;
          end
        else
          begin
             for (i=0;i<fifo_depth;i=i+1)
               begin
                  if (rdptr[i])
                    det_clkdomainX_read_data_mux <= det_clkdomainX_write_data_array[i];
               end
          end
     end

   assign data_out = det_clkdomainX_read_data_mux;

   // wrptr and rdptr generation
   assign start_ptr = 1;
   
   always@(posedge write_clk or negedge reset_ckWr)
     if(!reset_ckWr)
       wrptr <= start_ptr << separation;
     else
       wrptr <= {wrptr[(fifo_depth - 2):0], wrptr[(fifo_depth - 1)]};

   always@(posedge read_clk or negedge reset_ckRd)
     if(!reset_ckRd)
       rdptr <= start_ptr;
     else
       rdptr <= {rdptr[(fifo_depth - 2):0], rdptr[(fifo_depth - 1)]};

endmodule // det_clkdomainX


`ip2211ringpll_ASYNC_RST_2MSFF_META(rstoutsync1b,1'b1,clkin1,rstb)
`ip2211ringpll_ASYNC_RST_2MSFF_META(rstoutsync2b,1'b1,clkin2,rstb)

`ip2211ringpll_ASYNC_RST_2MSFF_META(sync1_out,sync1_in,clkin1,rstoutsync1b)
`ip2211ringpll_ASYNC_RST_2MSFF_META(sync1_out_sel, sync1_out,clkin1,rstoutsync1b)

`ip2211ringpll_ASYNC_RST_2MSFF_META(sync2_out,sync2_in,clkin2,rstoutsync2b)
`ip2211ringpll_ASYNC_RST_2MSFF_META(sync2_out_sel,sync2_out,clkin2,rstoutsync2b)


`ip2211ringpll_MAKE_CLK_GLITCHFREE_MUX(clkout, clkin1, clkin2, sync1_out, sync2_out)

endmodule // async_clock_mux


`define ASYNC_CLK_MUX(mclkout,mclkin1,mclkin2,mselect1,mrstb)                                 \
async_clock_mux \``iasync_clock_mux_``mclkout (                                               \
                                  .select1  (mselect1),                                       \
                                  .clkin1  (mclkin1),                                         \
                                  .clkin2  (mclkin2),                                         \
                                  .rstb    (mrstb),                                           \
                                  .clkout  (mclkout)                                          \
                                );
 -----/\----- EXCLUDED -----/\----- */




`endif //  `ifndef ip2211ringpll_SOC_CLOCK_MACROS_VH  



/*******************************************************************************************************************
*
 *  MACROS NOT BEING USED BY ANYONE ELSE -  for
   *  ISSUES 
*  
*******************************************************************************************************************/



//`define MAKE_CLK_DELAY4(clkd4out,clkd4clkin,clkd4in0,clkd4in1,clkd4in2)    \
//clk4delay \``clk4delay_``clkd4out (                                          \
//                                    .clk4delayout (clkd4out),              \
//                                    .clk4delayin (clkd4clkin),             \
//                                    .clk4in0 (clkd4in0),                   \
//                                    .clk4in1 (clkd4in1),                   \
//                                    .clk4in2 (clkd4in2)                    \
//                                );
//
//`define LIB_clk4delay(clk4delayout,clk4delayin,clk4in0,clk4in1,clk4in2) \
//  vl0dcc04ln0a0 ck2(.o(clk4delayout),.clk(clk4delayin),.rsel0(clk4in0),.rsel1(clk4in1),.rsel2(clk4in2)); \
//
//module clk4delay (clk4delayout,clk4delayin,clk4in0,clk4in1,clk4in2);
//output clk4delayout;
//input clk4delayin;
//input clk4in0;
//input clk4in1;
//input clk4in2;
//wire clk4delayout,clk4delayin,clk4in0,clk4in1,clk4in2;
//`ifdef INTC_DC
//     `LIB_clk4delay(clk4delayout,clk4delayin,clk4in0,clk4in1,clk4in2) 
// `else
//assign clk4delayout = clk4delayin;
//`endif
//endmodule
//
//
//`define MAKE_CLK_DELAY8(clkd8out,clkd8clkin,clkd8in0,clkd8in1,clkd8in2,clkd8in3,clkd8in4,clkd8in5,clkd8in6)    \
//clk8delay \``clk8delay_``clkd8out (                                                         \
//                                    .clk8delayout (clkd8out),                             \
//                                    .clk8delayin (clkd8clkin),                            \
//                                    .clk8in0 (clkd8in0),                                  \
//                                    .clk8in1 (clkd8in1),                                  \
//                                    .clk8in2 (clkd8in2),                                  \
//                                    .clk8in3 (clkd8in3),                                  \
//                                    .clk8in4 (clkd8in4),                                  \
//                                    .clk8in5 (clkd8in5),                                  \
//                                    .clk8in6 (clkd8in6)                                   \
//                                );
//
//
//`define LIB_clk8delay(clk8delayout,clk8delayin,clk8in0,clk8in1,clk8in2,clk8in3,clk8in4,clk8in5,clk8in6) \
//  vl0dcc08ln0a0 ck2(.o(clk8delayout),.clk(clk8delayin),.rsel0(clk8in0),.rsel1(clk8in1),.rsel2(clk8in2),.rsel3(clk8in3),.rsel4(clk8in4),.rsel5(clk8in5),.rsel6(clk8in6)); \
//
//module clk8delay (clk8delayout,clk8delayin,clk8in0,clk8in1,clk8in2,clk8in3,clk8in4,clk8in5,clk8in6);
//output clk8delayout;
//input clk8delayin;
//input clk8in0;
//input clk8in1;
//input clk8in2;
//input clk8in3;
//input clk8in4;
//input clk8in5;
//input clk8in6;
//wire clk8delayout,clk8delayin,clk8in0,clk8in1,clk8in2,clk8in3,clk8in4,clk8in5,clk8in6;
//`ifdef INTC_DC
//     `LIB_clk8delay(clk8delayout,clk8delayin,clk8in0,clk8in1,clk8in2,clk8in3,clk8in4,clk8in5,clk8in6) 
// `else
//assign clk8delayout = clk8delayin;
//`endif
//endmodule
//
//
//`define MAKE_CLK_DIV2SHIFT(ckdiv2shftout,ipinckdiv2shftin,usyncdiv2shft)      \
// clk2div2shft \``clk_div2shift_``ckdiv2shftout (                                             \
//                                              .div2shftckdiv2shftout (ckdiv2shftout),      \
//                                              .div2shftipinckdiv2shftin (ipinckdiv2shftin),\
//                                              .div2shftusyncdiv2shft (usyncdiv2shft)       \
//                                             );
//
//module clk2div2shft (div2shftckdiv2shftout,div2shftipinckdiv2shftin,div2shftusyncdiv2shft);
//output div2shftckdiv2shftout;
//input div2shftipinckdiv2shftin;
//input div2shftusyncdiv2shft;
//reg div2shftckdiv2shftout;
//wire div2shftipinckdiv2shftin,div2shftusyncdiv2shft;
// reg ckdiv2shftout_ffout;                                                          
//  wire ckdiv2shftout_invout,ckdiv2shftout_andout,ckdiv2shftout_ckinvout;        
//  always_ff @(posedge div2shftipinckdiv2shftin)                                               
//      begin                                                                           
//       ckdiv2shftout_ffout   <= div2shftusyncdiv2shft;                                      
//      end  
//  assign ckdiv2shftout_invout = ~ckdiv2shftout_ffout;       
//  ip2211ringpll_clkinv clkinvdiv2shft (
//                         .clkout (ckdiv2shftout_ckinvout),
//                         .clkin (div2shftipinckdiv2shftin)
//                        );
//  assign  ckdiv2shftout_andout = (ckdiv2shftout_invout) & (~div2shftckdiv2shftout);     
//  clockdivff clockdivff_ckdiv2shftout (                                            
//                                   .ffout(div2shftckdiv2shftout),                             
//                                   .ffin(ckdiv2shftout_andout),                     
//                                   .clockin(ckdiv2shftout_ckinvout)                 
//                                  );
//endmodule
//
//                                             
//
//
//
//
//
//`define MAKE_CLK_LOCAL_QUALDIV100(div100clkout, div100_base_clk, div100_reset_n, div100_byp_div, div100_clk_disable, div100_squash_div)        \
//   crp_sample_gen_common #(100) \``make_clk_qualdiv100_``div100clksample (                                           \
//                                                    .base_clk              (div100_base_clk),                \
//                                                    .byp_div               (div100_byp_div),                 \
//                                                    .reset_n               (div100_reset_n),                 \
//                                                    .clk_disable           (div100_clk_disable),             \
//                                                    .squash_div            (div100_squash_div),              \
//                                                    .clk_out               (div100clkout)                    \
//                                                    );
//
//`define MAKE_CLK_LOCAL_QUALDIV16(outclk,inclk,ipinck,inusync)             \
//clkqualdiv16_local \``clk_qualdiv4_local``outclk (                               \
//                                   .divckout (outclk),                      \
//                                   .divckin  (inclk),                       \
//                                   .divipinckin(ipinck),                      \
//                                   .divusync (inusync)                            \
//                                  );
//
///* lintra s-31500, s-33048, s-33050 */
//module clkqualdiv16_local (divckout,divckin,divipinckin,divusync);
//   output divckout;
//   input  divckin;
//   input  divipinckin;
//   input  divusync;
//   reg    divckout;
//   wire   divckin,divusync;
//   reg    ckdiv16out_pout;                                                
//   reg [3:0] ckdiv16out_rstffpst;                                      
//   wire [3:0] ckdiv16out_rstffnxt;
//   logic       temp1, usync;
//   always_latch                                                         
//     begin                                                          
//        if (~divipinckin) ckdiv16out_pout  <= divusync;        
//     end                                                            
//   always_ff @(posedge divipinckin)                                 
//     begin                                                          
//        if (ckdiv16out_pout) ckdiv16out_rstffpst  <= '0;
//        else ckdiv16out_rstffpst  <=  ckdiv16out_rstffnxt;     
//     end                                                            
//   assign ckdiv16out_rstffnxt = ckdiv16out_rstffpst  + 1 ;           
//   assign usync = &ckdiv16out_rstffpst;
//   
//   clockdivff clockdivff_ckdiv16out(                                 
//                                   .ffout(temp1),                      
//                                   .ffin(usync),              
//                                   .clockin(divckin)                      
//                                   );
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp1)
//
//endmodule
//
//`define MAKE_CLK_LOCAL_QUALDIV2(ckout,ckin,ipinckin,usync)         \
// clkqualdiv_local \``clk_qualdiv2_``ckout (                         \
//                                         .divckout(ckout),       \
//                                         .divckin(ckin) ,        \
//                                         .divipinckin(ipinckin), \
//                                         .divusync(usync)          \
//                                         );
//
//
//
///* lintra s-31500, s-33048, s-33050 */
//`define MAKE_CLK_LOCAL_QUALDIV4(ckout2,ckin2,ipinckin2,usync2)            \
//clkqualdiv4_local \``clk_qualdiv4_local``ckout2 (                                \
//                                   .divckout (ckout2),             \
//                                   .divckin  (ckin2),              \
//                                   .divipinckin(ipinckin2),        \
//                                   .divusync (usync2)                \
//                                  );
//
//`define MAKE_CLK_LOCAL_QUALDIV600(div600clkout, div600_base_clk, div600_reset_n, div600_byp_div, div600_clk_disable, div600_squash_div)        \
//   crp_sample_gen_common #(600) \``make_clk_qualdiv600_``div600clksample (                                           \
//                                                    .base_clk              (div600_base_clk),                \
//                                                    .reset_n               (div600_reset_n),                 \
//                                                    .byp_div               (div600_byp_div),                 \
//                                                    .clk_disable           (div600_clk_disable),             \
//                                                    .squash_div            (div600_squash_div),              \
//                                                    .clk_out               (div600clkout)                    \
//                                                    );
//
//module crp_sample_gen_common  #(parameter dWidth = 3) 
//                     (
//                      input                  base_clk,       // Pre or Post CTS based on Physical Design
//                      input                  reset_n,        // Must be pre-stinkronized to base_clk input
//                      input                  byp_div,        // PMU Register input
//                      input                  clk_disable,    // PMU Register input
//                      input [(dWidth - 1):0] squash_div,     // PMU Register input
//                      output                 clk_out
//                      );
//
//   reg [(dWidth - 1):0]    count;
//   reg                     clk_sample_fe;
//   wire                    clk_sample;
//
//   // Standard up-down counter with some extras
//   always @(posedge base_clk or negedge reset_n )
//     if (~reset_n)
//       count         <= 'b0;     // Divider initial 1 or 0
//     else if (clk_disable || (squash_div == 0))
//       count         <= 'b0;
//     else if (count < squash_div)
//       count         <= count + 1;
//     else
//       count         <= 'b0;
//
//   // Falling edge used to clock forward the sample signal
//   always @(negedge base_clk or negedge reset_n )
//     if (~reset_n)
//       clk_sample_fe <= 'b0;     
//     else if (clk_disable)    // I1 control
//       clk_sample_fe <= 'b0;
//     else if ( count == 0 )
//       clk_sample_fe <= 'b1;
//     else
//       clk_sample_fe <= 'b0;
//
//   assign  clk_sample = byp_div ? 1'b1 : clk_sample_fe;
//
//   ip2211ringpll_soc_rbe_clk \``soc_rbe_clk_``clk_out (clk_out,base_clk,clk_sample);
//endmodule // clk_sample_gen
//
//
//`define MAKE_CLK_LOCAL_QUALDIV8(ckout2,ckin2,ipinckin2,usync2)            \
//clkqualdiv8_local \``clk_qualdiv4_local``ckout2 (                                \
//                                   .divckout (ckout2),             \
//                                  .divckin  (ckin2),              \
//                                   .divipinckin(ipinckin2),        \
//                                   .divusync (usync2)                \
//                                  );
///* lintra s-31500, s-33048, s-33050 */
//module clkqualdiv8_local (divckout,divckin,divipinckin,divusync);
//   output divckout;
//   input  divckin;
//   input  divipinckin;
//   input  divusync;
//   reg    divckout;
//   wire   divckin,divusync;
//   reg    ckdiv8out_pout;                                                
//   reg [2:0] ckdiv8out_rstffpst;                                      
//   wire [2:0] ckdiv8out_rstffnxt;
//   logic       temp1, temp2, usync;
//   always_latch                                                         
//     begin                                                          
//        if (~divipinckin) ckdiv8out_pout  <= divusync;        
//     end                                                            
//   always_ff @(posedge divipinckin)                                 
//     begin                                                          
//        if (ckdiv8out_pout) ckdiv8out_rstffpst  <= '0;          
//        else ckdiv8out_rstffpst  <=  ckdiv8out_rstffnxt;     
//     end                                                            
//   assign ckdiv8out_rstffnxt = ckdiv8out_rstffpst  + 1 ;           
//   assign usync = &ckdiv8out_rstffpst;
//   
//   clockdivff clockdivff_ckdiv8out(                                 
//                                   .ffout(temp1),                      
//                                   .ffin(usync),              
//                                   .clockin(divckin)                      
//                                   );
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp1)
//endmodule
//                                  
//
//`define MAKE_CLK_LOCAL_QUALDIV8_ADJ(ckout2,ckin2,ipinckin2,usync2, ratiosel2)            \
//clkqualdiv8_local_adj \``clk_qualdiv4_local_adj``ckout2 (                                \
//                                   .divckout (ckout2),             \
//                                   .divckin  (ckin2),              \
//                                   .divipinckin(ipinckin2),        \
//                                   .divusync (usync2),               \
//                                   .ratiosel (ratiosel2)                \
//                                  );
///* lintra s-31500, s-33048, s-33050 */
//module clkqualdiv8_local_adj (divckout,divckin,divipinckin,divusync,ratiosel);
//   output divckout;
//   input  divckin;
//   input  divipinckin;
//   input  divusync;
//   input [2:0] ratiosel;
//   reg    divckout;
///   wire   divckin,divusync;
//   reg    ckdiv8out_pout;                                                
//   reg [2:0] ckdiv8out_rstffpst;                                      
//   wire [2:0] ckdiv8out_rstffnxt;
//   logic       temp1, usync;
//
//   `ip2211ringpll_LATCH_P_DESKEW(ckdiv8out_pout, divusync, divipinckin)           
//   assign ckdiv8out_rstffnxt = ckdiv8out_rstffpst  + 1 ;
//   `ip2211ringpll_RST_MSFF(ckdiv8out_rstffpst, ckdiv8out_rstffnxt, divipinckin, ckdiv8out_pout)                   
//
//   always_comb
//     case(ratiosel)
//       3'b000 : usync = &ckdiv8out_rstffpst[2:0]; // div 8
//       3'b001 : usync = &ckdiv8out_rstffpst[1:0]; // div 4
//       3'b011 : usync = ckdiv8out_rstffpst[0];    // div 2
//       3'b111 : usync = 1'b1;                     // div 1
//       default: usync = 1'b1;
//     endcase // case(ratiosel)
//       
//   clockdivff clockdivff_ckdiv8out(                                 
//                                   .ffout(temp1),                      
//                                   .ffin(usync),              
//                                   .clockin(divckin)                      
//                                   );
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp1)
//endmodule
//
//// original MAKE_CLK_QUALDIV2 need to comment out after iosf is inplace
//`define MAKE_CLK_QUALDIV2(ckout,ckin,ipinckin,qual)         \
// clkqualdiv \``clk_qualdiv2_``ckout (                         \
//                                    .divckout(ckout),       \
//                                    .divckin(ckin) ,        \
//                                    .divipinckin(ipinckin), \
//                                    .divqual(qual)          \
//                                   );
//module clkqualdiv_local (divckout,divckin,divipinckin,divusync);
//output divckout;
//input divckin;
//input divipinckin;
//input divusync;
//   logic temp, temp1, temp2, temp3;
//    wire ckout_tmp1, ckout_tmp2, ckout_tmp, ckout_invclk;                                 
//   `ip2211ringpll_LATCH_P(temp, divusync, divipinckin)
//   `ip2211ringpll_MSFF(temp1, temp2, divipinckin)
//   assign temp2 = ~temp1 & ~temp;
//   `ip2211ringpll_MSFF(temp3, temp1, divckin)
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp3)
// 
//     /* lintra s-31500 */
//endmodule
//
//// original MAKE_CLK_QUALDIV4 - need to comment out after iosf in place
//`define MAKE_CLK_QUALDIV4(ckout2,ckin2,ipinckin2,qual2)            \
//clkqualdiv \``clk_qualdiv4_``ckout2 (                                \
//                                   .divckout (ckout2),             \
//                                   .divckin  (ckin2),              \
//                                   .divipinckin(ipinckin2),        \
//                                   .divqual (qual2)                \
//                                  );
//
//
//`define MAKE_QUAL_LOCAL_QUALDIV2(qual_out, inclk, inusync, inqualovrd)     \
// qualdiv2_local \``qualdiv2_``qual_out (                                         \
//                                         .qualifier_out(qual_out),       \
//                                         .ipinclk(inclk) ,                  \
//                                         .usync(inusync),                       \
//                                         .qualovrd(inqualovrd)                  \
//                                         );
//
///* lintra s-31500, s-33048, s-33050 */
//module qualdiv2_local (qualifier_out,ipinclk,usync,qualovrd);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
// 
//  logic usync_lat, qual_staged;
//  logic nxt, pst;
// 
//  `ip2211ringpll_LATCH_P(usync_lat, usync, ipinclk)
//  assign nxt = pst + 1;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_lat)
//  `ip2211ringpll_MSFF(qual_staged, pst, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule
// 
//`define MAKE_QUAL_LOCAL_QUALDIV4(qual_out, inclk, inusync, inqualovrd)     \
// qualdiv4_local \``qualdiv4_``qual_out (                                         \
//                                         .qualifier_out(qual_out),       \
//                                         .ipinclk(inclk) ,                  \
//                                         .usync(inusync),                       \
//                                         .qualovrd(inqualovrd)                  \
//                                         );
///* lintra s-31500, s-33048, s-33050 */
//module clkqualdiv4_local (divckout,divckin,divipinckin,divusync);
//   output divckout;
//   input  divckin;
//   input  divipinckin;
//   input  divusync;
//   reg    divckout;
//   wire   divckin,divusync;
//   reg    ckdiv4out_pout;                                                
//   reg [1:0] ckdiv4out_rstffpst;                                      
//   wire [1:0] ckdiv4out_rstffnxt;
//   logic       temp1, usync;
//   always_latch                                                         
//     begin                                                          
//        if (~divipinckin) ckdiv4out_pout  <= divusync;        
//     end                                                            
//   always_ff @(posedge divipinckin)                                 
//     begin                                                          
//        if (ckdiv4out_pout) ckdiv4out_rstffpst  <= '0;          
//        else ckdiv4out_rstffpst  <=  ckdiv4out_rstffnxt;     
//     end                                                            
//   assign ckdiv4out_rstffnxt = ckdiv4out_rstffpst  + 1 ;           
//   assign usync = &ckdiv4out_rstffpst;
//   
//   clockdivff clockdivff_ckdiv4out(                                 
//                                   .ffout(temp1),                      
//                                   .ffin(usync),              
//                                   .clockin(divckin)                      
//                                   );
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp1)
//endmodule
//
//// origianl clkqualdiv - need to remove after iosf is in place
//module clkqualdiv (divckout,divckin,divipinckin,divqual);
//output divckout;
//input divckin;
//input divipinckin;
//input divqual;
//wire divckout,divckin,divipinckin,divqual;
//`ifdef INTC_DC                                                                                         
//    wire ckout_tmp1, ckout_tmp2, ckout_tmp, ckout_invclk;                                 
//    `LIB_clkqualdiv(divckout,divckin,divipinckin,divqual) 
//`else                                                                                             
//reg ckout_qualout, ckout_qual1out;                                                            
// always @(negedge divipinckin)                                                                       
//   begin                                                                                          
//      ckout_qual1out = divqual; /* lintra s-60028 */
//   end                                                                                            
// always @(negedge divipinckin)                                                                       
//  begin                                                                                           
//      ckout_qualout  = ckout_qual1out; /* lintra s-60028 */
//   end                                                                                            
//   assign divckout = ckout_qualout & divckin;                                                     
//`endif     /* lintra s-31500 */
//endmodule
//
//
//                                        
//`define MAKE_QUAL_LOCAL_QUALDIV8(qual_out, inclk, inusync, inqualovrd)     \
// qualdiv8_local \``qualdiv8_``qual_out (                                         \
//                                        .qualifier_out(qual_out),       \
//                                         .ipinclk(inclk) ,                  \
//                                         .usync(inusync),                       \
//                                        .qualovrd(inqualovrd)                  \
//                                         );
//
///* lintra s-31500, s-33048, s-33050 */
//module qualdiv8_local (qualifier_out,ipinclk,usync,qualovrd);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
// 
//  logic usync_lat, qual_staged, qual;
//  logic [2:0] nxt;
//  logic [2:0] pst;
// 
//  `ip2211ringpll_LATCH_P(usync_lat, usync, ipinclk)
//  assign nxt = pst + 1;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_lat)
//  assign qual = (&(pst));
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule
//
//*****ANY USES OF MAKE_QUAL_LOCAL_QUALDIV8_ADJ SHOULD EVENTUALLY BE REPLACED BY 
//*****MAKE_QUAL_LOCAL_QUALDIV1TO8_ADJ WE CAN'T JUST CHANGE THIS MACRO AS IT WOULD CAUSE FAILS
// ML_FIX : Eventually need to remove this define and module
//`define MAKE_QUAL_LOCAL_QUALDIV8_ADJ(qual_out, inclk, inusync, inqualovrd, inratiosel)     \
// qualdiv8_adj_local \``qualdiv8adj_``qual_out (                                                   \
//                                         .qualifier_out(qual_out),                     \
//                                         .ipinclk(inclk) ,                                \
//                                         .usync(inusync),                                     \
//                                         .qualovrd(inqualovrd),                                \
//                                         .ratiosel(inratiosel)                                \
//                                         );
//
///* lintra s-31500, s-33048, s-33050 */
//module qualdiv8_adj_local (qualifier_out,ipinclk,usync,qualovrd,ratiosel);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
//  input [2:0] ratiosel;
// 
//  logic usync_lat, qual_staged, qual;
//  logic [2:0] nxt;
//  logic [2:0] pst;
// 
//  `ip2211ringpll_LATCH_P_DESKEW(usync_lat, usync, ipinclk)
//  assign nxt = pst + 1;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_lat)
//  always_comb begin
//    casex(ratiosel)
//      3'b000 : qual = &pst[2:0]; // div 8
//      3'b001 : qual = &pst[1:0]; // div 4
//      3'b011 : qual = pst[0];    // div 2
//      3'b111 : qual = 1'b1;      // div 1
//      default: qual = 1'b1;
//    endcase // case(ratiosel)
//  end
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule // qualdiv8_adj_local
//
//`define CLK_FF_INV(ckdiv2routb,ckdiv2rin,ckdiv2clkin,ckdiv2resetin)                       \
//clockdivffreset_inv \``clockdivffreset_inv_``ckdiv2routb (                                \
//                                                         .ffoutresetb(ckdiv2routb),       \
//                                                         .ffinreset(ckdiv2rin),           \
//                                                         .clockinreset(ckdiv2clkin),      \
//                                                         .resetckdivff(ckdiv2resetin)     \
//                                                        );
//
//module clockdivffreset_inv (ffoutresetb, ffinreset, clockinreset,resetckdivff);    
//output ffoutresetb;
//input ffinreset;
//input clockinreset;
//input resetckdivff;
//reg ffoutresetb;
//wire ffinreset, clockinreset, resetckdivff;
//`ifdef INTC_DC
//     `LIB_clockdivffreset(ffoutresetb, ffinreset, clockinreset,resetckdivff) 
//`else 
//always @(negedge (resetckdivff) or posedge clockinreset)
//begin
//  if (~(resetckdivff))
//    ffoutresetb = 1'b0; /* lintra s-60028 */
//  else
//    ffoutresetb = ~(ffinreset); /* lintra s-60028 */
//end
//`endif
//endmodule
//
//
//`define CLK_GATE_HF(o, clk, a)                                                               \
// soc_rbe_clk_hf \``soc_rbe_clk_hf_``o (                                                      \
//                                       .ckrcbxpn  (o),                                       \
//                                       .ckgridxpn (clk),                                     \
//                                       .latrcben  (a)                                        \
//                                      );
//module soc_rbe_clk_hf (output logic ckrcbxpn, input logic ckgridxpn, latrcben);  //lintra s-51506
//
//`ifdef INTC_DC
//     `LIB_soc_rbe_clk_hf(ckrcbxpn,ckgridxpn,latrcben) 
//`else
//   logic latrcbenl; // rce state element
//  
//  `ip2211ringpll_LATCH_P(latrcbenl, latrcben, ckgridxpn) //lintra s-51552
//  `ip2211ringpll_CLKAND(ckrcbxpn,ckgridxpn,latrcbenl)
//`endif
//endmodule // soc_rbe_clk_hf
//
////CLKBF_GLITCH_GLOB is a clkbuf used to remove glitches
////It is coded as a buffer, but this doesnot match the schematics.
////NEED TO CHECK IF INTC_SYNTHESIS ISNT REPLACING THE CELL WITH A BUFFER
//`define CLKBF_GLITCH_GLOB(clkout, clkin)                          \
//`ifdef INTC_DC                                                         \
//   `LIB_CLKBF_GLITCH_GLOB(clkout,clkin)                           \
//`else                                                             \
//   assign clkout = clkin;                                         \
//`endif
//
//`define CLKDIVFF(iffout, iffin, iclockin)             \
//clockdivff \``clockdivff_``iffout (                   \
//                                   .ffout(iffout),    \
//                                   .ffin(iffin),      \
//                                   .clockin(iclockin) \
//);
//
//// creating FF module to be used by clock macros below
//module clockdivff (ffout, ffin, clockin);    
//output ffout;
//input ffin;
//input clockin;
//reg ffout;
//wire ffin, clockin;
//`ifdef INTC_DC 
//     wire ffin_b;
//     assign ffin_b = ~ffin;
//     `LIB_clockdivff(ffout, ffin_b, clockin) 
//`else                                                                         
// always @(posedge clockin)                                                
//      begin                                                                  
//         ffout = ffin; /* lintra s-60028 */
//      end 
//`endif
//endmodule
//
//`define MAKE_CLK_GATE_TRUNK(igatedclk, iipclk, iusync, iresetb, iclken, idfx_scan_dbg_mode) \
//   clk_gate_trunk \``clk_gate_trunk_``igatedclk (                                           \
//                                                 .gatedclk(igatedclk),                      \
//                                                 .ipclk(iipclk),                            \
//                                                 .usync(iusync),                            \
//                                                 .resetb(iresetb),                          \
//                                                 .clken(iclken),                            \
//                                                 .dfx_scan_dbg_mode(idfx_scan_dbg_mode)     \
//                                                );
//
//module clk_gate_trunk(output logic gatedclk,
//                      input logic ipclk,
//                      input logic usync,
//                      input logic resetb,
//                      input logic clken,
//                      input logic dfx_scan_dbg_mode);
//logic clken_qual_in, clken_qual_out;
//logic qual_or_ovrd;
//assign clken_qual_in = usync ? clken : clken_qual_out;
//`ip2211ringpll_SET_MSFF(clken_qual_out, clken_qual_in, ipclk, ~resetb)
//assign qual_or_ovrd = clken_qual_out | dfx_scan_dbg_mode;
//`CLK_GATE_HF(gatedclk, ipclk, qual_or_ovrd)
//endmodule
//                                                
//











//`define MAKE_CLK_LOCAL_QUALDIV1TO16_ADJ(qual_out,inclk,inusync,inqualovrd,inratiosel)     \
//clk_qualdiv1to16_adj_local \``clk_qualdiv1to16_adj_local_``qual_out (                           \
//                                                                  .qualclk_out(qual_out),    \
//                                                                  .clk(inclk),               \
//                                                                  .usync(inusync),           \
//                                                                  .qualovrd(inqualovrd),     \
//                                                                  .ratiosel(inratiosel)     \
//                                                                 ); /* lintra s-51500, s-53048, s-53050 */
//
//module clk_qualdiv1to16_adj_local(qualclk_out, clk, usync, qualovrd, ratiosel);
//  output qualclk_out;
//  input clk;
//  input usync;
//  input qualovrd;
//  input [3:0] ratiosel;
//  logic qual_out;
//  `MAKE_QUAL_LOCAL_QUALDIV1TO8_ADJ(qual_out, clk, usync, qualovrd, ratiosel)        
//  `ip2211ringpll_CLK_GATE(qualclk_out, clk,  qual_out)
//endmodule
//
//
//
//`define MAKE_CLK_LOCAL_QUALDIV1TO8_ADJ(qual_out,inclk,inusync,inqualovrd,inratiosel)     \
//clk_qualdiv1to8_adj_local \``clk_qualdiv1to8_adj_local_``qual_out (                           \
//                                                                  .qualclk_out(qual_out),    \
//                                                                  .clk(inclk),               \
//                                                                  .usync(inusync),           \
//                                                                  .qualovrd(inqualovrd),     \
//                                                                  .ratiosel(inratiosel)     \
//                                                                 ); /* lintra s-51500, s-53048, s-53050 */
//module clk_qualdiv1to8_adj_local(qualclk_out, clk, usync, qualovrd, ratiosel);
//  output qualclk_out;
//  input clk;
//  input usync;
//  input qualovrd;
//  input [2:0] ratiosel;
//  logic qual_out;
//  `MAKE_QUAL_LOCAL_QUALDIV1TO8_ADJ(qual_out, clk, usync, qualovrd, ratiosel)        
//  `ip2211ringpll_CLK_GATE(qualclk_out, clk,  qual_out) //lintra s-51557, s-51552
//endmodule
//
//`define MAKE_CLK_NOREN(cknorenout,cknorenckin,cknorenenin)              \
//clknoren \``clknoren_``cknorenout (                                     \
//                              .clknorenout (cknorenout),                \
//                              .clknorenckin (cknorenckin),              \
//                              .clknorenenin (cknorenenin)               \
//                             );
//
//module clknoren(clknorenout,clknorenckin,clknorenenin);
//output clknorenout;
//input clknorenckin;
//input clknorenenin;
//wire clknorenout,clknorenckin,clknorenenin;
//`ifdef INTC_DC
//     `LIB_clknoren(clknorenout,clknorenckin,clknorenenin) 
//`else
//assign clknorenout = ~(clknorenckin|clknorenenin);
//`endif
//endmodule
//



//
//`define MAKE_QUAL_LOCAL_QUALDIV16(qual_out, inclk, inusync, inqualovrd)          \
// qualdiv16_local \``qualdiv16_``qual_out (                                       \
//                                         .qualifier_out(qual_out),               \
//                                         .ipinclk(inclk) ,                       \
//                                         .usync(inusync),                        \
//                                         .qualovrd(inqualovrd)                   \
//                                         );
//module qualdiv16_local (qualifier_out,ipinclk,usync,qualovrd);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
// 
//  logic usync_lat, qual_staged, qual;
//  logic [3:0] nxt;
//  logic [3:0] pst;
// 
//  `ip2211ringpll_LATCH_P_DESKEW(usync_lat, usync, ipinclk)
//  assign nxt = pst + 4'b0001;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_lat)
//  assign qual = (&(pst));
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule
//
//`define MAKE_QUAL_LOCAL_QUALDIV1TO16_ADJ(qual_out, inclk, inusync, inqualovrd, inratiosel)     \
// qualdiv1to16_adj_local \``qualdiv1to16adj_``qual_out (                                         \
//                                                    .qualifier_out(qual_out),                 \
//                                                    .ipinclk(inclk) ,                         \
//                                                    .usync(inusync),                          \
//                                                    .qualovrd(inqualovrd),                    \
//                                                    .ratiosel(inratiosel)                     \
//                                                    );
///* lintra s-51500, s-53048, s-53050 */
//module qualdiv1to16_adj_local (qualifier_out,ipinclk,usync,qualovrd,ratiosel);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
//  input [3:0] ratiosel;
// 
//  logic usync_or_qual_lat, usync_or_qual, qual_staged, qual;
//  logic [3:0] ratiosel_muxed_staged, ratiosel_muxed;
//  logic [3:0] nxt;
//  logic [3:0] pst;
// 
//  //Whenever a qual or usync comes through we reset the counter
//  assign usync_or_qual = usync | qual;
//
//  `ip2211ringpll_LATCH_P_DESKEW(usync_or_qual_lat, usync_or_qual, ipinclk)
//  assign nxt = pst + 4'b0001;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_or_qual_lat)
//
//  //only grab ratiosel on usync boundary
//  assign ratiosel_muxed = usync ? ratiosel : ratiosel_muxed_staged;
//  `ip2211ringpll_MSFF(ratiosel_muxed_staged, ratiosel_muxed, ipinclk)
//
//  //Once we've reached the count that matches the ratiosel we're dividing by
//  //Set the qual indicator and reset the count
//  assign qual = (pst == ratiosel_muxed_staged);
//
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule // qualdiv1to16_adj_local
//
//`define MAKE_QUAL_LOCAL_QUALDIV1TO8_ADJ_WEN(qual_out, inclk, inusync, inqualovrd, inratiosel, inenable)     \
// qualdiv1to8_adj_wen_local \``qualdiv1to8adjwen_``qual_out (                                         \
//                                                    .qualifier_out(qual_out),                 \
//                                                    .ipinclk(inclk) ,                         \
//                                                    .usync(inusync),                          \
//                                                    .qualovrd(inqualovrd),                    \
//                                                    .ratiosel(inratiosel),                    \
//                                                    .enable(inenable)                         \
//                                                    );
///* lintra s-51500, s-53048, s-53050 */
//module qualdiv1to8_adj_wen_local (qualifier_out,ipinclk,usync,qualovrd,ratiosel,enable);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
//  input [2:0] ratiosel;
//  input enable;
// 
//  logic usync_or_qual_lat, usync_or_qual, qual_staged, qual;
//  logic [2:0] ratiosel_muxed_staged, ratiosel_muxed;
//  logic [2:0] nxt;
//  logic [2:0] pst;
// 
//  //Whenever a qual or usync comes through we reset the counter
//  assign usync_or_qual = usync | qual;
//
//  `ip2211ringpll_LATCH_P_DESKEW(usync_or_qual_lat, usync_or_qual, ipinclk)
//  assign nxt = pst + 1;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_or_qual_lat)
//
//  //only grab ratiosel on usync boundary
//  assign ratiosel_muxed = usync ? ratiosel : ratiosel_muxed_staged;
//  `ip2211ringpll_MSFF(ratiosel_muxed_staged, ratiosel_muxed, ipinclk)
//
//  //Once we've reached the count that matches the ratiosel we're dividing by
//  //Set the qual indicator and reset the count
//  assign qual = (pst == ratiosel_muxed_staged);
//
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = (qual_staged & enable) | qualovrd;
//endmodule // qualdiv1to8_adj_wen_local
//
//
////module qual_5_2(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [2:0]           count;
//
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 3'b000;
//     else
//       count <= (count + 3'b001) & {3{~(count == 4)}};
//
//   assign              fast_qual = (count == 0  ||
//                                    count == 3);
//   assign              slow_qual = 1'b1;
//endmodule //qual_5_2
//
//
//module qual_1_1(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//  
//   assign              fast_qual = 1'b1;
//   assign              slow_qual = 1'b1;
//endmodule // qual_1_1
//
//module qual_4_3(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [1:0]           count;
//
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//
//   assign              fast_qual = ~(count == 2);
//   assign              slow_qual = 1'b1;
//endmodule // qual_4_3
//
//module qual_8_5(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [2:0]           count;
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//   assign              fast_qual = (count == 0 ||
//                                    count == 2 ||
//                                    count == 3 ||
//                                    count == 5 ||
//                                    count == 6);
//   assign              slow_qual = 1'b1;
//endmodule // qual_8_5
//
//module qual_2_1(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg                 count;
//
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//
//   assign              fast_qual = count == 0;

/* -----\/----- EXCLUDED -----\/-----
//This macro has a decrementing counter and hence we would see a low phase on
//the output clock when get the usync.
`define MAKE_CLK_DIV2OR4(idivoutclk, iipinclk, iusync, iseldiv2)     \
clkdiv2or4 \``clk_div_2or4_``idivoutclk (                            \
                                          .divoutclk(idivoutclk),    \
                                          .ipinclk(iipinclk),        \
                                          .usync(iusync),            \
                                          .seldiv2(iseldiv2)         \
                                        );

module clkdiv2or4 (divoutclk, ipinclk, usync, seldiv2);
output divoutclk;
input  ipinclk;
input  usync;
input  seldiv2;

logic [1:0] nxt;
logic [1:0] pst;
logic usync_lat;
logic divinclk;
logic divinclk_b;
`LATCH_P_DESKEW(usync_lat, usync, ipinclk)
`SET_MSFF(pst, nxt, ipinclk, usync_lat)
assign nxt = ~(|(pst))? 2'b11:(pst - 1);
assign divinclk_b = seldiv2? pst[0] : pst[1];
assign divinclk  = ~divinclk_b; 
clockdivff clockdivff_clkdiv2or4(
                                  .ffout(divoutclk),
                                  .ffin(divinclk),
                                  .clockin(ipinclk)
                                );
endmodule


`define MAKE_CLK_DIV8(ckdiv8out,ipinckdiv8in,usyncdiv8in)        \
clkdiv8 \``clk_div8_``ckdiv8out (                                \
                               .div8ckdiv8out (ckdiv8out),       \
                               .div8ipinckdiv8in (ipinckdiv8in), \
                               .div8usyncdiv8in (usyncdiv8in)    \
                              );

module clkdiv8 (div8ckdiv8out,div8ipinckdiv8in,div8usyncdiv8in);
output div8ckdiv8out;
input div8ipinckdiv8in;
input div8usyncdiv8in;
reg div8ckdiv8out;
wire div8ipinckdiv8in,div8usyncdiv8in;
reg ckdiv8out_pout;                                                
reg [2:0] ckdiv8out_rstffpst;                                      
wire [2:0] ckdiv8out_rstffnxt;                                     
wire ckdiv8out_invout;                                             
always_latch                                                         
      begin                                                          
         if (~div8ipinckdiv8in) ckdiv8out_pout  = div8usyncdiv8in; /-* lintra s-60028 *-/
      end                                                            
   always_ff @(posedge div8ipinckdiv8in)                                 
      begin                                                          
         if (ckdiv8out_pout) ckdiv8out_rstffpst  <= '0;          
         else ckdiv8out_rstffpst  <=  ckdiv8out_rstffnxt;     
      end                                                            
 assign ckdiv8out_rstffnxt = ckdiv8out_rstffpst  + 1 ;           
assign ckdiv8out_invout = ~ckdiv8out_rstffpst[2];                
clockdivff clockdivff_ckdiv8out (                                 
                             .ffout(div8ckdiv8out),                      
                             .ffin(ckdiv8out_invout),              
                             .clockin(div8ipinckdiv8in)                      
                            );
endmodule



`define MAKE_CLK_DIV4(ckdiv4out,ipinckdiv4in,usyncdiv4in)        \
clkdiv4 \``clk_div4_``ckdiv4out (                                \
                               .div4ckdiv4out (ckdiv4out),       \
                               .div4ipinckdiv4in (ipinckdiv4in), \
                               .div4usyncdiv4in (usyncdiv4in)    \
                              );


module clkdiv4 (div4ckdiv4out,div4ipinckdiv4in,div4usyncdiv4in);
output div4ckdiv4out;
input div4ipinckdiv4in;
input div4usyncdiv4in;
reg div4ckdiv4out;
wire div4ipinckdiv4in,div4usyncdiv4in;
reg ckdiv4out_pout;                                                
reg [1:0] ckdiv4out_rstffpst;                                      
wire [1:0] ckdiv4out_rstffnxt;                                     
wire ckdiv4out_invout;                                             
always_latch                                                         
      begin                                                          
         if (~div4ipinckdiv4in) ckdiv4out_pout  = div4usyncdiv4in; /-* lintra s-60028 *-/
      end                                                            
   always_ff @(posedge div4ipinckdiv4in)                                 
      begin                                                          
         if (ckdiv4out_pout) ckdiv4out_rstffpst  <= '0;          
         else ckdiv4out_rstffpst  <=  ckdiv4out_rstffnxt;     
      end                                                            
 assign ckdiv4out_rstffnxt = ckdiv4out_rstffpst  + 1 ;           
assign ckdiv4out_invout = ~ckdiv4out_rstffpst[1];                
clockdivff clockdivff_ckdiv4out (                                 
                             .ffout(div4ckdiv4out),                      
                             .ffin(ckdiv4out_invout),              
                             .clockin(div4ipinckdiv4in)                      
                            );
endmodule
 -----/\----- EXCLUDED -----/\----- */


/*
`define ip2211ringpll_MAKE_CLK_GLITCHFREE_MUX(clkout, clka, clkb, sela, selb)             	 \
ip2211ringpll_clk_glitchfree_mux_part \clk_glitchfree_mux_part_``clkout (                      \
                                                            .clk_out(clkout),    \
                                                            .clk_a(clka),        \
                                                            .clk_b(clkb),        \
                                                            .sel_a(sela),        \
                                                            .sel_b(selb)         \
                                                          );               

module ip2211ringpll_clk_glitchfree_mux_part (clk_out, clk_a, clk_b, sel_a, sel_b);
output clk_out;
input clk_a;
input clk_b;
input sel_a;
input sel_b;
logic sel_a_l, sel_b_l;

//`ifdef INTC_DC
        //  `LIB_clk_glitchfree_mux_part(clk_out, clk_a, clk_b, sel_a, sel_b)
//    ctech_lib_clk_mux_2to1_glitchfree ctech_lib_clk_mux_2to1_glitchfree(.clkout(clk_out),.clk1(clk_a),.clk2(clk_b),.s1(sel_a),.s2(sel_b));
//`else
  `ip2211ringpll_LATCH_P(sel_a_l, sel_a, clk_a)
  `ip2211ringpll_LATCH_P(sel_b_l, sel_b, clk_b)
  assign clk_out = (clk_a & sel_a_l) | (clk_b & sel_b_l);
//`endif
endmodule
*/
// New clock buffer macro only for SIPs that use thick gate library cells as are RTC in VLV

/* -----\/----- EXCLUDED -----\/-----
`define TG_CLKBF(clkbufout,clkbufin)                                                           \
//`ifdef INTC_DC                                                                                   \
//     `LIB_TG_CLKBF_SOC(clkbufout,clkbufin)                                                     \
// `else                                                                                      \
  `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                    \
                                                                                            \
   `endif                                                                                   \
     assign clkbufout =  (~(~(clkbufin)));                                                  \
// `endif
 -----/\----- EXCLUDED -----/\----- */


/* -----\/----- EXCLUDED -----\/-----
//programmable divider with usync, divivalonehot can one have one of the 10 bits high
//0000000001 is for div1 to 1000000000 is for div 10

`define MAKE_CLK_DIV_1_TO_10_USYNC(clkout, divvalonehot, clkin, usync, asyncrstb )      	\
div1to10macro_usync \div1to10macro_usync_``clkout (                      			\
                                                            .clk_out(clkout),    		\
                                                            .div_val_onehot(divvalonehot),      \
                                                            .clk_in(clkin),        		\
                                                            .usync_in(usync),        		\
                                                            .asyncrst_in(asyncrstb)         	\
                                                          );

module div1to10macro_usync (clk_out, div_val_onehot, clk_in, usync_in, asyncrst_in);
         input logic clk_in, usync_in,asyncrst_in;
         input logic [9:0] div_val_onehot;
         output logic clk_out;

         logic clk_in_b;

         logic usync_lat;
         logic divclk, divclk_p1,divclkout;
         logic divodd;
         logic [3:0] divsel_flop;

         logic div1, div2, div3, div4, div5, div6, div7, div8, div9, div10;
         logic q0,q1,q2,q3,q4;
         logic q1_or_fb,q2_or_fb,q3_or_fb,q4_or_fb,q5in;
         logic div1_b;

         logic q0in;
         logic q1in;
         logic q2in;
         logic q3in;
         logic q4in;
         
         // Generate clk_in_b
         `ip2211ringpll_MAKE_CLK_INV(clk_in_b,clk_in)

         // Latch the incoming usync to prevent min-vio
         `ip2211ringpll_LATCH_P_DESKEW(usync_lat, usync_in, clk_in)
         
         //Flop hte div-sel based on usync_lat
         // Capture new value on usync_lat, else keep the old value
         always_ff @(posedge clk_in or negedge asyncrst_in)
         begin
                 if(asyncrst_in == 1'b0)
                 begin
                          div1 <= 0;
                          div2 <= 0;
                          div3 <= 0;
                          div4 <= 0;
                          div5 <= 0;
                          div6 <= 0;
                          div7 <= 0;
                          div8 <= 0;
                          div9 <= 0;
                          div10 <= 0;
                 end
                 else     
                 if(usync_lat)
                 begin    
                          div1 <= div_val_onehot[0];
                          div2 <= div_val_onehot[1];
                          div3 <= div_val_onehot[2];
                          div4 <= div_val_onehot[3];
                          div5 <= div_val_onehot[4];
                          div6 <= div_val_onehot[5];
                          div7 <= div_val_onehot[6];
                          div8 <= div_val_onehot[7];
                          div9 <= div_val_onehot[8];
                          div10 <= div_val_onehot[9];
                 end
         end



                 // Shift-reg based counter
                 
                 assign fb = divodd ?~(q0|q1):~q0;
                 

                 //If the divsel value is invalue, do a div1

                 assign div3or4 = div3 | div4;
                 assign div5or6 = div5 | div6;
                 assign div7or8 = div7 | div8;
                 assign div9or10 = div9 | div10;
                 assign divodd = div3 | div5 | div7 | div9 ;        
                 
                 //the feedback point is selected based on the div-value
                 assign q1_or_fb = div2?fb:q1;
                 assign q2_or_fb = div3or4?fb:q2;
                 assign q3_or_fb = div5or6?fb:q3;
                 assign q4_or_fb = div7or8?fb:q4;
                 assign q5in = div9or10 & fb;

                 assign q0in = usync_lat ?1'b0:q1_or_fb;
                 assign q1in = usync_lat ?1'b0:q2_or_fb;
                 assign q2in = usync_lat ?1'b0:q3_or_fb;
                 assign q3in = usync_lat ?1'b0:q4_or_fb;
                 assign q4in = usync_lat ?1'b0:q5in;
                 

                 `ip2211ringpll_CLK_FF(q0,q0in,clk_in,asyncrst_in)
                 `ip2211ringpll_CLK_FF(q1,q1in,clk_in,asyncrst_in)
                 `ip2211ringpll_CLK_FF(q2,q2in,clk_in,asyncrst_in)
                 `ip2211ringpll_CLK_FF(q3,q3in,clk_in,asyncrst_in)
                 `ip2211ringpll_CLK_FF(q4,q4in,clk_in,asyncrst_in)
         
                 
                 //If it is div1, then just send out the input clock
                 assign divinclk = div1?1'b0:fb;   



                 `ip2211ringpll_CLK_FF(divclk,divinclk,clk_in,asyncrst_in)
                 //`ip2211ringpll_CLK_FF(divclk_p1,(divodd & divclk),~clk_in,asyncrst_in)
                 `ip2211ringpll_CLK_FF(divclk_p1,(divodd & divclk),clk_in_b,asyncrst_in)

                 assign divclkout = divodd?(divclk | divclk_p1):divclk;
                 
                 //assign clkout = div1?clk_in:divclk_out;
                 //clkmux_glitchfree iclkmx(.clka(clk_in),.clkb(divclkout),.sela(div1),.clkout(clk_out));
                assign div1_b = ~div1;

                 `ip2211ringpll_MAKE_CLK_GLITCHFREE_MUX(clk_out,clk_in,divclkout,div1,~div1)

                 
endmodule
 -----/\----- EXCLUDED -----/\----- */



/* -----\/----- EXCLUDED -----\/-----
//programmable divider  divivalonehot can one have one of the 10 bits high
//0000000001 is for div1 to 1000000000 is for div 10

`define MAKE_CLK_DIV_1_TO_10(clkout, divvalonehot, clkin, asyncrstb)             		\
div1to10macro \div1to10macro_``clkout (                      					\
                                                            .clk_out(clkout),    		\
                                                            .div_val_onehot(divvalonehot),      \
                                                            .clk_in(clkin),        		\
                                                            .asyncrst_in(asyncrstb)         	\
                                                          );

module div1to10macro (clk_out, div_val_onehot, clk_in, asyncrst_in);
                    input logic clk_in, asyncrst_in;
                    input logic [9:0] div_val_onehot;
                    output logic clk_out;

                    logic clk_in_b;

                    logic usync_lat;
                    logic divclk, divclk_p1,divclkout;
                    logic divodd;
                    logic [3:0] divsel_flop;

                    logic div1, div2, div3, div4, div5, div6, div7, div8, div9, div10;
                   logic div1_b;
                    logic q0,q1,q2,q3,q4;
                    logic q1_or_fb,q2_or_fb,q3_or_fb,q4_or_fb,q5in;

                    logic q0in;
                    logic q1in;
                    logic q2in;
                    logic q3in;
                    logic q4in;

                                        // Generate clk_in_b
                                        `ip2211ringpll_MAKE_CLK_INV(clk_in_b,clk_in)

                                        // Shift-reg based counter
                                        
                                        assign fb = divodd?~(q0|q1):~q0;
                                        

                                        //If the divsel value is invalue, do a div1

                                        assign div3or4 = div_val_onehot[2] | div_val_onehot[3];
                                        assign div5or6 = div_val_onehot[4] | div_val_onehot[5];
                                        assign div7or8 = div_val_onehot[6] | div_val_onehot[7];
                                        assign div9or10 = div_val_onehot[8] | div_val_onehot[9];
                                        assign divodd = div_val_onehot[2] | div_val_onehot[4] | div_val_onehot[6] | div_val_onehot[8] ;     
                                        
                                        //the feedback point is selected based on the div-value

                                        assign q0in = div_val_onehot[1]?fb:q1;
                                        assign q1in = div3or4?fb:q2;
                                        assign q2in = div5or6?fb:q3;
                                        assign q3in = div7or8?fb:q4;
                                        assign q4in = div9or10 & fb;

                                        `ip2211ringpll_CLK_FF(q0,q0in,clk_in,asyncrst_in)
                                        `ip2211ringpll_CLK_FF(q1,q1in,clk_in,asyncrst_in)
                                        `ip2211ringpll_CLK_FF(q2,q2in,clk_in,asyncrst_in)
                                        `ip2211ringpll_CLK_FF(q3,q3in,clk_in,asyncrst_in)
                                        `ip2211ringpll_CLK_FF(q4,q4in,clk_in,asyncrst_in)
                    
                                        
                                        //If it is div1, then just send out the input clock
                                        assign divinclk = div_val_onehot[0]?1'b0:fb; 



                                        `ip2211ringpll_CLK_FF(divclk,divinclk,clk_in,asyncrst_in)
                                        //`ip2211ringpll_CLK_FF(divclk_p1,(divodd & divclk),~clk_in,asyncrst_in)
                                        `ip2211ringpll_CLK_FF(divclk_p1,(divodd & divclk),clk_in_b,asyncrst_in)

                                        assign divclkout = divodd?(divclk | divclk_p1):divclk;
                                        
//                                       clkmux_glitchfree iclkmx(.clka(clk_in),.clkb(divclkout),.sela(div_val_onehot[0]),.clkout(clk_out));
                                      assign div1 =  div_val_onehot[0];
                                      assign div1_b =  ~div_val_onehot[0];

                                         `ip2211ringpll_MAKE_CLK_GLITCHFREE_MUX(clk_out, clk_in, divclkout, div1, div1_b)  
                                          
endmodule


   
module ip2211ringpll_clockdiv4ffreset (clk_in, reset_in, clk_out);
output clk_out;
input clk_in; 
input reset_in;
wire counter_0, counter_0_b, xor_out, nand_out, and_out, nor_out;
`ip2211ringpll_MAKE_CLK_INV(counter_0_b,counter_0) 
`ip2211ringpll_CLK_FF(counter_0,counter_0_b,clk_in,reset_in)
`ip2211ringpll_CLK_FF(clk_out,xor_out,clk_in,reset_in)
`ip2211ringpll_CLK_NAND(nand_out,counter_0,clk_out)
`ip2211ringpll_MAKE_CLK_INV(and_out,nand_out)    
`ip2211ringpll_MAKE_CLKNOR(nor_out,counter_0,clk_out)
`ip2211ringpll_MAKE_CLKNOR(xor_out,nor_out,and_out)
endmodule





/-* novas s-51500, s-53048, s-53050 *-/
module qualdiv1to8_adj_local (qualifier_out,ipinclk,usync,qualovrd,ratiosel);
  output qualifier_out;
  input ipinclk;
  input usync;
  input qualovrd;
  input [2:0] ratiosel;
 
  logic usync_or_qual_lat, usync_or_qual, qual_staged, qual;
  logic [2:0] ratiosel_muxed_staged, ratiosel_muxed;
  logic [2:0] nxt;
  logic [2:0] pst;
 
  //Whenever a qual or usync comes through we reset the counter
  assign usync_or_qual = usync | qual;

  `ip2211ringpll_LATCH_P_DESKEW(usync_or_qual_lat, usync_or_qual, ipinclk)
  assign nxt = pst + 3'b001;
  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_or_qual_lat)

  //only grab ratiosel on usync boundary
  assign ratiosel_muxed = usync ? ratiosel : ratiosel_muxed_staged;
  `ip2211ringpll_MSFF(ratiosel_muxed_staged, ratiosel_muxed, ipinclk)

  //Once we've reached the count that matches the ratiosel we're dividing by
  //Set the qual indicator and reset the count
  assign qual = (pst == ratiosel_muxed_staged);

  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
  assign qualifier_out = qual_staged | qualovrd;
endmodule // qualdiv1to8_adj_local
 -----/\----- EXCLUDED -----/\----- */

/* -----\/----- EXCLUDED -----\/-----
`define MAKE_QUAL_LOCAL_QUALDIV1TO8_ADJ(qual_out, inclk, inusync, inqualovrd, inratiosel)     \
 qualdiv1to8_adj_local \``qualdiv1to8adj_``qual_out (                                         \
                                                    .qualifier_out(qual_out),                 \
                                                    .ipinclk(inclk),                          \
                                                    .usync(inusync),                          \
                                                    .qualovrd(inqualovrd),                    \
                                                    .ratiosel(inratiosel)                     \
                                                    );



//this macro will divide the clk with output qualified with the period of the clk coming in//
//ratio stting for dividering is://
//Raiosel(2) ratiosel(1) ratiosel(0)//
//000 div1//
//001 div2//
//010 div3//
//011 div4//
//100 div5//
//101 div6//
//110 div7//
//111 div8//

module clk_qualdiv1to8_adj_local(xqualclk_out, xclk, xusync, xqualovrd, xratiosel);
  output xqualclk_out;
  input xclk;
  input xusync;
  input xqualovrd;
  input [2:0] xratiosel;
  logic xqual_out;
  `MAKE_QUAL_LOCAL_QUALDIV1TO8_ADJ(xqual_out, xclk, xusync, xqualovrd, xratiosel)        
  `ip2211ringpll_CLK_GATE(xqualclk_out, xclk,  xqual_out) //novas s-51557, s-51552
endmodule

`define CLK_QUALDIV1TO8_ADJ_LOCAL(qualclk_out, clk, usync, qualovrd, ratiosel )                 \
clk_qualdiv1to8_adj_local \``clk_qualdiv1to8_adj_local_``qualclk_out (                          \
                                                            .xqualclk_out(qualclk_out),         \
                                                            .xclk(clk),                         \
                                                            .xusync(usync),                     \
                                                            .xqualovrd(qualovrd),               \
                                                            .xratiosel(ratiosel)                \
                                                          );




module async_clock_mux
  (
   input logic select1,
   input logic clkin1,
   input logic clkin2,
   input logic rstb,
   output logic clkout
   );


logic sync1_in, sync2_in, sync1_out,sync2_out, rstoutsync1b, rstoutsync2b;
logic sync1_out_sel , sync2_out_sel;
assign sync1_in =  select1 & ~sync2_out_sel;
assign sync2_in = ~select1 & ~sync1_out_sel;



`ip2211ringpll_ASYNC_RST_2MSFF_META(rstoutsync1b,1'b1,clkin1,rstb)
`ip2211ringpll_ASYNC_RST_2MSFF_META(rstoutsync2b,1'b1,clkin2,rstb)

`ip2211ringpll_ASYNC_RST_2MSFF_META(sync1_out,sync1_in,clkin1,rstoutsync1b)
`ip2211ringpll_ASYNC_RST_2MSFF_META(sync1_out_sel, sync1_out,clkin1,rstoutsync1b)

`ip2211ringpll_ASYNC_RST_2MSFF_META(sync2_out,sync2_in,clkin2,rstoutsync2b)
`ip2211ringpll_ASYNC_RST_2MSFF_META(sync2_out_sel,sync2_out,clkin2,rstoutsync2b)


`ip2211ringpll_MAKE_CLK_GLITCHFREE_MUX(clkout, clkin1, clkin2, sync1_out, sync2_out)

endmodule // async_clock_mux


`define ASYNC_CLK_MUX(mclkout,mclkin1,mclkin2,mselect1,mrstb)                                 \
async_clock_mux \``iasync_clock_mux_``mclkout (                                               \
                                  .select1  (mselect1),                                       \
                                  .clkin1  (mclkin1),                                         \
                                  .clkin2  (mclkin2),                                         \
                                  .rstb    (mrstb),                                           \
                                  .clkout  (mclkout)                                          \
                                );
 -----/\----- EXCLUDED -----/\----- */




//`endif //  `ifndef ip2211ringpll_SOC_CLOCK_MACROS_VH  



/*******************************************************************************************************************
*
 *  MACROS NOT BEING USED BY ANYONE ELSE -  for
   *  ISSUES 
*  
*******************************************************************************************************************/



//`define MAKE_CLK_DELAY4(clkd4out,clkd4clkin,clkd4in0,clkd4in1,clkd4in2)    \
//clk4delay \``clk4delay_``clkd4out (                                          \
//                                    .clk4delayout (clkd4out),              \
//                                    .clk4delayin (clkd4clkin),             \
//                                    .clk4in0 (clkd4in0),                   \
//                                    .clk4in1 (clkd4in1),                   \
//                                    .clk4in2 (clkd4in2)                    \
//                                );
//
//`define LIB_clk4delay(clk4delayout,clk4delayin,clk4in0,clk4in1,clk4in2) \
//  vl0dcc04ln0a0 ck2(.o(clk4delayout),.clk(clk4delayin),.rsel0(clk4in0),.rsel1(clk4in1),.rsel2(clk4in2)); \
//
//module clk4delay (clk4delayout,clk4delayin,clk4in0,clk4in1,clk4in2);
//output clk4delayout;
//input clk4delayin;
//input clk4in0;
//input clk4in1;
//input clk4in2;
//wire clk4delayout,clk4delayin,clk4in0,clk4in1,clk4in2;
//`ifdef INTC_DC
//     `LIB_clk4delay(clk4delayout,clk4delayin,clk4in0,clk4in1,clk4in2) 
// `else
//assign clk4delayout = clk4delayin;
//`endif
//endmodule
//
//
//`define MAKE_CLK_DELAY8(clkd8out,clkd8clkin,clkd8in0,clkd8in1,clkd8in2,clkd8in3,clkd8in4,clkd8in5,clkd8in6)    \
//clk8delay \``clk8delay_``clkd8out (                                                         \
//                                    .clk8delayout (clkd8out),                             \
//                                    .clk8delayin (clkd8clkin),                            \
//                                    .clk8in0 (clkd8in0),                                  \
//                                    .clk8in1 (clkd8in1),                                  \
//                                    .clk8in2 (clkd8in2),                                  \
//                                    .clk8in3 (clkd8in3),                                  \
//                                    .clk8in4 (clkd8in4),                                  \
//                                    .clk8in5 (clkd8in5),                                  \
//                                    .clk8in6 (clkd8in6)                                   \
//                                );
//
//
//`define LIB_clk8delay(clk8delayout,clk8delayin,clk8in0,clk8in1,clk8in2,clk8in3,clk8in4,clk8in5,clk8in6) \
//  vl0dcc08ln0a0 ck2(.o(clk8delayout),.clk(clk8delayin),.rsel0(clk8in0),.rsel1(clk8in1),.rsel2(clk8in2),.rsel3(clk8in3),.rsel4(clk8in4),.rsel5(clk8in5),.rsel6(clk8in6)); \
//
//module clk8delay (clk8delayout,clk8delayin,clk8in0,clk8in1,clk8in2,clk8in3,clk8in4,clk8in5,clk8in6);
//output clk8delayout;
//input clk8delayin;
//input clk8in0;
//input clk8in1;
//input clk8in2;
//input clk8in3;
//input clk8in4;
//input clk8in5;
//input clk8in6;
//wire clk8delayout,clk8delayin,clk8in0,clk8in1,clk8in2,clk8in3,clk8in4,clk8in5,clk8in6;
//`ifdef INTC_DC
//     `LIB_clk8delay(clk8delayout,clk8delayin,clk8in0,clk8in1,clk8in2,clk8in3,clk8in4,clk8in5,clk8in6) 
// `else
//assign clk8delayout = clk8delayin;
//`endif
//endmodule
//
//
//`define MAKE_CLK_DIV2SHIFT(ckdiv2shftout,ipinckdiv2shftin,usyncdiv2shft)      \
// clk2div2shft \``clk_div2shift_``ckdiv2shftout (                                             \
//                                              .div2shftckdiv2shftout (ckdiv2shftout),      \
//                                              .div2shftipinckdiv2shftin (ipinckdiv2shftin),\
//                                              .div2shftusyncdiv2shft (usyncdiv2shft)       \
//                                             );
//
//module clk2div2shft (div2shftckdiv2shftout,div2shftipinckdiv2shftin,div2shftusyncdiv2shft);
//output div2shftckdiv2shftout;
//input div2shftipinckdiv2shftin;
//input div2shftusyncdiv2shft;
//reg div2shftckdiv2shftout;
//wire div2shftipinckdiv2shftin,div2shftusyncdiv2shft;
// reg ckdiv2shftout_ffout;                                                          
//  wire ckdiv2shftout_invout,ckdiv2shftout_andout,ckdiv2shftout_ckinvout;        
//  always_ff @(posedge div2shftipinckdiv2shftin)                                               
//      begin                                                                           
//       ckdiv2shftout_ffout   <= div2shftusyncdiv2shft;                                      
//      end  
//  assign ckdiv2shftout_invout = ~ckdiv2shftout_ffougmake run RUN_OPTS="-ucli -do vcs-fsdb.do"t;       
//  ip2211ringpll_clkinv clkinvdiv2shft (
//                         .clkout (ckdiv2shftout_ckinvout),
//                         .clkin (div2shftipinckdiv2shftin)
//                        );
//  assign  ckdiv2shftout_andout = (ckdiv2shftout_invout) & (~div2shftckdiv2shftout);     
//  clockdivff clockdivff_ckdiv2shftout (                                            
//                                   .ffout(div2shftckdiv2shftout),                             
//                                   .ffin(ckdiv2shftout_andout),                     
//                                   .clockin(ckdiv2shftout_ckinvout)                 
//                                  );
//endmodule
//
//                                             
//
//
//
//
//
//`define MAKE_CLK_LOCAL_QUALDIV100(div100clkout, div100_base_clk, div100_reset_n, div100_byp_div, div100_clk_disable, div100_squash_div)        \
//   crp_sample_gen_common #(100) \``make_clk_qualdiv100_``div100clksample (                                           \
//                                                    .base_clk              (div100_base_clk),                \
//                                                    .byp_div               (div100_byp_div),                 \
//                                                    .reset_n               (div100_reset_n),                 \
//                                                    .clk_disable           (div100_clk_disable),             \
//                                                    .squash_div            (div100_squash_div),              \
//                                                    .clk_out               (div100clkout)                    \
//                                                    );
//
//`define MAKE_CLK_LOCAL_QUALDIV16(outclk,inclk,ipinck,inusync)             \
//clkqualdiv16_local \``clk_qualdiv4_local``outclk (                               \
//                                   .divckout (outclk),                      \
//                                   .divckin  (inclk),                       \
//                                   .divipinckin(ipinck),                      \
//                                   .divusync (inusync)                            \
//                                  );
//
///* lintra s-31500, s-33048, s-33050 */
//module clkqualdiv16_local (divckout,divckin,divipinckin,divusync);
//   output divckout;
//   input  divckin;
//   input  divipinckin;
//   input  divusync;
//   reg    divckout;
//   wire   divckin,divusync;
//   reg    ckdiv16out_pout;                                                
//   reg [3:0] ckdiv16out_rstffpst;                                      
//   wire [3:0] ckdiv16out_rstffnxt;
//   logic       temp1, usync;
//   always_latch                                                         
//     begin                                                          
//        if (~divipinckin) ckdiv16out_pout  <= divusync;        
//     end                                                            
//   always_ff @(posedge divipinckin)                                 
//     begin                                                          
//        if (ckdiv16out_pout) ckdiv16out_rstffpst  <= '0;
//        else ckdiv16out_rstffpst  <=  ckdiv16out_rstffnxt;     
//     end                                                            
//   assign ckdiv16out_rstffnxt = ckdiv16out_rstffpst  + 1 ;           
//   assign usync = &ckdiv16out_rstffpst;
//   
//   clockdivff clockdivff_ckdiv16out(                                 
//                                   .ffout(temp1),                      
//                                   .ffin(usync),              
//                                   .clockin(divckin)                      
//                                   );
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp1)
//
//endmodule
//
//`define MAKE_CLK_LOCAL_QUALDIV2(ckout,ckin,ipinckin,usync)         \
// clkqualdiv_local \``clk_qualdiv2_``ckout (                         \
//                                         .divckout(ckout),       \
//                                         .divckin(ckin) ,        \
//                                         .divipinckin(ipinckin), \
//                                         .divusync(usync)          \
//                                         );
//
//
//
///* lintra s-31500, s-33048, s-33050 */
//`define MAKE_CLK_LOCAL_QUALDIV4(ckout2,ckin2,ipinckin2,usync2)            \
//clkqualdiv4_local \``clk_qualdiv4_local``ckout2 (                                \
//                                   .divckout (ckout2),             \
//                                   .divckin  (ckin2),              \
//                                   .divipinckin(ipinckin2),        \
//                                   .divusync (usync2)                \
//                                  );
//
//`define MAKE_CLK_LOCAL_QUALDIV600(div600clkout, div600_base_clk, div600_reset_n, div600_byp_div, div600_clk_disable, div600_squash_div)        \
//   crp_sample_gen_common #(600) \``make_clk_qualdiv600_``div600clksample (                                           \
//                                                    .base_clk              (div600_base_clk),                \
//                                                    .reset_n               (div600_reset_n),                 \
//                                                    .byp_div               (div600_byp_div),                 \
//                                                    .clk_disable           (div600_clk_disable),             \
//                                                    .squash_div            (div600_squash_div),              \
//                                                    .clk_out               (div600clkout)                    \
//                                                    );
//
//module crp_sample_gen_common  #(parameter dWidth = 3) 
//                     (
//                      input                  base_clk,       // Pre or Post CTS based on Physical Design
//                      input                  reset_n,        // Must be pre-stinkronized to base_clk input
//                      input                  byp_div,        // PMU Register input
//                      input                  clk_disable,    // PMU Register input
//                      input [(dWidth - 1):0] squash_div,     // PMU Register input
//                      output                 clk_out
//                      );
//
//   reg [(dWidth - 1):0]    count;
//   reg                     clk_sample_fe;
//   wire                    clk_sample;
//
//   // Standard up-down counter with some extras
//   always @(posedge base_clk or negedge reset_n )
//     if (~reset_n)
//       count         <= 'b0;     // Divider initial 1 or 0
//     else if (clk_disable || (squash_div == 0))
//       count         <= 'b0;
//     else if (count < squash_div)
//       count         <= count + 1;
//     else
//       count         <= 'b0;
//
//   // Falling edge used to clock forward the sample signal
//   always @(negedge base_clk or negedge reset_n )
//     if (~reset_n)
//       clk_sample_fe <= 'b0;     
//     else if (clk_disable)    // I1 control
//       clk_sample_fe <= 'b0;
//     else if ( count == 0 )
//       clk_sample_fe <= 'b1;
//     else
//       clk_sample_fe <= 'b0;
//
//   assign  clk_sample = byp_div ? 1'b1 : clk_sample_fe;
//
//   ip2211ringpll_soc_rbe_clk \``soc_rbe_clk_``clk_out (clk_out,base_clk,clk_sample);
//endmodule // clk_sample_gen
//
//
//`define MAKE_CLK_LOCAL_QUALDIV8(ckout2,ckin2,ipinckin2,usync2)            \
//clkqualdiv8_local \``clk_qualdiv4_local``ckout2 (                                \
//                                   .divckout (ckout2),             \
//                                  .divckin  (ckin2),              \
//                                   .divipinckin(ipinckin2),        \
//                                   .divusync (usync2)                \
//                                  );
///* lintra s-31500, s-33048, s-33050 */
//module clkqualdiv8_local (divckout,divckin,divipinckin,divusync);
//   output divckout;
//   input  divckin;
//   input  divipinckin;
//   input  divusync;
//   reg    divckout;
//   wire   divckin,divusync;
//   reg    ckdiv8out_pout;                                                
//   reg [2:0] ckdiv8out_rstffpst;                                      
//   wire [2:0] ckdiv8out_rstffnxt;
//   logic       temp1, temp2, usync;
//   always_latch                                                         
//     begin                                                          
//        if (~divipinckin) ckdiv8out_pout  <= divusync;        
//     end                                                            
//   always_ff @(posedge divipinckin)                                 
//     begin                                                          
//        if (ckdiv8out_pout) ckdiv8out_rstffpst  <= '0;          
//        else ckdiv8out_rstffpst  <=  ckdiv8out_rstffnxt;     
//     end                                                            
//   assign ckdiv8out_rstffnxt = ckdiv8out_rstffpst  + 1 ;           
//   assign usync = &ckdiv8out_rstffpst;
//   
//   clockdivff clockdivff_ckdiv8out(                                 
//                                   .ffout(temp1),                      
//                                   .ffin(usync),              
//                                   .clockin(divckin)                      
//                                   );
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp1)
//endmodule
//                                  
//
//`define MAKE_CLK_LOCAL_QUALDIV8_ADJ(ckout2,ckin2,ipinckin2,usync2, ratiosel2)            \
//clkqualdiv8_local_adj \``clk_qualdiv4_local_adj``ckout2 (                                \
//                                   .divckout (ckout2),             \
//                                   .divckin  (ckin2),              \
//                                   .divipinckin(ipinckin2),        \
//                                   .divusync (usync2),               \
//                                   .ratiosel (ratiosel2)                \
//                                  );
///* lintra s-31500, s-33048, s-33050 */
//module clkqualdiv8_local_adj (divckout,divckin,divipinckin,divusync,ratiosel);
//   output divckout;
//   input  divckin;
//   input  divipinckin;
//   input  divusync;
//   input [2:0] ratiosel;
//   reg    divckout;
///   wire   divckin,divusync;
//   reg    ckdiv8out_pout;                                                
//   reg [2:0] ckdiv8out_rstffpst;                                      
//   wire [2:0] ckdiv8out_rstffnxt;
//   logic       temp1, usync;
//
//   `ip2211ringpll_LATCH_P_DESKEW(ckdiv8out_pout, divusync, divipinckin)           
//   assign ckdiv8out_rstffnxt = ckdiv8out_rstffpst  + 1 ;
//   `ip2211ringpll_RST_MSFF(ckdiv8out_rstffpst, ckdiv8out_rstffnxt, divipinckin, ckdiv8out_pout)                   
//
//   always_comb
//     case(ratiosel)
//       3'b000 : usync = &ckdiv8out_rstffpst[2:0]; // div 8
//       3'b001 : usync = &ckdiv8out_rstffpst[1:0]; // div 4
//       3'b011 : usync = ckdiv8out_rstffpst[0];    // div 2
//       3'b111 : usync = 1'b1;                     // div 1
//       default: usync = 1'b1;
//     endcase // case(ratiosel)
//       
//   clockdivff clockdivff_ckdiv8out(                                 
//                                   .ffout(temp1),                      
//                                   .ffin(usync),              
//                                   .clockin(divckin)                      
//                                   );
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp1)
//endmodule
//
//// original MAKE_CLK_QUALDIV2 need to comment out after iosf is inplace
//`define MAKE_CLK_QUALDIV2(ckout,ckin,ipinckin,qual)         \
// clkqualdiv \``clk_qualdiv2_``ckout (                         \
//                                    .divckout(ckout),       \
//                                    .divckin(ckin) ,        \
//                                    .divipinckin(ipinckin), \
//                                    .divqual(qual)          \
//                                   );
//module clkqualdiv_local (divckout,divckin,divipinckin,divusync);
//output divckout;
//input divckin;
//input divipinckin;
//input divusync;
//   logic temp, temp1, temp2, temp3;
//    wire ckout_tmp1, ckout_tmp2, ckout_tmp, ckout_invclk;                                 
//   `ip2211ringpll_LATCH_P(temp, divusync, divipinckin)
//   `ip2211ringpll_MSFF(temp1, temp2, divipinckin)
//   assign temp2 = ~temp1 & ~temp;
//   `ip2211ringpll_MSFF(temp3, temp1, divckin)
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp3)
// 
//     /* lintra s-31500 */
//endmodule
//
//// original MAKE_CLK_QUALDIV4 - need to comment out after iosf in place
//`define MAKE_CLK_QUALDIV4(ckout2,ckin2,ipinckin2,qual2)            \
//clkqualdiv \``clk_qualdiv4_``ckout2 (                                \
//                                   .divckout (ckout2),             \
//                                   .divckin  (ckin2),              \
//                                   .divipinckin(ipinckin2),        \
//                                   .divqual (qual2)                \
//                                  );
//
//
//`define MAKE_QUAL_LOCAL_QUALDIV2(qual_out, inclk, inusync, inqualovrd)     \
// qualdiv2_local \``qualdiv2_``qual_out (                                         \
//                                         .qualifier_out(qual_out),       \
//                                         .ipinclk(inclk) ,                  \
//                                         .usync(inusync),                       \
//                                         .qualovrd(inqualovrd)                  \
//                                         );
//
///* lintra s-31500, s-33048, s-33050 */
//module qualdiv2_local (qualifier_out,ipinclk,usync,qualovrd);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
// 
//  logic usync_lat, qual_staged;
//  logic nxt, pst;
// 
//  `ip2211ringpll_LATCH_P(usync_lat, usync, ipinclk)
//  assign nxt = pst + 1;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_lat)
//  `ip2211ringpll_MSFF(qual_staged, pst, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule
// 
//`define MAKE_QUAL_LOCAL_QUALDIV4(qual_out, inclk, inusync, inqualovrd)     \
// qualdiv4_local \``qualdiv4_``qual_out (                                         \
//                                         .qualifier_out(qual_out),       \
//                                         .ipinclk(inclk) ,                  \
//                                         .usync(inusync),                       \
//                                         .qualovrd(inqualovrd)                  \
//                                         );
///* lintra s-31500, s-33048, s-33050 */
//module clkqualdiv4_local (divckout,divckin,divipinckin,divusync);
//   output divckout;
//   input  divckin;
//   input  divipinckin;
//   input  divusync;
//   reg    divckout;
//   wire   divckin,divusync;
//   reg    ckdiv4out_pout;                                                
//   reg [1:0] ckdiv4out_rstffpst;                                      
//   wire [1:0] ckdiv4out_rstffnxt;
//   logic       temp1, usync;
//   always_latch                                               `ifndef ip2211ringpll_SOC_CLOCK_MACROS_VH          
//     begin                                                          
//        if (~divipinckin) ckdiv4out_pout  <= divusync;        
//     end                                                            
//   always_ff @(posedge divipinckin)                                 
//     begin                                                          
//        if (ckdiv4out_pout) ckdiv4out_rstffpst  <= '0;          
//        else ckdiv4out_rstffpst  <=  ckdiv4out_rstffnxt;     
//     end                                                            
//   assign ckdiv4out_rstffnxt = ckdiv4out_rstffpst  + 1 ;           
//   assign usync = &ckdiv4out_rstffpst;
//   
//   clockdivff clockdivff_ckdiv4out(                                 
//                                   .ffout(temp1),                      
//                                   .ffin(usync),              
//                                   .clockin(divckin)                      
//                                   );
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp1)
//endmodule
//
//// origianl clkqualdiv - need to remove after iosf is in place
//module clkqualdiv (divckout,divckin,divipinckin,divqual);
//output divckout;
//input divckin;
//input divipinckin;
//input divqual;
//wire divckout,divckin,divipinckin,divqual;
//`ifdef INTC_DC                                                                                         
//    wire ckout_tmp1, ckout_tmp2, ckout_tmp, ckout_invclk;                                 
//    `LIB_clkqualdiv(divckout,divckin,divipinckin,divqual) 
//`else                                                                                             
//reg ckout_qualout, ckout_qual1out;                                                            
// always @(negedge divipinckin)                                                                       
//   begin                                                                                          
//      ckout_qual1out = divqual; /* lintra s-60028 */
//   end                                                                                            
// always @(negedge divipinckin)                                                                       
//  begin                                                                                           
//      ckout_qualout  = ckout_qual1out; /* lintra s-60028 */
//   end                                                                                            
//   assign divckout = ckout_qualout & divckin;                                                     
//`endif     /* lintra s-31500 */
//endmodule
//
//
//                                        
//`define MAKE_QUAL_LOCAL_QUALDIV8(qual_out, inclk, inusync, inqualovrd)     \
// qualdiv8_local \``qualdiv8_``qual_out (                                         \
//                                        .qualifier_out(qual_out),       \
//                                         .ipinclk(inclk) ,                  \
//                                         .usync(inusync),                       \
//                                        .qualovrd(inqualovrd)                  \
//                                         );
//
///* lintra s-31500, s-33048, s-33050 */
//module qualdiv8_local (qualifier_out,ipinclk,usync,qualovrd);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
// 
//  logic usync_lat, qual_staged, qual;
//  logic [2:0] nxt;
//  logic [2:0] pst;
// 
//  `ip2211ringpll_LATCH_P(usync_lat, usync, ipinclk)
//  assign nxt = pst + 1;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_lat)
//  assign qual = (&(pst));
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule
//
//*****ANY USES OF MAKE_QUAL_LOCAL_QUALDIV8_ADJ SHOULD EVENTUALLY BE REPLACED BY 
//*****MAKE_QUAL_LOCAL_QUALDIV1TO8_ADJ WE CAN'T JUST CHANGE THIS MACRO AS IT WOULD CAUSE FAILS
// ML_FIX : Eventually need to remove this define and module
//`define MAKE_QUAL_LOCAL_QUALDIV8_ADJ(qual_gmake run RUN_OPTS="-ucli -do vcs-fsdb.do"out, inclk, inusync, inqualovrd, inratiosel)     \
// qualdiv8_adj_local \``qualdiv8adj_``qual_out (                                                   \
//                                         .qualifier_out(qual_out),                     \
//                                         .ipinclk(inclk) ,                                \
//                                         .usync(inusync),                                     \
//                                         .qualovrd(inqualovrd),                                \
//                                         .ratiosel(inratiosel)                                \
//                                         );
//
///* lintra s-31500, s-33048, s-33050 */
//module qualdiv8_adj_local (qualifier_out,ipinclk,usync,qualovrd,ratiosel);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
//  input [2:0] ratiosel;
// 
//  logic usync_lat, qual_staged, qual;
//  logic [2:0] nxt;
//  logic [2:0] pst;
// 
//  `ip2211ringpll_LATCH_P_DESKEW(usync_lat, usync, ipinclk)
//  assign nxt = pst + 1;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_lat)
//  always_comb begin
//    casex(ratiosel)
//      3'b000 : qual = &pst[2:0]; // div 8
//      3'b001 : qual = &pst[1:0]; // div 4
//      3'b011 : qual = pst[0];    // div 2
//      3'b111 : qual = 1'b1;      // div 1
//      default: qual = 1'b1;
//    endcase // case(ratiosel)
//  end
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule // qualdiv8_adj_local
//
//`define CLK_FF_INV(ckdiv2routb,ckdiv2rin,ckdiv2clkin,ckdiv2resetin)                       \
//clockdivffreset_inv \``clockdivffreset_inv_``ckdiv2routb (                                \
//                                                         .ffoutresetb(ckdiv2routb),       \
//                                                         .ffinreset(ckdiv2rin),           \
//                                                         .clockinreset(ckdiv2clkin),      \
//                                                         .resetckdivff(ckdiv2resetin)     \
//                                                        );
//
//module clockdivffreset_inv (ffoutresetb, ffinreset, clockinreset,resetckdivff);    
//output ffoutresetb;
//input ffinreset;
//input clockinreset;
//input resetckdivff;
//reg ffoutresetb;
//wire ffinreset, clockinreset, resetckdivff;
//`ifdef INTC_DC
//     `LIB_clockdivffreset(ffoutresetb, ffinreset, clockinreset,resetckdivff) 
//`else 
//always @(negedge (resetckdivff) or posedge clockinreset)
//begin
//  if (~(resetckdivff))
//    ffoutresetb = 1'b0; /* lintra s-60028 */
//  else
//    ffoutresetb = ~(ffinreset); /* lintra s-60028 */
//end
//`endif
//endmodule
//
//
//`define CLK_GATE_HF(o, clk, a)                                                               \
// soc_rbe_clk_hf \``soc_rbe_clk_hf_``o (                                                      \
//                                       .ckrcbxpn  (o),                                       \
//                                       .ckgridxpn (clk),                                     \
//                                       .latrcben  (a)                                        \
//                                      );
//module soc_rbe_clk_hf (output logic ckrcbxpn, input logic ckgridxpn, latrcben);  //lintra s-51506
//
//`ifdef INTC_DC
//     `LIB_soc_rbe_clk_hf(ckrcbxpn,ckgridxpn,latrcben) 
//`else
//   logic latrcbenl; // rce state element
//  
//  `ip2211ringpll_LATCH_P(latrcbenl, latrcben, ckgridxpn) //lintra s-51552
//  `ip2211ringpll_CLKAND(ckrcbxpn,ckgridxpn,latrcbenl)
//`endif
//endmodule // soc_rbe_clk_hf
//
////CLKBF_GLITCH_GLOB is a clkbuf used to remove glitches
////It is coded as a buffer, but this doesnot match the schematics.
////NEED TO CHECK IF INTC_SYNTHESIS ISNT REPLACING THE CELL WITH A BUFFER
//`define CLKBF_GLITCH_GLOB(clkout, clkin)                          \
//`ifdef INTC_DC                                                         \
//   `LIB_CLKBF_GLITCH_GLOB(clkout,clkin)                           \
//`else                                                             \
//   assign clkout = clkin;                                         \
//`endif
//
//`define CLKDIVFF(iffout, iffin, iclockin)             \
//clockdivff \``clockdivff_``iffout (                   \
//                                   .ffout(iffout),    \
//                                   .ffin(iffin),      \
//                                   .clockin(iclockin) \
//);
//
//// creating FF module to be used by clock macros below
//module clockdivff (ffout, ffin, clockin);    
//output ffout;
//input ffin;
//input clockin;
//reg ffout;
//wire ffin, clockin;
//`ifdef INTC_DC 
//     wire ffin_b;
//     assign ffin_b = ~ffin;
//     `LIB_clockdivff(ffout, ffin_b, clockin) 
//`else                                                                         
// always @(posedge clockin)                                                
//      begin                                                                  
//         ffout = ffin; /* lintra s-60028 */
//      end 
//`endif
//endmodule
//
//`define MAKE_CLK_GATE_TRUNK(igatedclk, iipclk, iusync, iresetb, iclken, idfx_scan_dbg_mode) \
//   clk_gate_trunk \``clk_gate_trunk_``igatedclk (                                           \
//                                                 .gatedclk(igatedclk),                      \
//                                                 .ipclk(iipclk),                            \
//                                                 .usync(iusync),                            \
//                                                 .resetb(iresetb),                          \
//                                                 .clken(iclken),                            \
//                                                 .dfx_scan_dbg_mode(idfx_scan_dbg_mode)     \
//                                                );
//
//module clk_gate_trunk(output logic gatedclk,
//                      input logic ipclk,
//                      input logic usync,
//                      input logic resetb,
//                      input logic clken,
//                      input logic dfx_scan_dbg_mode);
//logic clken_qual_in, clken_qual_out;
//logic qual_or_ovrd;
//assign clken_qual_in = usync ? clken : clken_qual_out;
//`ip2211ringpll_SET_MSFF(clken_qual_out, clken_qual_in, ipclk, ~resetb)
//assign qual_or_ovrd = clken_qual_out | dfx_scan_dbg_mode;
//`CLK_GATE_HF(gatedclk, ipclk, qual_or_ovrd)
//endmodule
//                                                
//











//`define MAKE_CLK_LOCAL_QUALDIV1TO16_ADJ(qual_out,inclk,inusync,inqualovrd,inratiosel)     \
//clk_qualdiv1to16_adj_local \``clk_qualdiv1to16_adj_local_``qual_out (                           \
//                                                                  .qualclk_out(qual_out),    \
//                                                                  .clk(inclk),               \
//                                                                  .usync(inusync),           \
//                                                                  .qualovrd(inqualovrd),     \
//                                                                  .ratiosel(inratiosel)     \
//                                                                 ); /* lintra s-51500, s-53048, s-53050 */
//
//module clk_qualdiv1to16_adj_local(qualclk_out, clk, usync, qualovrd, ratiosel);
//  output qualclk_out;
//  input clk;
//  input usync;
//  input qualovrd;
//  input [3:0] ratiosel;
//  logic qual_out;
//  `MAKE_QUAL_LOCAL_QUALDIV1TO8_ADJ(qual_out, clk, usync, qualovrd, ratiosel)        
//  `ip2211ringpll_CLK_GATE(qualclk_out, clk,  qual_out)
//endmodule
//
//
//
//`define MAKE_CLK_LOCAL_QUALDIV1TO8_ADJ(qual_out,inclk,inusync,inqualovrd,inratiosel)     \
//clk_qualdiv1to8_adj_local \``clk_qualdiv1to8_adj_local_``qual_out (                           \
//                                                                  .qualclk_out(qual_out),    \
//                                                                  .clk(inclk),               \
//                                                                  .usync(inusync),           \
//                                                                  .qualovrd(inqualovrd),     \
//                                                                  .ratiosel(inratiosel)     \
//                                                                 ); /* lintra s-51500, s-53048, s-53050 */
//module clk_qualdiv1to8_adj_local(qualclk_out, clk, usync, qualovrd, ratiosel);
//  output qualclk_out;
//  input clk;
//  input usync;
//  input qualovrd;
//  input [2:0] ratiosel;
//  logic qual_out;
//  `MAKE_QUAL_LOCAL_QUALDIV1TO8_ADJ(qual_out, clk, usync, qualovrd, ratiosel)        
//  `ip2211ringpll_CLK_GATE(qualclk_out, clk,  qual_out) //lintra s-51557, s-51552
//endmodule
//
//`define MAKE_CLK_NOREN(cknorenout,cknorenckin,cknorenenin)              \
//clknoren \``clknoren_``cknorenout (                                     \
//                              .clknorenout (cknorenout),                \
//                              .clknorenckin (cknorenckin),              \
//                              .clknorenenin (cknorenenin)               \
//                             );
//
//module clknoren(clknorenout,clknorenckin,clknorenenin);
//output clknorenout;
//input clknorenckin;
//input clknorenenin;
//wire clknorenout,clknorenckin,clknorenenin;
//`ifdef INTC_DC
//     `LIB_clknoren(clknorenout,clknorenckin,clknorenenin) 
//`else
//assign clknorenout = ~(clknorenckin|clknorenenin);
//`endif
//endmodule
//



//
//`define MAKE_QUAL_LOCAL_QUALDIV16(qual_out, inclk, inusync, inqualovrd)          \
// qualdiv16_local \``qualdiv16_``qual_out (                                       \
//                                         .qualifier_out(qual_out),               \
//                                         .ipinclk(inclk) ,                       \
//                                         .usync(inusync),                        \
//                                         .qualovrd(inqualovrd)                   \
//                                         );
//module qualdiv16_local (qualifier_out,ipinclk,usync,qualovrd);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
// 
//  logic usync_lat, qual_staged, qual;
//  logic [3:0] nxt;
//  logic [3:0] pst;
// 
//  `ip2211ringpll_LATCH_P_DESKEW(usync_lat, usync, ipinclk)
//  assign nxt = pst + 4'b0001;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_lat)
//  assign qual = (&(pst));
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule
//
//`define MAKE_QUAL_LOCAL_QUALDIV1TO16_ADJ(qual_out, inclk, inusync, inqualovrd, inratiosel)     \
// qualdiv1to16_adj_local \``qualdiv1to16adj_``qual_out (                                         \
//                                                    .qualifier_out(qual_out),                 \
//                                                    .ipinclk(inclk) ,                         \
//                                                    .usync(inusync),                          \
//                                                    .qualovrd(inqualovrd),                    \
//                                                    .ratiosel(inratiosel)                     \
//                                                    );
///* lintra s-51500, s-53048, s-53050 */
//module qualdiv1to16_adj_local (qualifier_out,ipinclk,usync,qualovrd,ratiosel);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
//  input [3:0] ratiosel;
// 
//  logic usync_or_qual_lat, usync_or_qual, qual_staged, qual;
//  logic [3:0] ratiosel_muxed_staged, ratiosel_muxed;
//  logic [3:0] nxt;
//  logic [3:0] pst;
// 
//  //Whenever a qual or usync comes through we reset the counter
//  assign usync_or_qual = usync | qual;
//
//  `ip2211ringpll_LATCH_P_DESKEW(usync_or_qual_lat, usync_or_qual, ipinclk)
//  assign nxt = pst + 4'b0001;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_or_qual_lat)
//
//  //only grab ratiosel on usync boundary
//  assign ratiosel_muxed = usync ? ratiosel : ratiosel_muxed_staged;
//  `ip2211ringpll_MSFF(ratiosel_muxed_staged, ratiosel_muxed, ipinclk)
//
//  //Once we've reached the count that matches the ratiosel we're dividing by
//  //Set the qual indicator and reset the count
//  assign qual = (pst == ratiosel_muxed_staged);
//
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule // qualdiv1to16_adj_local
//
//`define MAKE_QUAL_LOCAL_QUALDIV1TO8_ADJ_WEN(qual_out, inclk, inusync, inqualovrd, inratiosel, inenable)     \
// qualdiv1to8_adj_wen_local \``qualdiv1to8adjwen_``qual_out (                                         \
//                                                    .qualifier_out(qual_out),                 \
//                                                    .ipinclk(inclk) ,                         \
//                                                    .usync(inusync),                          \
//                                                    .qualovrd(inqualovrd),                    \
//                                                    .ratiosel(inratiosel),                    \
//                                                    .enable(inenable)                         \
//                                                    );
///* lintra s-51500, s-53048, s-53050 */
//module qualdiv1to8_adj_wen_local (qualifier_out,ipinclk,usync,qualovrd,ratiosel,enable);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
//  input [2:0] ratiosel;
//  input enable;
// 
//  logic usync_or_qual_lat, usync_or_qual, qual_staged, qual;
//  logic [2:0] ratiosel_muxed_staged, ratiosel_muxed;
//  logic [2:0] nxt;
//  logic [2:0] pst;
// 
//  //Whenever a qual or usync comes through we reset the counter
//  assign usync_or_qual = usync | qual;
//
//  `ip2211ringpll_LATCH_P_DESKEW(usync_or_qual_lat, usync_or_qual, ipinclk)
//  assign nxt = pst + 1;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_or_qual_lat)
//
//  //only grab ratiosel on usync boundary
//  assign ratiosel_muxed = usync ? ratiosel : ratiosel_muxed_staged;
//  `ip2211ringpll_MSFF(ratiosel_muxed_staged, ratiosel_muxed, ipinclk)
//
//  //Once we've reached the count that matches the ratiosel we're dividing by
//  //Set the qual indicator and reset the count
//  assign qual = (pst == ratiosel_muxed_staged);
//
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = (qual_staged & enable) | qualovrd;
//endmodule // qualdiv1to8_adj_wen_local
//
//
////module qual_5_2(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [2:0]           count;
//
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 3'b000;
//     else
//       count <= (count + 3'b001) & {3{~(count == 4)}};
//
//   assign              fast_qual = (count == 0  ||
//                                    count == 3);
//   assign              slow_qual = 1'b1;
//endmodule //qual_5_2
//
//
//module qual_1_1(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//  
//   assign              fast_qual = 1'b1;
//   assign              slow_qual = 1'b1;
//endmodule // qual_1_1
//
//module qual_4_3(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [1:0]           count;
//
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//
//   assign              fast_qual = ~(count == 2);
//   assign              slow_qual = 1'b1;
//endmodule // qual_4_3
//
//module qual_8_5(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [2:0]           count;
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//   assign              fast_qual = (count == 0 ||
//                                    count == 2 ||
//                                    count == 3 ||
//                                    count == 5 ||
//                                    count == 6);
//   assign              slow_qual = 1'b1;
//endmodule // qual_8_5
//
//module qual_2_1(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg                 count;
//
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//
//   assign              fast_qual = count == 0;
//   assign              slow_qual = 1'b1;
//endmodule // qual_2_1
//
//module qual_16_7(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [3:0]           count;
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//   assign              fast_qual = (count == 0  ||
//                                    count == 2  ||
//                                    count == 5  ||
//                                    count == 7  ||
//                                    count == 9  ||
//                                    count == 11 ||
//                                    count == 14);
//   assign              slow_qual = 1'b1;
//endmodule // qual_16_7
//
//module qual_8_3(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [2:0]           count;
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//   assign              fast_qual = (count == 0 ||
//                                    count == 3 ||
//                                    count == 5);
//   assign              slow_qual = 1'b1;
//endmodule // qual_8_3
//
//module qual_16_5(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [3:0]           count;
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//   assign              fast_qual = (count == 0  ||
//                                    count == 3  ||
//                                    count == 6  ||
//                                    count == 10 ||
//                                    count == 13);
//   assign              slow_qual = 1'b1;
//endmodule // qual_16_5
//
//module qual_4_1(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [1:0]           count;
//
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//
//   assign              fast_qual = count == 0;
//   assign              slow_qual = 1'b1;
//endmodule // qual_4_1
//
//module qual_5_3(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [2:0]           count;
//
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= (count + 1) & {3{~(count == 4)}};
//
//   assign              fast_qual = (count == 1  ||
//                                    count == 2  ||
//                                    count == 4);
//   assign              slow_qual = 1'b1;
//endmodule // qual_5_3
//
//
//
//module det_clkdomainX_with_usync #(parameter dWidth = 32, parameter fifo_depth = 10, parameter separation = 2) 
////  for synchronization that's done between two clocks that are derived from the same reference clock and use separation 1,
//// this synchronizer must initiate it's rd/wr pointers at usync and not at reset!
//// otherwise separation is not ensured.
//// module det_clkdomainX must be abandoned and only this module det_clkdomainX_with_usync must be used.
//                     (
//                      input reset_ckRd,
//                      input reset_ckWr,
//                      input ckWr,
//                      input ckRd,
//                      input qualWr,
//                      input qualRd,
//                    input first_usyncWr,
//                    input first_usyncRd,
//                      input [dWidth-1:0] data_in,
//                      output [dWidth-1:0] data_out
//                      );
//
//   logic [dWidth-1:0] det_clkdomainX_write_data_array[fifo_depth - 1:0];
//   logic [dWidth-1:0] det_clkdomainX_read_data_mux;
//   logic [fifo_depth - 1:0] wrptr;
//   logic [fifo_depth - 1:0] rdptr;
//   logic [fifo_depth - 1:0] start_ptr;
//   logic write_clk;
//   logic read_clk;
//
//   `ip2211ringpll_CLK_GATE(write_clk, ckWr, qualWr)
//   `ip2211ringpll_CLK_GATE(read_clk, ckRd, qualRd)
//  
//   // data path generation
//   always@(posedge write_clk or negedge reset_ckWr)
//     begin: write_clk_scope
//        integer i;
//        if (~reset_ckWr)
//          begin
//             for (i=0;i<fifo_depth;i=i+1)
//               begin
//                  det_clkdomainX_write_data_array[i] <= 0;
//               end
//          end
//        else
//          begin
//             for (i=0;i<fifo_depth;i=i+1)
//               begin
//                  if (wrptr[i])
//                    det_clkdomainX_write_data_array[i] <= data_in;
//               end
//          end
//     end
//
//   always@(posedge read_clk or negedge reset_ckRd)
//     begin: read_clk_scope
//        integer i;
//        if (~reset_ckRd)
//          begin
//             det_clkdomainX_read_data_mux <= 0;
//          end
//        else
//          begin
//             for (i=0;i<fifo_depth;i=i+1)
//               begin
//                  if (rdptr[i])
//                    det_clkdomainX_read_data_mux <= det_clkdomainX_write_data_array[i];
//               end
//          end
//     end
//
//   assign data_out = det_clkdomainX_read_data_mux;
//
//   // wrptr and rdptr generation
//   assign start_ptr = 1;
//   
//   always@(posedge write_clk or negedge reset_ckWr)
//     if(!reset_ckWr)
//       wrptr <= start_ptr << separation;
//     else if (first_usyncWr)
//       wrptr <= start_ptr << separation;
//     else
//       wrptr <= {wrptr[(fifo_depth - 2):0], wrptr[(fifo_depth - 1)]};
//
//   always@(posedge read_clk or negedge reset_ckRd)
//     if(!reset_ckRd)
//       rdptr <= start_ptr;
//     else if (first_usyncRd)
//       rdptr <= start_ptr;
//     else
//       rdptr <= {rdptr[(fifo_depth - 2):0], rdptr[(fifo_depth - 1)]};
//
//endmodule // det_clkdomainX_with_usync
//

`ifndef ip2211ringpll_SOC_POWER_MACROS_VH
`define ip2211ringpll_SOC_POWER_MACROS_VH

////`include "vlv_macro_tech_map.vh"

`ifdef INTC_EXPERIMENTAL_POWER_INTENT 
 //`include "sppowerintent.vh"
`endif

///============================================================================================
///
/// Firewall
///
///============================================================================================


//SAME as ip2211ringpll_FIREWALL_AND from soc_macros.sv but created seperate version
//for different checking on clocks. Still same library cell though.
`define ip2211ringpll_FIREWALL_AND_CLK(out,data,enable)                                           \
`ifdef INTC_EXPERIMENTAL_POWER_INTENT                                                          \
fw_and_bus #(.BW($bits(out))) \``fw_and_\``out   (.fwout(out),.fwdata(data),.fwenable(enable)); \
`else										    \
 `ifdef INTC_DC                                                                           \
  `LIB_FIREWALL_AND(out,data,enable)                                               \
 `else \
	 assign out = data & {$bits(out){enable}}; /* lintra s-35000, s-35006 */          \
 `endif \
`endif
	   	 

	   
	 
//SAME as ip2211ringpll_LS_WITH_AND_FW from soc_macros.sv but created seperate version
//for different checking on clocks. Still same library cell though.
`define ip2211ringpll_LS_WITH_AND_FW_CLK(o, pro, a, vcc_in, en)                                                 \
`ifdef INTC_EXPERIMENTAL_POWER_INTENT                                                          \
	   fw_ls_and_bus_ck #(.BW($bits(o))) \``fw_ls_and_\``o   (.lspro(pro),.fwout(o),.lsvcc_in(vcc_in),.fwdata(a),.fwenable(en)); \
`elsif INTC_DC                                                                                         \
  `LIB_LS_WITH_AND_FW_CLK(o, pro, a, vcc_in, en)                                                   \
`else \
       	assign o = a & {$bits(o){en}}; \
`endif \


//Needed for sVID GPIO clk pin (added on request by Chad Coburn)
`define ip2211ringpll_LS_WITH_OR_FW_CLK(o, pro, a, vcc_in, en)                                 \
`ifdef INTC_DC                                                                        \
     `LIB_LS_WITH_OR_FW(o, pro, a, vcc_in, en)                                   \
`else                                                                            \
     `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                      \
                                                                                 \
     `endif                                                                      \
     assign o = a | ~{$bits(o){en}};        /* lintra s-35019 */                 \
`endif

	  
   `define ip2211ringpll_FIREWALL_AND(out,data,enable)                                               \
   `ifdef INTC_EXPERIMENTAL_POWER_INTENT                                                          \
       fw_and_bus #(.BW($bits(out))) \``fw_and_\``out   (.fwout(out),.fwdata(data),.fwenable(enable)); \
   `else										    \
    `ifdef INTC_DC                                                                           \
	 `LIB_FIREWALL_AND(out,data,enable)                                               \
    `else \
	  assign out = data & {$bits(out){enable}}; /* lintra s-35000, s-35006 */          \
    `endif \
   `endif
	    									
	    
			
   `define ip2211ringpll_FIREWALL_OR(out,data,enable)                                                \
   `ifdef INTC_EXPERIMENTAL_POWER_INTENT  \
	    fw_or_bus  #(.BW($bits(out))) \``fw_or_\``out    (.fwout(out),.fwdata(data),.fwenable(enable)); \
    `else \
     `ifdef INTC_DC                                                                           \
	      `LIB_FIREWALL_OR(out,data,enable)                                                \
     `else \
	     assign out = data | ~{$bits(out){enable}}; /* lintra s-35000, s-35006 */ \
     `endif \
    `endif
	       
///============================================================================================
///
/// Voltage Level Shifters
///
///============================================================================================



//Signal Description
//outb       Level shifter output, 
//ipro       Output supply domain name (example: vccxxxvidsi0gt_1p05), 
// ib        Input signal to be level shifted,
//iwrite_en  Level shifter firewall enable. Should come from the output supply domain.
//Note: Input supply domain is implicit vcc!

`define ip2211ringpll_LS_LATCH_DN(outb,ipro,ib,iwrite_en)                                               \
`ifdef INTC_DC                                                                                 \
     `LIB_LS_LATCH_DN(outb,iwrite_en,ipro,ib)                                             \
`else                                                                                     \
   `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                 \
                                                                                          \
   `endif                                                                                 \
   always_latch                                                                           \
      begin                                                                               \
         if (iwrite_en) outb <= ~ib;   /* lintra s-30529, s-30518, s-31501, s-35006 */    \
      end                                                                                 \
/* lintra s-30500, s-30543 */                                                             \
`endif


  


  
//Signal Description
//outb       Level shifter output, 
//ipro       Output supply domain name (example: vccxxxvidsi0gt_1p05), 
//ib         Input signal to be level shifted,
//vccin      Input supply domain name (example: vccxxxvidsi0_1p05),
//iwrite_en  Level shifter firewall enable. Should come from the output supply domain.

`define ip2211ringpll_LS_LATCH_PWR_PN(outb, ipro, ib, vccin, iwrite_en )                                  \
  `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                    \
                                                                                            \
  `endif                                                                                    \
  always_latch                                                                              \
      begin                                                                                 \
         if (iwrite_en) outb <= ~ib; /* lintra s-30529, s-30518, s-35006 */                 \
      end   

  
  
//Signal Description
//outb       Level shifter output,
//ib         Input signal to be level shifted,
//ipro       Input supply domain name (example: vccxxxvidsi0gt_1p05), 
//iwrite_en  Level shifter firewall enable. Should come from the output supply domain.
//Note: Output supply domain is implicit vcc!

`define ip2211ringpll_LS_LATCH_UP(outb,ib,ipro,iwrite_en)                                               \
`ifdef INTC_DC                                                                                 \
     `LIB_LS_LATCH_UP(outb,iwrite_en,ipro,ib)                                             \
`else                                                                                     \
   `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                 \
                                                                                          \
   `endif                                                                                 \
   always_latch                                                                           \
      begin                                                                               \
         if (iwrite_en) outb <= ~ib;   /* lintra s-30529, s-30518, s-31501, s-35006 */    \
      end                                                                                 \
/* lintra s-30500, s-30543 */                                                             \
`endif

  
/* lintra s-30500, s-30543 */

//Signal Desctiption
//o       Level shifter output,
//pro     Output supply domain name (example: vccxxxvidsi0gt_1p05),
//a       Input signal to be level shifted,
//vcc_in  Input supply domain name (example: vccxxxvidsi0_1p05),
//en      Level shifter firewall enable. Should come from the output supply domain.
//To code level shifters with no firewall enable, please use ip2211ringpll_LS_WITH_AND_FW macro with en tied to the output supply domain.

`define ip2211ringpll_LS_WITH_AND_FW(o, pro, a, vcc_in, en)                                                     \
   `ifdef INTC_EXPERIMENTAL_POWER_INTENT                                                          \
 fw_ls_and_bus #(.BW($bits(o))) \``fw_ls_and_\``o   (.lspro(pro),.fwout(o),.lsvcc_in(vcc_in),.fwdata(a),.fwenable(en)); \
   `elsif INTC_DC                                                                                         \
     `LIB_LS_WITH_AND_FW(o, pro, a, vcc_in, en)                                                   \
   `else  \
	    assign o = a & {$bits(o){en}};   /* lintra s-35019 */                                        \
   `endif \
	      
	      
	      

     
       

//Signal Description
//o       Level shifter output,
//pro     Output supply domain name (example: vccxxxvidsi0gt_1p05),
//a       Input signal to be level shifted,
//vcc_in  Input supply domain name (example: vccxxxvidsi0_1p05),
//en      Level shifter firewall enable. Should come from the output supply domain.
   `define ip2211ringpll_LS_WITH_OR_FW(o, pro, a, vcc_in, en) \
   `ifdef INTC_EXPERIMENTAL_POWER_INTENT                                                          \
	      fw_ls_or_bus #(.BW($bits(o))) \``fw_ls_or_\``o   (.lspro(pro),.fwout(o),.lsvcc_in(vcc_in),.fwdata(a),.fwenable(en)); \
  `else \
  `ifdef INTC_DC                                                                                         \
    `LIB_LS_WITH_OR_FW(o, pro, a, vcc_in, en)                                                    \
   `else \
	 assign o = a | ~{$bits(o){en}};   /* lintra s-35019 */                                       \
   `endif \
  `endif   
    
	   
  
// New always ON inverter macro for Mihir
// Usage is only for the other power plane (Non-Vnn power plane)
`define ip2211ringpll_POWER_INVERTER_D(powerenout, powerenin, vcc_in)                                          \
`ifdef INTC_DC                                                                                        \
     `LIB_POWER_INVERTER_D(powerenout, powerenin, vcc_in)                                        \
`else                                                                                            \
  `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                         \
                                                                                                 \
  `endif                                                                                         \
  assign powerenout = ~powerenin ;     /* lintra s-35000, s-35006 */                             \
`endif 

    
///============================================================================================
///
/// Power Switch
///
///============================================================================================



//`define ip2211ringpll_POWERSWITCH(pwren_out, vcc_out, pwren_in, vcc_in, vss_in)  \
//   assign vcc_out   = ~pwren_in ? vcc_in : 1'bz ;                  \
//   assign pwren_out = ~(~(pwren_in)); /* lintra s-35022 */         \

//// new FW macro proposed by Bradley Erwin
`define ip2211ringpll_POWERSWITCH(pwren_out, vcc_out, pwren_in, vcc_in, vss_in)                                         \
`ifdef INTC_DC                                                                                                 \
    `LIB_POWERSWITCH(pwren_out, vcc_out, pwren_in, vcc_in, vss_in)                                       \
`else                                                                                                    \
 `ifdef INTC_EXPERIMENTAL_POWER_INTENT                                                          \
          `LIB_POWERSWITCH(pwren_out, vcc_out, pwren_in, vcc_in, vss_in)                                       \
 `else \
	 assign vcc_out = ~pwren_in ? vcc_in : 1'bz; /* lintra s-30505 */                                       \
	   assign pwren_out = ~(~(pwren_in)); /* lintra s-35022 */                                                \
 `endif \
`endif
	     
	   
	     
     
    

//Signal Description
//o                    Level shifter output,
//vccout            Output supply domain name (example: vccxxxvidsi0gt_1p05),
//a                    Input signal to be level shifted,
//vccin              Input supply domain name (example: vccxxxvidsi0_1p05),
//THIS MACRO SHOULD ONLY BE USED GOING FROM ALWAYS ON SUPPLIES TO COLLAPSIBLE SUPPLIES
 
`define ip2211ringpll_LS_WITH_NO_FW(o, vccout, a, vccin)                                                                \
`ifdef INTC_DC                                                                                                 \
`else                                                                                                     \
     `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                               \
         (* macro_attribute = `"LS_WITH_NO_FW(o``,vccout``,a``,vccin``)`" *)                              \
     `endif                                                                                               \
     assign o = a;   /* lintra s-35000, s-35019 */                                                        \
`endif                                                                                                    
       
//Adding this macro after approval from Raboul. 
//Email notes from Quddus, Wasim: We need a MACRO to instantiate LS going from rtc_well to sus_well.
//I talked with Rabiul, he suggested to use a different name, i.e. ip2211ringpll_LS_WITH_NO_FW_TG.
//We want the b12sirblnx20tg cell to implement the LS from TG library.

//
`define ip2211ringpll_LS_WITH_NO_FW_TG(o, vccout, a, vccin)                                                             \
`ifdef INTC_DC                                                                                                 \
       `LIB_LS_WITH_NO_FW_TG(o, pro, a, vcc_in)                                                                \
`else                                                                                                     \
 `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                               \
         (* macro_attribute = `"LS_WITH_NO_FW_TG(o``,vccout``,a``,vccin``)`" *)                           \
     `endif                                                                                               \
	   assign o = a;   /* lintra s-35000, s-35019 */                                                        \
    `endif
	     
	     
      

//New dual power switch macro ---- Added by Nasim Uddin
//dual power switch macro had not been tested out yet
`define ip2211ringpll_POWERSWITCH_DUAL(pwren1_out, pwren2_out, vcc_out, pwren1_in, pwren2_in, vcc_in, vss_in)           \
`ifdef INTC_DC                                                                                                 \
     `LIB_POWERSWITCH_DUAL(pwren1_out,  pwren2_out, vcc_out, pwren1_in, pwren2_in, vcc_in, vss_in)        \
`else                                                                                                     \
   `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                                 \
                                                                                                          \
   `endif                                                                                                 \
   assign vcc_out = ~pwren1_in | ~pwren2_in ? vcc_in : 1'bz; /* lintra s-30505 */                         \
   assign pwren1_out = ~(~(pwren1_in)); /* lintra s-35022 */                                              \
   assign pwren2_out = ~(~(pwren2_in)); /* lintra s-35022 */                                              \
  `endif                                                             \
 

 `endif //  `ifndef ip2211ringpll_SOC_POWER_MACROS_VH
     
     

/*******************************************************************************************************************
*
 *  MACROS NOT BEING USED BY ANYONE ELSE -  for
   *  ISSUES 
*  
*******************************************************************************************************************/



//`define MAKE_CLK_DELAY4(clkd4out,clkd4clkin,clkd4in0,clkd4in1,clkd4in2)    \
//clk4delay \``clk4delay_``clkd4out (                                          \
//                                    .clk4delayout (clkd4out),              \
//                                    .clk4delayin (clkd4clkin),             \
//                                    .clk4in0 (clkd4in0),                   \
//                                    .clk4in1 (clkd4in1),                   \
//                                    .clk4in2 (clkd4in2)                    \
//                                );
//
//`define LIB_clk4delay(clk4delayout,clk4delayin,clk4in0,clk4in1,clk4in2) \
//  vl0dcc04ln0a0 ck2(.o(clk4delayout),.clk(clk4delayin),.rsel0(clk4in0),.rsel1(clk4in1),.rsel2(clk4in2)); \
//
//module clk4delay (clk4delayout,clk4delayin,clk4in0,clk4in1,clk4in2);
//output clk4delayout;
//input clk4delayin;
//input clk4in0;
//input clk4in1;
//input clk4in2;
//wire clk4delayout,clk4delayin,clk4in0,clk4in1,clk4in2;
//`ifdef INTC_DC
//     `LIB_clk4delay(clk4delayout,clk4delayin,clk4in0,clk4in1,clk4in2) 
// `else
//assign clk4delayout = clk4delayin;
//`endif
//endmodule
//
//
//`define MAKE_CLK_DELAY8(clkd8out,clkd8clkin,clkd8in0,clkd8in1,clkd8in2,clkd8in3,clkd8in4,clkd8in5,clkd8in6)    \
//clk8delay \``clk8delay_``clkd8out (                                                         \
//                                    .clk8delayout (clkd8out),                             \
//                                    .clk8delayin (clkd8clkin),                            \
//                                    .clk8in0 (clkd8in0),                                  \
//                                    .clk8in1 (clkd8in1),                                  \
//                                    .clk8in2 (clkd8in2),                                  \
//                                    .clk8in3 (clkd8in3),                                  \
//                                    .clk8in4 (clkd8in4),                                  \
//                                    .clk8in5 (clkd8in5),                                  \
//                                    .clk8in6 (clkd8in6)                                   \
//                                );
//
//
//`define LIB_clk8delay(clk8delayout,clk8delayin,clk8in0,clk8in1,clk8in2,clk8in3,clk8in4,clk8in5,clk8in6) \
//  vl0dcc08ln0a0 ck2(.o(clk8delayout),.clk(clk8delayin),.rsel0(clk8in0),.rsel1(clk8in1),.rsel2(clk8in2),.rsel3(clk8in3),.rsel4(clk8in4),.rsel5(clk8in5),.rsel6(clk8in6)); \
//
//module clk8delay (clk8delayout,clk8delayin,clk8in0,clk8in1,clk8in2,clk8in3,clk8in4,clk8in5,clk8in6);
//output clk8delayout;
//input clk8delayin;
//input clk8in0;
//input clk8in1;
//input clk8in2;
//input clk8in3;
//input clk8in4;
//input clk8in5;
//input clk8in6;
//wire clk8delayout,clk8delayin,clk8in0,clk8in1,clk8in2,clk8in3,clk8in4,clk8in5,clk8in6;
//`ifdef INTC_DC
//     `LIB_clk8delay(clk8delayout,clk8delayin,clk8in0,clk8in1,clk8in2,clk8in3,clk8in4,clk8in5,clk8in6) 
// `else
//assign clk8delayout = clk8delayin;
//`endif
//endmodule
//
//
//`define MAKE_CLK_DIV2SHIFT(ckdiv2shftout,ipinckdiv2shftin,usyncdiv2shft)      \
// clk2div2shft \``clk_div2shift_``ckdiv2shftout (                                             \
//                                              .div2shftckdiv2shftout (ckdiv2shftout),      \
//                                              .div2shftipinckdiv2shftin (ipinckdiv2shftin),\
//                                              .div2shftusyncdiv2shft (usyncdiv2shft)       \
//                                             );
//
//module clk2div2shft (div2shftckdiv2shftout,div2shftipinckdiv2shftin,div2shftusyncdiv2shft);
//output div2shftckdiv2shftout;
//input div2shftipinckdiv2shftin;
//input div2shftusyncdiv2shft;
//reg div2shftckdiv2shftout;
//wire div2shftipinckdiv2shftin,div2shftusyncdiv2shft;
// reg ckdiv2shftout_ffout;                                                          
//  wire ckdiv2shftout_invout,ckdiv2shftout_andout,ckdiv2shftout_ckinvout;        
//  always_ff @(posedge div2shftipinckdiv2shftin)                                               
//      begin                                                                           
//       ckdiv2shftout_ffout   <= div2shftusyncdiv2shft;                                      
//      end  
//  assign ckdiv2shftout_invout = ~ckdiv2shftout_ffout;       
//  ip2211ringpll_clkinv clkinvdiv2shft (
//                         .clkout (ckdiv2shftout_ckinvout),
//                         .clkin (div2shftipinckdiv2shftin)
//                        );
//  assign  ckdiv2shftout_andout = (ckdiv2shftout_invout) & (~div2shftckdiv2shftout);     
//  clockdivff clockdivff_ckdiv2shftout (                                            
//                                   .ffout(div2shftckdiv2shftout),                             
//                                   .ffin(ckdiv2shftout_andout),                     
//                                   .clockin(ckdiv2shftout_ckinvout)                 
//                                  );
//endmodule
//
//                                             
//
//
//
//
//
//`define MAKE_CLK_LOCAL_QUALDIV100(div100clkout, div100_base_clk, div100_reset_n, div100_byp_div, div100_clk_disable, div100_squash_div)        \
//   crp_sample_gen_common #(100) \``make_clk_qualdiv100_``div100clksample (                                           \
//                                                    .base_clk              (div100_base_clk),                \
//                                                    .byp_div               (div100_byp_div),                 \
//                                                    .reset_n               (div100_reset_n),                 \
//                                                    .clk_disable           (div100_clk_disable),             \
//                                                    .squash_div            (div100_squash_div),              \
//                                                    .clk_out               (div100clkout)                    \
//                                                    );
//
//`define MAKE_CLK_LOCAL_QUALDIV16(outclk,inclk,ipinck,inusync)             \
//clkqualdiv16_local \``clk_qualdiv4_local``outclk (                               \
//                                   .divckout (outclk),                      \
//                                   .divckin  (inclk),                       \
//                                   .divipinckin(ipinck),                      \
//                                   .divusync (inusync)                            \
//                                  );
//
///* lintra s-31500, s-33048, s-33050 */
//module clkqualdiv16_local (divckout,divckin,divipinckin,divusync);
//   output divckout;
//   input  divckin;
//   input  divipinckin;
//   input  divusync;
//   reg    divckout;
//   wire   divckin,divusync;
//   reg    ckdiv16out_pout;                                                
//   reg [3:0] ckdiv16out_rstffpst;                                      
//   wire [3:0] ckdiv16out_rstffnxt;
//   logic       temp1, usync;
//   always_latch                                                         
//     begin                                                          
//        if (~divipinckin) ckdiv16out_pout  <= divusync;        
//     end                                                            
//   always_ff @(posedge divipinckin)                                 
//     begin                                                          
//        if (ckdiv16out_pout) ckdiv16out_rstffpst  <= '0;
//        else ckdiv16out_rstffpst  <=  ckdiv16out_rstffnxt;     
//     end                                                            
//   assign ckdiv16out_rstffnxt = ckdiv16out_rstffpst  + 1 ;           
//   assign usync = &ckdiv16out_rstffpst;
//   
//   clockdivff clockdivff_ckdiv16out(                                 
//                                   .ffout(temp1),                      
//                                   .ffin(usync),              
//                                   .clockin(divckin)                      
//                                   );
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp1)
//
//endmodule
//
//`define MAKE_CLK_LOCAL_QUALDIV2(ckout,ckin,ipinckin,usync)         \
// clkqualdiv_local \``clk_qualdiv2_``ckout (                         \
//                                         .divckout(ckout),       \
//                                         .divckin(ckin) ,        \
//                                         .divipinckin(ipinckin), \
//                                         .divusync(usync)          \
//                                         );
//
//
//
///* lintra s-31500, s-33048, s-33050 */
//`define MAKE_CLK_LOCAL_QUALDIV4(ckout2,ckin2,ipinckin2,usync2)            \
//clkqualdiv4_local \``clk_qualdiv4_local``ckout2 (                                \
//                                   .divckout (ckout2),             \
//                                   .divckin  (ckin2),              \
//                                   .divipinckin(ipinckin2),        \
//                                   .divusync (usync2)                \
//                                  );
//
//`define MAKE_CLK_LOCAL_QUALDIV600(div600clkout, div600_base_clk, div600_reset_n, div600_byp_div, div600_clk_disable, div600_squash_div)        \
//   crp_sample_gen_common #(600) \``make_clk_qualdiv600_``div600clksample (                                           \
//                                                    .base_clk              (div600_base_clk),                \
//                                                    .reset_n               (div600_reset_n),                 \
//                                                    .byp_div               (div600_byp_div),                 \
//                                                    .clk_disable           (div600_clk_disable),             \
//                                                    .squash_div            (div600_squash_div),              \
//                                                    .clk_out               (div600clkout)                    \
//                                                    );
//
//module crp_sample_gen_common  #(parameter dWidth = 3) 
//                     (
//                      input                  base_clk,       // Pre or Post CTS based on Physical Design
//                      input                  reset_n,        // Must be pre-stinkronized to base_clk input
//                      input                  byp_div,        // PMU Register input
//                      input                  clk_disable,    // PMU Register input
//                      input [(dWidth - 1):0] squash_div,     // PMU Register input
//                      output                 clk_out
//                      );
//
//   reg [(dWidth - 1):0]    count;
//   reg                     clk_sample_fe;
//   wire                    clk_sample;
//
//   // Standard up-down counter with some extras
//   always @(posedge base_clk or negedge reset_n )
//     if (~reset_n)
//       count         <= 'b0;     // Divider initial 1 or 0
//     else if (clk_disable || (squash_div == 0))
//       count         <= 'b0;
//     else if (count < squash_div)
//       count         <= count + 1;
//     else
//       count         <= 'b0;
//
//   // Falling edge used to clock forward the sample signal
//   always @(negedge base_clk or negedge reset_n )
//     if (~reset_n)
//       clk_sample_fe <= 'b0;     
//     else if (clk_disable)    // I1 control
//       clk_sample_fe <= 'b0;
//     else if ( count == 0 )
//       clk_sample_fe <= 'b1;
//     else
//       clk_sample_fe <= 'b0;
//
//   assign  clk_sample = byp_div ? 1'b1 : clk_sample_fe;
//
//   ip2211ringpll_soc_rbe_clk \``soc_rbe_clk_``clk_out (clk_out,base_clk,clk_sample);
//endmodule // clk_sample_gen
//
//
//`define MAKE_CLK_LOCAL_QUALDIV8(ckout2,ckin2,ipinckin2,usync2)            \
//clkqualdiv8_local \``clk_qualdiv4_local``ckout2 (                                \
//                                   .divckout (ckout2),             \
//                                  .divckin  (ckin2),              \
//                                   .divipinckin(ipinckin2),        \
//                                   .divusync (usync2)                \
//                                  );
///* lintra s-31500, s-33048, s-33050 */
//module clkqualdiv8_local (divckout,divckin,divipinckin,divusync);
//   output divckout;
//   input  divckin;
//   input  divipinckin;
//   input  divusync;
//   reg    divckout;
//   wire   divckin,divusync;
//   reg    ckdiv8out_pout;                                                
//   reg [2:0] ckdiv8out_rstffpst;                                      
//   wire [2:0] ckdiv8out_rstffnxt;
//   logic       temp1, temp2, usync;
//   always_latch                                                         
//     begin                                                          
//        if (~divipinckin) ckdiv8out_pout  <= divusync;        
//     end                                                            
//   always_ff @(posedge divipinckin)                                 
//     begin                                                          
//        if (ckdiv8out_pout) ckdiv8out_rstffpst  <= '0;          
//        else ckdiv8out_rstffpst  <=  ckdiv8out_rstffnxt;     
//     end                                                            
//   assign ckdiv8out_rstffnxt = ckdiv8out_rstffpst  + 1 ;           
//   assign usync = &ckdiv8out_rstffpst;
//   
//   clockdivff clockdivff_ckdiv8out(                                 
//                                   .ffout(temp1),                      
//                                   .ffin(usync),              
//                                   .clockin(divckin)                      
//                                   );
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp1)
//endmodule
//                                  
//
//`define MAKE_CLK_LOCAL_QUALDIV8_ADJ(ckout2,ckin2,ipinckin2,usync2, ratiosel2)            \
//clkqualdiv8_local_adj \``clk_qualdiv4_local_adj``ckout2 (                                \
//                                   .divckout (ckout2),             \
//                                   .divckin  (ckin2),              \
//                                   .divipinckin(ipinckin2),        \
//                                   .divusync (usync2),               \
//                                   .ratiosel (ratiosel2)                \
//                                  );
///* lintra s-31500, s-33048, s-33050 */
//module clkqualdiv8_local_adj (divckout,divckin,divipinckin,divusync,ratiosel);
//   output divckout;
//   input  divckin;
//   input  divipinckin;
//   input  divusync;
//   input [2:0] ratiosel;
//   reg    divckout;
///   wire   divckin,divusync;
//   reg    ckdiv8out_pout;                                                
//   reg [2:0] ckdiv8out_rstffpst;                                      
//   wire [2:0] ckdiv8out_rstffnxt;
//   logic       temp1, usync;
//
//   `ip2211ringpll_LATCH_P_DESKEW(ckdiv8out_pout, divusync, divipinckin)           
//   assign ckdiv8out_rstffnxt = ckdiv8out_rstffpst  + 1 ;
//   `ip2211ringpll_RST_MSFF(ckdiv8out_rstffpst, ckdiv8out_rstffnxt, divipinckin, ckdiv8out_pout)                   
//
//   always_comb
//     case(ratiosel)
//       3'b000 : usync = &ckdiv8out_rstffpst[2:0]; // div 8
//       3'b001 : usync = &ckdiv8out_rstffpst[1:0]; // div 4
//       3'b011 : usync = ckdiv8out_rstffpst[0];    // div 2
//       3'b111 : usync = 1'b1;                     // div 1
//       default: usync = 1'b1;
//     endcase // case(ratiosel)
//       
//   clockdivff clockdivff_ckdiv8out(                                 
//                                   .ffout(temp1),                      
//                                   .ffin(usync),              
//                                   .clockin(divckin)                      
//                                   );
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp1)
//endmodule
//
//// original MAKE_CLK_QUALDIV2 need to comment out after iosf is inplace
//`define MAKE_CLK_QUALDIV2(ckout,ckin,ipinckin,qual)         \
// clkqualdiv \``clk_qualdiv2_``ckout (                         \
//                                    .divckout(ckout),       \
//                                    .divckin(ckin) ,        \
//                                    .divipinckin(ipinckin), \
//                                    .divqual(qual)          \
//                                   );
//module clkqualdiv_local (divckout,divckin,divipinckin,divusync);
//output divckout;
//input divckin;
//input divipinckin;
//input divusync;
//   logic temp, temp1, temp2, temp3;
//    wire ckout_tmp1, ckout_tmp2, ckout_tmp, ckout_invclk;                                 
//   `ip2211ringpll_LATCH_P(temp, divusync, divipinckin)
//   `ip2211ringpll_MSFF(temp1, temp2, divipinckin)
//   assign temp2 = ~temp1 & ~temp;
//   `ip2211ringpll_MSFF(temp3, temp1, divckin)
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp3)
// 
//     /* lintra s-31500 */
//endmodule
//
//// original MAKE_CLK_QUALDIV4 - need to comment out after iosf in place
//`define MAKE_CLK_QUALDIV4(ckout2,ckin2,ipinckin2,qual2)            \
//clkqualdiv \``clk_qualdiv4_``ckout2 (                                \
//                                   .divckout (ckout2),             \
//                                   .divckin  (ckin2),              \
//                                   .divipinckin(ipinckin2),        \
//                                   .divqual (qual2)                \
//                                  );
//
//
//`define MAKE_QUAL_LOCAL_QUALDIV2(qual_out, inclk, inusync, inqualovrd)     \
// qualdiv2_local \``qualdiv2_``qual_out (                                         \
//                                         .qualifier_out(qual_out),       \
//                                         .ipinclk(inclk) ,                  \
//                                         .usync(inusync),                       \
//                                         .qualovrd(inqualovrd)                  \
//                                         );
//
///* lintra s-31500, s-33048, s-33050 */
//module qualdiv2_local (qualifier_out,ipinclk,usync,qualovrd);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
// 
//  logic usync_lat, qual_staged;
//  logic nxt, pst;
// 
//  `ip2211ringpll_LATCH_P(usync_lat, usync, ipinclk)
//  assign nxt = pst + 1;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_lat)
//  `ip2211ringpll_MSFF(qual_staged, pst, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule
// 
//`define MAKE_QUAL_LOCAL_QUALDIV4(qual_out, inclk, inusync, inqualovrd)     \
// qualdiv4_local \``qualdiv4_``qual_out (                                         \
//                                         .qualifier_out(qual_out),       \
//                                         .ipinclk(inclk) ,                  \
//                                         .usync(inusync),                       \
//                                         .qualovrd(inqualovrd)                  \
//                                         );
///* lintra s-31500, s-33048, s-33050 */
//module clkqualdiv4_local (divckout,divckin,divipinckin,divusync);
//   output divckout;
//   input  divckin;
//   input  divipinckin;
//   input  divusync;
//   reg    divckout;
//   wire   divckin,divusync;
//   reg    ckdiv4out_pout;                                                
//   reg [1:0] ckdiv4out_rstffpst;                                      
//   wire [1:0] ckdiv4out_rstffnxt;
//   logic       temp1, usync;
//   always_latch                                                         
//     begin                                                          
//        if (~divipinckin) ckdiv4out_pout  <= divusync;        
//     end                                                            
//   always_ff @(posedge divipinckin)                                 
//     begin                                                          
//        if (ckdiv4out_pout) ckdiv4out_rstffpst  <= '0;          
//        else ckdiv4out_rstffpst  <=  ckdiv4out_rstffnxt;     
//     end                                                            
//   assign ckdiv4out_rstffnxt = ckdiv4out_rstffpst  + 1 ;           
//   assign usync = &ckdiv4out_rstffpst;
//   
//   clockdivff clockdivff_ckdiv4out(                                 
//                                   .ffout(temp1),                      
//                                   .ffin(usync),              
//                                   .clockin(divckin)                      
//                                   );
//   `ip2211ringpll_CLK_GATE(divckout, divckin, temp1)
//endmodule
//
//// origianl clkqualdiv - need to remove after iosf is in place
//module clkqualdiv (divckout,divckin,divipinckin,divqual);
//output divckout;
//input divckin;
//input divipinckin;
//input divqual;
//wire divckout,divckin,divipinckin,divqual;
//`ifdef INTC_DC                                                                                         
//    wire ckout_tmp1, ckout_tmp2, ckout_tmp, ckout_invclk;                                 
//    `LIB_clkqualdiv(divckout,divckin,divipinckin,divqual) 
//`else                                                                                             
//reg ckout_qualout, ckout_qual1out;                                                            
// always @(negedge divipinckin)                                                                       
//   begin                                                                                          
//      ckout_qual1out = divqual; /* lintra s-60028 */
//   end                                                                                            
// always @(negedge divipinckin)                                                                       
//  begin                                                                                           
//      ckout_qualout  = ckout_qual1out; /* lintra s-60028 */
//   end                                                                                            
//   assign divckout = ckout_qualout & divckin;                                                     
//`endif     /* lintra s-31500 */
//endmodule
//
//
//                                        
//`define MAKE_QUAL_LOCAL_QUALDIV8(qual_out, inclk, inusync, inqualovrd)     \
// qualdiv8_local \``qualdiv8_``qual_out (                                         \
//                                        .qualifier_out(qual_out),       \
//                                         .ipinclk(inclk) ,                  \
//                                         .usync(inusync),                       \
//                                        .qualovrd(inqualovrd)                  \
//                                         );
//
///* lintra s-31500, s-33048, s-33050 */
//module qualdiv8_local (qualifier_out,ipinclk,usync,qualovrd);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
// 
//  logic usync_lat, qual_staged, qual;
//  logic [2:0] nxt;
//  logic [2:0] pst;
// 
//  `ip2211ringpll_LATCH_P(usync_lat, usync, ipinclk)
//  assign nxt = pst + 1;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_lat)
//  assign qual = (&(pst));
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule
//
//*****ANY USES OF MAKE_QUAL_LOCAL_QUALDIV8_ADJ SHOULD EVENTUALLY BE REPLACED BY 
//*****MAKE_QUAL_LOCAL_QUALDIV1TO8_ADJ WE CAN'T JUST CHANGE THIS MACRO AS IT WOULD CAUSE FAILS
// ML_FIX : Eventually need to remove this define and module
//`define MAKE_QUAL_LOCAL_QUALDIV8_ADJ(qual_out, inclk, inusync, inqualovrd, inratiosel)     \
// qualdiv8_adj_local \``qualdiv8adj_``qual_out (                                                   \
//                                         .qualifier_out(qual_out),                     \
//                                         .ipinclk(inclk) ,                                \
//                                         .usync(inusync),                                     \
//                                         .qualovrd(inqualovrd),                                \
//                                         .ratiosel(inratiosel)                                \
//                                         );
//
///* lintra s-31500, s-33048, s-33050 */
//module qualdiv8_adj_local (qualifier_out,ipinclk,usync,qualovrd,ratiosel);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
//  input [2:0] ratiosel;
// 
//  logic usync_lat, qual_staged, qual;
//  logic [2:0] nxt;
//  logic [2:0] pst;
// 
//  `ip2211ringpll_LATCH_P_DESKEW(usync_lat, usync, ipinclk)
//  assign nxt = pst + 1;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_lat)
//  always_comb begin
//    casex(ratiosel)
//      3'b000 : qual = &pst[2:0]; // div 8
//      3'b001 : qual = &pst[1:0]; // div 4
//      3'b011 : qual = pst[0];    // div 2
//      3'b111 : qual = 1'b1;      // div 1
//      default: qual = 1'b1;
//    endcase // case(ratiosel)
//  endip2211ringpll_soc_rbe_clk
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule // qualdiv8_adj_local
//
//`define CLK_FF_INV(ckdiv2routb,ckdiv2rin,ckdiv2clkin,ckdiv2resetin)                       \
//clockdivffreset_inv \``clockdivffreset_inv_``ckdiv2routb (                                \
//                                                         .ffoutresetb(ckdiv2routb),       \
//                                                         .ffinreset(ckdiv2rin),           \
//                                                         .clockinreset(ckdiv2clkin),      \
//                                                         .resetckdivff(ckdiv2resetin)     \
//                                                        );
//
//module clockdivffreset_inv (ffoutresetb, ffinreset, clockinreset,resetckdivff);    
//output ffoutresetb;
//input ffinreset;
//input clockinreset;
//input resetckdivff;
//reg ffoutresetb;
//wire ffinreset, clockinreset, resetckdivff;
//`ifdef INTC_DC
//     `LIB_clockdivffreset(ffoutresetb, ffinreset, clockinreset,resetckdivff) 
//`else 
//always @(negedge (resetckdivff) or posedge clockinreset)
//begin
//  if (~(resetckdivff))
//    ffoutresetb = 1'b0; /* lintra s-60028 */
//  else
//    ffoutresetb = ~(ffinreset); /* lintra s-60028 */
//end
//`endif
//endmodule
//
//
//`define CLK_GATE_HF(o, clk, a)                                                               \
// soc_rbe_clk_hf \``soc_rbe_clk_hf_``o (                                                      \
//                                       .ckrcbxpn  (o),                                       \
//                                       .ckgridxpn (clk),                                     \
//                                       .latrcben  (a)                                        \
//                                      );
//module soc_rbe_clk_hf (output logic ckrcbxpn, input logic ckgridxpn, latrcben);  //lintra s-51506
//
//`ifdef INTC_DC
//     `LIB_soc_rbe_clk_hf(ckrcbxpn,ckgridxpn,latrcben) 
//`else
//   logic latrcbenl; // rce state element
//  
//  `ip2211ringpll_LATCH_P(latrcbenl, latrcben, ckgridxpn) //lintra s-51552
//  `ip2211ringpll_CLKAND(ckrcbxpn,ckgridxpn,latrcbenl)
//`endif
//endmodule // soc_rbe_clk_hf
//
////CLKBF_GLITCH_GLOB is a clkbuf used to remove glitches
////It is coded as a buffer, but this doesnot match the schematics.
////NEED TO CHECK IF INTC_SYNTHESIS ISNT REPLACING THE CELL WITH A BUFFER
//`define CLKBF_GLITCH_GLOB(clkout, clkin)                          \
//`ifdef INTC_DC                                                         \
//   `LIB_CLKBF_GLITCH_GLOB(clkout,clkin)                           \
//`else                                                             \
//   assign clkout = clkin;                                         \
//`endif
//
//`define CLKDIVFF(iffout, iffin, iclockin)             \
//clockdivff \``clockdivff_``iffout (                   \
//                                   .ffout(iffout),    \
//                                   .ffin(iffin),      \
//                                   .clockin(iclockin) \
//);
//
//// creating FF module to be used by clock macros below
//module clockdivff (ffout, ffin, clockin);    
//output ffout;
//input ffin;
//input clockin;
//reg ffout;
//wire ffin, clockin;
//`ifdef INTC_DC 
//     wire ffin_b;
//     assign ffin_b = ~ffin;
//     `LIB_clockdivff(ffout, ffin_b, clockin) 
//`else                                                                         
// always @(posedge clockin)                                                
//      begin                                                                  
//         ffout = ffin; /* lintra s-60028 */
//      end 
//`endif
//endmodule
//
//`define MAKE_CLK_GATE_TRUNK(igatedclk, iipclk, iusync, iresetb, iclken, idfx_scan_dbg_mode) \
//   clk_gate_trunk \``clk_gate_trunk_``igatedclk (                                           \
//                                                 .gatedclk(igatedclk),                      \
//                                                 .ipclk(iipclk),                            \
//                                                 .usync(iusync),                            \
//                                                 .resetb(iresetb),                          \
//                                                 .clken(iclken),                            \
//                                                 .dfx_scan_dbg_mode(idfx_scan_dbg_mode)     \
//                                                );
//
//module clk_gate_trunk(output logic gatedclk,
//                      input logic ipclk,
//                      input logic usync,
//                      input logic resetb,
//                      input logic clken,
//                      input logic dfx_scan_dbg_mode);
//logic clken_qual_in, clken_qual_out;
//logic qual_or_ovrd;
//assign clken_qual_in = usync ? clken : clken_qual_out;
//`ip2211ringpll_SET_MSFF(clken_qual_out, clken_qual_in, ipclk, ~resetb)
//assign qual_or_ovrd = clken_qual_out | dfx_scan_dbg_mode;
//`CLK_GATE_HF(gatedclk, ipclk, qual_or_ovrd)
//endmodule
//                                                
//











//`define MAKE_CLK_LOCAL_QUALDIV1TO16_ADJ(qual_out,inclk,inusync,inqualovrd,inratiosel)     \
//clk_qualdiv1to16_adj_local \``clk_qualdiv1to16_adj_local_``qual_out (                           \
//                                                                  .qualclk_out(qual_out),    \
//                                                                  .clk(inclk),               \
//                                                                  .usync(inusync),           \
//                                                                  .qualovrd(inqualovrd),     \
//                                                                  .ratiosel(inratiosel)     \
//                                                                 ); /* lintra s-51500, s-53048, s-53050 */
//
//module clk_qualdiv1to16_adj_local(qualclk_out, clk, usync, qualovrd, ratiosel);
//  output qualclk_out;
//  input clk;
//  input usync;
//  input qualovrd;
//  input [3:0] ratiosel;
//  logic qual_out;
//  `MAKE_QUAL_LOCAL_QUALDIV1TO8_ADJ(qual_out, clk, usync, qualovrd, ratiosel)        
//  `ip2211ringpll_CLK_GATE(qualclk_out, clk,  qual_out)
//endmodule
//
//
//
//`define MAKE_CLK_LOCAL_QUALDIV1TO8_ADJ(qual_out,inclk,inusync,inqualovrd,inratiosel)     \
//clk_qualdiv1to8_adj_local \``clk_qualdiv1to8_adj_local_``qual_out (                           \
//                                                                  .qualclk_out(qual_out),    \
//                                                                  .clk(inclk),               \
//                                                                  .usync(inusync),           \
//                                                                  .qualovrd(inqualovrd),     \
//                                                                  .ratiosel(inratiosel)     \
//                                                                 ); /* lintra s-51500, s-53048, s-53050 */
//module clk_qualdiv1to8_adj_local(qualclk_out, clk, usync, qualovrd, ratiosel);
//  output qualclk_out;
//  input clk;
//  input usync;
//  input qualovrd;
//  input [2:0] ratiosel;
//  logic qual_out;
//  `MAKE_QUAL_LOCAL_QUALDIV1TO8_ADJ(qual_out, clk, usync, qualovrd, ratiosel)        
//  `ip2211ringpll_CLK_GATE(qualclk_out, clk,  qual_out) //lintra s-51557, s-51552
//endmodule
//
//`define MAKE_CLK_NOREN(cknorenout,cknorenckin,cknorenenin)              \
//clknoren \``clknoren_``cknorenout (                                     \
//                              .clknorenout (cknorenout),                \
//                              .clknorenckin (cknorenckin),              \
//                              .clknorenenin (cknorenenin)               \
//                             );
//
//module clknoren(clknorenout,clknorenckin,clknorenenin);
//output clknorenout;
//input clknorenckin;
//input clknorenenin;
//wire clknorenout,clknorenckin,clknoreneninip2211ringpll_SOC_CLOCK_MACROS_VH;
//`ifdef INTC_DC
//     `LIB_clknoren(clknorenout,clknorenckin,clknorenenin) 
//`else
//assign clknorenout = ~(clknorenckin|clknorenenin);
//`endif
//endmodule
//



//
//`define MAKE_QUAL_LOCAL_QUALDIV16(qual_out, inclk, inusync, inqualovrd)          \
// qualdiv16_local \``qualdiv16_``qual_out (                                       \
//                                         .qualifier_out(qual_out),               \
//                                         .ipinclk(inclk) ,                       \
//                                         .usync(inusync),                        \
//                                         .qualovrd(inqualovrd)                   \
//                                         );
//module qualdiv16_local (qualifier_out,ipinclk,usync,qualovrd);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
// 
//  logic usync_lat, qual_staged, qual;
//  logic [3:0] nxt;
//  logic [3:0] pst;
// 
//  `ip2211ringpll_LATCH_P_DESKEW(usync_lat, usync, ipinclk)
//  assign nxt = pst + 4'b0001;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_lat)
//  assign qual = (&(pst));
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule
//
//`define MAKE_QUAL_LOCAL_QUALDIV1TO16_ADJ(qual_out, inclk, inusync, inqualovrd, inratiosel)     \
// qualdiv1to16_adj_local \``qualdiv1to16adj_``qual_out (                                         \
//                                                    .qualifier_out(qual_out),                 \
//                                                    .ipinclk(inclk) ,                         \
//                                                    .usync(inusync),                          \
//                                                    .qualovrd(inqualovrd),                    \
//                                                    .ratiosel(inratiosel)                     \
//                                                    );
///* lintra s-51500, s-53048, s-53050 */
//module qualdiv1to16_adj_local (qualifier_out,ipinclk,usync,qualovrd,ratiosel);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
//  input [3:0] ratiosel;
// 
//  logic usync_or_qual_lat, usync_or_qual, qual_staged, qual;
//  logic [3:0] ratiosel_muxed_staged, ratiosel_muxed;
//  logic [3:0] nxt;
//  logic [3:0] pst;
// 
//  //Whenever a qual or usync comes through we reset the counter
//  assign usync_or_qual = usync | qual;
//
//  `ip2211ringpll_LATCH_P_DESKEW(usync_or_qual_lat, usync_or_qual, ipinclk)
//  assign nxt = pst + 4'b0001;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_or_qual_lat)
//
//  //only grab ratiosel on usync boundary
//  assign ratiosel_muxed = usync ? ratiosel : ratiosel_muxed_staged;
//  `ip2211ringpll_MSFF(ratiosel_muxed_staged, ratiosel_muxed, ipinclk)
//
//  //Once we've reached the count that matches the ratiosel we're dividing by
//  //Set the qual indicator and reset the count
//  assign qual = (pst == ratiosel_muxed_staged);
//
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = qual_staged | qualovrd;
//endmodule // qualdiv1to16_adj_local
//
//`define MAKE_QUAL_LOCAL_QUALDIV1TO8_ADJ_WEN(qual_out, inclk, inusync, inqualovrd, inratiosel, inenable)     \
// qualdiv1to8_adj_wen_local \``qualdiv1to8adjwen_``qual_out (                                         \
//                                                    .qualifier_out(qual_out),                 \
//                                                    .ipinclk(inclk) ,                         \
//                                                    .usync(inusync),                          \
//                                                    .qualovrd(inqualovrd),                    \
//                                                    .ratiosel(inratiosel),                    \
//                                                    .enable(inenable)                         \
//                                                    );
///* lintra s-51500, s-53048, s-53050 */
//module qualdiv1to8_adj_wen_local (qualifier_out,ipinclk,usync,qualovrd,ratiosel,enable);
//  output qualifier_out;
//  input ipinclk;
//  input usync;
//  input qualovrd;
//  input [2:0] ratiosel;
//  input enable;
// 
//  logic usync_or_qual_lat, usync_or_qual, qual_staged, qual;
//  logic [2:0] ratiosel_muxed_staged, ratiosel_muxed;
//  logic [2:0] nxt;
//  logic [2:0] pst;
// 
//  //Whenever a qual or usync comes through we reset the counter
//  assign usync_or_qual = usync | qual;
//
//  `ip2211ringpll_LATCH_P_DESKEW(usync_or_qual_lat, usync_or_qual, ipinclk)
//  assign nxt = pst + 1;
//  `ip2211ringpll_RST_MSFF(pst, nxt, ipinclk, usync_or_qual_lat)
//
//  //only grab ratiosel on usync boundary
//  assign ratiosel_muxed = usync ? ratiosel : ratiosel_muxed_staged;
//  `ip2211ringpll_MSFF(ratiosel_muxed_staged, ratiosel_muxed, ipinclk)
//
//  //Once we've reached the count that matches the ratiosel we're dividing by
//  //Set the qual indicator and reset the count
//  assign qual = (pst == ratiosel_muxed_staged);
//
//  `ip2211ringpll_MSFF(qual_staged, qual, ipinclk)
//  assign qualifier_out = (qual_staged & enable) | qualovrd;
//endmodule // qualdiv1to8_adj_wen_local
//
//
////module qual_5_2(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [2:0]           count;
//
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 3'b000;
//     else
//       count <= (count + 3'b001) & {3{~(count == 4)}};
//
//   assign              fast_qual = (count == 0  ||
//                                    count == 3);
//   assign              slow_qual = 1'b1;
//endmodule //qual_5_2
//
//
//module qual_1_1(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//  
//   assign              fast_qual = 1'b1;
//   assign              slow_qual = 1'b1;
//endmodule // qual_1_1
//
//module qual_4_3(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [1:0]           count;
//
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//
//   assign              fast_qual = ~(count == 2);
//   assign              slow_qual = 1'b1;
//endmodule // qual_4_3
//
//module qual_8_5(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [2:0]           count;
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//   assign              fast_qual = (count == 0 ||
//                                    count == 2 ||
//                                    count == 3 ||
//                                    count == 5 ||
//                                    count == 6);
//   assign              slow_qual = 1'b1;
//endmodule // qual_8_5
//
//module qual_2_1(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg                 count;
//
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//
//   assign              fast_qual = count == 0;
//   assign              slow_qual = 1'b1;
//endmodule // qual_2_1
//
//module qual_16_7(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [3:0]           count;
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//   assign              fast_qual = (count == 0  ||
//                                    count == 2  ||
//                                    count == 5  ||
//                                    count == 7  ||
//                                    count == 9  ||
//                                    count == 11 ||
//                                    count == 14);
//   assign              slow_qual = 1'b1;
//endmodule // qual_16_7
//
//module qual_8_3(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [2:0]           count;
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//   assign              fast_qual = (count == 0 ||
//                                    count == 3 ||
//                                    count == 5);
//   assign              slow_qual = 1'b1;
//endmodule // qual_8_3
//
//module qual_16_5(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [3:0]           count;
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//   assign              fast_qual = (count == 0  ||
//                                    count == 3  ||
//                                    count == 6  ||
//                                    count == 10 ||
//                                    count == 13);
//   assign              slow_qual = 1'b1;
//endmodule // qual_16_5
//
//module qual_4_1(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [1:0]           count;
//
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= count + 1;
//
//   assign              fast_qual = count == 0;
//   assign              slow_qual = 1'b1;
//endmodule // qual_4_1
//
//module qual_5_3(
//                input usync_fast_clk,
//                input fast_clk,
//                output fast_qual,
//                output slow_qual
//                );
//   reg [2:0]           count;
//
//   always@(posedge fast_clk)
//     if(usync_fast_clk)
//       count <= 0;
//     else
//       count <= (count + 1) & {3{~(count == 4)}};
//
//   assign              fast_qual = (count == 1  ||
//                                    count == 2  ||
//                                    count == 4);
//   assign              slow_qual = 1'b1;
//endmodule // qual_5_3
//
//
//
//module det_clkdomainX_with_usync #(parameter dWidth = 32, parameter fifo_depth = 10, parameter separation = 2) 
////  for synchronization that's done between two clocks that are derived from the same reference clock and use separation 1,
//// this synchronizer must initiate it's rd/wr pointers at usync and not at reset!
//// otherwise separation is not ensured.
//// module det_clkdomainX must be abandoned and only this module det_clkdomainX_with_usync must be used.
//                     (
//                      input reset_ckRd,
//                      input reset_ckWr,
//                      input ckWr,
//                      input ckRd,
//                      input qualWr,
//                      input qualRd,
//                    input first_usyncWr,
//                    input first_usyncRd,
//                      input [dWidth-1:0] data_in,
//                      output [dWidth-1:0] data_out
//                      );
//
//   logic [dWidth-1:0] det_clkdomainX_write_data_array[fifo_depth - 1:0];
//   logic [dWidth-1:0] det_clkdomainX_read_data_mux;
//   logic [fifo_depth - 1:0] wrptr;
//   logic [fifo_depth - 1:0] rdptr;
//   logic [fifo_depth - 1:0] start_ptr;
//   logic write_clk;
//   logic read_clk;
//
//   `ip2211ringpll_CLK_GATE(write_clk, ckWr, qualWr)
//   `ip2211ringpll_CLK_GATE(read_clk, ckRd, qualRd)
//  
//   // data path generation
//   always@(posedge write_clk or negedge reset_ckWr)
//     begin: write_clk_scope
//        integer i;
//        if (~reset_ckWr)
//          begin
//             for (i=0;i<fifo_depth;i=i+1)
//               begin
//                  det_clkdomainX_write_data_array[i] <= 0;
//               end
//          end
//        else
//          begin
//             for (i=0;i<fifo_depth;i=i+1)
//               begin
//                  if (wrptr[i])
//                    det_clkdomainX_write_data_array[i] <= data_in;
//               end
//          end
//     end
//
//   always@(posedge read_clk or negedge reset_ckRd)
//     begin: read_clk_scope
//        integer i;
//        if (~reset_ckRd)
//          begin
//             det_clkdomainX_read_data_mux <= 0;
//          end
//        else
//          begin
//             for (i=0;i<fifo_depth;i=i+1)
//               begin
//                  if (rdptr[i])
//                    det_clkdomainX_read_data_mux <= det_clkdomainX_write_data_array[i];
//               end
//          end
//     end
//
//   assign data_out = det_clkdomainX_read_data_mux;
//
//   // wrptr and rdptr generation
//   assign start_ptr = 1;
//   
//   always@(posedge write_clk or negedge reset_ckWr)
//     if(!reset_ckWr)
//       wrptr <= start_ptr << separation;
//     else if (first_usyncWr)
//       wrptr <= start_ptr << separation;
//     else
//       wrptr <= {wrptr[(fifo_depth - 2):0], wrptr[(fifo_depth - 1)]};
//
//   always@(posedge read_clk or negedge reset_ckRd)
//     if(!reset_ckRd)
//       rdptr <= start_ptr;
//     else if (first_usyncRd)
//       rdptr <= start_ptr;
//     else
//       rdptr <= {rdptr[(fifo_depth - 2):0], rdptr[(fifo_depth - 1)]};
//
//endmodule // det_clkdomainX_with_usync
//
`ifndef ip2211ringpll_INTEL_CHECKERS_VS
`define ip2211ringpll_INTEL_CHECKERS_VS

`ifndef INTC_SVA_LIB_SVA2009
`define ip2211ringpll_SVA_LIB_SVA2005
`endif

/*
### VER 7.0 ###

There are three files representing the library templates: 

intel_checkers_core.vs: Core Library templates.
intel_checkers_ext.vs: Project specific Library extensions.
intel_checkers_coverg_ext.vs: Covergroups library extensions.

Blocking the extensions part is done by defining the compiler directive:
 INTC_SVA_LIB_CORE.

*/



`ifndef ip2211ringpll_SVA_LIB_SVA2005
   `ifdef INTC_SVA_LIB_FINAL_SEMANTICS
        `define ip2211ringpll_FINAL final
   `else  
        `define ip2211ringpll_FINAL #0
   `endif 
`else
   `define ip2211ringpll_FINAL final
`endif

`ifndef ip2211ringpll_SVA_LIB_SVA2005
   `define ip2211ringpll_default_clk $inferred_clock
   `define ip2211ringpll_SYS_CLK $global_clock
`else
   `ifndef ip2211ringpll_NO_VCSSIM
      `define ip2211ringpll_default_clk null
   `else
      `define ip2211ringpll_default_clk $default_clk
   `endif
`endif



// === === ===  macro definitions for error reporting

`define ip2211ringpll_MSG $psprintf
`define ip2211ringpll_ERR_MSG else $error
`define ip2211ringpll_ERR `ip2211ringpll_ERR_MSG()
`define ip2211ringpll_ERR_MSG_VARG else $error
`define ip2211ringpll_WARNING_MSG else $warning
`define ip2211ringpll_WARN `ip2211ringpll_WARNING_MSG()
`define ip2211ringpll_FATAL_MSG else $fatal
`define ip2211ringpll_FATAL `ip2211ringpll_FATAL_MSG(2,"")
`define ip2211ringpll_INFO_MSG else $info

// The following mechanism is to allow the project to control printing the 'cover message'
// generated information to stdout. When using cover properties, the messages
// generated by the simulator/emulator may slow down the runtime significantly.
// It is used by some tools (JemHW) during compilation time without any impact on
// performance.
// The following mechanism enables several control modes:
//      1) Basic compile-time expression, such as 1'b0.  (Recommended)
//      2) Runtime global/local expression: users can implement/define dedicated 
//         signal/signals to cover message information. They may choose a global
//         signal to represent the whole design or several signals defined across 
//         the design hierarchies. These signals should be driven either during
//         simulation (CTE injection / do file / use $test$plusargs()/ ... ) or
//         in the design itself.
// 
`ifdef INTC_SVA_LIB_ENABLE_COVER_STDOUT
    `ifdef INTC_SVA_LIB_COVER_STDOUT_EXPR
        `define ip2211ringpll_COVER_MSG if(`INTC_SVA_LIB_COVER_STDOUT_EXPR) $info 
    `else
        `define ip2211ringpll_COVER_MSG $info
    `endif
`else
     `define ip2211ringpll_COVER_MSG if(1'b0) $info
`endif


`define ip2211ringpll_ERR_GLITCH_MSG(text, glitch_ns) $info("assertion is up"); \
  else $error("%s Not sensitive to glitch less than %d ns", (text), (glitch_ns))


// === === === Implementation for the templates

//`include "intel_checkers_core.vs"

// --- --- --- --- --- --- --- --- --- --- ----


`ifndef INTC_SVA_LIB_CORE

//`include "intel_checkers_ext.vs"
//`include "intel_checkers_coverg_ext.vs"

`endif


`endif // ip2211ringpll_INTEL_CHECKERS_VS


`ifndef ip2211ringpll_INTEL_CHECKERS_CORE_VS
`define ip2211ringpll_INTEL_CHECKERS_CORE_VS

/*                                                                             
There are two kinds of core entities, sequential and combinational.            
The combinational entities do not use a sampling clock and are implemented     
on top of deferred assertions.                                                 
The sequential entities require a clock for sampling the design signals and    
are implemented on top of concurrent assertions.                               

The sequential entities can infer the clock from its context if not specified  
explicitly in the entity instance. The clk is inherited either from the        
enclosing always procedure (with posedge/negedge control) or from the default  
clocking. The reset has a default value of 1'b0. Therefore, if an actual       
argument for rst is omitted, the assertion is always enabled.                  

Both kinds of entities can be instantiated in procedural and in concurrent     
(structural) contexts. Both positional and named association between the       
formal and the actual arguments is supported.                                  
The combinational entities start with ASSERTC, The sequential entities start   
with ASSERTS. The legacy format used by SNB is also supported.                 

Stability assertions: there are two sets of sequential entities:               
Those checking also between specified clock ticks, and those which check only  
on specified clock ticks.                                                      

Note 1:  the first operate on system clock that samples the design clock, clk, 
and the design signals. Those entities start with ASSERTS_G... . These entities
trigger on both edges of the system clock.                                     

Note2: The system-clock based entites come in two varieties,  event based      
checkers and signal based.  They are distinguished by the suffixes in the names.
For the second  group only the clock name or its complement must be provided as
the  actual argument, i.e., there should be no edge specifier.                 



Examples:                                                                      
=========                                                                      

Combinational entity:                                                          
    `ip2211ringpll_ASSERTC_MUTEXED(name, myBusEnables, `ip2211ringpll_ERR_MSG("I have error"));            

Sequential entity:                                                             
    `ip2211ringpll_ASSERTS_TRIGGER(name, x, y, posedge clk, rst, `ip2211ringpll_ERR_MSG("I have error"));  

Usage Examples:                                                                
    // declare default clock if so desired                                     
    default clocking def_clk @(posedge clk);                                   
    endclocking                                                                

    Positional association:                                                    
       // clk inferred either from always or def_clk, rst is 0                 
       `ip2211ringpll_ASSERTS_TRIGGER(name, x, y, , , `ip2211ringpll_ERR_MSG("I have error"))              
       // clk inferred either from always or def_clk,                          
       `ip2211ringpll_ASSERTS_TRIGGER(name, x, y, , rst, `ip2211ringpll_ERR_MSG("I have error"))           
       // default rst of 0                                                     
       `ip2211ringpll_ASSERTS_TRIGGER(name, x, y, posedge clk, , `ip2211ringpll_ERR_MSG("I have error"))   
       // no default or inference                                              
       `ip2211ringpll_ASSERTS_TRIGGER(name, x, y, posedge clk, rst, `ip2211ringpll_ERR_MSG("I have error"))

    Named associations:                                                        
        // clk inferred either from always or def_clk, rst is 0                
       `ip2211ringpll_ASSERTS_TRIGGER(name, .en(x), .ev(y), .prop(z), `ip2211ringpll_ERR_MSG("I have error"))

*/                                                                             






// === === === Implementation for the templates                                

//`include "intel_checkers_core_imp.vs"                                          

// --- --- --- --- --- --- --- --- --- --- ----                                



// ****************************************************************************************** //
// Common arguments:                                                           
//      clk     event       Clock event. Default: $inferred_clock.             
//      rst     Boolean     Reset signal.                                      
//      name    string      Assertion label.                                   
//      ip2211ringpll_MSG     string      Error message.                                     
//                                                                             
// ------------------------------------------------------------------------------------------ //

// --- --- --- Immediate Templates --- --- --- //                              


// ****************************************************************************************** //
// Name:   mutexed                                                             
// Category: Combinational                                                     
// Description:                                                                
//       At most one bit of 'sig' is high. x and z values are counted, which means that at most
//       one bit can be high or x or z.                                        
// Arguments:                                                                  
//       - sig    Bit-vector  At most one bit of <sig> is high. Limitation: 'sig' must be a packed
//       array                                                                 
// Comments:                                                                   
//       - MUTEXED is equivalent to AT_MOST_BITS_HIGH where 'n' is equal to 1. 
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//       - The pass or failure of an immediate assertion inside an always_ff block would be delayed
//         by one sampling edge compared to when the assertion is in an always_comb or in
//         structural context.                                                 
// Related:                                                                    
//       ONE_HOT                                                               
//       AT_MOST_BITS_HIGH                                                     
//       BITS_HIGH                                                             
// Example:                                                                    
//       The following will fail | @VIEW@(001x);                               
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_MUTEXED(sig, rst)                                                \
    assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_mutexed(sig))  /* novas s-2050,s-2056 */             

`define ip2211ringpll_ASSUME_MUTEXED(sig, clk, rst)                                           \
    assume property(p_mutexed(sig, clk, rst))                                  

`define ip2211ringpll_COVER_MUTEXED(sig, clk, rst)                                            \
    cover property(p_cover_mutexed(sig, clk, rst))                             

`define ip2211ringpll_NOT_MUTEXED_COVER(sig, clk ,rst)                                        \
    cover property(p_not_mutexed_covered(sig, clk, rst))                       

`endif                                                                         


`define ip2211ringpll_ASSERTC_MUTEXED(name, sig, rst, ip2211ringpll_MSG)                                    \
    name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_mutexed(sig)) /* novas s-2050,s-2056 */   ip2211ringpll_MSG  

`define ip2211ringpll_ASSUMEC_MUTEXED(name, sig, rst, ip2211ringpll_MSG)                                    \
    name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_mutexed(sig)) /* novas s-2050,s-2056 */   ip2211ringpll_MSG  


`define ip2211ringpll_ASSERTS_MUTEXED(name, sig, clk, rst, ip2211ringpll_MSG)                               \
    name: assert property(p_mutexed(sig, clk, rst)) ip2211ringpll_MSG                        

`define ip2211ringpll_ASSUMES_MUTEXED(name, sig, clk, rst, ip2211ringpll_MSG)                               \
    name: assume property(p_mutexed(sig, clk, rst)) ip2211ringpll_MSG                        


`define ip2211ringpll_COVERC_MUTEXED(name, sig, rst, ip2211ringpll_MSG)                                     \
    `ifndef INTC_SVA_LIB_COVER_ENABLE                                                \
        typedef bit t_``name                                                    \
    `else                                                                       \
        name: cover `ip2211ringpll_FINAL (!(rst) && `ip2211ringpll_l_mutexed(sig)) /* novas s-2050,s-2056 */  ip2211ringpll_MSG \
    `endif                                                                     

`define ip2211ringpll_COVERS_MUTEXED(name, sig, clk, rst, ip2211ringpll_MSG)                                \
    `ifndef INTC_SVA_LIB_COVER_ENABLE                                                \
        typedef bit t_``name                                                    \
    `else                                                                       \
        name: cover property(p_cover_mutexed(sig, clk, rst)) ip2211ringpll_MSG                \
    `endif                                                                     



`define ip2211ringpll_NOT_MUTEXED_COVERC(name, sig, rst, ip2211ringpll_MSG)                                 \
    `ifndef INTC_SVA_LIB_COVER_ENABLE                                                \
        typedef bit t_``name                                                    \
    `else                                                                       \
        name: cover `ip2211ringpll_FINAL (!(rst) && ! `ip2211ringpll_l_mutexed(sig)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG  \
    `endif                                                                     


`define ip2211ringpll_NOT_MUTEXED_COVERS(name, sig, clk, rst, ip2211ringpll_MSG)                            \
    `ifndef INTC_SVA_LIB_COVER_ENABLE                                                \
        typedef bit t_``name                                                    \
    `else                                                                       \
        name: cover property(p_not_mutexed_covered(sig, clk, rst)) ip2211ringpll_MSG          \
    `endif                                                                     

// ****************************************************************************************** //



// --- --- ---                                                                 



// ****************************************************************************************** //
// Name:   one hot                                                             
// Category: Combinational                                                     
// Description:                                                                
//       Exactly one bit of 'sig' is high, other bits are low, and there are no x and z values
//       in 'sig'.                                                             
// Arguments:                                                                  
//       - sig    Bit-vector  Exactly one bit of 'sig' is high.                
// Comments:                                                                   
//       - ONE_HOT is equivalent to BITS_HIGH where 'n' is equal to 1.         
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//         The pass or failure of an immediate assertion inside an always_ff block would be delayed
//         by one sampling edge compared to when the assertion is in an always_comb or in structural
//         context.                                                            
// Related:                                                                    
//       MUTEXED                                                               
//       AT_MOST_BITS_HIGH                                                     
//       BITS_HIGH                                                             
// Example:                                                                    
//       The following will fail | @VIEW@(001x);                               
//                                                                             
// ------------------------------------------------------------------------------------------ //


`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_ONE_HOT(sig, rst)                                                \
   assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_one_hot(sig))      /* novas s-2050,s-2056 */       

`define ip2211ringpll_ASSUME_ONE_HOT(sig, clk, rst)                                           \
   assume property(p_one_hot(sig, clk, rst))                                   

`define ip2211ringpll_COVER_ONE_HOT(sig, clk, rst)                                            \
   cover property(p_cover_one_hot(sig, clk, rst))                              

`define ip2211ringpll_NOT_ONE_HOT_COVER(sig, clk, rst)                                        \
   cover property(p_not_one_hot_cover(sig, clk, rst))                          

`endif                                                                         



`define ip2211ringpll_ASSERTC_ONE_HOT(name, sig, rst, ip2211ringpll_MSG)                                    \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_one_hot(sig)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG     

`define ip2211ringpll_ASSUMEC_ONE_HOT(name, sig, rst, ip2211ringpll_MSG)                                    \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_one_hot(sig)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG     



`define ip2211ringpll_ASSERTS_ONE_HOT(name, sig, clk, rst, ip2211ringpll_MSG)                               \
   name: assert property(p_one_hot(sig, clk, rst)) ip2211ringpll_MSG                         

`define ip2211ringpll_ASSUMES_ONE_HOT(name, sig, clk, rst, ip2211ringpll_MSG)                               \
   name: assume property(p_one_hot(sig, clk, rst)) ip2211ringpll_MSG                         



`define ip2211ringpll_COVERC_ONE_HOT(name, sig, rst, ip2211ringpll_MSG)                                     \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && `ip2211ringpll_l_one_hot(sig)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif

`define ip2211ringpll_COVERS_ONE_HOT(name, sig, clk, rst, ip2211ringpll_MSG)                                \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_cover_one_hot(sig, clk, rst)) ip2211ringpll_MSG                 \
   `endif



`define ip2211ringpll_NOT_ONE_HOT_COVERC(name, sig, rst, ip2211ringpll_MSG)                                 \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && !`ip2211ringpll_l_one_hot(sig)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif

`define ip2211ringpll_NOT_ONE_HOT_COVERS(name, sig, clk, rst, ip2211ringpll_MSG)                            \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_not_one_hot_cover(sig, clk, rst)) ip2211ringpll_MSG             \
   `endif



// ****************************************************************************************** //



// --- --- ---                                                                 



// ****************************************************************************************** //
// Name:   same bits                                                           
// Category: Combinational                                                     
// Description:                                                                
//       All bits of 'sig' have the same value: high or low.                   
// Arguments:                                                                  
//       - sig    Bit-vector    All bits of 'sig' have the same value: high or low. 
// Comments:                                                                   
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//       - The pass or failure of an immediate assertion inside an always_ff block would be
//         delayed by one sampling edge compared to when the assertion is in an always_comb or
//         in structural context.                                              
// Related:                                                                    
//       None                                                                  
// Example:                                                                    
//       The following will fail | @VIEW@(000x);                               
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_SAME_BITS(sig, rst)                                              \
   assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_same_bits(sig))        /* novas s-2050,s-2056 */      

`define ip2211ringpll_ASSUME_SAME_BITS(sig, clk, rst)                                         \
   assume property(p_same_bits(sig, clk, rst))                                 

`define ip2211ringpll_COVER_SAME_BITS(sig, clk, rst)                                          \
   cover property(p_cover_same_bits(sig, clk, rst))                            

`define ip2211ringpll_NOT_SAME_BITS_COVER(sig, clk, rst)                                      \
   cover property(p_not_same_bits_cover(sig, clk, rst))                        

`endif                                                                         



`define ip2211ringpll_ASSERTC_SAME_BITS(name, sig, rst, ip2211ringpll_MSG)                                  \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_same_bits(sig)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG                      

`define ip2211ringpll_ASSUMEC_SAME_BITS(name, sig, rst, ip2211ringpll_MSG)                                  \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_same_bits(sig)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG                      



`define ip2211ringpll_ASSERTS_SAME_BITS(name, sig, clk, rst, ip2211ringpll_MSG)                             \
   name: assert property(p_same_bits(sig, clk, rst)) ip2211ringpll_MSG                       

`define ip2211ringpll_ASSUMES_SAME_BITS(name, sig, clk, rst, ip2211ringpll_MSG)                             \
   name: assume property(p_same_bits(sig, clk, rst)) ip2211ringpll_MSG                       



`define ip2211ringpll_COVERC_SAME_BITS(name, sig, rst, ip2211ringpll_MSG)                                   \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && `ip2211ringpll_l_same_bits(sig)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif

`define ip2211ringpll_COVERS_SAME_BITS(name, sig, clk, rst, ip2211ringpll_MSG)                              \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_cover_same_bits(sig, clk, rst)) ip2211ringpll_MSG               \
   `endif



`define ip2211ringpll_NOT_SAME_BITS_COVERS(name, sig, clk, rst, ip2211ringpll_MSG)                          \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_not_same_bits_cover(sig, clk, rst)) ip2211ringpll_MSG           \
   `endif

`define ip2211ringpll_NOT_SAME_BITS_COVERC(name, sig, rst, ip2211ringpll_MSG)                               \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && ! `ip2211ringpll_l_same_bits(sig)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  range                                                                
// Category: Combinational                                                     
// Description:                                                                
//       Signal 'sig' must always be in the range [low, high], inclusive of both the range
//       values.                                                               
// Arguments:                                                                  
//       - sig    Bit-vector  Signal to be monitored for its value to be within a specified range.
//       - low    Number>=0   Lower bound on 'sig'.                            
//       - high   Number>=0   Upper bound on 'sig'.                            
// Comments:                                                                   
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//       - The pass or failure of an immediate assertion inside an always_ff block would be
//         delayed by one sampling edge compared to when the assertion is in an always_comb or
//         in structural context.                                              
// Related:                                                                    
//       ONE_OF                                                                
//       MIN                                                                   
//       MAX                                                                   
// Example:                                                                    
//       Valid port number is 5 to 10 | @VIEW@(port, 5, 10);                   
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_RANGE(sig, low, high, rst)                                       \
   assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_range(sig, low, high))     /* novas s-2050,s-2056,s-0393 */  

`define ip2211ringpll_ASSUME_RANGE(sig, low, high, clk, rst)                                  \
   assume property(p_range(sig, low, high, clk, rst))                          

`define ip2211ringpll_COVER_RANGE(sig, low, high, clk, rst)                                   \
   cover property(p_cover_range(sig, low, high, clk, rst))                     

`define ip2211ringpll_NOT_RANGE_COVER(sig, low, high, clk ,rst)                               \
   cover property(p_not_range_cover(sig, low, high, clk, rst))                 

`endif                                                                         


`define ip2211ringpll_ASSERTC_RANGE(name, sig, low, high, rst, ip2211ringpll_MSG)                           \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_range(sig, low, high)) /* novas s-2050,s-2056,s-0393 */ ip2211ringpll_MSG               

`define ip2211ringpll_ASSUMEC_RANGE(name, sig, low, high, rst, ip2211ringpll_MSG)                           \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_range(sig, low, high)) /* novas s-2050,s-2056,s-0393 */ ip2211ringpll_MSG             



`define ip2211ringpll_ASSERTS_RANGE(name, sig, low, high, clk, rst, ip2211ringpll_MSG)                      \
   name: assert property(p_range(sig, low, high, clk, rst)) ip2211ringpll_MSG                

`define ip2211ringpll_ASSUMES_RANGE(name, sig, low, high, clk, rst, ip2211ringpll_MSG)                      \
   name: assume property(p_range(sig, low, high, clk, rst)) ip2211ringpll_MSG                



`define ip2211ringpll_COVERC_RANGE(name, sig, low, high, rst, ip2211ringpll_MSG)                            \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && `ip2211ringpll_l_range(sig, low, high)) /* novas s-2050,s-2056,s-0393 */ ip2211ringpll_MSG \
   `endif

`define ip2211ringpll_COVERS_RANGE(name, sig, low, high, clk, rst, ip2211ringpll_MSG)                       \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property (p_cover_range(sig, low, high, clk, rst)) ip2211ringpll_MSG       \
   `endif



`define ip2211ringpll_NOT_RANGE_COVERS(name, sig, low, high, clk ,rst, ip2211ringpll_MSG)                   \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_not_range_cover(sig, low, high, clk, rst)) ip2211ringpll_MSG    \
   `endif

`define ip2211ringpll_NOT_RANGE_COVERC(name, sig, low, high, rst, ip2211ringpll_MSG)                        \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && ! `ip2211ringpll_l_range(sig, low, high)) /* novas s-2050,s-2056,s-0393 */ ip2211ringpll_MSG \
   `endif



// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  at most bits high                                                    
// Category: Combinational                                                     
// Description:                                                                
//       At most 'n' bits in 'sig' are high. x and z values are counted as high for this
//       calculation.                                                          
// Arguments:                                                                  
//       - sig    Bit-vector    At most 'n' bits in 'sig' can be high. Limitation: 'sig' must be
//                              a packed array.                                
//       - n      Number>=0     The maximum number of bits in 'sig' that are allowed to be high.
// Comments:                                                                   
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//       - The pass or failure of an immediate assertion inside an always_ff block would be
//         delayed by one sampling edge compared to when the assertion is in an always_comb or
//         in structural context.                                              
// Related:                                                                    
//       BITS_HIGH                                                             
//       MUTEXED                                                               
//       ONE_HOT                                                               
// Example:                                                                    
//       The following will fail | @VIEW@(001x, 1);                            
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_AT_MOST_BITS_HIGH(sig, n, rst)                                   \
   assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_at_most_bits_high(sig, n))     /* novas s-2050,s-2056 */

`define ip2211ringpll_ASSUME_AT_MOST_BITS_HIGH(sig, n, clk, rst)                              \
   assume property(p_at_most_bits_high(sig, n, clk, rst))                      

`define ip2211ringpll_COVER_AT_MOST_BITS_HIGH(sig, n, clk, rst)                               \
   cover property(p_cover_at_most_bits_high(sig, n, clk, rst))                 

`define ip2211ringpll_NOT_AT_MOST_BITS_HIGH_COVER(sig, n, clk, rst)                           \
   cover property(p_not_at_most_bits_high_cover(sig, n, clk, rst))             

`endif                                                                         



`define ip2211ringpll_ASSERTC_AT_MOST_BITS_HIGH(name, sig, n, rst, ip2211ringpll_MSG)                       \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_at_most_bits_high(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG

`define ip2211ringpll_ASSUMEC_AT_MOST_BITS_HIGH(name, sig, n, rst, ip2211ringpll_MSG)                       \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_at_most_bits_high(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG



`define ip2211ringpll_ASSERTS_AT_MOST_BITS_HIGH(name, sig, n, clk, rst, ip2211ringpll_MSG)                  \
   name: assert property(p_at_most_bits_high(sig, n, clk, rst)) ip2211ringpll_MSG            

`define ip2211ringpll_ASSUMES_AT_MOST_BITS_HIGH(name, sig, n, clk, rst, ip2211ringpll_MSG)                  \
   name: assume property(p_at_most_bits_high(sig, n, clk, rst)) ip2211ringpll_MSG            



`define ip2211ringpll_COVERC_AT_MOST_BITS_HIGH(name, sig, n, rst, ip2211ringpll_MSG)                        \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && `ip2211ringpll_l_at_most_bits_high(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif

`define ip2211ringpll_COVERS_AT_MOST_BITS_HIGH(name, sig, n, clk, rst, ip2211ringpll_MSG)                   \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_cover_at_most_bits_high(sig, n, clk, rst)) ip2211ringpll_MSG    \
   `endif



`define ip2211ringpll_NOT_AT_MOST_BITS_HIGH_COVERS(name, sig, n, clk, rst, ip2211ringpll_MSG)               \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_not_at_most_bits_high_cover(sig, n, clk, rst)) ip2211ringpll_MSG \
   `endif

`define ip2211ringpll_NOT_AT_MOST_BITS_HIGH_COVERC(name ,sig, n, rst, ip2211ringpll_MSG)                    \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && ! `ip2211ringpll_l_at_most_bits_high(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  bits high                                                            
// Category: Combinational                                                     
// Description:                                                                
//       Exactly 'n' bits of 'sig' are high, other bits are low, and there are no x or z
//       values in 'sig'.                                                      
// Arguments:                                                                  
//       - sig    Bit-vector   Exactly 'n' bits in 'sig' are high.             
//       - n      Number>=0    The number of bits in 'sig' that are high.      
// Comments:                                                                   
//       - BITS_HIGH where 'n' is equal to 1 is equivalent to ONE_HOT.         
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//       - The pass or failure of an immediate assertion inside an always_ff block would be
//         delayed by one sampling edge compared to when the assertion is in an always_comb or
//         in structural context.                                              
// Related:                                                                    
//       AT_MOST_BITS_HIGH                                                     
//       REMAIN_HIGH                                                           
//       BITS_LOW                                                              
//       ONE_HOT                                                               
// Example:                                                                    
//       The following will fail | @VIEW@(001x, 1);                            
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_BITS_HIGH(sig, n, rst)                                           \
   assert `ip2211ringpll_FINAL (( (|(rst)) | `ip2211ringpll_l_bits_high(sig, n)))     /* novas s-2050,s-2056 */   

`define ip2211ringpll_ASSUME_BITS_HIGH(sig, n, clk, rst)                                      \
   assume property(p_bits_high(sig, n, clk, rst))                              

`define ip2211ringpll_COVER_BITS_HIGH(sig, n, clk, rst)                                       \
   cover property(p_cover_bits_high(sig, n, clk, rst))                         

`define ip2211ringpll_NOT_BITS_HIGH_COVER(sig, n, clk, rst)                                   \
   cover property(p_not_bits_high_cover(sig, n, clk, rst))                     

`endif                                                                         



`define ip2211ringpll_ASSERTC_BITS_HIGH(name, sig, n, rst, ip2211ringpll_MSG)                               \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_bits_high(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG

`define ip2211ringpll_ASSUMEC_BITS_HIGH(name, sig, n, rst, ip2211ringpll_MSG)                               \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_bits_high(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG



`define ip2211ringpll_ASSERTS_BITS_HIGH(name, sig, n, clk, rst, ip2211ringpll_MSG)                          \
   name: assert property(p_bits_high(sig, n, clk, rst)) ip2211ringpll_MSG                    

`define ip2211ringpll_ASSUMES_BITS_HIGH(name, sig, n, clk, rst, ip2211ringpll_MSG)                          \
   name: assume property(p_bits_high(sig, n, clk, rst)) ip2211ringpll_MSG                    



`define ip2211ringpll_COVERS_BITS_HIGH(name, sig, n, clk, rst, ip2211ringpll_MSG)                           \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_cover_bits_high(sig, n, clk, rst)) ip2211ringpll_MSG            \
   `endif

`define ip2211ringpll_COVERC_BITS_HIGH(name, sig, n, rst, ip2211ringpll_MSG)                                \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && `ip2211ringpll_l_bits_high(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif



`define ip2211ringpll_NOT_BITS_HIGH_COVERS(name, sig, n, clk, rst, ip2211ringpll_MSG)                       \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_not_bits_high_cover(sig, n, clk, rst)) ip2211ringpll_MSG        \
   `endif

`define ip2211ringpll_NOT_BITS_HIGH_COVERC(name ,sig, n, rst, ip2211ringpll_MSG)                            \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && ! `ip2211ringpll_l_bits_high(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  one of                                                               
// Category: Combinational                                                     
// Description:                                                                
//      Signal 'sig' must be equal to one of the values listed.                
// Arguments:                                                                  
//       - sig    Bit-vector   Signal to be monitored for its value to be one of the values listed.
//       - set    Number>=0    Comma separated set of integers.                
// Comments:                                                                   
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//       - The pass or failure of an immediate assertion inside an always_ff block would be delayed
//         by one sampling edge compared to when the assertion is in an always_comb or in
//         structural context.                                                 
//       - set of elements is currently not supported in let statments         
//       - Sequential views are not supported for this macro.                  
// Related:                                                                    
//       RANGE                                                                 
//       MIN                                                                   
//       MAX                                                                   
// Example:                                                                    
//       TBD |                                                                 
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_ONE_OF(sig, set, rst)                                            \
   assert `ip2211ringpll_FINAL ((|(rst)) | ((sig) inside set) & `ip2211ringpll_SVA_LIB_KNOWN(sig))  /* novas s-2050,s-2056 */

// `define ASSUME_ONE_OF(sig, set, clk, rst)                                    \
//    assume property(p_one_of(sig, set, clk, rst))                            

// `define COVER_ONE_OF(sig, sig, clk, rst)                                     \
//    cover property(p_cover_one_of(sig, set, clk, rst))                       

// `define NOT_ONE_OF_COVER(sig, sig, clk, rst)                                 \
//    cover property(p_not_one_of_cover(sig, set, clk, rst))                   

`endif                                                                         


`define ip2211ringpll_ASSERTC_ONE_OF(name, sig, set, rst, ip2211ringpll_MSG)                                \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | (((sig) inside set) & `ip2211ringpll_SVA_LIB_KNOWN(sig))) /* novas s-2050,s-2056 */ ip2211ringpll_MSG

`define ip2211ringpll_ASSUMEC_ONE_OF(name, sig, set, rst, ip2211ringpll_MSG)                                \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | (((sig) inside set) & `ip2211ringpll_SVA_LIB_KNOWN(sig))) /* novas s-2050,s-2056 */ ip2211ringpll_MSG



// `define ASSUMES_ONE_OF(name, sig, set, clk, rst, ip2211ringpll_MSG)                        \
//    name: `ASSUME_ONE_OF(sig, set, clk, rst) ip2211ringpll_MSG                             

// `define ASSERTS_ONE_OF(name, sig, set, clk, rst, ip2211ringpll_MSG)                        \
//    name: assert property(p_one_of(sig, set, clk, rst)) ip2211ringpll_MSG                  



// `define COVERS_ONE_OF(name, sig, set, clk, rst, ip2211ringpll_MSG)                         \
//    name: `COVER_ONE_OF(sig, set, clk, rst) ip2211ringpll_MSG                              

`define ip2211ringpll_COVERC_ONE_OF(name, sig, set, rst, ip2211ringpll_MSG)                                 \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && ((sig) inside set)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif



// `define NOT_ONE_OF_COVERS(name, sig, set, clk, rst, ip2211ringpll_MSG)                     \
//    name: `NOT_ONE_OF_COVER(sig, set, clk, rst) ip2211ringpll_MSG                          

`define ip2211ringpll_NOT_ONE_OF_COVERC(name ,sig, set, rst, ip2211ringpll_MSG)                             \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && !((sig) inside set)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:   known driven                                                        
// Category: Combinational                                                     
// Description:                                                                
//       All bits of 'sig' are both known (not X) and driven (not Z). This property passes
//       vacuously in formal verification since signals in formal verification have concrete
//       (known) values (0 or 1).                                              
// Arguments:                                                                  
//       - sig    Bit-vector    Signal to check.                               
// Comments:                                                                   
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//       - The pass or failure of an immediate assertion inside an always_ff block would be delayed
//         by one sampling edge compared to when the assertion is in an always_comb or in structural
//         context.                                                            
// Related:                                                                    
//       None                                                                  
// Example:                                                                    
//       Not relevant|                                                         
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_KNOWN_DRIVEN(sig, rst)                                           \
   assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_known_driven(sig))     /* novas s-2050,s-2056 */     

`define ip2211ringpll_ASSUME_KNOWN_DRIVEN(sig, clk, rst)                                      \
   assume property(p_known_driven(sig, clk, rst))                              

`define ip2211ringpll_COVER_KNOWN_DRIVEN(sig, clk ,rst)                                       \
   cover property(p_cover_known_driven(sig, clk, rst))                         

`define ip2211ringpll_NOT_KNOWN_DRIVEN_COVER(sig, clk ,rst)                                   \
   cover property(p_not_known_driven_cover(sig, clk, rst))                     

`endif                                                                         


`define ip2211ringpll_ASSERTC_KNOWN_DRIVEN(name, sig, rst, ip2211ringpll_MSG)                               \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_known_driven(sig)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG

`define ip2211ringpll_ASSUMEC_KNOWN_DRIVEN(name, sig, rst, ip2211ringpll_MSG)                               \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_known_driven(sig)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG



`define ip2211ringpll_ASSERTS_KNOWN_DRIVEN(name, sig, clk, rst, ip2211ringpll_MSG)                          \
   name: assert property(p_known_driven(sig, clk, rst)) ip2211ringpll_MSG                    

`define ip2211ringpll_ASSUMES_KNOWN_DRIVEN(name, sig, clk, rst, ip2211ringpll_MSG)                          \
   name: assume property(p_known_driven(sig, clk, rst)) ip2211ringpll_MSG                    



`define ip2211ringpll_COVERS_KNOWN_DRIVEN(name, sig, clk, rst, ip2211ringpll_MSG)                           \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_cover_known_driven(sig, clk, rst)) ip2211ringpll_MSG            \
   `endif

`define ip2211ringpll_COVERC_KNOWN_DRIVEN(name, sig, rst, ip2211ringpll_MSG)                                \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && `ip2211ringpll_l_known_driven(sig)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif



`define ip2211ringpll_NOT_KNOWN_DRIVEN_COVERS(name, sig, clk, rst, ip2211ringpll_MSG)                       \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_not_known_driven_cover(sig, clk, rst)) ip2211ringpll_MSG        \
   `endif

`define ip2211ringpll_NOT_KNOWN_DRIVEN_COVERC(name, sig, rst, ip2211ringpll_MSG)                            \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && ! `ip2211ringpll_l_known_driven(sig)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif


// ****************************************************************************************** //



// --- --- ---                                                                 

// ****************************************************************************************** //
// Name:   same                                                                
// Category: Combinational                                                     
// Description:                                                                
//       The vectors have same value . The checker compares 2 input vectors - 'siga' has the
//       same value as 'sigb'.                                                 
// Arguments:                                                                  
//       - siga    Bit-vector    First vector to be checked.                   
//       - sigb    Bit-vector    Second vector to be checked.                  
// Comments:                                                                   
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//       - The pass or failure of an immediate assertion inside an always_ff block would be
//         delayed by one sampling edge compared to when the assertion is in an always_comb or
//         in structural context.                                              
// Related:                                                                    
//       SAME_BITS                                                             
// Example:                                                                    
//       Not relevant. |                                                       
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_SAME(siga, sigb, rst)                                            \
    assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_same(siga, sigb))    /* novas s-2050,s-2056 */       

`define ip2211ringpll_ASSUME_SAME(siga, sigb, clk, rst)                                       \
    assume property(p_same(siga, sigb, clk, rst))                              

`define ip2211ringpll_COVER_SAME(siga, sigb, clk, rst)                                        \
    cover property(p_cover_same(siga, sigb, clk, rst))                         

`define ip2211ringpll_NOT_SAME_COVER(siga, sigb, clk, rst)                                    \
    cover property(p_not_same_cover(siga, sigb, clk, rst))                     

`endif                                                                         



`define ip2211ringpll_ASSERTC_SAME(name, siga, sigb, rst, ip2211ringpll_MSG)                                \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_same(siga, sigb)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG 

`define ip2211ringpll_ASSUMEC_SAME(name, siga, sigb, rst, ip2211ringpll_MSG)                                \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_same(siga, sigb)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG 



`define ip2211ringpll_ASSERTS_SAME(name, siga, sigb, clk, rst, ip2211ringpll_MSG)                           \
   name: assert property(p_same(siga, sigb, clk, rst)) ip2211ringpll_MSG                     

`define ip2211ringpll_ASSUMES_SAME(name, siga, sigb, clk, rst, ip2211ringpll_MSG)                           \
   name: assume property(p_same(siga, sigb, clk, rst)) ip2211ringpll_MSG                     



`define ip2211ringpll_COVERC_SAME(name, siga, sigb, rst, ip2211ringpll_MSG)                                 \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && `ip2211ringpll_l_same(siga, sigb)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif

`define ip2211ringpll_COVERS_SAME(name, siga, sigb, clk, rst, ip2211ringpll_MSG)                            \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_cover_same(siga, sigb, clk ,rst)) ip2211ringpll_MSG             \
   `endif



`define ip2211ringpll_NOT_SAME_COVERC(name, siga, sigb, rst, ip2211ringpll_MSG)                             \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && !(`ip2211ringpll_l_same(siga, sigb))) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif

`define ip2211ringpll_NOT_SAME_COVERS(name, siga, sigb, clk, rst, ip2211ringpll_MSG)                        \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_not_same_cover(siga, sigb, clk, rst)) ip2211ringpll_MSG         \
   `endif


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:   must                                                                
// Category: Combinational                                                     
// Description:                                                                
//       Boolean condition 'prop' must always be true.                         
// Arguments:                                                                  
//       - prop    Boolean  The boolean condition that must always be true.    
// Comments:                                                                   
//       - The condition must be a boolean.                                    
//       - When the condition is boolean and clocked, ip2211ringpll_ASSERTS_MUST is equivalent to ip2211ringpll_ASSERTS_VERIFY.
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//       - The pass or failure of an immediate assertion inside an always_ff block would be delayed by 
//         one sampling edge compared to when the assertion is in an always_comb or in structural
//         context.                                                            
// Related:                                                                    
//       VERIFY                                                                
//       FORBIDDEN                                                             
//       NEVER                                                                 
// Example:                                                                    
//       N/A |                                                                 
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_MUST(prop, rst)                                                  \
   assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_must(prop))            /* novas s-2050,s-2056 */      

`define ip2211ringpll_ASSUME_MUST(prop, clk, rst)                                             \
   assume property(p_must(prop, clk, rst))                                     

`endif                                                                         


`define ip2211ringpll_ASSERTC_MUST(name, prop, rst, ip2211ringpll_MSG)                                      \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_must(prop)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG       

`define ip2211ringpll_ASSUMEC_MUST(name, prop, rst, ip2211ringpll_MSG)                                      \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_must(prop)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG       



`define ip2211ringpll_ASSUMES_MUST(name, prop, clk, rst, ip2211ringpll_MSG)                                 \
   name: assume property(p_must(prop, clk, rst)) ip2211ringpll_MSG                           

`define ip2211ringpll_ASSERTS_MUST(name, prop, clk, rst, ip2211ringpll_MSG)                                 \
   name: assert property(p_must(prop, clk, rst)) ip2211ringpll_MSG                           


// ****************************************************************************************** //



// --- --- ---                                                                 



// ****************************************************************************************** //
// Name:   forbidden                                                           
// Category: Combinational                                                     
// Description:                                                                
//       Boolean condition 'cond' must never occur.                            
// Arguments:                                                                  
//       - cond    Boolean   The boolean condition that must never occur.      
// Comments:                                                                   
//       - The condition must be a boolean.                                    
//       - When the condition is boolean and clocked, ip2211ringpll_ASSERTS_FORBIDDEN is equivalent to
//       - ip2211ringpll_ASSERTS_NEVER.                                                      
//       - The difference between ip2211ringpll_ASSERTS_NEVER and ip2211ringpll_ASSERTS_FORBIDDEN is that with
//         ip2211ringpll_ASSERTS_FORBIDDEN the condition must be boolean, whereas with ip2211ringpll_ASSERTS_NEVER the
//         condition may also span over time (i.e. be sequential).             
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//       - The pass or failure of an immediate assertion inside an always_ff block would be
//         delayed by one sampling edge compared to when the assertion is in an always_comb or
//         in structural context.                                              
// Related:                                                                    
//       VERIFY                                                                
//       FORBIDDEN                                                             
//       NEVER                                                                 
// Example:                                                                    
//       N/A |                                                                 
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_FORBIDDEN(cond, rst)                                             \
   assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_forbidden(cond))       /* novas s-2050,s-2056 */      

`define ip2211ringpll_ASSUME_FORBIDDEN(cond, clk, rst)                                        \
   assume property(p_forbidden(cond, clk, rst))                                

`endif                                                                         


`define ip2211ringpll_ASSERTC_FORBIDDEN(name, cond, rst, ip2211ringpll_MSG)                                 \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_forbidden(cond)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG       

`define ip2211ringpll_ASSUMEC_FORBIDDEN(name, cond, rst, ip2211ringpll_MSG)                                 \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_forbidden(cond)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG   



`define ip2211ringpll_ASSUMES_FORBIDDEN(name, cond, clk, rst, ip2211ringpll_MSG)                            \
   name: assume property(p_forbidden(cond, clk, rst)) ip2211ringpll_MSG                      

`define ip2211ringpll_ASSERTS_FORBIDDEN(name, cond, clk, rst, ip2211ringpll_MSG)                            \
   name: assert property(p_forbidden(cond, clk, rst)) ip2211ringpll_MSG                      


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:   min                                                                 
// Category: Combinational                                                     
// Description:                                                                
//       The value of 'sig' must be no less than 'min_val'. It may be equal to 'min_val'.
// Arguments:                                                                  
//       - sig        Bit-vector  Signal to be monitored for its value to be no lower than
//                                'min_val'.                                   
//       - min_val    Number>=0   The minimum value that 'sig' can have.       
// Comments:                                                                   
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//       - The pass or failure of an immediate assertion inside an always_ff block would be
//         delayed by one sampling edge compared to when the assertion is in an always_comb or
//         in structural context.                                              
// Related:                                                                    
//       MAX                                                                   
//       RANGE                                                                 
//       ONE_OF                                                                
// Example:                                                                    
//       Valid port number is no less than 5 | @VIEW@(port, 5);                
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_MIN(sig, min_val, rst)                                           \
   assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_min_value(sig, min_val))       /* novas s-2050,s-2056 */

`define ip2211ringpll_ASSUME_MIN(sig, min_val, clk, rst)                                      \
   assume property(p_min_value(sig, min_val, clk, rst))                        

`define ip2211ringpll_COVER_MIN(sig, min_val, clk, rst)                                       \
   cover property(p_cover_min_value(sig, min_val, clk, rst))                   

`define ip2211ringpll_NOT_MIN_COVER(sig, min_val, clk, rst)                                   \
   cover property(p_not_min_value_cover(sig, min_val, clk, rst))               

`endif                                                                         


`define ip2211ringpll_ASSERTC_MIN(name, sig, min_val, rst, ip2211ringpll_MSG)                               \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_min_value(sig, min_val)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG

`define ip2211ringpll_ASSUMEC_MIN(name, sig, min_val, rst, ip2211ringpll_MSG)                               \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_min_value(sig, min_val)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG



`define ip2211ringpll_ASSUMES_MIN(name, sig, min_val, clk, rst, ip2211ringpll_MSG)                          \
   name: assume property(p_min_value(sig, min_val, clk, rst)) ip2211ringpll_MSG              

`define ip2211ringpll_ASSERTS_MIN(name, sig, min_val, clk, rst, ip2211ringpll_MSG)                          \
   name: assert property(p_min_value(sig, min_val, clk, rst)) ip2211ringpll_MSG              



`define ip2211ringpll_COVERS_MIN(name, sig, min_val, clk, rst, ip2211ringpll_MSG)                           \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_cover_min_value(sig, min_val, clk, rst)) ip2211ringpll_MSG      \
   `endif

`define ip2211ringpll_COVERC_MIN(name, sig, min_val, rst, ip2211ringpll_MSG)                                \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL ((!(rst) && `ip2211ringpll_l_min_value(sig, min_val))) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif



`define ip2211ringpll_NOT_MIN_COVERS(name ,sig, min_val, clk, rst, ip2211ringpll_MSG)                       \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_not_min_value_cover(sig, min_val, clk, rst)) ip2211ringpll_MSG  \
   `endif

`define ip2211ringpll_NOT_MIN_COVERC(name, sig, min_val, rst, ip2211ringpll_MSG)                            \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && `ip2211ringpll_l_min_value(sig, min_val)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:   max                                                                 
// Category: Combinational                                                     
// Description:                                                                
//       The value of 'sig' must be no greater than 'max_val'. It may be equal to 'max_val'.
// Arguments:                                                                  
//       - sig        Bit-vector   Signal to be monitored for its value to be no greater than
//                                 'max_val'.                                  
//       - max_val    Number>=0    The maximum value that 'sig' can have.      
// Comments:                                                                   
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//       - The pass or failure of an immediate assertion inside an always_ff block would be delayed
//         by one sampling edge compared to when the assertion is in an always_comb or in structural
//         context.                                                            
// Related:                                                                    
//       MIN                                                                   
//       RANGE                                                                 
//       ONE_OF                                                                
// Example:                                                                    
//       Valid port number is no more than 5 | @VIEW@(port, 5);                
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_MAX(sig, max_val, rst)                                           \
   assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_max_value(sig, max_val))       /* novas s-2050,s-2056 */

`define ip2211ringpll_ASSUME_MAX(sig, max_val, clk, rst)                                      \
   assume property(p_max_value(sig, max_val, clk, rst))                        

`define ip2211ringpll_COVER_MAX(sig, max_val, clk, rst)                                       \
   cover property(p_cover_max_value(sig, max_val, clk, rst))                   

`define ip2211ringpll_NOT_MAX_COVER(sig, max_val, clk, rst)                                   \
   cover property(p_not_max_value_cover(sig, max_val, clk, rst))               

`endif                                                                         


`define ip2211ringpll_ASSERTC_MAX(name, sig, max_val, rst, ip2211ringpll_MSG)                               \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_max_value(sig, max_val)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG

`define ip2211ringpll_ASSUMEC_MAX(name, sig, max_val, rst, ip2211ringpll_MSG)                               \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_max_value(sig, max_val)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG



`define ip2211ringpll_ASSUMES_MAX(name, sig, max_val, clk, rst, ip2211ringpll_MSG)                          \
   name: assume property(p_max_value(sig, max_val, clk, rst)) ip2211ringpll_MSG              

`define ip2211ringpll_ASSERTS_MAX(name, sig, max_val, clk, rst, ip2211ringpll_MSG)                          \
   name: assert property(p_max_value(sig, max_val, clk, rst)) ip2211ringpll_MSG              



`define ip2211ringpll_COVERS_MAX(name, sig, max_val, clk, rst, ip2211ringpll_MSG)                           \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_cover_max_value(sig, max_val, clk, rst)) ip2211ringpll_MSG      \
   `endif

`define ip2211ringpll_COVERC_MAX(name, sig, max_val, rst, ip2211ringpll_MSG)                                \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL ((!(rst) && `ip2211ringpll_l_max_value(sig, max_val))) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif



`define ip2211ringpll_NOT_MAX_COVERS(name ,sig, max_val, clk, rst, ip2211ringpll_MSG)                       \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_not_max_value_cover(sig, max_val, clk, rst)) ip2211ringpll_MSG  \
   `endif

`define ip2211ringpll_NOT_MAX_COVERC(name, sig, max_val, rst, ip2211ringpll_MSG)                            \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && `ip2211ringpll_l_max_value(sig, max_val)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:   at most bits low                                                    
// Category: Combinational                                                     
// Description:                                                                
//       At most 'n' bits in 'sig' are low. x and z values are counted as low for this calculation.
// Arguments:                                                                  
//       - sig   Bit-vector    At most 'n' bits in 'sig' can be low. Limitation: 'sig' must be a
//                             packed array.                                   
//       - n     Number>=0     The maximum number of bits in 'sig' that are allowed to be low.
// Comments:                                                                   
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//       - The pass or failure of an immediate assertion inside an always_ff block would be delayed
//         by one sampling edge compared to when the assertion is in an always_comb or in structural
//         context.                                                            
// Related:                                                                    
//       AT_MOST_BITS_HIGH                                                     
//       BITS_LOW                                                              
// Example:                                                                    
//       The following will fail | @VIEW@(001x, 3);                            
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_AT_MOST_BITS_LOW(sig, n, rst)                                    \
   assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_at_most_bits_low(sig, n))      /* novas s-2050,s-2056 */

`define ip2211ringpll_ASSUME_AT_MOST_BITS_LOW(sig, n, clk, rst)                               \
   assume property(p_at_most_bits_low(sig, n, clk, rst))                       

`define ip2211ringpll_COVER_AT_MOST_BITS_LOW(sig, n, clk, rst)                                \
   cover property(p_cover_at_most_bits_low(sig, n, clk, rst))                  

`define ip2211ringpll_NOT_AT_MOST_BITS_LOW_COVER(sig, n, clk, rst)                            \
   cover property(p_not_at_most_bits_low_cover(sig, n, clk, rst))              

`endif                                                                         



`define ip2211ringpll_ASSERTC_AT_MOST_BITS_LOW(name, sig, n, rst, ip2211ringpll_MSG)                        \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_at_most_bits_low(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG

`define ip2211ringpll_ASSUMEC_AT_MOST_BITS_LOW(name, sig, n, rst, ip2211ringpll_MSG)                        \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_at_most_bits_low(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG



`define ip2211ringpll_ASSUMES_AT_MOST_BITS_LOW(name, sig, n, clk, rst, ip2211ringpll_MSG)                   \
   name: assume property(p_at_most_bits_low(sig, n, clk, rst)) ip2211ringpll_MSG             

`define ip2211ringpll_ASSERTS_AT_MOST_BITS_LOW(name, sig, n, clk, rst, ip2211ringpll_MSG)                   \
   name: assert property(p_at_most_bits_low(sig, n, clk, rst)) ip2211ringpll_MSG             



`define ip2211ringpll_COVERS_AT_MOST_BITS_LOW(name, sig, n, clk, rst, ip2211ringpll_MSG)                    \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_cover_at_most_bits_low(sig, n, clk, rst)) ip2211ringpll_MSG     \
   `endif

`define ip2211ringpll_COVERC_AT_MOST_BITS_LOW(name, sig, n, rst, ip2211ringpll_MSG)                         \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && `ip2211ringpll_l_at_most_bits_low(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif



`define ip2211ringpll_NOT_AT_MOST_BITS_LOW_COVERS(name, sig, n, clk, rst, ip2211ringpll_MSG)                \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_not_at_most_bits_low_cover(sig, n, clk, rst)) ip2211ringpll_MSG \
   `endif

`define ip2211ringpll_NOT_AT_MOST_BITS_LOW_COVERC(name ,sig, n, rst, ip2211ringpll_MSG)                     \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && ! `ip2211ringpll_l_at_most_bits_low(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:   bits low                                                            
// Category: Combinational                                                     
// Description:                                                                
//       Exactly 'n' bits of 'sig' are low, other bits are high, and there are no x or z
//       values in 'sig'.                                                      
// Arguments:                                                                  
//       - sig   Bit-vector   Exactly 'n' bits in 'sig' are low.               
//       - n     Number>=0    The number of bits in 'sig' that are low.        
// Comments:                                                                   
//       - ASSERTC view This is an immediate checker and can be used anywhere including functions.
//       - ASSUMES view This is temporal and recommended for formal verification users.
//       - The pass or failure of an immediate assertion inside an always_ff block would be
//         delayed by one sampling edge compared to when the assertion is in an always_comb or
//         in structural context.                                              
// Related:                                                                    
//       AT_MOST_BITS_LOW                                                      
//       BITS_HIGH                                                             
//       REMAIN_LOW                                                            
// Example:                                                                    
//       The following will fail | @VIEW@(001x, 2);                            
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_BITS_LOW(sig, n, rst)                                            \
   assert `ip2211ringpll_FINAL (( (|(rst)) | `ip2211ringpll_l_bits_low(sig, n)))      /* novas s-2050,s-2056 */   

`define ip2211ringpll_ASSUME_BITS_LOW(sig, n, clk, rst)                                       \
   assume property(p_bits_low(sig, n, clk, rst))                               

`define ip2211ringpll_COVER_BITS_LOW(sig, n, clk, rst)                                        \
   cover property(p_cover_bits_low(sig, n, clk, rst))                          

`define ip2211ringpll_NOT_BITS_LOW_COVER(sig, n, clk, rst)                                    \
   cover property(p_not_bits_low_cover(sig, n, clk, rst))                      

`endif                                                                         



`define ip2211ringpll_ASSERTC_BITS_LOW(name, sig, n, rst, ip2211ringpll_MSG)                                \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_bits_low(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG 

`define ip2211ringpll_ASSUMEC_BITS_LOW(name, sig, n, rst, ip2211ringpll_MSG)                                \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_bits_low(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG 



`define ip2211ringpll_ASSUMES_BITS_LOW(name, sig, n, clk, rst, ip2211ringpll_MSG)                           \
   name: assume property(p_bits_low(sig, n, clk, rst)) ip2211ringpll_MSG                     

`define ip2211ringpll_ASSERTS_BITS_LOW(name, sig, n, clk, rst, ip2211ringpll_MSG)                           \
   name: assert property(p_bits_low(sig, n, clk, rst)) ip2211ringpll_MSG                     



`define ip2211ringpll_COVERS_BITS_LOW(name, sig, n, clk, rst, ip2211ringpll_MSG)                            \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_cover_bits_low(sig, n, clk, rst)) ip2211ringpll_MSG             \
   `endif

`define ip2211ringpll_COVERC_BITS_LOW(name, sig, n, rst, ip2211ringpll_MSG)                                 \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && `ip2211ringpll_l_bits_low(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif



`define ip2211ringpll_NOT_BITS_LOW_COVERS(name, sig, n, clk, rst, ip2211ringpll_MSG)                        \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_not_bits_low_cover(sig, n, clk, rst)) ip2211ringpll_MSG         \
   `endif

`define ip2211ringpll_NOT_BITS_LOW_COVERC(name ,sig, n, rst, ip2211ringpll_MSG)                             \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover `ip2211ringpll_FINAL (!(rst) && ! `ip2211ringpll_l_bits_low(sig, n)) /* novas s-2050,s-2056 */ ip2211ringpll_MSG \
   `endif


// ****************************************************************************************** //


// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  cover                                                                
// Category: Cover                                                             
// Description:                                                                
//      Cover a sequence.                                                      
// Arguments:                                                                  
//      - seq  Sequence   Sequence to be covered.                              
// Comments:                                                                   
//      None.                                                                  
// Related:                                                                    
//      None                                                                   
// Example:                                                                    
//      TBD |                                                                  
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                     

`define ip2211ringpll_COVER(seq, clk, rst)                                                    \
   cover property(p_cover(seq, clk, rst))                                      

`endif                                                                         


`define ip2211ringpll_COVERS(name, prop, clk, rst, ip2211ringpll_MSG)                                        \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
       typedef bit t_``name                                                     \
   `else                                                                        \
       name: cover property(p_cover(prop, clk, rst)) ip2211ringpll_MSG                        \
   `endif


`define ip2211ringpll_COVERS_ENABLE(name, en, prop, clk, rst, ip2211ringpll_MSG)                            \
   `ifndef INTC_SVA_LIB_COVER_ENABLE                                                 \
      typedef bit t_``name                                                      \
   `else                                                                        \
      name: cover property(p_cover_enable(en, prop, clk, rst)) ip2211ringpll_MSG              \
   `endif




// ****************************************************************************************** //                                                                              

// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:   fire                                                                
// Category: Combinational                                                     
// Description:                                                                
//       Fire an error message whenever reached.                               
// Arguments:                                                                  
//       - sig    Bit-vector   At most one bit of <sig> is high. Limitation: 'sig' must be a
//                           packed array                                      
// Comments:                                                                   
//       - This checker has generic arguments only. It is only used to fire error messages.
//       - This template is mainly useful in default clauses of case statements.
// Related:                                                                    
//       None                                                                  
// Code sample:                                                                
//       always_comb                                                           
//         unique casex (1'b1)                                                 
//           iq_4flight_CM105H[0] : iq_instflight_CM105H[0] = 3'b100;          
//           iq_3flight_CM105H[0] : iq_instflight_CM105H[0] = 3'b011;          
//         default :                                                           
//           iq_instflight_CM105H[0] = 3'b000;                                 
//           `ip2211ringpll_ASSERTC_FIRE(R_IFU_iq_instflight, `ip2211ringpll_ERR_MSG("error in sva1"));    
//       endcase                                                               
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_FIRE                                                             \
   assert `ip2211ringpll_FINAL (1'b0)                                                        

`endif                                                                         


`define ip2211ringpll_ASSERTC_FIRE(name, ip2211ringpll_MSG)                                                 \
   name: assert `ip2211ringpll_FINAL (1'b0) ip2211ringpll_MSG                                              


// ****************************************************************************************** //





// --- --- --- Concurent Templates --- --- --- //                              


// ****************************************************************************************** //
// Name:  trigger                                                              
// Category: Antecedent/Consequence                                            
// Description:                                                                
//       When 'trig' occurs, 'prop' should occur.                              
// Arguments:                                                                  
//      - trig    Sequence   Triggering event. Checking begins each time the sequence 'trig' is
//                           matched. In the special case where the sequence is a Boolean, each
//                           time the Boolean is high.                         
//      - prop    Property   Property to be satisfied.                         
// Comments:                                                                   
//      - If sequence 'trig' occurs, then property 'prop' must hold at the completion of that
//        sequence. Can also be used for simple Boolean implication, i.e. if Boolean 'b1' holds,
//        then Boolean 'b2' holds as well.                                     
// Related:                                                                    
//      DELAYED_TRIGGER                                                        
//      RECUR_TRIGGERS                                                         
// Code sample:                                                                
//      sequence e;                                                            
//        sig1 ##1 !sig1 ##1 sig1;                                             
//      endsequence                                                            
//      sequence form;                                                         
//        sig2 ##1 !sig2 ##1 sig2[*2];                                         
//      endsequence                                                            
//      `ip2211ringpll_ASSERTS_TRIGGER(trigger_edge_clk, e, form, posedge clk, rst, `ip2211ringpll_ERR_MSG("Error!"));
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_TRIGGER(trig, prop, clk, rst)                                    \
   assert property(p_trigger(trig, prop, clk, rst))                            

`define ip2211ringpll_ASSUME_TRIGGER(trig, prop, clk, rst)                                    \
   assume property(p_trigger(trig, prop, clk, rst))                            

`endif                                                                         

`define ip2211ringpll_ASSERTC_TRIGGER(name, trig, sig, rst, ip2211ringpll_MSG)                              \
   name: assert `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_trigger(trig, sig))  /* novas s-2050 */  ip2211ringpll_MSG

`define ip2211ringpll_ASSERTS_TRIGGER(name, trig, prop, clk, rst, ip2211ringpll_MSG)                        \
   name: assert property(p_trigger(trig, prop, clk, rst)) ip2211ringpll_MSG                  

`define ip2211ringpll_ASSUMEC_TRIGGER(name, trig, sig, rst, ip2211ringpll_MSG)                         \
   name: assume `ip2211ringpll_FINAL ((|(rst)) | `ip2211ringpll_l_trigger(trig, sig))  /* novas s-2050 */  ip2211ringpll_MSG

`define ip2211ringpll_ASSUMES_TRIGGER(name, trig, prop, clk, rst, ip2211ringpll_MSG)                        \
   name: assume property(p_trigger(trig, prop, clk, rst)) ip2211ringpll_MSG                  


// ****************************************************************************************** //



// --- --- ---                                                                 



// ****************************************************************************************** //
// Name:  delayed trigger                                                      
// Category: Antecedent/Consequence                                            
// Description:                                                                
//      When 'trig' occurs, 'prop' should occur 'delay' clock ticks after the completion of
//      'trig'.                                                                
// Arguments:                                                                  
//      - trig    Sequence     Triggering event. Checking begins each time the sequence
//                             'trig' is matched. In the special case where the sequence is
//                             a Boolean, each time the Boolean is high.       
//      - delay   Number>0     Delay in clock ticks after the completion of 'trig'.
//      - prop    Property     The property that should occur.                 
// Comments:                                                                   
//      - This template no longer supports a delay of 0. To achieve this purpose, use TRIGGER.
//      - This template is expensive for a large 'delay'.                      
//      - If sequence 'trig' is satisfied, then property 'prop' must be satisfied 'delay' clock
//        ticks after the completion of 'trig'. Can also be used for simple Boolean implication,
//        i.e. if Boolean 'b1' holds, then after 'delay' clock ticks Boolean 'b2' holds as well.
// Related:                                                                    
//      TRIGGER                                                                
//      RECUR_TRIGGERS                                                         
// Code sample:                                                                
//      sequence e;                                                            
//        sig1 ##1 !sig1 ##1 sig1;                                             
//      endsequence                                                            
//      sequence form;                                                         
//        sig2 ##1 !sig2 ##1 sig2[*2];                                         
//      endsequence                                                            
//      `ip2211ringpll_ASSERTS_DELAYED_TRIGGER(delayed_name, e, 2, form, posedge clk, rst, `ip2211ringpll_ERR_MSG("Error"));
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_DELAYED_TRIGGER(trig, delay, prop, clk, rst)                     \
   assert property(p_delayed_trigger(trig, delay, prop, clk, rst))             

`define ip2211ringpll_ASSUME_DELAYED_TRIGGER(trig, delay, prop, clk, rst)                     \
   assume property(p_delayed_trigger(trig, delay, prop, clk, rst))             

`endif                                                                         

`define ip2211ringpll_ASSERTS_DELAYED_TRIGGER(name, trig, delay, prop, clk, rst, ip2211ringpll_MSG)         \
   name: assert property(p_delayed_trigger(trig, delay, prop, clk, rst)) ip2211ringpll_MSG   

`define ip2211ringpll_ASSUMES_DELAYED_TRIGGER(name, trig, delay, prop, clk, rst, ip2211ringpll_MSG)         \
   name: assume property(p_delayed_trigger(trig, delay, prop, clk, rst)) ip2211ringpll_MSG   


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  never                                                                
// Category: Data Checking                                                     
// Description:                                                                
//      The property 'prop' never occurs.                                      
// Arguments:                                                                  
//      - prop    Property  The property that should never occur.              
// Comments:                                                                   
//      - When the condition is boolean and clocked, ip2211ringpll_ASSERTS_FORBIDDEN is equivalent to 
//        ip2211ringpll_ASSERTS_NEVER. The difference between ip2211ringpll_ASSERTS_NEVER and ip2211ringpll_ASSERTS_FORBIDDEN is that with
//        ip2211ringpll_ASSERTS_FORBIDDEN the condition must be boolean, whereas with ip2211ringpll_ASSERTS_NEVER the 
//        condition may also span over time (i.e. be sequential).              
// Related:                                                                    
//      FORBIDDEN                                                              
//      MUST                                                                   
//      VERIFY                                                                 
// Example:                                                                    
//      N/A |                                                                  
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_NEVER(prop, clk, rst)                                            \
   assert property(p_never(prop, clk, rst))                                    

`define ip2211ringpll_ASSUME_NEVER(prop, clk, rst)                                            \
   assume property(p_never(prop, clk, rst))                                    

`endif                                                                         

`define ip2211ringpll_ASSERTS_NEVER(name, prop, clk, rst, ip2211ringpll_MSG)                                \
   name: assert property(p_never(prop, clk, rst)) ip2211ringpll_MSG                          

`define ip2211ringpll_ASSUMES_NEVER(name, prop, clk, rst, ip2211ringpll_MSG)                                \
   name: assume property(p_never(prop, clk, rst)) ip2211ringpll_MSG                          


// ****************************************************************************************** //



// --- --- ---                                                                 



// ****************************************************************************************** //
// Name:  eventually holds                                                     
// Category: Data Checking                                                     
// Description:                                                                
//      Once the enable 'en' is high, 'prop' should eventually hold (strong eventually relation).
//      There is no time bound.                                                
//      Thus, the property is violated if 'prop' never holds or if the clock stops ticking.
// Arguments:                                                                  
//      - en    Sequence   Enabling event. Checking begins each time the sequence 'en' is matched.
//                         In the special case where the sequence is a Boolean, each time the
//                         Boolean is high.                                    
//      - prop  Property   Property that should eventually hold.               
// Comments:                                                                   
//      - ip2211ringpll_ASSERT_EVENTUALLY_HOLDS is only useful for formal verification.      
// Related:                                                                    
//      NEXT_EVENT                                                             
//      REQ_GRANTED                                                            
//      UNTIL_STRONG                                                           
// Example:                                                                    
//      TBD |                                                                  
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_EVENTUALLY_HOLDS(en, prop, clk, rst)                             \
   assert property(p_eventually_holds(en, prop, clk, rst))                     

`define ip2211ringpll_ASSUME_EVENTUALLY_HOLDS(en, prop, clk, rst)                             \
   assume property(p_eventually_holds(en, prop, clk, rst))                     

`endif                                                                         

`define ip2211ringpll_ASSERTS_EVENTUALLY_HOLDS(name, en, prop, clk, rst, ip2211ringpll_MSG)                 \
   name: assert property(p_eventually_holds(en, prop, clk, rst)) ip2211ringpll_MSG           

`define ip2211ringpll_ASSUMES_EVENTUALLY_HOLDS(name, en, prop, clk, rst, ip2211ringpll_MSG)                 \
   name: assume property(p_eventually_holds(en, prop, clk, rst)) ip2211ringpll_MSG           


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  between                                                              
// Category: Stability , Events                                                
// Description:                                                                
//      'cond' holds at every sampling point between the two events 'start_ev' and 'end_ev'
//      inclusive. The end event may never occur, in which case 'cond' continues to hold forever.
// Arguments:                                                                  
//      - start_ev    Sequence   Start checking event. Checking begins each time the sequence
//                               'start_ev' is matched. In the special case where the sequence
//                               is a Boolean, each time the Boolean is high.  
//      - end_ev      Property   End event is when 'end_ev' is true.           
//      - cond        Property   A property that must be true between 'start_ev' and 'end_ev'.
// Comments:                                                                   
//      None.                                                                  
// Related:                                                                    
//      BETWEEN_TIME                                                           
//      BEFORE_EVENT                                                           
//      NEXT_EVENT                                                             
// Code sample:                                                                
//      sequence e;                                                            
//        sig1 ##1 !sig1 ##1 sig1;                                             
//      endsequence                                                            
//      `ip2211ringpll_ASSERTS_BETWEEN(between_posedge_clk, e, end_b, cond, posedge clk, rst, `ip2211ringpll_ERR_MSG("Bad"));
// Example:                                                                    
//      Success (start-time:195 and end-time:235) | | images/BETWEEN_1.png     
// Example:                                                                    
//      Failure (start-time:135 and end-time:175) | | images/BETWEEN_2.png     
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_BETWEEN(start_ev, end_ev, cond, clk, rst)                        \
   assert property(p_between(start_ev, end_ev, cond, clk, rst))                

`define ip2211ringpll_ASSUME_BETWEEN(start_ev, end_ev, cond, clk, rst)                        \
   assume property(p_between(start_ev, end_ev, cond, clk, rst))                

`endif                                                                         

`define ip2211ringpll_ASSERTS_BETWEEN(name, start_ev, end_ev, cond, clk, rst, ip2211ringpll_MSG)            \
   name: assert property(p_between(start_ev, end_ev, cond, clk, rst)) ip2211ringpll_MSG      

`define ip2211ringpll_ASSUMES_BETWEEN(name, start_ev, end_ev, cond, clk, rst, ip2211ringpll_MSG)            \
   name: assume property(p_between(start_ev, end_ev, cond, clk, rst)) ip2211ringpll_MSG      


// ****************************************************************************************** //



// --- --- ---                                                                 

// ****************************************************************************************** //
// Name:   between time                                                        
// Category: Stability , Events                                                
// Description:                                                                
//       After the triggering event 'trig', 'cond' holds continuously starting at time
//       'start_time' until time 'end_time' (inclusive). Start time 0 is at the last tick
//       of the event 'trig' (or simply at 'trig' if it is a Boolean). Start time 1 is a tick
//       after 'trig' etc. There are no restrictions on 'cond' outside the [start_time, end_time]
//       interval.                                                             
// Arguments:                                                                  
//      - trig        Sequence   Triggering event. Checking begins each time the sequence 'trig'
//                               is matched. In the special case where the sequence is a Boolean,
//                               each time the Boolean is high.                
//      - start_time  Number>=0  Starting time greater than or equal to zero.  
//      - end_time    Number>=0  Ending time greater than or equal to 'start_time'.
//      - cond        Property   A property that must true between 'start_time' and 'end_time'.
// Comments:                                                                   
//      - This template is expensive for large start or end times. Use BETWEEN if possible.
// Related:                                                                    
//      BETWEEN                                                                
//      BEFORE_EVENT                                                           
//      NEXT_EVENT                                                             
// Example:                                                                    
//       | | images/BETWEEN_TIME_1.png                                         
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_BETWEEN_TIME(trig, start_time, end_time, cond, clk, rst)         \
   assert property(p_between_time(trig, start_time, end_time, cond, clk, rst)) 

`define ip2211ringpll_ASSUME_BETWEEN_TIME(trig, start_time, end_time, cond, clk, rst)         \
   assume property(p_between_time(trig, start_time, end_time, cond, clk, rst)) 

`endif                                                                         

`define ip2211ringpll_ASSERTS_BETWEEN_TIME(name, trig, start_time, end_time, cond, clk, rst, ip2211ringpll_MSG) \
   name: assert property(p_between_time(trig, start_time, end_time, cond, clk, rst)) ip2211ringpll_MSG

`define ip2211ringpll_ASSUMES_BETWEEN_TIME(name, trig, start_time, end_time, cond, clk, rst, ip2211ringpll_MSG) \
   name: assume property(p_between_time(trig, start_time, end_time, cond, clk, rst)) ip2211ringpll_MSG


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:   next event                                                          
// Category: Events                                                            
// Description:                                                                
//      If 'en' is high, then the next time that 'ev' holds, property 'prop' must hold as well.
//      'ev' and 'en' can hold simultaneously. 'ev' may never hold.            
// Arguments:                                                                  
//      - en      Boolean     Enabler.                                         
//      - ev      Boolean     Sampling event.                                  
//      - prop    Property    Property to be checked.                          
// Comments:                                                                   
//      - This template is expensive for large start or end times. Use BETWEEN if possible.
// Related:                                                                    
//      BEFORE_EVENT                                                           
//      BETWEEN                                                                
//      UNTIL_STRONG                                                           
// Example:                                                                    
//      TBD |                                                                  
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_NEXT_EVENT(en, ev, prop, clk, rst)                               \
   assert property(p_next_event(en, ev, prop, clk, rst))                       

`define ip2211ringpll_ASSUME_NEXT_EVENT(en, ev, prop, clk, rst)                               \
   assume property(p_next_event(en, ev, prop, clk, rst))                       

`endif                                                                         

`define ip2211ringpll_ASSERTS_NEXT_EVENT(name, en, ev, prop, clk, rst, ip2211ringpll_MSG)                   \
   name: assert property(p_next_event(en, ev, prop, clk, rst)) ip2211ringpll_MSG             

`define ip2211ringpll_ASSUMES_NEXT_EVENT(name, en, ev, prop, clk, rst, ip2211ringpll_MSG)                   \
   name: assume property(p_next_event(en, ev, prop, clk, rst)) ip2211ringpll_MSG             


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:   before event                                                        
// Category: Events                                                            
// Description:                                                                
//      Whenever 'en' holds, 'first' must hold before 'second'. The earliest 'second' can hold
//      is one cycle after 'first' holds. 'first' is not required to hold, in which case 'second'
//      should never hold.                                                     
// Arguments:                                                                  
//      - en       Sequence   Enabling sequence. Checking begins each time the sequence 'en' is
//                            matched. In the special case where the sequence is a Boolean, each
//                            time the Boolean is high.                        
//      - first    Property   Must be true before 'second' holds. 'first' and 'en' can hold
//                            simutaneously.                                   
//      - second   Property   Cannot hold before 'first' is true.              
// Comments:                                                                   
//      None.                                                                  
// Related:                                                                    
//      NEXT_EVENT                                                             
//      BETWEEN                                                                
//      BETWEEN TIME                                                           
//      UNTIL_STRONG                                                           
// Example:                                                                    
//      TBD |                                                                  
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_BEFORE_EVENT(en, first, second, clk, rst)                        \
   assert property(p_before_event(en, first, second, clk, rst))                

`define ip2211ringpll_ASSUME_BEFORE_EVENT(en, first, second, clk, rst)                        \
   assume property(p_before_event(en, first, second, clk, rst))                

`endif                                                                         

`define ip2211ringpll_ASSERTS_BEFORE_EVENT(name, en, first, second, clk, rst, ip2211ringpll_MSG)            \
   name: assert property(p_before_event(en, first, second, clk, rst)) ip2211ringpll_MSG      

`define ip2211ringpll_ASSUMES_BEFORE_EVENT(name, en, first, second, clk, rst, ip2211ringpll_MSG)            \
   name: assume property(p_before_event(en, first, second, clk, rst)) ip2211ringpll_MSG      


// ****************************************************************************************** //



// --- --- ---                                                                 



// ****************************************************************************************** //
// Name:  remain high                                                          
// Category: Stability                                                         
// Description:                                                                
//      Whenever 'sig' rises, it remains high for 'n' additional clocks. The number of clocks 
//      'n' does not include the clock at which 'sig' changed. 'sig' must be high at the 'n'th
//      tick point. Values of 'sig' are only sampled at the clock ticks. The behavior of 'sig'
//      between the clock ticks is not checked.                                
// Arguments:                                                                  
//      - sig  Bit-vector  Signal to be checked.                               
//      - n    Number>0    The minimum number of cycles thoughtout which 'sig' must remain high.
// Comments:                                                                   
//      - This checker is expensive for a large 'n'. In this case use STABLE if possible (if the
//        signal retains its value between events, rather than throughout a time interval).
// Related:                                                                    
//      GREMAIN_HIGH                                                           
//      REMAIN_LOW                                                             
//      GREMAIN_LOW                                                            
// Example:                                                                    
//      In the following example, both sig 1 and sig 2 pass. | | images/REMAIN_HIGH_1.png
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_REMAIN_HIGH(sig, n, clk, rst)                                    \
   assert property(p_remain_high(sig, n, clk, rst))                            

`define ip2211ringpll_ASSUME_REMAIN_HIGH(sig, n, clk, rst)                                    \
   assume property(p_remain_high(sig, n, clk, rst))                            

`endif                                                                         

`define ip2211ringpll_ASSERTS_REMAIN_HIGH(name, sig, n, clk, rst, ip2211ringpll_MSG)                        \
   name: assert property(p_remain_high(sig, n, clk, rst)) ip2211ringpll_MSG                  

`define ip2211ringpll_ASSUMES_REMAIN_HIGH(name, sig, n, clk, rst, ip2211ringpll_MSG)                        \
   name: assume property(p_remain_high(sig, n, clk, rst)) ip2211ringpll_MSG                  


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  gremain high                                                         
// Category: Stability                                                         
// Description:                                                                
//      Whenever 'sig' rises, it remains high for 'n' additional clocks. The number of clocks
//      'n' does not include the clock at which 'sig' changed. 'sig' must also be high at the
//      'n'th tick point. Values of 'sig' are only sampled at the clock ticks. However, 'sig
//      is required to be high at all times during the 'n' clock ticks, even at the non-tick
//      points of the clock.                                                   
// Arguments:                                                                  
//      - sig  Bit-vector   Signal to be checked.                              
//      - n    Number>0     The minimum number of cycles throughout which 'sig' must remain high.
// Comments:                                                                   
//      - This checker is expensive for a large 'n'. In such cases, use GSTABLE if possible
//        (if the signal retains its value between events, rather than throughout a time interval).
// Related:                                                                    
//      REMAIN_HIGH                                                            
//      REMAIN_LOW                                                             
//      GREMAIN_LOW                                                            
// Example:                                                                    
//      In the following example, sig 1 passes, while sig 2 fails. | | images/GREMAIN_HIGH_1.png
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_GREMAIN_HIGH(sig, n, clk, rst)                                   \
   assert property(p_gremain_high(sig, n, clk, rst))                           

`define ip2211ringpll_ASSUME_GREMAIN_HIGH(sig, n, clk, rst)                                   \
   assume property(p_gremain_high(sig, n, clk, rst))                           

`endif                                                                         

`define ip2211ringpll_ASSERTS_GREMAIN_HIGH(name, sig, n, clk, rst, ip2211ringpll_MSG)                       \
   name: assert property(p_gremain_high(sig, n, clk, rst)) ip2211ringpll_MSG                 

`define ip2211ringpll_ASSUMES_GREMAIN_HIGH(name, sig, n, clk, rst, ip2211ringpll_MSG)                       \
   name: assume property(p_gremain_high(sig, n, clk, rst)) ip2211ringpll_MSG                 


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  remain low                                                           
// Category: Stability                                                         
// Description:                                                                
//      Whenever 'sig' falls, it remains low for 'n' additional clocks. The number of clocks 'n'
//       does not include the clock at which 'sig' changed. 'sig' must be low at the 'n'th tick
//       point. Values of 'sig' are only sampled at the clock ticks. The behavior of 'sig'
//       between the clock ticks is not checked.                               
// Arguments:                                                                  
//       - sig   Bit-vector   Signal to be checked.                            
//       - n     Number>0     The minimum number of cycles thoughtout which 'sig' must remain low.
// Comments:                                                                   
//       - This checker is expensive for a large 'n'. In such cases, use STABLE if possible
//         (if the signal retains its value between events, rather than throughout a time interval).
// Related:                                                                    
//       GREMAIN_LOW                                                           
//       REMAIN_HIGH                                                           
//       GREMAIN_HIGH                                                          
// Example:                                                                    
//       In the following example, both sig 1 and sig 2 pass.| | images/REMAIN_LOW_1.png
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_REMAIN_LOW(sig, n, clk, rst)                                     \
   assert property(p_remain_high(!(sig), n, clk, rst))                         

`define ip2211ringpll_ASSUME_REMAIN_LOW(sig, n, clk, rst)                                     \
   assume property(p_remain_high(!(sig), n, clk, rst))                         

`endif                                                                         

`define ip2211ringpll_ASSERTS_REMAIN_LOW(name, sig, n, clk, rst, ip2211ringpll_MSG)                         \
   name: assert property(p_remain_high(!(sig), n, clk, rst)) ip2211ringpll_MSG               

`define ip2211ringpll_ASSUMES_REMAIN_LOW(name, sig, n, clk, rst, ip2211ringpll_MSG)                         \
   name: assume property(p_remain_high(!(sig), n, clk, rst)) ip2211ringpll_MSG               


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  gremain low                                                          
// Category: Stability                                                         
// Description:                                                                
//       Whenever 'sig' falls, it remains low for 'n' additional clocks. The number of clocks
//       'n' does not include the clock at which 'sig' changed. 'sig' must also be low at the
//       'n'th tick point. Values of 'sig' are only sampled at the clock ticks. However, 'sig'
//       is required to be low at all times during the 'n' clock ticks, even at the non-tick
//       points of the clock.                                                  
// Arguments:                                                                  
//       - sig   Bit-vector   Signal to be checked.                            
//       - n     Number>0     The minimum number of cycles thoughtout which 'sig' must remain low.
// Comments:                                                                   
//       - This checker is expensive for a large 'n'. In such cases, use GSTABLE if possible
//         (if the signal retains its value between events, rather than throughout a time interval).
// Related:                                                                    
//       REMAIN_LOW                                                            
//       REMAIN_HIGH                                                           
//       GREMAIN_HIGH                                                          
// Example:                                                                    
//       In the following example, sig 1 passes, while sig 2 fails. | | images/GREMAIN_LOW_1.png
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_GREMAIN_LOW(sig, n, clk, rst)                                    \
   assert property(p_gremain_high(!(sig), n, clk, rst))                        

`define ip2211ringpll_ASSUME_GREMAIN_LOW(sig, n, clk, rst)                                    \
   assume property(p_gremain_high(!(sig), n, clk, rst))                        

`endif                                                                         

`define ip2211ringpll_ASSERTS_GREMAIN_LOW(name, sig, n, clk, rst, ip2211ringpll_MSG)                        \
   name: assert property(p_gremain_high(!(sig), n, clk, rst)) ip2211ringpll_MSG              

`define ip2211ringpll_ASSUMES_GREMAIN_LOW(name, sig, n, clk, rst, ip2211ringpll_MSG)                        \
   name: assume property(p_gremain_high(!(sig), n, clk, rst)) ip2211ringpll_MSG              


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  remain_high_at_most                                                  
// Category: Stability                                                         
// Description:                                                                
//      Whenever 'sig' rises, it remains high for at most 'n' additional clocks. The number 
//      of clocks 'n' does not include the clock at which 'sig' changed. Values of 'sig' are
//      only sampled at the clock ticks.                                       
// Arguments:                                                                  
//      - sig  Bit-vector   Signal to be checked.                              
//      - n    Number>=0    The maximal number of cycles thoughtout which 'sig' is allowed 
//                          to remain high.                                    
// Comments:                                                                   
//       - This checker is expensive for a large 'n'. In such cases, use GSTABLE if possible
//         (if the signal retains its value between events, rather than throughout a time interval).
// Related:                                                                    
//       REMAIN_LOW                                                            
//       GREMAIN_HIGH                                                          
//       REMAIN_HIGH                                                           
//       GREMAIN_HIGH                                                          
//       GREMAIN_HIGH_AT_MOST                                                  
// Example:                                                                    
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_REMAIN_HIGH_AT_MOST(sig, n, clk, rst)                            \
   assert property(p_remain_high_at_most(sig, n, clk, rst))                    

`define ip2211ringpll_ASSUME_REMAIN_HIGH_AT_MOST(sig, n, clk, rst)                            \
   assume property(p_remain_high_at_most(sig, n, clk, rst))                    


`define ip2211ringpll_ASSERTS_REMAIN_HIGH_AT_MOST(name, sig, n, clk, rst, ip2211ringpll_MSG)                \
   name: assert property(p_remain_high_at_most(sig, n, clk, rst)) ip2211ringpll_MSG          

`define ip2211ringpll_ASSUMES_REMAIN_HIGH_AT_MOST(name, sig, n, clk, rst, ip2211ringpll_MSG)                \
   name: assume property(p_remain_high_at_most(sig, n, clk, rst)) ip2211ringpll_MSG          

`endif                                                                         

// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:   gremain_high_at_most                                                
// Category: Stability                                                         
// Description:                                                                
//       Whenever 'sig' rises, it remains high for at most 'n' additional clocks, that is 'sig'
//       should fall in no more than 'n' clocks. The number of clocks 'n' does not include the 
//       clock at which 'sig' changed.                                         
//       Values of 'sig' are also checked between the clock ticks.             
// Arguments:                                                                  
//      - sig  Bit-vector   Signal to be checked.                              
//      - n    Number>=0    The maximal number of cycles thoughtout which 'sig' is allowed 
//                          to remain high.                                    
// Comments:                                                                   
//      - This checker is expensive for a large 'n'. In such cases, use GSTABLE if possible
//        (if the signal retains its value between events, rather than throughout a time interval).
// Related:                                                                    
//       REMAIN_LOW                                                            
//       GREMAIN_HIGH                                                          
//       REMAIN_HIGH                                                           
//       GREMAIN_HIGH                                                          
//       REMAIN_HIGH_AT_MOST                                                   
// Example:                                                                    
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_GREMAIN_HIGH_AT_MOST(sig, n, clk, rst)                           \
   assert property(p_gremain_high_at_most(sig, n, clk, rst))                   

`define ip2211ringpll_ASSUME_GREMAIN_HIGH_AT_MOST(sig, n, clk, rst)                           \
   assume property(p_gremain_high_at_most(sig, n, clk, rst))                   

`endif                                                                         

`define ip2211ringpll_ASSERTS_GREMAIN_HIGH_AT_MOST(name, sig, n, clk, rst, ip2211ringpll_MSG)               \
   name: assert property(p_gremain_high_at_most(sig, n, clk, rst)) ip2211ringpll_MSG         

`define ip2211ringpll_ASSUMES_GREMAIN_HIGH_AT_MOST(name, sig, n, clk, rst, ip2211ringpll_MSG)               \
   name: assume property(p_gremain_high_at_most(sig, n, clk, rst)) ip2211ringpll_MSG         


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  verify                                                               
// Category: Data Checking                                                     
// Description:                                                                
//      The property 'prop' must always be true.                               
// Arguments:                                                                  
//      - prop    Property    The property that must always be true.           
// Comments:                                                                   
//      - When the condition is boolean and clocked, ip2211ringpll_ASSERTS_MUST is equivalent to ip2211ringpll_ASSERTS_VERIFY.
// Related:                                                                    
//      MUST                                                                   
//      FORBIDDEN                                                              
//      NEVER                                                                  
// Example:                                                                    
//      N/A |                                                                  
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_VERIFY(prop, clk, rst)                                           \
   assert property(p_verify(prop, clk, rst))                                   

`define ip2211ringpll_ASSUME_VERIFY(prop, clk, rst)                                           \
   assume property(p_verify(prop, clk, rst))                                   

`endif                                                                         

`define ip2211ringpll_ASSERTS_VERIFY(name, prop, clk, rst, ip2211ringpll_MSG)                               \
   name: assert property(p_verify(prop, clk, rst)) ip2211ringpll_MSG                         

`define ip2211ringpll_ASSUMES_VERIFY(name, prop, clk, rst, ip2211ringpll_MSG)                               \
   name: assume property(p_verify(prop, clk, rst)) ip2211ringpll_MSG                         


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  req granted                                                          
// Category: Antecedent/Consequence                                            
// Description:                                                                
//       A request is eventually granted. A request is registered when 'req' rises and there
//       is no pending request, or when there is a 'gnt' followed by 'req'. As long as the
//       request is not satisfied, no new requests can be registered.          
// Arguments:                                                                  
//       - req   Boolean   Request signal.                                     
//       - gnt   Boolean   Grant signal.                                       
// Comments:                                                                   
//       - The property passes if the grant holds at the same time the request is made.
//       - There is no explicit bound by which the request must be granted.    
// Related:                                                                    
//       CONT_REQ_GRANTED                                                      
//       REQ_GRANTED_WITHIN                                                    
// Code sample:                                                                
//       `ip2211ringpll_ASSERTS_REQ_GRANTED(req_granted_clk, req, gnt, posedge clk, rst, `ip2211ringpll_ERR_MSG("Error"));
// Example:                                                                    
//       success (start-time:51 and end-time:81) | | images/REQ_GRANTED_1.png  
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_REQ_GRANTED(req, gnt, clk, rst)                                  \
   assert property(p_req_granted(req, gnt, clk, rst))                          

`define ip2211ringpll_ASSUME_REQ_GRANTED(req, gnt, clk, rst)                                  \
   assume property(p_req_granted(req, gnt, clk, rst))                          

`endif                                                                         

`define ip2211ringpll_ASSERTS_REQ_GRANTED(name, req, gnt, clk, rst, ip2211ringpll_MSG)                      \
   name: assert property(p_req_granted(req, gnt, clk, rst)) ip2211ringpll_MSG                

`define ip2211ringpll_ASSUMES_REQ_GRANTED(name, req, gnt, clk, rst, ip2211ringpll_MSG)                      \
   name: assume property(p_req_granted(req, gnt, clk, rst)) ip2211ringpll_MSG                


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  cont req granted                                                     
// Category: Data Checking , Antecedent/Consequence                            
// Description:                                                                
//       A continuous request is eventually granted. A request is registered when 'req' rises
//       and there is no pending request, or when there is a 'gnt' followed by 'req'. 'req'
//       should remain high as long as the request is not satisfied.           
// Arguments:                                                                  
//       - req  Boolean     Request signal.                                    
//       - gnt  Boolean     Grant signal.                                      
// Comments:                                                                   
//       - The property passes if the grant holds at the same time the request is made.
//       - There is no explicit bound by which the request must be granted.    
// Related:                                                                    
//       REQ_GRANTED                                                           
//       REQ_GRANTED_WITHIN                                                    
// Code sample:                                                                
//       `ip2211ringpll_ASSERTS_CONT_REQ_GRANTED(cont_req_granted, req, gnt, clk, rst, `ip2211ringpll_ERR_MSG("Error"));
// Example:                                                                    
//       failure (start-time:75 and end-time:111) | | images/CONT_REQ_GRANTED_1.png
// Example:                                                                    
//       success (start-time:27 and end-time:63) | | images/CONT_REQ_GRANTED_2.png
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_CONT_REQ_GRANTED(req, gnt, clk, rst)                             \
   assert property(p_cont_req_granted(req, gnt, clk, rst))                     

`define ip2211ringpll_ASSUME_CONT_REQ_GRANTED(req, gnt, clk, rst)                             \
   assume property(p_cont_req_granted(req, gnt, clk, rst))                     

`endif                                                                         

`define ip2211ringpll_ASSERTS_CONT_REQ_GRANTED(name, req, gnt, clk, rst, ip2211ringpll_MSG)                 \
   name: assert property(p_cont_req_granted(req, gnt, clk, rst)) ip2211ringpll_MSG           

`define ip2211ringpll_ASSUMES_CONT_REQ_GRANTED(name, req, gnt, clk, rst, ip2211ringpll_MSG)                 \
   name: assume property(p_cont_req_granted(req, gnt, clk, rst)) ip2211ringpll_MSG           


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  req granted within                                                   
// Category: Antecedent/Consequence                                            
// Description:                                                                
//       A request is granted at some sampling point between (and including) the m-th and n-th
//       sampling points after the current point. A single grant may satisfy more than one
//       request, as long as for each request the grant occurs within the m to n interval with
//       respect to that request.                                              
// Arguments:                                                                  
//       - req  Boolean     Request signal.                                    
//       - m    Number>=0   Starting sampling point.                           
//       - n    Number>0    Ending sampling point.                             
//       - gnt  Boolean     Grant signal.                                      
// Comments:                                                                   
//       - The request does not need to remain pending until it is granted.    
//       - This template is expensive for large 'm's or 'n's. Use REQ_GRANTED if possible.
// Related:                                                                    
//       REQ_GRANTED                                                           
//       CONT_REQ_GRANTED                                                      
// Code sample:                                                                
//       `ip2211ringpll_ASSERTS_REQ_GRANTED_WITHIN(reg_granted_within_check, req, 3, 6, gnt, clk, rst, `ip2211ringpll_ERR_MSG(""));
// Example:                                                                    
//       failure (start-time:33 and end-time:51) | | images/REQ_GRANTED_WITHIN_1.png
// Example:                                                                    
//       success (start-time:63 and end-time:87) | | images/REQ_GRANTED_WITHIN_2.png
// Example:                                                                    
//       failure (start-time:219 and end-time:261) | | images/REQ_GRANTED_WITHIN_3.png
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_REQ_GRANTED_WITHIN(req, min, max, gnt, clk, rst)                 \
   assert property(p_req_granted_within(req, min, max, gnt, clk, rst))         

`define ip2211ringpll_ASSUME_REQ_GRANTED_WITHIN(req, min, max, gnt, clk, rst)                 \
   assume property(p_req_granted_within(req, min, max, gnt, clk, rst))         

`endif                                                                         

`define ip2211ringpll_ASSERTS_REQ_GRANTED_WITHIN(name, req, min, max, gnt, clk, rst, ip2211ringpll_MSG)     \
   name: assert property(p_req_granted_within(req, min, max, gnt, clk, rst)) ip2211ringpll_MSG

`define ip2211ringpll_ASSUMES_REQ_GRANTED_WITHIN(name, req, min, max, gnt, clk, rst, ip2211ringpll_MSG)     \
   name: assume property(p_req_granted_within(req, min, max, gnt, clk, rst)) ip2211ringpll_MSG


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  until strong                                                         
// Category: Stability                                                         
// Description:                                                                
//       Whenever 'start_ev' is high, 'cond' must hold until 'end_ev' holds. 'end_ev' must
//       eventually hold. 'cond' is not required to hold at the time 'end_ev' holds.
// Arguments:                                                                  
//       - start_ev    Sequence   Enabling event. Occurs each time the sequence 'start_ev' is
//                                matched. In the special case where the sequence is a Boolean,
//                                each time the Boolean is high.               
//       - cond        Property   A property that must hold until 'end_ev' holds.
//       - end_ev      Property   End event is when the property 'end_ev' is true.
// Comments:                                                                   
//       - The property passes if 'end_ev' holds at the same time as 'start_ev'.
//       - There is no explicit bound by which 'end_ev' must occur.            
// Related:                                                                    
//       NEXT_EVENT                                                            
//       REQ_GRANTED                                                           
//       BETWEEN                                                               
//       UNTIL_WEAK                                                            
// Code sample:                                                                
//       `ip2211ringpll_ASSERTS_UNTIL_STRONG(until_strong_clk, start_bool, sig==8'h10, end_bool, posedge clk, rst, `ip2211ringpll_ERR_MSG(""));
// Example:                                                                    
//       success (start-time:33 and end-time:51) | | images/UNTIL_STRONG_1.png 
// Example:                                                                    
//       failure (start-time:201 and end-time:213) | | images/UNTIL_STRONG_2.png
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_UNTIL_STRONG(start_ev, cond, end_ev, clk, rst)                   \
   assert property(p_until_strong(start_ev, cond, end_ev, clk, rst))           

`define ip2211ringpll_ASSUME_UNTIL_STRONG(start_ev, cond, end_ev, clk, rst)                   \
   assume property(p_until_strong(start_ev, cond, end_ev, clk, rst))           

`endif                                                                         

`define ip2211ringpll_ASSERTS_UNTIL_STRONG(name, start_ev, cond, end_ev, clk, rst, ip2211ringpll_MSG)       \
   name: assert property(p_until_strong(start_ev, cond, end_ev, clk, rst)) ip2211ringpll_MSG 

`define ip2211ringpll_ASSUMES_UNTIL_STRONG(name, start_ev, cond, end_ev, clk, rst, ip2211ringpll_MSG)       \
   name: assume property(p_until_strong(start_ev, cond, end_ev, clk, rst)) ip2211ringpll_MSG 


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:   until weak                                                          
// Category: Stability                                                         
// Description:                                                                
//       Whenever 'start_ev' is high, formula 'cond' must hold until 'end_ev' holds.
//       Formula 'end_ev' is NOT required to eventually hold, that is, 'cond' may hold forever.
//       Formula 'cond' is not required to hold at the time 'end_ev' holds     
// Arguments:                                                                  
//       - start_ev    Sequence   Enabling event. Occurs each time the sequence 'start_ev' is
//                                matched. In the special case where the sequence is a Boolean,
//                                each time the Boolean is high.               
//       - cond        Property   A property that must hold until 'end_ev' holds.
//       - end_ev      Property   End event is when the property 'end_ev' is true.
// Comments:                                                                   
//       - The property passes if 'end_ev' holds at the same time as 'start_ev'.
//       - There is no explicit bound by which 'end_ev' must occur.            
// Related:                                                                    
//       NEXT_EVENT                                                            
//       REQ_GRANTED                                                           
//       BETWEEN                                                               
//       UNTIL_STRONG                                                          
// Code sample:                                                                
//       `ip2211ringpll_ASSERTS_UNTIL_WEAK(until_w_clk, start_bool, sig==8'h1, end_bool, posedge clk, rst, `ip2211ringpll_ERR_MSG(""));
// Example:                                                                    
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_UNTIL_WEAK(start_ev, cond, end_ev, clk, rst)                     \
   assert property(p_until_weak(start_ev, cond, end_ev, clk, rst))             

`define ip2211ringpll_ASSUME_UNTIL_WEAK(start_ev, cond, end_ev, clk, rst)                     \
   assume property(p_until_weak(start_ev, cond, end_ev, clk, rst))             

`endif                                                                         

`define ip2211ringpll_ASSERTS_UNTIL_WEAK(name, start_ev, cond, end_ev, clk, rst, ip2211ringpll_MSG)         \
   name: assert property(p_until_weak(start_ev, cond, end_ev, clk, rst)) ip2211ringpll_MSG   

`define ip2211ringpll_ASSUMES_UNTIL_WEAK(name, start_ev, cond, end_ev, clk, rst, ip2211ringpll_MSG)         \
   name: assume property(p_until_weak(start_ev, cond, end_ev, clk, rst)) ip2211ringpll_MSG   


// ****************************************************************************************** //



// --- --- ---                                                                 



// ****************************************************************************************** //
// Name:   recur triggers                                                      
// Category: Antecedent/Consequence                                            
// Description:                                                                
//       The Boolean 'cond' must hold after at most 'n' repetitions of the event 'trig'.
//       That is, the 'n'-th next time event 'event' occurs without 'cond' being satisfied,
//       'cond' must be satisfied at the completion of that event.             
// Arguments:                                                                  
//       - trig     Boolean    The Boolean that we count its repetitions.      
//       - n        Number>0   The number of repetitions counted.              
//       - cond     Boolean    The cond that should hold.                      
// Comments:                                                                   
//       None.                                                                 
// Related:                                                                    
// Example:                                                                    
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_RECUR_TRIGGERS(trig, n, cond, clk, rst)                          \
   assert property(p_recur_triggers(trig, n, cond, clk, rst))                  

`define ip2211ringpll_ASSUME_RECUR_TRIGGERS(trig, n, cond, clk, rst)                          \
   assume property(p_recur_triggers(trig, n, cond, clk, rst))                  

`endif                                                                         

`define ip2211ringpll_ASSERTS_RECUR_TRIGGERS(name, trig, n, cond, clk, rst, ip2211ringpll_MSG)              \
   name: assert property(p_recur_triggers(trig, n, cond, clk, rst)) ip2211ringpll_MSG        

`define ip2211ringpll_ASSUMES_RECUR_TRIGGERS(name, trig, n, cond, clk, rst, ip2211ringpll_MSG)              \
    name: assume property(p_recur_triggers(trig, n, cond, clk, rst)) ip2211ringpll_MSG       


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  data transfer                                                        
// Category: Data Checking                                                     
// Description:                                                                
//      Data is transferred correctly from 'start_ev' to 'end_ev'. That is, 'start_data' when
//      'start_ev' holds must be equal to 'end_data' when 'end_ev' holds. If 'start_ev' holds
//      multiple times before 'end_ev' holds, the value of 'start_data' at the occurrence of the
//      last 'start_ev' must match 'end_data' when 'end_ev' holds.             
// Arguments:                                                                  
//      - start_ev    Boolean     Signal denoting the beginning of the transaction.
//      - start_data  Bit-vector  Data at the beginning of transaction.        
//      - end_ev      Boolean     Signal denoting the end of the transaction.  
//      - end_data    Bit-vector  Data at the end of transaction.              
// Comments:                                                                   
//      None.                                                                  
// Related:                                                                    
//      None.                                                                  
// Example:                                                                    
//      TBD |                                                                  
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_DATA_TRANSFER(start_ev, start_data, end_ev, end_data, clk, rst)  \
   assert property(p_data_transfer(start_ev, start_data, end_ev, end_data, clk, rst))

`define ip2211ringpll_ASSUME_DATA_TRANSFER(start_ev, start_data, end_ev, end_data, clk, rst)  \
   assume property(p_data_transfer(start_ev, start_data, end_ev, end_data, clk, rst))

`endif                                                                         

`define ip2211ringpll_ASSERTS_DATA_TRANSFER(name, start_ev, start_data, end_ev, end_data, clk, rst, ip2211ringpll_MSG) \
   name: assert property(p_data_transfer(start_ev, start_data, end_ev, end_data, clk, rst)) ip2211ringpll_MSG

`define ip2211ringpll_ASSUMES_DATA_TRANSFER(name, start_ev, start_data, end_ev, end_data, clk, rst, ip2211ringpll_MSG) \
   name: assume property(p_data_transfer(start_ev, start_data, end_ev, end_data, clk, rst)) ip2211ringpll_MSG


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  gray code                                                            
// Category: Data Checking                                                     
// Description:                                                                
//      At most one bit in 'sig' can change between any two consecutive clock ticks.
// Arguments:                                                                  
//      - sig   Bit-vector   Signal to be checked.                             
// Comments:                                                                   
//      None.                                                                  
// Related:                                                                    
//      None                                                                   
// Example:                                                                    
//      TBD |                                                                  
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_GRAY_CODE(sig, clk, rst)                                         \
   assert property(p_gray_code(sig, clk, rst))                                 

`define ip2211ringpll_ASSUME_GRAY_CODE(sig, clk, rst)                                         \
   assume property(p_gray_code(sig, clk, rst))                                 

`endif                                                                         

`define ip2211ringpll_ASSERTS_GRAY_CODE(name, sig, clk, rst, ip2211ringpll_MSG)                             \
   name: assert property(p_gray_code(sig, clk, rst)) ip2211ringpll_MSG                       

`define ip2211ringpll_ASSUMES_GRAY_CODE(name, sig, clk, rst, ip2211ringpll_MSG)                             \
   name: assume property(p_gray_code(sig, clk, rst)) ip2211ringpll_MSG                       


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  clock ticking                                                        
// Category: Clocks and Resets                                                 
// Description:                                                                
//      The clock 'clock' is ticking. The clock is only required to tick repeatedly. This
//      template requires $global_clock.                                       
// Arguments:                                                                  
// Comments:                                                                   
//      - There is no specific pattern the clock is required to follow.        
// Related:                                                                    
//      None                                                                   
// Example:                                                                    
//      TBD |                                                                  
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_CLOCK_TICKING(clk)                                               \
   assert property(p_clock_ticking(clk))                                       

`define ip2211ringpll_ASSUME_CLOCK_TICKING(clk)                                               \
   assume property(p_clock_ticking(clk))                                       

`endif                                                                         

`define ip2211ringpll_ASSERTS_CLOCK_TICKING(name, clk, ip2211ringpll_MSG)                                   \
   name: assert property(p_clock_ticking(clk)) ip2211ringpll_MSG                             

`define ip2211ringpll_ASSUMES_CLOCK_TICKING(name, clk, ip2211ringpll_MSG)                                   \
   name: assume property(p_clock_ticking(clk)) ip2211ringpll_MSG                             


// ****************************************************************************************** //



// --- --- --- Stability Templates --- --- --- //                              


// ****************************************************************************************** //
// Name:  rigid                                                                
// Category: Stability                                                         
// Description:                                                                
//      Signal 'sig' is considered to be rigid if the first value of 'sig' is determined when
//      the reset becomes low and maintains that value as long as the reset is low.
//      Pay attention, the reset for this template behaves as a lock; when the reset is high,
//      the signal can change its value freely.                                
// Arguments:                                                                  
//      - sig    Bit-vector  The signal that should fulfill rigid constraint.  
// Comments:                                                                   
//      - If no 'rst' signal is passed, the default value will be used, and then 'sig' must 
//        retain its value all the time.                                       
// Related:                                                                    
//      None                                                                   
// Example:                                                                    
//      TBD |//                                                                
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_RIGID(sig, clk, rst)                                             \
   assert property(p_rigid(sig, clk, rst))                                     

`define ip2211ringpll_ASSUME_RIGID(sig, clk, rst)                                             \
   assume property(p_rigid(sig, clk, rst))                                     

`endif                                                                         

`define ip2211ringpll_ASSERTS_RIGID(name, sig, clk, rst, ip2211ringpll_MSG)                                 \
   name: assert property(p_rigid(sig, clk, rst)) ip2211ringpll_MSG                           

`define ip2211ringpll_ASSUMES_RIGID(name, sig, clk, rst, ip2211ringpll_MSG)                                 \
   name: assume property(p_rigid(sig, clk, rst)) ip2211ringpll_MSG                           


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  stable                                                               
// Category: Stability                                                         
// Description:                                                                
//      Signal 'sig' is stable between the two events 'start_ev' and 'end_ev'. The behavior
//      of 'sig' between the clk ticks *is not* checked.                       
// Arguments:                                                                  
//      - sig         Bit-vector  Signal that should remain stable.            
//      - start_ev    Sequence    Start checking event. Checking begins each time the sequence
//                                'start_ev' is matched. In the special case where the sequence
//                                is a Boolean, each time the Boolean is high. 
//      - end_ev      Property    End event is when 'end_ev' is true.          
// Comments:                                                                   
//      - This template checks the behavior of 'sig' only on specified clock ticks. To check
//        the behavior of 'sig' also between specified clock ticks, use GSTABLE.
// Related:                                                                    
//      GSTABLE                                                                
//      STABLE_POSEDGE                                                         
//      STABLE_NEGEDGE                                                         
//      STABLE_EDGE                                                            
// Example:                                                                    
//       | | images/STABLE_1a.png                                              
// Code sample:                                                                
//      `ip2211ringpll_ASSERTS_STABLE(stable_clk, sig, write, stop_write, posedge clk, rst, `ip2211ringpll_ERR_MSG("Bad!"));
// Example:                                                                    
//      Success (start-time:33 and end-time:51) | | images/STABLE_1.png        
// Example:                                                                    
//      Failure (start-stime:111 and end-time:135)  | | images/STABLE_2.png    
// Code sample:                                                                
//     `ip2211ringpll_ASSERTS_STABLE(stable_edge_clk, sig, write, stop_write, clk, rst, `ip2211ringpll_ERR_MSG("Bad!"));
// Example:                                                                    
//     Failure (start-time:1746 and end-time:1770) | | images/STABLE_3.png     
// Example:                                                                    
//     Failure (start-time:1404 and end-time:1458) | | images/STABLE_4.png     
// Code sample:                                                                
//    `ip2211ringpll_ASSERTS_STABLE(stable_posedge_clk, sig, write, write_stop, posedge clk, rst, `ip2211ringpll_ERR_MSG("Bad!"));
// Example:                                                                    
//      Success (start-time:3798 and end-time:3942) | | images/STABLE_5.png    
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_STABLE(sig, start_ev, end_ev, clk, rst)                          \
   assert property(p_stable(sig, start_ev, end_ev, clk, rst))                  

`define ip2211ringpll_ASSUME_STABLE(sig, start_ev, end_ev, clk, rst)                          \
   assume property(p_stable(sig, start_ev, end_ev, clk, rst))                  

`endif                                                                         

`define ip2211ringpll_ASSERTS_STABLE(name, sig, start_ev, end_ev, clk, rst, ip2211ringpll_MSG)              \
   name: assert property(p_stable(sig, start_ev, end_ev, clk, rst)) ip2211ringpll_MSG        

`define ip2211ringpll_ASSUMES_STABLE(name, sig, start_ev, end_ev, clk, rst, ip2211ringpll_MSG)              \
   name: assume property(p_stable(sig, start_ev, end_ev, clk, rst)) ip2211ringpll_MSG        


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  gstable                                                              
// Category: Stability                                                         
// Description:                                                                
//      Signal 'sig' is stable between the two events 'start_ev' and 'end_ev'. The behavior of
//      'sig' between the clk ticks *is not* checked.                          
// Arguments:                                                                  
//      - sig        Bit-vector  Signal that should remain stable.             
//      - start_ev   Sequence    Start checking event. Checking begins each time the sequence
//                               'start_ev' is matched. In the special case where the sequence
//                               is a Boolean, each time the Boolean is high.  
//      - end_ev     Property    End event is when 'end_ev' is true.           
// Comments:                                                                   
//      - To use this checker, the global clocking should be defined.          
//      - GSTABLE works correctly only when each clock tick is at least two global clock ticks.
//      - The lint assertion associated with GSTABLE checks this condition.    
//      - To get same functionality using a clock that is represented by a Boolean signal,
//        use STABLE_POSEDGE, STABLE_NEGEDGE, or STABLE_EDGE.                  
//      - For formal verification this template is also useful as an assumption, since it is
//        easier to debug a counter-example when the signals are stable between user-given events.
// Related:                                                                    
//      STABLE                                                                 
//      STABLE_POSEDGE                                                         
//      STABLE_NEGEDGE                                                         
//      STABLE_EDGE                                                            
// Example:                                                                    
//       | | images/GSTABLE_1.png                                              
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_GSTABLE(sig, start_ev, end_ev, clk, rst)                         \
   assert property(p_gstable_ev(sig, start_ev, end_ev, clk, rst))              

`define ip2211ringpll_ASSUME_GSTABLE(sig, start_ev, end_ev, clk, rst)                         \
   assume property(p_gstable_ev(sig, start_ev, end_ev, clk, rst))              

`endif                                                                         

`define ip2211ringpll_ASSERTS_GSTABLE(name, sig, start_ev, end_ev, clk, rst, ip2211ringpll_MSG)             \
   name: assert property(p_gstable_ev(sig, start_ev, end_ev, clk, rst)) ip2211ringpll_MSG    

`define ip2211ringpll_ASSUMES_GSTABLE(name, sig, start_ev, end_ev, clk, rst, ip2211ringpll_MSG)             \
   name: assume property(p_gstable_ev(sig, start_ev, end_ev, clk, rst)) ip2211ringpll_MSG    


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  stable posedge                                                       
// Category: Stability                                                         
// Description:                                                                
//      Signal 'sig' is stable between the two events 'start_ev' and 'end_ev'. The behavior of
//      'sig' between the clk ticks is checked. The clock argument of this template must be a
//      Boolean signal. This template regards the POSEDGE of 'clk' as the clock tick. This is
//      a global-clock based property.                                         
// Arguments:                                                                  
//      - sig         Bit-vector  Signal that should remain stable.            
//      - start_ev    Sequence    Start checking event. Checking begins each time the sequence
//                                'start_ev' is matched. In the special case where the sequence
//                                is a Boolean, each time the Boolean is high. 
//      - end_ev      Property    End event is when 'end_ev' is true.          
// Comments:                                                                   
//      - To use this checker, the global clocking should be defined.          
//      - To get same functionality using a clock that is represented by an event, use GSTABLE
//      - For formal verification this template is also useful as an assumption, since it is
//        easier to debug a counter-example when the signals are stable between user-given 
//        events.                                                              
// Related:                                                                    
//      GSTABLE                                                                
//      STABLE_NEGEDGE                                                         
//      STABLE_EDGE                                                            
// Example:                                                                    
//       | | images/STABLE_POSEDGE_1.png                                       
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`ifndef ip2211ringpll_SVA_LIB_SVA2005                                                        

`define ip2211ringpll_ASSERT_STABLE_POSEDGE(sig, start_ev, end_ev, clk, rst)                  \
   `ip2211ringpll_ASSERT_GSTABLE(sig, start_ev, end_ev, posedge (clk), rst)                  

`define ip2211ringpll_ASSUME_STABLE_POSEDGE(sig, start_ev, end_ev, clk, rst)                  \
   `ip2211ringpll_ASSUME_GSTABLE(sig, start_ev, end_ev, posedge (clk), rst)                  

`else                                                                          

`define ip2211ringpll_ASSERT_STABLE_POSEDGE(sig, start_ev, end_ev, clk, rst)                  \
   assert property(p_gstable_sig_posedge(sig, start_ev, end_ev, clk, rst))     

`define ip2211ringpll_ASSUME_STABLE_POSEDGE(sig, start_ev, end_ev, clk, rst)                  \
   assume property(p_gstable_sig_posedge(sig, start_ev, end_ev, clk, rst))     

`endif                                                                         

`endif                                                                         

// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  stable negedge                                                       
// Category: Stability                                                         
// Description:                                                                
//      Signal 'sig' is stable between the two events 'start_ev' and 'end_ev'. The behavior of
//      'sig' between the clk ticks is checked. The clock argument of this template must be a
//      Boolean signal. This template regards the NEGEDGE of 'clk' as the clock tick. This is
//      a global-clock based property.                                         
// Arguments:                                                                  
//      - sig        Bit-vector  Signal that should remain stable.             
//      - start_ev   Sequence    Start checking event. Checking begins each time the sequence
//                               'start_ev' is matched. In the special case where the sequence
//                               is a Boolean, each time the Boolean is high.  
//      - end_ev     Property    End event is when 'end_ev' is true.           
// Comments:                                                                   
//      - To use this checker, the global clocking should be defined.          
//      - To get same functionality using a clock that is represented by an event, use GSTABLE
//      - For formal verification this template is also useful as an assumption, since it is
//        easier to debug a counter-example when the signals are stable between user-given events.
// Related:                                                                    
//      GSTABLE                                                                
//      STABLE_POSEDGE                                                         
//      STABLE_EDGE                                                            
// Example:                                                                    
//       | | images/STABLE_NEGEDGE_1.png                                       
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`ifndef ip2211ringpll_SVA_LIB_SVA2005                                                        

`define ip2211ringpll_ASSERT_STABLE_NEGEDGE(sig, start_ev, end_ev, clk, rst)                  \
   `ip2211ringpll_ASSERT_GSTABLE(sig, start_ev, end_ev, negedge (clk), rst)                   \

`define ip2211ringpll_ASSUME_STABLE_NEGEDGE(sig, start_ev, end_ev, clk, rst)                  \
   `ip2211ringpll_ASSUME_GSTABLE(sig, start_ev, end_ev, negedge (clk), rst)                   \

`else                                                                          

`define ip2211ringpll_ASSERT_STABLE_NEGEDGE(sig, start_ev, end_ev, clk, rst)                  \
   assert property(p_gstable_sig_negedge(sig, start_ev, end_ev, clk, rst))      

`define ip2211ringpll_ASSUME_STABLE_NEGEDGE(sig, start_ev, end_ev, clk, rst)                  \
   assume property(p_gstable_sig_negedge(sig, start_ev, end_ev, clk, rst))     

`endif                                                                         

`endif                                                                         

// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  stable edge                                                          
// Category: Stability                                                         
// Description:                                                                
//      Signal 'sig' is stable between the two events 'start_ev' and 'end_ev'. The behavior of
//      'sig' between the clk ticks is checked. The clock argument of this template must be a
//      Boolean signal. This template regards every change of 'clk' as a clock tick. This is a
//      global-clock based property.                                           
// Arguments:                                                                  
//      - sig        Bit-vector  Signal that should remain stable.             
//      - start_ev   Sequence    Start checking event. Checking begins each time the sequence
//                               'start_ev' is matched. In the special case where the sequence
//                               is a Boolean, each time the Boolean is high.  
//      - end_ev     Property    End event is when 'end_ev' is true.           
// Comments:                                                                   
//      - To use this checker, the global clocking should be defined.          
//      - To get same functionality using a clock that is represented by an event, use GSTABLE
// Related:                                                                    
//      GSTABLE                                                                
//      STABLE_POSEDGE                                                         
//      STABLE_NEGEDGE                                                         
// Example:                                                                    
//       | | images/STABLE_EDGE_1.png                                          
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`ifndef ip2211ringpll_SVA_LIB_SVA2005                                                        

`define ip2211ringpll_ASSERT_STABLE_EDGE(sig, start_ev, end_ev, clk, rst)                     \
   `ip2211ringpll_ASSERT_GSTABLE(sig, start_ev, end_ev, clk, rst)                             \

`define ip2211ringpll_ASSUME_STABLE_EDGE(sig, start_ev, end_ev, clk, rst)                     \
   `ip2211ringpll_ASSUME_GSTABLE(sig, start_ev, end_ev, clk, rst)                             \

`else                                                                          

`define ip2211ringpll_ASSERT_STABLE_EDGE(sig, start_ev, end_ev, clk, rst)                     \
   assert property(p_gstable_sig_edge(sig, start_ev, end_ev, clk, rst))        

`define ip2211ringpll_ASSUME_STABLE_EDGE(sig, start_ev, end_ev, clk, rst)                     \
   assume property(p_gstable_sig_edge(sig, start_ev, end_ev, clk, rst))       

`endif                                                                         

`endif                                                                         

// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  stable window                                                        
// Category: Stability                                                         
// Description:                                                                
//      Whenever 'sample' is high, 'sig' must keep its value for 'clks_after' additional clocks
//      after the sampling point, and 'clks_before' clocks before the sampling point. 'sig' is
//      not required to remain stable between the clock ticks.                 
// Arguments:                                                                  
//      - sample      Boolean         Sampling signal.                         
//      - sig         Bit-vector      Signal that should remain stable.        
//      - clks_before Number>=0       Number of cycles before the sampling point during which
//                                    'sig' must keep its value.               
//      - clks_after  Number>=0       Number of cycles after the sampling point during which
//                                    'sig' must keep its value.               
// Comments:                                                                   
//      - This checker is *not* backward compatible. The previous implementation effectively used
//        'clks_before' -1, and required that 'clks_before' be strongly positive.
//      - This template checks the value of 'sig' only on clock ticks; 'sig' is not required to
//        remain stable between the clock ticks.                               
//      - When 'clks_before' is equal to 0, this template is equivalent to STABLE_AFTER.
// Related:                                                                    
//      GSTABLE_WINDOW                                                         
//      STABLE_AFTER                                                           
//      BETWEEN_TIME                                                           
// Example:                                                                    
//       | | images/STABLE_WINDOW_1.png                                        
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_STABLE_WINDOW(sample, sig, clks_before, clks_after, clk, rst)    \
   assert property(p_stable_window(sample, sig, clks_before, clks_after, clk, rst))

`define ip2211ringpll_ASSUME_STABLE_WINDOW(sample, sig, clks_before, clks_after, clk, rst)    \
   assume property(p_stable_window(sample, sig, clks_before, clks_after, clk, rst))

`endif                                                                         

`define ip2211ringpll_ASSERTS_STABLE_WINDOW(name, sample, sig, clks_before, clks_after, clk, rst, ip2211ringpll_MSG) \
   name: assert property(p_stable_window(sample, sig, clks_before, clks_after, clk, rst)) ip2211ringpll_MSG

`define ip2211ringpll_ASSUMES_STABLE_WINDOW(name, sample, sig, clks_before, clks_after, clk, rst, ip2211ringpll_MSG) \
   name: assume property(p_stable_window(sample, sig, clks_before, clks_after, clk, rst)) ip2211ringpll_MSG


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  gstable window                                                       
// Category: Stability                                                         
// Description:                                                                
//      Whenever 'sample' is high, 'sig' must be stable 'clks_after' additional clocks
//      (including) after the sampling point and 'clks_before' clocks (including) before the
//      sampling point. 'sig' must be stable between the clock ticks as well.  
// Arguments:                                                                  
//      - sample      Boolean         Sampling signal.                         
//      - sig         Bit-vector      Signal that should remain stable.        
//      - clks_before Number>=0       Number of cycles before the sampling point during which
//                                    'sig' must keep its value.               
//      - clks_after  Number>=0       Number of cycles after the sampling point during which
//                                    'sig' must keep its value.               
// Comments:                                                                   
//      - To use this checker, the global clocking should be defined.          
//        GSTABLE_WINDOW works correctly only when each clock tick is at least two global clock
//        ticks. This template checks the value of 'sig' only on clock ticks; 'sig' is required
//      - to remain stable between the clock ticks. When 'clks_before' is equal to 0, this template
//        is equivalent to GSTABLE_AFTER.                                      
// Related:                                                                    
//      STABLE_WINDOW                                                          
//      GSTABLE_AFTER                                                          
// Example:                                                                    
//       | | images/GSTABLE_WINDOW_1.png                                       
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_GSTABLE_WINDOW(sample, sig, clks_before, clks_after, clk, rst)   \
   assert property(p_gstable_window(sample, sig, clks_before, clks_after, clk, rst))

`define ip2211ringpll_ASSUME_GSTABLE_WINDOW(sample, sig, clks_before, clks_after, clk, rst)   \
   assume property(p_gstable_window(sample, sig, clks_before, clks_after, clk, rst))

`endif                                                                         

`define ip2211ringpll_ASSERTS_GSTABLE_WINDOW(name, sample, sig, clks_before, clks_after, clk, rst, ip2211ringpll_MSG) \
   name: assert property(p_gstable_window(sample, sig, clks_before, clks_after, clk, rst)) ip2211ringpll_MSG

`define ip2211ringpll_ASSUMES_GSTABLE_WINDOW(name, sample, sig, clks_before, clks_after, clk, rst, ip2211ringpll_MSG) \
   name: assume property(p_gstable_window(sample, sig, clks_before, clks_after, clk, rst)) ip2211ringpll_MSG


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  stable for                                                           
// Category: Stability                                                         
// Description:                                                                
//      Whenever 'sig' changes, it must keep its value for n additional clocks. The number of
//      clocks n does not include the clock at which 'sig' changed. 'sig' must be stable at the
//      'n'th tick point. Values of 'sig' are only sampled at the ticks of 'clk'. The change of
//      'sig' should be from one clock tick to another. The behavior of 'sig' between the clock
//      ticks *is not* checked                                                 
// Arguments:                                                                  
//      - sig     Bit-vector  Signal that should remain stable.                
//      - n       Number>0    The minimum number of cycles throughout which 'sig' keeps its value.
// Comments:                                                                   
//      - This checker is expensive for a large n. In this case use, STABLE if possible (if the
//        signal retains its value between events, rather than during a time interval).
// Related:                                                                    
//      REMAIN_HIGH                                                            
//      REMAIN_LOW                                                             
//      BETWEEN_TIME                                                           
//      GSTABLE_FOR                                                            
// Example:                                                                    
//       | | images/STABLE_FOR_1.png                                           
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_STABLE_FOR(sig, n, clk, rst)                                     \
   assert property(p_stable_for(sig, n, clk, rst))                             

`define ip2211ringpll_ASSUME_STABLE_FOR(sig, n, clk, rst)                                     \
   assume property(p_stable_for(sig, n, clk, rst))                             

`endif                                                                         

`define ip2211ringpll_ASSERTS_STABLE_FOR(name, sig, n, clk, rst, ip2211ringpll_MSG)                         \
   name: assert property(p_stable_for(sig, n, clk, rst)) ip2211ringpll_MSG                   

`define ip2211ringpll_ASSUMES_STABLE_FOR(name, sig, n, clk, rst, ip2211ringpll_MSG)                         \
   name: assume property(p_stable_for(sig, n, clk, rst)) ip2211ringpll_MSG                   


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  gstable for                                                          
// Category: Stability                                                         
// Description:                                                                
//      Whenever 'sig' changes, it must keep its value for n additional clocks. The number of
//      clocks n does not include the clock at which 'sig' changed. 'sig' must be stable at the
//      n-th tick point. Values of 'sig' are only sampled at the ticks of 'clk'. The change of
//      'sig' should be from one clock tick to another. However, 'sig' *is* required to be stable
//      at all times during the n clock ticks, even at the non-tick points of the clock.
// Arguments:                                                                  
//      - sig     Bit-vector  Signal that should remain stable.                
//      - n       Number>0    The minimum number of cycles throughout which 'sig' keeps its value.
// Comments:                                                                   
//      - To use this checker, the global clocking should be defined.          
//      - This checker is expensive for a large n. In this case use GSTABLE if possible (if the
//        signal retains its value between events, rather than during a time interval).
//      - In formal verification, although the value of 'sig' may be irrelevant between the tick
//        points of 'clk', it is more convenient to examine the counter-example when it is stable.
// Related:                                                                    
//      STABLE_AFTER                                                           
//      GSTABLE_WINDOW                                                         
//      STABLE_FOR                                                             
// Example:                                                                    
//       | | images/GSTABLE_FOR_1.png                                          
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_GSTABLE_FOR(sig, n, clk, rst)                                    \
   assert property(p_gstable_for(sig, n, clk, rst))                            

`define ip2211ringpll_ASSUME_GSTABLE_FOR(sig, n, clk, rst)                                    \
   assume property(p_gstable_for(sig, n, clk, rst))                            

`endif                                                                         

`define ip2211ringpll_ASSERTS_GSTABLE_FOR(name, sig, n, clk, rst, ip2211ringpll_MSG)                        \
   name: assert property(p_gstable_for(sig, n, clk, rst)) ip2211ringpll_MSG                  

`define ip2211ringpll_ASSUMES_GSTABLE_FOR(name, sig, n, clk, rst, ip2211ringpll_MSG)                        \
   name: assume property(p_gstable_for(sig, n, clk, rst)) ip2211ringpll_MSG                  


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  stable after                                                         
// Category: Stability                                                         
// Description:                                                                
//      Whenever sample is high, 'sig' must keep its value for 'clks_after' additional clocks
//      after the sampling point. The behavior of 'sig' between the clock ticks *is* checked.
// Arguments:                                                                  
//      - sample      Sequence    Sampling event. Sampling begins each time the sequence
//                                'sample' is matched. In the special case where the
//                                sequence is a Boolean, each time the Boolean is high.
//      - sig         Bit-vector  Signal that should remain stable.            
//      - clks_after  Number>0    Number of additional cycles after the sampling point
//                                during which 'sig' must keep its value.      
// Comments:                                                                   
//      None.                                                                  
// Related:                                                                    
//      GSTABLE_AFTER                                                          
//      STABLE_WINDOW                                                          
//      STABLE_FOR                                                             
// Example:                                                                    
//       | | images/STABLE_AFTER_1.png                                         
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_STABLE_AFTER(sample, sig, clks_after, clk, rst)                  \
   assert property(p_stable_after(sample, sig, clks_after, clk, rst))          

`define ip2211ringpll_ASSUME_STABLE_AFTER(sample, sig, clks_after, clk, rst)                  \
   assume property(p_stable_after(sample, sig, clks_after, clk, rst))          

`endif                                                                         

`define ip2211ringpll_ASSERTS_STABLE_AFTER(name, sample, sig, clks_after, clk, rst, ip2211ringpll_MSG)      \
   name: assert property(p_stable_after(sample, sig, clks_after, clk, rst)) ip2211ringpll_MSG

`define ip2211ringpll_ASSUMES_STABLE_AFTER(name, sample, sig, clks_after, clk, rst, ip2211ringpll_MSG)      \
   name: assume property(p_stable_after(sample, sig, clks_after, clk, rst)) ip2211ringpll_MSG


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  gstable after                                                        
// Category: Stability                                                         
// Description:                                                                
//      Whenever sample is high, 'sig' must keep its value for 'clks_after' additional clocks
//      after the sampling point. The behavior of 'sig' between the clock ticks *is* checked.
// Arguments:                                                                  
//      - sample      Sequence    Sampling event. Sampling begins each time the sequence
//                                'sample' is matched. In the special case where the sequence
//                                is a Boolean, each time the Boolean is high. 
//      - sig         Bit-vector  Signal that should remain stable.            
//      - clks_after  Number>0    Number of additional cycles after the sampling point during
//                                which 'sig' must keep its value.             
// Comments:                                                                   
//      None.                                                                  
// Related:                                                                    
//      TBD                                                                    
// Example:                                                                    
//       | | images/GSTABLE_AFTER_1.png                                        
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_GSTABLE_AFTER(sample, sig, clks_after, clk, rst)                 \
   assert property(p_gstable_after(sample, sig, clks_after, clk, rst))         

`define ip2211ringpll_ASSUME_GSTABLE_AFTER(sample, sig, clks_after, clk, rst)                 \
   assume property(p_gstable_after(sample, sig, clks_after, clk, rst))         

`endif                                                                         

`define ip2211ringpll_ASSERTS_GSTABLE_AFTER(name, sample, sig, clks_after, clk, rst, ip2211ringpll_MSG)     \
   name: assert property(p_gstable_after(sample, sig, clks_after, clk, rst)) ip2211ringpll_MSG

`define ip2211ringpll_ASSUMES_GSTABLE_AFTER(name, sample, sig, clks_after, clk, rst, ip2211ringpll_MSG)     \
   name: assume property(p_gstable_after(sample, sig, clks_after, clk, rst)) ip2211ringpll_MSG


// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  gstable between ticks                                                
// Category: Stability                                                         
// Description:                                                                
//      Signal 'sig' is stable between every two clock events. The value of 'sig' can only
//      change at a clock event (i.e. when 'sig' is sampled). The value of 'sig' at event 'i'
//      should hold until event 'i+1' (exclusively). The clock argument of this template must
//      be an event (e.g. a signal with an edge specifier).                    
//      This is a global-clock based property.                                 
// Arguments:                                                                  
//      - sig     Bit-vector  Signal that should remain stable.                
// Comments:                                                                   
//      - To use this checker, the global clocking should be defined.          
//      - To get same functionality using a clock that is represented by a Boolean signal, use
//        STABLE_BETWEEN_TICKS_POSEDGE, STABLE_BETWEEN_TICKS_NEGEDGE, or STABLE_BETWEEN_TICKS_EDGE.
//      - For formal verification this template is also useful as an assumption, since it is easier
//        to debug a counter-example when the signals are stable between clock ticks.
//      - Pay attention: A clock tick is needed in order to start checking, i.e, the signal is 
//        not checked for stability starting from point where the reset becomes in-active, until
//        the first clock tick.                                                
// Related:                                                                    
//      STABLE                                                                 
//      GSTABLE_BETWEEN_TICKS                                                  
//      STABLE_BETWEEN_TICKS_POSEDGE                                           
//      STABLE_BETWEEN_TICKS_NEGEDGE                                           
//      STABLE_BETWEEN_TICKS_EDGE                                              
// Example:                                                                    
//      TBD |                                                                  
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`define ip2211ringpll_ASSERT_GSTABLE_BETWEEN_TICKS(sig, clk, rst)                             \
   assert property(p_gstable_between_ticks_ev(sig, clk, rst)) /* novas s-70517 */

`define ip2211ringpll_ASSUME_GSTABLE_BETWEEN_TICKS(sig, clk, rst)                             \
   assume property(p_gstable_between_ticks_ev(sig, clk, rst)) /* novas s-70517 */

`endif                                                                         

`define ip2211ringpll_ASSERTS_GSTABLE_BETWEEN_TICKS(name, sig, clk, rst, ip2211ringpll_MSG)                 \
   name: assert property(p_gstable_between_ticks_ev(sig, clk, rst)) /* novas s-70517 */ ip2211ringpll_MSG        

`define ip2211ringpll_ASSUMES_GSTABLE_BETWEEN_TICKS(name, sig, clk, rst, ip2211ringpll_MSG)                 \
   name: assume property(p_gstable_between_ticks_ev(sig, clk, rst)) /* novas s-70517 */ ip2211ringpll_MSG        


// ****************************************************************************************** //



// --- --- ---                                                                 



// ****************************************************************************************** //
// Name:  stable between ticks posedge                                         
// Category: Stability                                                         
// Description:                                                                
//      Signal 'sig' is stable between every two 'clk' ticks. The value of 'sig' can only
//      change at a 'clk' tick (i.e. when 'sig' is sampled). The value of 'sig' at tick 'i'
//      should hold until tick 'i+1' (exclusively). The clock argument of this template must be
//      a Boolean signal. This version regards the POSEDGE of 'clk' as the clock tick. This is
//      a global-clock based property.                                         
// Arguments:                                                                  
//      - sig     Bit-vector  Signal that should remain stable.                
//      - clk     Boolean     clk is treated as regular signal.                
// Comments:                                                                   
//      - To use this checker, the global clocking should be defined.          
//      - To get same functionality using a clock that is represented by an event use
//        GSTABLE_BETWEEN_TICKS. For formal verification this template is also useful as an assumption,
//        since it is easier to debug a counter-example when the signals are stable between clock ticks.
//      - This template immitates the clock behaviour by itself.               
// Related:                                                                    
//      STABLE                                                                 
//      GSTABLE_BETWEEN_TICKS                                                  
//      STABLE_BETWEEN_TICKS_NEGEDGE                                           
//      STABLE_BETWEEN_TICKS_EDGE                                              
// Example:                                                                    
//      TBD |                                                                  
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`ifndef ip2211ringpll_SVA_LIB_SVA2005                                                        

`define ip2211ringpll_ASSERT_STABLE_BETWEEN_TICKS_POSEDGE(sig, clk, rst)                      \
   `ip2211ringpll_ASSERT_GSTABLE_BETWEEN_TICKS(sig, posedge (clk), rst)                      

`define ip2211ringpll_ASSUME_STABLE_BETWEEN_TICKS_POSEDGE(sig, clk, rst)                      \
   `ip2211ringpll_ASSUME_GSTABLE_BETWEEN_TICKS(sig, posedge (clk), rst)                      

`else                                                                          

`define ip2211ringpll_ASSERT_STABLE_BETWEEN_TICKS_POSEDGE(sig, clk, rst)                      \
   assert property(p_gstable_between_ticks_sig_posedge(sig, clk, rst)) /* novas s-70517 */

`define ip2211ringpll_ASSUME_STABLE_BETWEEN_TICKS_POSEDGE(sig, clk, rst)                      \
   assume property(p_gstable_between_ticks_sig_posedge(sig, clk, rst)) /* novas s-70517 */

`endif                                                                         

`endif                                                                         

// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  stable between ticks negedge                                         
// Category: Stability                                                         
// Description:                                                                
//      Signal 'sig' is stable between every two 'clk' ticks. The value of 'sig' can only change
//      at a 'clk' tick (i.e. when 'sig' is sampled). The value of 'sig' at tick 'i' should hold
//      until tick 'i+1' (exclusively). The clock argument of this template must be a Boolean
//      signal. This version regards the NEGEDGE of 'clk' as the clock tick. This is a global-clock
//      based property.                                                        
// Arguments:                                                                  
//      - sig     Bit-vector  Signal that should remain stable.                
//      - clk     Boolean     clk is treated as regular signal.                
// Comments:                                                                   
//      - To use this checker, the global clocking should be defined.          
//      - To get same functionality using a clock that is represented by an event use
//        GSTABLE_BETWEEN_TICKS. For formal verification this template is also useful as an
//        assumption, since it is easier to debug a counter-example when the signals are stable
//        between clock ticks. This template immitates the clock behaviour by itself.
// Related:                                                                    
//      STABLE                                                                 
//      GSTABLE_BETWEEN_TICKS                                                  
//      STABLE_BETWEEN_TICKS_POSEDGE                                           
//      STABLE_BETWEEN_TICKS_EDGE                                              
// Example:                                                                    
//      TBD |                                                                  
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`ifndef ip2211ringpll_SVA_LIB_SVA2005                                                        

`define ip2211ringpll_ASSERT_STABLE_BETWEEN_TICKS_NEGEDGE(sig, clk, rst)                      \
   `ip2211ringpll_ASSERT_GSTABLE_BETWEEN_TICKS(sig, negedge (clk), rst)                      

`define ip2211ringpll_ASSUME_STABLE_BETWEEN_TICKS_NEGEDGE(sig, clk, rst)                      \
   `ip2211ringpll_ASSUME_GSTABLE_BETWEEN_TICKS(sig, negedge (clk), rst)                      


`else                                                                          

`define ip2211ringpll_ASSERT_STABLE_BETWEEN_TICKS_NEGEDGE(sig, clk, rst)                      \
   assert property(p_gstable_between_ticks_sig_negedge(sig, clk, rst)) /* novas s-70517 */ 

`define ip2211ringpll_ASSUME_STABLE_BETWEEN_TICKS_NEGEDGE(sig, clk, rst)                      \
   assume property(p_gstable_between_ticks_sig_negedge(sig, clk, rst)) /* novas s-70517 */

`endif                                                                         

`endif                                                                         

// ****************************************************************************************** //



// --- --- ---                                                                 


// ****************************************************************************************** //
// Name:  stable between ticks edge                                            
// Category: Stability                                                         
// Description:                                                                
//      Signal 'sig' is stable between every two 'clk' ticks. The value of 'sig' can only change
//      at a 'clk' tick (i.e. when 'sig' is sampled). The value of 'sig' at tick 'i' should hold
//      until tick 'i+1' (exclusively). The clock argument of this template must be a Boolean
//      signal. This template regards every change of 'clk' as a clock tick. This is a global-clock
//      based property.                                                        
// Arguments:                                                                  
//      - sig     Bit-vector  Signal that should remain stable.                
//      - clk     Boolean     clk is treated as regular signal.                
// Comments:                                                                   
//      - To use this checker, the global clocking should be defined.          
//      - To get same functionality using a clock that is represented by an event use
//        GSTABLE_BETWEEN_TICKS. For formal verification this template is also useful as an
//        assumption, since it is easier to debug a counter-example when the signals are stable
//        between clock ticks. This template immitates the clock behaviour by itself.
// Related:                                                                    
//      STABLE                                                                 
//      GSTABLE_BETWEEN_TICKS                                                  
//      STABLE_BETWEEN_TICKS_POSEDGE                                           
//      STABLE_BETWEEN_TICKS_NEGEDGE                                           
// Example:                                                                    
//      TBD |                                                                  
//                                                                             
// ------------------------------------------------------------------------------------------ //

`ifdef INTC_SVA_LIB_OLD_FORMAT                                                      

`ifndef ip2211ringpll_SVA_LIB_SVA2005                                                        

`define ip2211ringpll_ASSERT_STABLE_BETWEEN_TICKS_EDGE(sig, clk, rst)                         \
   `ip2211ringpll_ASSERT_GSTABLE_BETWEEN_TICKS(sig, clk, rst)                                

`define ip2211ringpll_ASSUME_STABLE_BETWEEN_TICKS_EDGE(sig, clk, rst)                         \
   `ip2211ringpll_ASSUME_GSTABLE_BETWEEN_TICKS(sig, clk, rst)                                

`else                                                                          

`define ip2211ringpll_ASSERT_STABLE_BETWEEN_TICKS_EDGE(sig, clk, rst)                         \
   assert property(p_gstable_between_ticks_sig_edge(sig, clk, rst)) /* novas s-70517 */ 

`define ip2211ringpll_ASSUME_STABLE_BETWEEN_TICKS_EDGE(sig, clk, rst)                         \
   assume property(p_gstable_between_ticks_sig_edge(sig, clk, rst)) /* novas s-70517 */

`endif                                                                         

`endif                                                                         

// ****************************************************************************************** //



// --- --- ---                                                                 


// ***********Currently not supported******************************************************** //
// Name:   transaction length                                                  
// Description:                                                                
//       Check that a transaction delimited by start_ev and end_ev lasts at least min cycles
//       and at most max cycles.                                               
// Arguments:                                                                  
//       start_ev   Formula                                                    
//       end_ev     Boolean                                                    
//       min        Signal or constant                                         
//       max        Signal or constant                                         
// Comments:                                                                   
// Related:                                                                    
// Example:                                                                    
//                                                                             
// ------------------------------------------------------------------------------------------ //
//                                                                             
//`define ASSERT_TRANSACTION_LENGTH (start_ev, end_ev, min , max, clk , rst)    \
//   assert property(p_transaction_length(start_ev, end_ev, min , max, clk , rst)
//                                                                             
//`define ASSUME_TRANSACTION_LENGTH (start_ev, end_ev, min , max, clk , rst)    \
//   assume property(p_transaction_length(start_ev, end_ev, min , max, clk , rst)
//                                                                             
//`ifndef INTC_SVA_LIB_OLD_FORMAT                                                   
//                                                                             
//`define ASSERTS_TRANSACTION_LENGTH (name, start_ev, end_ev, min , max, clk , rst, ip2211ringpll_MSG) \
//   name: `ASSERT_TRANSACTION_LENGTH (start_ev, end_ev, min , max, clk , rst) ip2211ringpll_MSG
//                                                                             
//`define ASSUMES_TRANSACTION_LENGTH (name, start_ev, end_ev, min , max, clk , rst, ip2211ringpll_MSG) \
//   name: `ASSUME_TRANSACTION_LENGTH (start_ev, end_ev, min , max, clk , rst) ip2211ringpll_MSG
//                                                                             
//`endif                                                                       
//                                                                             
// ****************************************************************************************** //



// --- --- ---                                                                 


// **********Currently not supported********************************************************** //
// Name:   tagged request granted                                              
// Description:                                                                
//       A tagged request is eventually granted with a signal having same tag. 
//       The request does not need to remain pending until it is granted       
// Arguments:                                                                  
//       req       Formula                                                     
//       gnt       Formula                                                     
//       req_tag   Bit-vector                                                  
//       gnt_tag   Bit-vector                                                  
//                                                                             
// ------------------------------------------------------------------------------------------ //
//                                                                             
//`define ASSERT_TAGGED_REQ_GRANTED(req, req_tag, gnt, gnt_tag, clk, rst)       \
//   assert property(tagged_req_granted(req, req_tag, gnt, gnt_tag, clk, rst)) 
//                                                                             
//`define ASSUME_TAGGED_REQ_GRANTED(req, req_tag, gnt, gnt_tag, clk, rst)       \
//   assume property(tagged_req_granted(req, req_tag, gnt, gnt_tag, clk, rst)) 
//                                                                             
//`ifndef INTC_SVA_LIB_OLD_FORMAT                                                   
//                                                                             
//`define ASSERTS_TAGGED_REQ_GRANTED(name, req, req_tag, gnt, gnt_tag, clk, rst, ip2211ringpll_MSG) \
//   name:  `ASSERT_TAGGED_REQ_GRANTED(req, req_tag, gnt, gnt_tag, clk, rst) ip2211ringpll_MSG
//                                                                             
//`define ASSUMES_TAGGED_REQ_GRANTED(name, req, req_tag, gnt, gnt_tag, clk, rst, ip2211ringpll_MSG) \
//   name:  `ASSUME_TAGGED_REQ_GRANTED(req, req_tag, gnt, gnt_tag, clk, rst) ip2211ringpll_MSG
//                                                                             
//`endif                                                                       
//                                                                             
// ****************************************************************************************** //

`endif // ip2211ringpll_INTEL_CHECKERS_CORE_VS



`ifndef ip2211ringpll_INTEL_CHECKERS_CORE_IMP_VS
`define ip2211ringpll_INTEL_CHECKERS_CORE_IMP_VS

// X/Z checking 
`ifndef INTC_SVA_LIB_IGNOREXZ
    `define ip2211ringpll_SVA_LIB_KNOWN(sig) (!($isunknown({>>{sig}})))
    `define ip2211ringpll_SVA_LIB_SAME(siga,sigb) ((siga)==(sigb))
`else
    `define ip2211ringpll_SVA_LIB_KNOWN(sig) (1'b1)
    `define ip2211ringpll_SVA_LIB_SAME(siga,sigb) ((siga)===(sigb))
`endif

`ifndef ip2211ringpll_SVA_LIB_SVA2005

    let ip2211ringpll_l_mutexed(sig) = $onehot0({>>{sig}}) && `ip2211ringpll_SVA_LIB_KNOWN(sig);
    `define ip2211ringpll_l_mutexed(sig) ip2211ringpll_l_mutexed(sig)
    let ip2211ringpll_l_at_most_bits_high(sig, n) = ($countones({>>{sig}}) <= n) && `ip2211ringpll_SVA_LIB_KNOWN(sig);
    `define ip2211ringpll_l_at_most_bits_high(sig, n) ip2211ringpll_l_at_most_bits_high(sig, n)
    let ip2211ringpll_l_at_most_bits_low(sig, n) = ($countones({>>{~sig}}) <= n) && `ip2211ringpll_SVA_LIB_KNOWN(sig);
    `define ip2211ringpll_l_at_most_bits_low(sig, n) ip2211ringpll_l_at_most_bits_low(sig, n)
    let ip2211ringpll_l_bits_high(sig, n) = ($countones({>>{sig}}) == n) && `ip2211ringpll_SVA_LIB_KNOWN(sig);
    `define ip2211ringpll_l_bits_high(sig, n) ip2211ringpll_l_bits_high(sig, n)
    let ip2211ringpll_l_bits_low(sig, n) = ($countones({>>{~sig}}) == n) && `ip2211ringpll_SVA_LIB_KNOWN(sig);
    `define ip2211ringpll_l_bits_low(sig, n) ip2211ringpll_l_bits_low(sig, n)
    let ip2211ringpll_l_same_bits(sig) = (&(sig)) || !(|(sig)) && `ip2211ringpll_SVA_LIB_KNOWN(sig);
    `define ip2211ringpll_l_same_bits(sig) ip2211ringpll_l_same_bits(sig)
    let ip2211ringpll_l_one_hot(sig) = $onehot({>>{sig}}) && `ip2211ringpll_SVA_LIB_KNOWN(sig);
    `define ip2211ringpll_l_one_hot(sig) ip2211ringpll_l_one_hot(sig)
    let ip2211ringpll_l_known_driven(sig) = `ip2211ringpll_SVA_LIB_KNOWN(sig);
    `define ip2211ringpll_l_known_driven(sig) ip2211ringpll_l_known_driven(sig)
    let ip2211ringpll_l_forbidden(cond) = !(cond);
    `define ip2211ringpll_l_forbidden(cond) ip2211ringpll_l_forbidden(cond)
    let ip2211ringpll_l_must(prop) = (prop);
    `define ip2211ringpll_l_must(prop) ip2211ringpll_l_must(prop)
    let ip2211ringpll_l_trigger(trig_sig, prop_sig) = (trig_sig -> prop_sig);
    `define ip2211ringpll_l_trigger(trig_sig, prop_sig) ip2211ringpll_l_trigger(trig_sig, prop_sig)
    let ip2211ringpll_l_range(sig, low, high) = (((sig) >=(low)) & ((sig) <=(high)));
    `define ip2211ringpll_l_range(sig, low, high) ip2211ringpll_l_range(sig, low, high)
    let ip2211ringpll_l_max_value(sig, max_val) = ((sig) <= (max_val));
    `define ip2211ringpll_l_max_value(sig, max_val) ip2211ringpll_l_max_value(sig, max_val)
    let ip2211ringpll_l_min_value(sig, min_val) = ((sig) >= (min_val));
    `define ip2211ringpll_l_min_value(sig, min_val) ip2211ringpll_l_min_value(sig, min_val)
    let ip2211ringpll_l_same(siga, sigb) = `ip2211ringpll_SVA_LIB_SAME(siga,sigb);
    `define ip2211ringpll_l_same(siga, sigb) ip2211ringpll_l_same(siga, sigb)

`else

    `define ip2211ringpll_l_mutexed(sig)  ($onehot0({>>{sig}}) && `ip2211ringpll_SVA_LIB_KNOWN(sig))
    `define ip2211ringpll_l_at_most_bits_high(sig, n)  (($countones({>>{sig}}) <= n) && `ip2211ringpll_SVA_LIB_KNOWN(sig))
    `define ip2211ringpll_l_at_most_bits_low(sig, n)  (($countones({>>{~sig}}) <= n) && `ip2211ringpll_SVA_LIB_KNOWN(sig))
    `define ip2211ringpll_l_bits_high(sig, n)  (($countones({>>{sig}}) == n) && `ip2211ringpll_SVA_LIB_KNOWN(sig))
    `define ip2211ringpll_l_bits_low(sig, n)  (($countones({>>{~sig}}) == n) && `ip2211ringpll_SVA_LIB_KNOWN(sig))
    `define ip2211ringpll_l_same_bits(sig)  ((&(sig)) || !(|(sig)) && `ip2211ringpll_SVA_LIB_KNOWN(sig))
    `define ip2211ringpll_l_one_hot(sig)  ($onehot({>>{sig}}) && `ip2211ringpll_SVA_LIB_KNOWN(sig))
    `define ip2211ringpll_l_known_driven(sig)  `ip2211ringpll_SVA_LIB_KNOWN(sig)
    `define ip2211ringpll_l_forbidden(cond)  (!(cond))
    `define ip2211ringpll_l_must(prop)  (prop)
    `define ip2211ringpll_l_trigger(trig_sig, prop_sig) (trig_sig -> prop_sig)
    `define ip2211ringpll_l_range(sig, low, high)  (((sig) >=(low)) & ((sig) <=(high)))
    `define ip2211ringpll_l_max_value(sig, max_val)  ((sig) <= (max_val))
    `define ip2211ringpll_l_min_value(sig, min_val)  ((sig) >= (min_val))
    `define ip2211ringpll_l_same(siga, sigb)  `ip2211ringpll_SVA_LIB_SAME(siga,sigb)

`endif





// --- --- Assumption Properties --- --- //

property p_max_value(sig, max_val, clk=`ip2211ringpll_default_clk, rst=1'b0);
     @(clk) disable iff(rst) `ip2211ringpll_l_max_value(sig, max_val);
endproperty : p_max_value

property p_min_value(sig, min_val, clk=`ip2211ringpll_default_clk, rst=1'b0);
     @(clk) disable iff(rst) `ip2211ringpll_l_min_value(sig, min_val);
endproperty : p_min_value

property p_mutexed(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
     @(clk) disable iff(rst) `ip2211ringpll_l_mutexed(sig) ;
endproperty : p_mutexed

property p_one_hot(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
     @(clk) disable iff(rst) `ip2211ringpll_l_one_hot(sig);
endproperty : p_one_hot

property p_same_bits(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
     @(clk) disable iff(rst) `ip2211ringpll_l_same_bits(sig);
endproperty : p_same_bits

property p_range(sig, low, high, clk=`ip2211ringpll_default_clk, rst=1'b0);
     @(clk) disable iff(rst) `ip2211ringpll_l_range(sig, low, high);
endproperty : p_range

property p_at_most_bits_high(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
     @(clk) disable iff(rst) `ip2211ringpll_l_at_most_bits_high(sig, n);
endproperty : p_at_most_bits_high

property p_at_most_bits_low(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
     @(clk) disable iff(rst) `ip2211ringpll_l_at_most_bits_low(sig, n);
endproperty : p_at_most_bits_low

property p_bits_high(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
     @(clk) disable iff(rst) `ip2211ringpll_l_bits_high(sig, n);
endproperty : p_bits_high

property p_forbidden(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
  @(clk) disable iff(rst) `ip2211ringpll_l_forbidden(sig);
endproperty : p_forbidden

property p_must(prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
  @(clk) disable iff(rst) `ip2211ringpll_l_must(prop);
endproperty : p_must

property p_known_driven(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
  @(clk) disable iff(rst) `ip2211ringpll_l_known_driven(sig);
endproperty : p_known_driven

property p_same(siga, sigb, clk=`ip2211ringpll_default_clk, rst=1'b0);
  @(clk) disable iff(rst) `ip2211ringpll_l_same(siga, sigb);
endproperty : p_same

property p_bits_low(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk disable iff(rst) `ip2211ringpll_l_bits_low(sig, n);
endproperty : p_bits_low

//   --- --- --- Currently not supported in let statements --- --- --- //

//property one_of(sig, set, clk=`ip2211ringpll_default_clk, rst=1'b0);
//     @(clk) disable iff(rst) ((sig) inside set);
//endproperty : p_one_of

//property one_of(sig, set, clk=`ip2211ringpll_default_clk, rst=1'b0);
//     @(clk) disable iff(rst) one_of(sig, set);
//endproperty : p_one_of

// --- --- --- --- --- --- --- --- --- --- --- --- --- --- --- --- --- //




// --- --- ---Cover Properties --- --- --- //


property p_cover_mutexed(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) && `ip2211ringpll_l_mutexed(sig);
endproperty : p_cover_mutexed

property p_not_mutexed_covered(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) && !(`ip2211ringpll_l_mutexed(sig));
endproperty : p_not_mutexed_covered

property p_cover_one_hot(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) && `ip2211ringpll_l_one_hot(sig);
endproperty : p_cover_one_hot

property p_not_one_hot_cover(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) && !(`ip2211ringpll_l_one_hot(sig));
endproperty : p_not_one_hot_cover

property p_cover_same_bits(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk  !(rst) && `ip2211ringpll_l_same_bits(sig);
endproperty : p_cover_same_bits

property p_not_same_bits_cover(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk  !(rst) && !(`ip2211ringpll_l_same_bits(sig));
endproperty : p_not_same_bits_cover

property p_cover_range(sig, low, high, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk  !(rst) && `ip2211ringpll_l_range(sig, low, high);
endproperty : p_cover_range

property p_not_range_cover(sig, low, high, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk  !(rst) && !(`ip2211ringpll_l_range(sig, low, high));
endproperty : p_not_range_cover

property p_cover_at_most_bits_high(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk  !(rst) &&  `ip2211ringpll_l_at_most_bits_high(sig, n);
endproperty : p_cover_at_most_bits_high

property p_not_at_most_bits_high_cover(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk  !(rst) &&  !(`ip2211ringpll_l_at_most_bits_high(sig, n));
endproperty : p_not_at_most_bits_high_cover

property p_cover_at_most_bits_low(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk  !(rst) &&  `ip2211ringpll_l_at_most_bits_low(sig, n);
endproperty : p_cover_at_most_bits_low

property p_not_at_most_bits_low_cover(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk  !(rst) &&  !(`ip2211ringpll_l_at_most_bits_low(sig, n));
endproperty : p_not_at_most_bits_low_cover

property p_cover_bits_high(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) && `ip2211ringpll_l_bits_high(sig, n);
endproperty : p_cover_bits_high

property p_not_bits_high_cover(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) && !(`ip2211ringpll_l_bits_high(sig, n));
endproperty : p_not_bits_high_cover

property p_cover_known_driven(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) && `ip2211ringpll_l_known_driven(sig);
endproperty : p_cover_known_driven

property p_not_known_driven_cover(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) && !(`ip2211ringpll_l_known_driven(sig));
endproperty : p_not_known_driven_cover

property p_cover_same(siga, sigb, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) && `ip2211ringpll_l_same(siga, sigb);
endproperty : p_cover_same

property p_not_same_cover(siga, sigb, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) && !(`ip2211ringpll_l_same(siga, sigb));
endproperty : p_not_same_cover

property p_cover_max_value(sig, max_val, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) &&  `ip2211ringpll_l_max_value(sig, max_val);
endproperty : p_cover_max_value

property p_not_max_value_cover(sig, max_val, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) && !(`ip2211ringpll_l_max_value(sig, max_val));
endproperty : p_not_max_value_cover

property p_cover_min_value(sig, min_val, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) &&  `ip2211ringpll_l_min_value(sig, min_val);
endproperty : p_cover_min_value

property p_not_min_value_cover(sig, min_val, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) && !(`ip2211ringpll_l_min_value(sig, min_val));
endproperty : p_not_min_value_cover

property p_cover_bits_low(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) && `ip2211ringpll_l_bits_low(sig, n);
endproperty : p_cover_bits_low

property p_not_bits_low_cover(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk !(rst) &&  !(`ip2211ringpll_l_bits_low(sig, n));
endproperty : p_not_bits_low_cover


//   --- --- --- Currently not supported in let statements --- --- --- //

//property cover_one_of(sig, set, clk=`ip2211ringpll_default_clk, rst=1'b0);
//  @clk !(rst) && l_one_of(sig, set);
//endproperty : p_cover_one_of


//property not_one_of_cover(sig, set, clk=`ip2211ringpll_default_clk, rst=1'b0);
//  @clk !(rst) && !(l_one_of(sig, set));
//endproperty : p_not_one_of_cover

// --- --- --- --- --- --- --- --- --- --- --- --- --- --- --- --- --- //






// --- --- Sequential Properties --- --- //


property p_trigger(trig, prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) trig |-> prop;
endproperty : p_trigger


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_delayed_trigger(trig, delay, prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) trig |-> nexttime[delay] prop;
endproperty : p_delayed_trigger

`else

property p_delayed_trigger(trig, delay, prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) trig ##delay 1'b1 |->  prop;
endproperty : p_delayed_trigger

`endif


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_never(prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) not(strong(prop));
endproperty : p_never

`else

property p_never(prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) not(prop);
endproperty : p_never

`endif


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_eventually_holds(en, prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) en |-> s_eventually prop;
endproperty : p_eventually_holds

`else

property p_eventually_holds(en, prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) en |-> ##[0:$] prop;
endproperty : p_eventually_holds

`endif


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_between(start_ev, end_ev, cond, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) start_ev |-> cond until_with end_ev;
endproperty : p_between

`else

property p_between(start_ev, end_ev, cond, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) start_ev ##0 !(end_ev && cond)[*1:$] |-> cond;
endproperty : p_between

`endif


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_between_time(trig, start_time, end_time, cond, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) trig |-> always [start_time:end_time] cond;
endproperty : p_between_time

`else

property p_between_time(trig, start_time, end_time, cond, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst)
        trig |-> ##start_time (cond[*(end_time-start_time+1)]);
endproperty : p_between_time

`endif


// --- --- ---


property p_next_event(en, ev, prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) en ##0 ev[->1] |-> prop;
endproperty : p_next_event


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_before_event(en, first, second, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) en |-> (not strong(second)) until_with first;
endproperty : p_before_event

`else

property p_before_event(en, first, second, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) en ##0 (!first[*1:$] or first[->1]) |-> not second;
endproperty : p_before_event

`endif


// --- --- ---


property p_remain_high(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) !sig ##1 sig |=> sig[*n];
endproperty : p_remain_high


// --- --- ---


property p_remain_high_at_most(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) !sig ##1 sig |=> sig[*0:n] ##1 !sig;
endproperty : p_remain_high_at_most


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_gremain_high(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk disable iff(rst) !sig ##1 sig |=> reject_on(!sig) 1'b1[*n];
endproperty : p_gremain_high

`else

property p_gremain_high(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) 1;
endproperty : p_gremain_high

`endif


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_gremain_high_at_most(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
   @clk disable iff(rst) !sig ##1 sig |=> accept_on(!sig) ##n !sig;
endproperty : p_gremain_high_at_most

`else

property p_gremain_high_at_most(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) 1;
endproperty : p_gremain_high_at_most

`endif


// --- --- ---


property p_verify(prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) prop;
endproperty : p_verify


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_req_granted(req, gnt, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) (gnt || !req) ##1 req |-> s_eventually (gnt);
endproperty : p_req_granted

`else

property p_req_granted(req, gnt, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff (rst)
    (gnt || !req) ##1 req |-> gnt[->1];
endproperty : p_req_granted

`endif


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_cont_req_granted(req, gnt, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst)
    (gnt || !req) ##1 req |-> strong(req throughout gnt[->1]);
endproperty : p_cont_req_granted

`else

property p_cont_req_granted(req, gnt, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff (rst)
    (gnt || !req) ##1 req |-> req throughout gnt[->1];
endproperty : p_cont_req_granted

`endif


// --- --- ---


property p_req_granted_within(req, min, max, gnt, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst)
    (gnt || !req) ##1 req |-> !gnt[*min:max] ##1 gnt;
endproperty : p_req_granted_within


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_until_strong(start_ev, cond, end_ev, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst)
    start_ev |-> cond s_until end_ev;
endproperty : p_until_strong

`else

property p_until_strong(start_ev, cond, end_ev, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff (rst)
    start_ev |-> cond[*0:$] ##1 end_ev;
endproperty : p_until_strong

`endif


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_until_weak(start_ev, cond, end_ev, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disablintel_checkers_core_imp.vse iff(rst)
    start_ev |-> cond until end_ev;
endproperty : p_until_weak

`else

property p_until_weak(start_ev, cond, end_ev, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff (rst)
    start_ev ##0 (!cond || end_ev)[->1] |-> end_ev;
endproperty : p_until_weak

`endif


// --- --- ---


property p_recur_triggers(trig, n, cond, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst)
     not( !cond throughout (trig ##1 trig[->(n-1)]) );
endproperty : p_recur_triggers


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_gray_code(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst)  nexttime $onehot0(sig ^ $past(sig));
endproperty : p_gray_code

`else

property p_gray_code(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst)  ##1 $onehot0(sig ^ $past(sig));
endproperty : p_gray_code

`endif


// --- --- ---


property p_rigid(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
  @(clk) disable iff(rst) ##1 $stable(sig);
endproperty : p_rigid


// --- --- ---


property p_data_transfer(start_ev, start_data, end_ev, end_data, clk=`ip2211ringpll_default_clk, rst=1'b0);
    logic [$bits(start_data)-1:0] local_data;
    @(clk) disable iff(rst)
    (start_ev, local_data = start_data) ##0
      (end_ev or (!end_ev ##1 (!start_ev throughout end_ev[->1])))
             |-> (local_data == end_data);
endproperty : p_data_transfer



// --- --- ---


property p_cover(prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) prop;
endproperty : p_cover


// --- --- ---

`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_cover_enable(en, prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) en #-# prop;
endproperty : p_cover_enable

`else

property p_cover_enable(en, prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) 1'b0;
endproperty : p_cover_enable

`endif

// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_clock_ticking(clk);
    @($global_clock) s_eventually $changing_gclk(clk);
endproperty : p_clock_ticking

`else

`ifdef ip2211ringpll_SYS_CLK

property p_clock_ticking(clk);
    @(`ip2211ringpll_SYS_CLK) !$stable(clk)[->1];
endproperty : p_clock_ticking

`else

property p_clock_ticking(clk);
    @(clk) 1;
endproperty : p_clock_ticking

`endif

`endif

// --- --- ---


// --- --- --- Stability Properties --- --- --- //


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_stable(sig, start_ev, end_ev, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) start_ev |=> $stable(sig) until_with end_ev;
endproperty : p_stable

`else

property p_stable(sig, start_ev, end_ev, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst)
        start_ev
        ##1 !(end_ev && $stable(sig))[*1:$]
              |-> $stable(sig);
endproperty : p_stable

`endif


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_gstable_ev(sig, start_ev, end_ev, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) start_ev |->
        @($global_clock) nexttime reject_on($changed_gclk(sig)) @clk 1'b1 until_with end_ev;
endproperty : p_gstable_ev

`else

property p_gstable_ev(sig, start_ev, end_ev, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) 1;
endproperty : p_gstable_ev

`endif


// --- --- ---

`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_gstable_sig_posedge(sig, start_ev, end_ev, clk, rst=1'b0);
   @(clk) 1;
endproperty : p_gstable_sig_posedge


property p_gstable_sig_negedge(sig, start_ev, end_ev, clk, rst=1'b0);
   @(clk) 1;
endproperty : p_gstable_sig_negedge


property p_gstable_sig_edge(sig, start_ev, end_ev, clk, rst=1'b0);
   @(clk) 1;
endproperty : p_gstable_sig_edge


`else

`ifdef ip2211ringpll_SYS_CLK


property p_gstable_sig(sig, start_ev, end_ev, clk, rst=1'b0);
    start_ev ##1 clk
     ##1
       (!(clk && $past(end_ev) && ($past(sig)==$past(sig,2)))[*1:$])
             |-> ($past(sig)==$past(sig,2));
endproperty : p_gstable_sig


property p_gstable_sig_posedge(sig, start_ev, end_ev, clk, rst=1'b0);
    @(`ip2211ringpll_SYS_CLK) disable iff(rst) 
        p_gstable_sig(sig, start_ev, end_ev, $rose(clk), rst);
endproperty : p_gstable_sig_posedge


property p_gstable_sig_negedge(sig, start_ev, end_ev, clk, rst=1'b0);
    @(`ip2211ringpll_SYS_CLK) disable iff(rst) 
        p_gstable_sig(sig, start_ev, end_ev, $fell(clk), rst);
endproperty : p_gstable_sig_negedge


property p_gstable_sig_edge(sig, start_ev, end_ev, clk, rst=1'b0);
    @(`ip2211ringpll_SYS_CLK) disable iff(rst) 
        p_gstable_sig(sig, start_ev, end_ev, !$stable(clk), rst);
endproperty : p_gstable_sig_edge


`else 


property p_gstable_sig_posedge(sig, start_ev, end_ev, clk, rst=1'b0);
   @(clk) 1;
endproperty : p_gstable_sig_posedge


property p_gstable_sig_negedge(sig, start_ev, end_ev, clk, rst=1'b0);
   @(clk) 1;
endproperty : p_gstable_sig_negedge


property p_gstable_sig_edge(sig, start_ev, end_ev, clk, rst=1'b0);
   @(clk) 1;
endproperty : p_gstable_sig_edge


`endif

`endif


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_stable_window(sample, sig, win_start, win_end, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) nexttime[win_start] sample implies ##1 $stable(sig)[*win_end + win_start];
endproperty : p_stable_window

`else

sequence stable_before_s(sig, clks_before, clk);
    @(clk) ##1 $stable(sig)[*clks_before-1];
endsequence : stable_before_s

property p_stable_window(sample, sig, clks_before, clks_after, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) ##clks_before sample
        |-> stable_before_s(sig, clks_before, clk).ended ##1
                ($stable(sig)[*clks_after]);
endproperty : p_stable_window

`endif


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_gstable_window(sample, sig, win_start, win_end, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @clk disable iff(rst) nexttime[win_start] sample implies
        @($global_clock) nexttime[1] reject_on($changed_gclk(sig)) @clk 1'b1[*win_end + win_start];
endproperty : p_gstable_window

`else

property p_gstable_window(sample, sig, win_start, win_end, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) 1;
endproperty : p_gstable_window

`endif


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005


property p_stable_for(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) ##1 $changed(sig) |=> $stable(sig)[*n];
endproperty : p_stable_for

`else

property p_stable_for(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) ##1 !$stable(sig) |=> $stable(sig)[*n];
endproperty : p_stable_for

`endif


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_gstable_for(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) ##1 $changed(sig) |->
            @($global_clock) nexttime reject_on($changed_gclk(sig)) @(clk) 1'b1[*n];
endproperty : p_gstable_for

`else

property p_gstable_for(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) 1;
endproperty : p_gstable_for

`endif


// --- --- ---


property p_stable_after(sample, sig, clks_after, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) sample |=> $stable(sig)[*clks_after];
endproperty : p_stable_after


// --- --- ---


`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_gstable_after(sample, sig, clks_after, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) sample |->
        @($global_clock) nexttime reject_on($changed_gclk(sig)) @(clk) 1'b1[*clks_after];
endproperty : p_gstable_after

`else

property p_gstable_after(sample, sig, clks_after, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) 1;
endproperty : p_gstable_after

`endif


// --- --- ---



`ifndef ip2211ringpll_SVA_LIB_SVA2005

property p_gstable_between_ticks_ev(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
    @(clk) disable iff(rst) 1'b1 |-> @($global_clock) nexttime[2]
        reject_on($changed_gclk(sig)) @(clk) 1'b1;
endproperty : p_gstable_between_ticks_ev


`else

property p_gstable_between_ticks_ev(sig, clk, rst=1'b0);
    @(clk) 1;
endproperty : p_gstable_between_ticks_ev

`endif


// --- --- ---


`ifdef ip2211ringpll_SYS_CLK

property p_gstable_between_ticks_sig_posedge(sig, clk, rst=1'b0);
    @(`ip2211ringpll_SYS_CLK) disable iff(rst) ##1 !$stable(sig) |-> $rose(clk);
endproperty : p_gstable_between_ticks_sig_posedge


property p_gstable_between_ticks_sig_negedge(sig, clk, rst=1'b0);
    @(`ip2211ringpll_SYS_CLK) disable iff(rst) ##1 !$stable(sig) |-> $fell(clk);
endproperty : p_gstable_between_ticks_sig_negedge


property p_gstable_between_ticks_sig_edge(sig, clk, rst=1'b0);
    @(`ip2211ringpll_SYS_CLK) disable iff(rst) ##1 !$stable(sig) |-> !$stable(clk);
endproperty : p_gstable_between_ticks_sig_edge

`else

property p_gstable_between_ticks_sig_posedge(sig, clk, rst=1'b0);
    @(clk) 1;
endproperty : p_gstable_between_ticks_sig_posedge


property p_gstable_between_ticks_sig_negedge(sig, clk, rst=1'b0);
    @(clk) 1;
endproperty : p_gstable_between_ticks_sig_negedge


property p_gstable_between_ticks_sig_edge(sig, clk, rst=1'b0);
    @(clk) 1;
endproperty : p_gstable_between_ticks_sig_edge


`endif


//
// DEPRECATED NON-'p_' PROPERTIES
// These are only kept because some projects hard-coded internal library 
// property names from sva_lib 4.4.  Please avoid using them.
//

property req_granted(req, gnt, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_req_granted(req, gnt, clk, rst);
endproperty

property one_hot(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_one_hot(sig,clk,rst);
endproperty

property stable_window(sample, sig, win_start, win_end, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_stable_window(sample,sig,win_start,win_end,clk,rst);
endproperty

property at_most_bits_high(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_at_most_bits_high(sig, n, clk, rst);
endproperty

property delayed_trigger(trig, delay, prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_delayed_trigger(trig, delay, prop, clk, rst);
endproperty

property never(prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_never(prop,clk,rst);
endproperty

property cont_req_granted(req, gnt, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_cont_req_granted(req, gnt, clk, rst);
endproperty

property trigger(trig, prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_trigger(trig, prop, clk, rst);
endproperty

property verify(prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_verify(prop, clk, rst);
endproperty

property forbidden(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_forbidden(sig, clk, rst);
endproperty

property between(start_ev, end_ev, cond, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_between(start_ev, end_ev, cond, clk, rst);
endproperty

property stable(sig, start_ev, end_ev, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_stable(sig, start_ev, end_ev, clk, rst);
endproperty

property mutexed(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_mutexed(sig, clk, rst);
endproperty

property must(prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_must(prop, clk, rst);
endproperty

property remain_high(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_remain_high(sig, n, clk, rst);
endproperty

property remain_low(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_remain_high(!sig, n, clk, rst);
endproperty

property stable_for(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_stable_for(sig, n, clk, rst);
endproperty

property req_granted_within(req, min, max, gnt, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_req_granted_within(req, min, max, gnt, clk, rst);
endproperty

property recur_triggers(trig, n, cond, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_recur_triggers(trig, n, cond, clk, rst);
endproperty

property clock_ticking(clk);
    p_clock_ticking(clk);
endproperty

property same_bits(sig, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_same_bits(sig, clk, rst);
endproperty

property range(sig, low, high, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_range(sig, low, high, clk, rst);
endproperty

property bits_high(sig, n, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_bits_high(sig, n, clk, rst);
endproperty

property between_time(trig, start_time, end_time, cond, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_between_time(trig, start_time, end_time, cond, clk, rst);
endproperty

property next_event(en, ev, prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_next_event(en, ev, prop, clk, rst);
endproperty

property before_event(en, first, second, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_before_event(en, first, second, clk, rst);
endproperty

property cov_seq(seq, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_cover(seq, clk, rst);
endproperty

property eventually_holds(en, prop, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_eventually_holds(en, prop, clk, rst);
endproperty

property stable_after(sample, sig, clks_after, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_stable_after(sample, sig, clks_after, clk, rst);
endproperty

property until_strong(start_ev, cond, end_ev, clk=`ip2211ringpll_default_clk, rst=1'b0);
    p_until_strong(start_ev, cond, end_ev, clk, rst);
endproperty

`endif	// ip2211ringpll_INTEL_CHECKERS_CORE_IMP_VS

`ifndef ip2211ringpll_INTEL_CHECKERS_EXT_VS
`define ip2211ringpll_INTEL_CHECKERS_EXT_VS

`define ip2211ringpll_FPV_RESTRICT

`ifdef INTC_SVA_LIB_OLD_FORMAT


`define ip2211ringpll_ASSERT_MUTEXED_HW(fire, label, sig, rst)        \
	assert(1);					\
	fire = ~((rst) || `ip2211ringpll_SVA_LIB_ONEHOT0({>>{sig}}));	         \
	label``_hw: `ip2211ringpll_ASSERT_MUTEXED(sig, rst) 
    
`endif

`define ip2211ringpll_ASSERTH_MUTEXED(fire, label, sig, rst, ip2211ringpll_MSG)        \
	fire = ~((rst) || `ip2211ringpll_SVA_LIB_ONEHOT0({>>{sig}}));	         \
	`ip2211ringpll_ASSERTC_MUTEXED(label``_hw, sig, rst, ip2211ringpll_MSG)


`ifdef INTC_SVA_LIB_OLD_FORMAT

`define ip2211ringpll_ASSERT_ONE_HOT_HW(fire, label, sig, rst)	\
	assert(1);					\
	fire = ~((rst) || `ip2211ringpll_SVA_LIB_ONEHOT({>>{sig}}));		\
	label``_hw: `ip2211ringpll_ASSERT_ONE_HOT(sig,rst) 

`endif

`define ip2211ringpll_ASSERTH_ONE_HOT(fire, label, sig, rst, ip2211ringpll_MSG)	\
	fire = ~((rst) || `ip2211ringpll_SVA_LIB_ONEHOT({>>{sig}}));		\
	`ip2211ringpll_ASSERTC_ONE_HOT(label``_hw, sig, rst, ip2211ringpll_MSG)
    

`ifdef INTC_SVA_LIB_OLD_FORMAT

`define ip2211ringpll_ASSERT_SAME_BITS_HW(fire, label, sig, rst)		\
	assert(1);					\
	fire = ~((rst) || ((&(sig)) || !(|(sig))) );	\
	label``_hw: `ip2211ringpll_ASSERT_SAME_BITS(sig,rst)  

`endif

`define ip2211ringpll_ASSERTH_SAME_BITS(fire, label, sig, rst, ip2211ringpll_MSG)		\
	fire = ~((rst) || ((&(sig)) || !(|(sig))) );	\
        `ip2211ringpll_ASSERTC_SAME_BITS(label``_hw, sig, rst, ip2211ringpll_MSG)


`ifdef INTC_SVA_LIB_OLD_FORMAT

`define ip2211ringpll_ASSERT_AT_MOST_BITS_HIGH_HW(fire, label, sig, n, rst) \
	assert(1);						\
	fire = ~((rst) || (`ip2211ringpll_SVA_LIB_COUNTONES({>>{sig}}) <= n));	      \
	label``_hw: `ip2211ringpll_ASSERT_AT_MOST_BITS_HIGH(sig, n, rst) 
    
`endif
 
`define ip2211ringpll_ASSERTH_AT_MOST_BITS_HIGH(fire, label, sig, n, rst, ip2211ringpll_MSG) \
	fire = ~((rst) || (`ip2211ringpll_SVA_LIB_COUNTONES({>>{sig}}) <= n));	      \
	`ip2211ringpll_ASSERTC_AT_MOST_BITS_HIGH(label``_hw, sig, n, rst, ip2211ringpll_MSG)


`ifdef INTC_SVA_LIB_OLD_FORMAT

`define ip2211ringpll_ASSERT_BITS_HIGH_HW(fire, label, sig, n, rst )		\
	assert(1);						\
	fire = ~((rst) || (`ip2211ringpll_SVA_LIB_COUNTONES({>>{sig}}) == n));	\
	label``_hw: `ip2211ringpll_ASSERT_BITS_HIGH(sig, n, rst) 

`endif

`define ip2211ringpll_ASSERTH_BITS_HIGH(fire, label, sig, n, rst, ip2211ringpll_MSG)	\
	fire = ~((rst) || (`ip2211ringpll_SVA_LIB_COUNTONES({>>{sig}}) == n));	\
	`ip2211ringpll_ASSERTC_BITS_HIGH(label``_hw, sig, n, rst, ip2211ringpll_MSG)


`ifdef INTC_SVA_LIB_OLD_FORMAT

`define ip2211ringpll_ASSERT_FORBIDDEN_HW(fire, label, prop, rst) \
	assert (1);				\
	fire = ~((rst) || !(prop));	    \
	label``_hw: `ip2211ringpll_ASSERT_FORBIDDEN(prop, rst) 

`endif

`define ip2211ringpll_ASSERTH_FORBIDDEN(fire, label, prop, rst, ip2211ringpll_MSG) \
	fire = ~((rst) || !(prop));	    \
    `ip2211ringpll_ASSERTC_FORBIDDEN(label``_hw, prop, rst, ip2211ringpll_MSG)


`ifdef INTC_SVA_LIB_OLD_FORMAT

`define ip2211ringpll_ASSERT_MUST_HW(fire, label,  prop, rst)			\
	assert(1);						\
	fire = ~((rst) || (prop));				\
	label``_hw: `ip2211ringpll_ASSERT_MUST(prop, rst) 

`endif

`define ip2211ringpll_ASSERTH_MUST(fire, label, prop, rst, ip2211ringpll_MSG)			\
	fire = ~((rst) || (prop));				\
    `ip2211ringpll_ASSERTC_MUST(label``_hw, prop, rst, ip2211ringpll_MSG)


`ifdef INTC_SVA_LIB_OLD_FORMAT

`define ip2211ringpll_ASSERT_SAME_HW(fire, label, siga, sigb, rst)		\
	assert(1);						\
	fire = ~((rst) || ((siga) == (sigb)));		\
	label``_hw: `ip2211ringpll_ASSERT_SAME(siga, sigb, rst) 

`endif

`define ip2211ringpll_ASSERTH_SAME(fire, label, siga, sigb, rst, ip2211ringpll_MSG)		\
	fire = ~((rst) || ((siga) == (sigb)));		\
	`ip2211ringpll_ASSERTC_SAME(label``_hw, siga, sigb, rst, ip2211ringpll_MSG)



//ip2211ringpll_MCP Assertions
// these macros assume that the user adds manually the ip2211ringpll_ERR_MSG. 
//
`define ip2211ringpll_ASSERT_SIGNAL_IS_PH2(clk,sig,constr_name) \
  `ifdef INTC_FEV \
     always \
  lira_transimply_``constr_name: $transimply("$rising",clk,"$unchanging",sig);\
  `endif \
  `ip2211ringpll_ASSERTS_GSTABLE_BETWEEN_TICKS(sva_``constr_name, sig, negedge clk, 1'b0, $info("")); 


`define ip2211ringpll_ASSERT_SIGNAL_IS_PH1(clk,sig,constr_name) \
  `ifdef INTC_FEV \
     always \
  lira_transimply_``constr_name: $transimply("$falling",clk,"$unchanging",sig);\
  `endif \
  `ip2211ringpll_ASSERTS_GSTABLE_BETWEEN_TICKS(sva_``constr_name, sig, posedge clk, 1'b0, $info(""));



`ifndef INTC_SVA_LIB_DONT_SYNTHESIZE_BOOL_SF
    `define ip2211ringpll_SVA_LIB_ONEHOT    f_onehot
    `define ip2211ringpll_SVA_LIB_ONEHOT0   f_onehot0
    `define ip2211ringpll_SVA_LIB_COUNTONES f_countones 
`else
    `define ip2211ringpll_SVA_LIB_ONEHOT    $onehot
    `define ip2211ringpll_SVA_LIB_ONEHOT0   $onehot0
    `define ip2211ringpll_SVA_LIB_COUNTONES $countones 
`endif


`ifndef INTC_SVA_LIB_DONT_SYNTHESIZE_BOOL_SF

// VCS / LIRA today handle $onehot / $countones also in constraints
// RLS flow probably uses different synthesis tool, which doesn't compile
// $onehot / $countones.
// The goal of the separation is not to lose optimizations that are done 
// in the tools.

function automatic bit [2:0] f_countones_4 (input bit [3:0] i);
begin
	unique casez (i)
		4'b0001 : f_countones_4=3'b001;
		4'b0010 : f_countones_4=3'b001;
		4'b0011 : f_countones_4=3'b010;
		4'b0100 : f_countones_4=3'b001;
		4'b0101 : f_countones_4=3'b010;
		4'b0110 : f_countones_4=3'b010;
		4'b0111 : f_countones_4=3'b011;
		4'b1000 : f_countones_4=3'b001;
		4'b1001 : f_countones_4=3'b010;
		4'b1010 : f_countones_4=3'b010;
		4'b1011 : f_countones_4=3'b011;
		4'b1100 : f_countones_4=3'b010;
		4'b1101 : f_countones_4=3'b011;
		4'b1110 : f_countones_4=3'b011;
		4'b1111 : f_countones_4=3'b100;
		default : f_countones_4=3'b000;
	endcase;
end
endfunction

function automatic bit [3:0] f_countones_8 (input bit [7:0] i);
begin
	f_countones_8=f_countones_4(i[7:4])+f_countones_4(i[3:0]); // lintra s-0393
end
endfunction

function automatic bit [4:0] f_countones_16 (input bit [15:0] i);
begin
	f_countones_16=f_countones_8(i[15:8])+f_countones_8(i[7:0]); // lintra s-0393
end
endfunction

function automatic bit [5:0] f_countones_32 (input bit [31:0] i);
begin
	f_countones_32=f_countones_16(i[31:16])+f_countones_16(i[15:0]); // lintra s-0393
end
endfunction

function automatic bit [6:0] f_countones_64 (input bit [63:0] i);
begin
	f_countones_64=f_countones_32(i[63:32])+f_countones_32(i[31:0]); // lintra s-0393
end
endfunction

function automatic bit [7:0] f_countones_128 (input bit [127:0] i);
begin
	f_countones_128=f_countones_64(i[127:64])+f_countones_64(i[63:0]); // lintra s-0393
end
endfunction

function automatic bit [8:0] f_countones (input bit [255:0] i);
begin
	f_countones=f_countones_128(i[255:128])+f_countones_128(i[127:0]); // lintra s-0393
end
endfunction

function automatic bit [1:0] f_onehot_8 (input bit [7:0] i);
begin
	unique casez (i)
		8'b00000000 : f_onehot_8=2'b00;
		8'b10000000 : f_onehot_8=2'b01;
		8'b01000000 : f_onehot_8=2'b01;
		8'b00100000 : f_onehot_8=2'b01;
		8'b00010000 : f_onehot_8=2'b01;
		8'b00001000 : f_onehot_8=2'b01;
		8'b00000100 : f_onehot_8=2'b01;
		8'b00000010 : f_onehot_8=2'b01;
		8'b00000001 : f_onehot_8=2'b01;
		default     : f_onehot_8=2'b11;
	endcase;
end
endfunction

function automatic bit [1:0] f_onehot_adder (input bit [1:0] i1,i2);
begin
	unique casez ({i1,i2})
		4'b0000 : f_onehot_adder=2'b00;
		4'b0001 : f_onehot_adder=2'b01;
		4'b0100 : f_onehot_adder=2'b01;
		default : f_onehot_adder=2'b11;
	endcase;
end
endfunction

function automatic bit [1:0] f_onehot_16 (input bit [15:0] i);
begin
	f_onehot_16=f_onehot_adder(f_onehot_8(i[15:8]),f_onehot_8(i[7:0]));
end
endfunction

function automatic bit [1:0] f_onehot_32 (input bit [31:0] i);
begin
	f_onehot_32=f_onehot_adder(f_onehot_16(i[31:16]),f_onehot_16(i[15:0]));
end
endfunction

function automatic bit [1:0] f_onehot_64 (input bit [63:0] i);
begin
	f_onehot_64=f_onehot_adder(f_onehot_32(i[63:32]),f_onehot_32(i[31:0]));
end
endfunction

function automatic bit [1:0] f_onehot_128 (input bit [127:0] i);
begin
	f_onehot_128=f_onehot_adder(f_onehot_64(i[127:64]),f_onehot_64(i[63:0]));
end
endfunction

function automatic bit f_onehot (input bit [255:0] i);
begin
	bit [1:0] t;
	t=f_onehot_adder(f_onehot_128(i[255:128]),f_onehot_128(i[127:0]));
	f_onehot=((~t[1]) && t[0]);
end
endfunction

function automatic bit f_onehot0 (input bit [255:0] i);
begin
	bit [1:0] t;
	t=f_onehot_adder(f_onehot_128(i[255:128]),f_onehot_128(i[127:0]));
	f_onehot0=~t[1];
end
endfunction

`endif



// --- --- ---
//
//
// This macro was added by SKL FPV to supply eventually check in simulation
//
// ******************************************************************************************
//
// Name:   eventually holds FV - DV
// Description:
//     This assertion has diff meanings depending on environment FV or DV.
//     1. FV mode - the macro calls to the "regular" eventually macro ip2211ringpll_ASSERTS_EVENTUALLY_HOLDS and
//              checks that if a req came than eventually an ack will come
//     2. DV mode - because a simulation cannot check if sometime in the future an ack will come, 
//              this assertion checks that if a req came than an ack came in the time window of
//              0 cycles to timeout_for_dv cycles.
//              If an ack didn't came until timeout_for_dv, the assertion will fail.
//              Pay attention: when 'req' comes the assertion waits for an 'ack' to come, and 
//              ignores comming 'req' until ack comes.
//
// Arguments:
//     req              Boolean          Indication that a request is submitted.
//     ack              Boolean          Indication that an ack has been recieved.
//     timeout_for_dv   Natural-Number   timeout time.
//     
//
// Comments:
//     short description of implementation:
//         As long as the request hasn't received an ack, the request is in progress. The macro 
//         has a counter which counts all the cycles where the request is in progress.
//         if this counter reaches the value of timeout_for_dv, than the assertion fails.
//     BKM's to debug in simulation:
//         In case you want to see the counter of the macro, you have to:
//         1. Go to the call to the macro (definition of your assertion) and press "m", 
//            this will expand the macro to its implementation.
//         2. The name of the counter is "InProgressCnt". 
//            2.1 in case the assertion is not used in a loop click ctrl +w to load to wave form
//            2,2 in case it is used in a loop, you have to sepiciy which instance you want to see:
//                2.2.1 click "x" to see values of signals
//                2.2.2 right click on the index variable and choode "Specify array index"
//                2.2.3 choose a value
//                2.2.4 ctrl +w on the counter name to load it to waveform 
// Related:
//       EVENTUALLY_HOLDS
//
// Example:
//    `ip2211ringpll_ASSERTS_EVENTUALLY_HOLDS_FV_AND_DV(P_Request_will_eventully_Get_An_Ack, 
//                  req, ack, 9'b111110100, clk, rst,
//    `ip2211ringpll_ERR_MSG("FV: Req didn't received an ack back, DV: No ack during time-out of 500 cycles"));
//
// ------------------------------------------------------------------------------------------
//
//


`ifndef ip2211ringpll_FPV_RESTRICT    

`define ip2211ringpll_ASSERTS_EVENTUALLY_HOLDS_DV(name, request, acknowledge, timeout_for_dv ,clock, reset) \
    ip2211ringpll_eventually_module #(.BITS($bits(timeout_for_dv)), .TIMEOUT(timeout_for_dv))    \
    name(.ack(acknowledge), .req(request), .rst(reset),.clk(clock))

`endif

`ifdef ip2211ringpll_FPV_RESTRICT 
  `define ip2211ringpll_ASSERTS_EVENTUALLY_HOLDS_FV_AND_DV(name, req, ack, timeout_for_dv, clk, rst ,ip2211ringpll_MSG ) \
       `ip2211ringpll_ASSERTS_EVENTUALLY_HOLDS(name, req, ack, clk, rst, ip2211ringpll_MSG) 
`else
  `define ip2211ringpll_ASSERTS_EVENTUALLY_HOLDS_FV_AND_DV( name, req , ack , timeout_for_dv ,clk , rst ,ip2211ringpll_MSG ) \
       `ip2211ringpll_ASSERTS_EVENTUALLY_HOLDS_DV(name, req, ack, timeout_for_dv, clk, rst) 
`endif


// ***************************************************************************************** //
`ifndef ip2211ringpll_FPV_RESTRICT
module ip2211ringpll_eventually_module 
      #(parameter BITS = 5, parameter TIMEOUT = 32) 
      (input bit req, input bit ack, input wire clk, input bit rst);

bit             InProgress      ;
bit [BITS -1:0] InProgressCnt   ;
      
always_ff @(posedge clk or posedge rst)
begin
    if (rst || ack) 
       begin
          InProgressCnt = {BITS{1'b0}}; 
          InProgress = 1'b0;
       end
      else
       begin
          if (req)
            begin        
               InProgress = 1'b1;
            end
          InProgressCnt = InProgressCnt + InProgress;
       end
end

`ip2211ringpll_ASSERTS_NEVER(assertion_name, InProgressCnt == TIMEOUT, clk, rst, 
`ip2211ringpll_ERR_MSG("eventually_module ip2211ringpll_ERR ip2211ringpll_MSG: an ack didn't follow the req during %d cycles", TIMEOUT));

endmodule

`endif

`endif	// `ifdef ip2211ringpll_INTEL_CHECKERS_EXT_VS

`ifndef ip2211ringpll_INTEL_CHECKERS_COVERG_EXT_VS
`define ip2211ringpll_INTEL_CHECKERS_COVERG_EXT_VS

/*
 * Coverg is an SVA_LIB extension which contains covergroup-based macros.
 *
 * The SystemVerilog language provides a rich set of features for creating and
 * defining coverage specs through the utilization of the SVA cover property and
 * covergroup constructs. Although the language allows the creation of complex
 * scenarios to cover, the syntax of these constructs is often non-trivial and 
 * requires a higher-than-basic level of expertise. The coverg extension aims 
 * to provide simpler, more concise and easy-to-learn coverage spec constructs
 * that are sufficient for the vast majority of coding needs.
 *
 * These macros, when processed by any SystemVerilog-capable tool, expand to
 * standard covergroup specifications. They are not tailored to any specific
 * tool or flow, but rather are general and designed to work in any flow that
 * supports coverage collection using covergroups. Unlike the coverage macros
 * supplied in the core library, the macros supplied by this extension are 
 * covergroup-based and generally non-synthesizable by EDA tools. They are
 * handled natively by simulation tools and are synthesizable for emulation by
 * the DTS tool Jem. When code utilizing these macros is fed into FPV and
 * synthesis tools other than Jem, this extension should be disabled (as it is
 * today by default).
 *
 * Generally speaking, a coverage specification consists of a set of coverage
 * conditions. 
 * All coverage conditions are synchronized to a clocking event. 
 * The term 'coverage condition hit' refers to a specific moment in time when
 * a coverage condition is determined to be true. The tool collecting coverage
 * internally manages counters (also called bins) that accumulate the number of
 * coverage condition hits during a test execution. A specific coverage condition 
 * hits count may be incremented only at its associated clocking event.
 *
 * One of the parameters of the macros defined in this extension is
 * 'int_expr'. If the user passes a Boolean expression, then coverage conditions
 * may evaluate to either true or false, and result in a single bin being used 
 * during execution to accumulate the condition hits. On the other hand, integral
 * conditions (such as those with values of type int, packed array/struct, etc.)
 * may evaluate to multiple (integral) values, and may have one or more bins 
 * created, depending on the condition specification. Thus, for example, for an
 * enumerated variable "opcode", a single coverage condition specification may
 * be coded to separately cover the cases when it has the value OP_ADD and OP_SUB.
 *
 * The macros can be used at the module scope level, in generate constructs,
 * or in procedural initial blocks. They cannot be used inside always procedural
 * blocks.
 *
 * All extension macros may be globally enabled or disabled at compile-time, as
 * controlled by the INTC_SVA_LIB_COVERG_ENABLE macro. When compiling code that uses
 * covergroup macros, it is required to define INTC_SVA_LIB_COVERG_ENABLE for the macros
 * to take effect. This is typically done with the +define or -D command line options
 * of SystemVerilog simulators/emulator compilers. If the INTC_SVA_LIB_COVERG_ENABLE 
 * macro is not defined during compilation, all coverg extension macros expand
 * to empty text.
 *
 */


`ifndef INTC_SVA_LIB_COVER_ENABLE
  `ifdef INTC_SVA_LIB_COVERG_ENABLE
`undef  INTC_SVA_LIB_COVERG_ENABLE
`endif
`endif



// ****************************************************************************************** //
// Name:   all_values                                                             
// Category: CoverGroups                                                     
// Description:                                                                
//       Separately cover all values of an integral expression. Each possible value of the 
//       expression results with a separate bin.
// Arguments:   
//       - int_exp  expression  combinational expression of which are covered (Packed Datatype).
// Comments:                                                                   
//       - In order to clarify, the difference between ONE_OF and ALL_VALUES is as follows:
//           - ONE_OF is implemented as a cover property and covers the case where the expression 
//             has one of the values passed as an argument.
//           - ALL_VALUES is implemented as a covergroup, and the tool collecting coverage will 
//             automatically create a bin for each possible value. Coverage is collected per bin.
//       - For this macro, the 'name' argument is used as the base name of the condition. 
//         If the covered integral expression is of an enumerated type, each created bin will be
//         named <name>.val.auto[<enum_value>]. Otherwise, each created bin will be named 
//         <name>.val.auto[<integral_value>].
// Related:                                                                    
//       ONE_OF                                                               
//       ALL_VALUES_WITH_IGNORE
//       VALUES
//       VALUES_WITH_IGNORE
// Example:                                                                    
//       The following example separately covers all the values of variable imph.GfxTileTypeU267H 
//       of an enumerated type with the following possible values: TILE_LINEAR, TILE_X, TILE_Y, 
//       GTT, IOBAR. A total of five bins will be created, one per possible value of the variable,
//       which will be named imph_gfx_tile_type_hit_gtlb.val.auto[TILE_LINEAR], 
//       imph_gfx_tile_type_hit_gtlb.val.auto[TILE_X], and so on.
// 
// Code sample:
//         `ip2211ringpll_COVERG_ALL_VALUES(
//               imph_gfx_tilen_type_hit_gtlb,
//               imph.GfxTileTypeU267H,
//               posedge imph.Uclk,
//               imph.mpcohtrk.NCRadecspwrgoodU002H);
//                                     
// ------------------------------------------------------------------------------------------ //


`define ip2211ringpll_COVERG_ALL_VALUES(name, int_expr, clk, rst, DESC)                   \
    `ifndef INTC_SVA_LIB_COVERG_ENABLE                                               \
        typedef bit t_``name                                                    \
    `else                                                                       \
        (* cover_lib_macro = "COVERG_ALL_VALUES" *)                             \
        covergroup cg``name @(clk);                                                 \
            option.comment = DESC;                                              \
            name: coverpoint (int_expr) iff (!(rst));                           \
        endgroup                                                                \
        cg``name name = new                                                     \
    `endif


// ****************************************************************************************** //



// --- --- ---   



// ****************************************************************************************** //
// Name:   all_values_with_ignore                                                             
// Category: CoverGroups                                                     
// Description:                                                                
//       Separately cover all values of an integral expression, with the exception of some 
//       explicitly specified ignored values. Each possible non-ignored value is covered 
//       with a separate bin.
// Arguments:   
//       - int_exp         expression     Combinational expression values of which are covered.  
//       - ignored_values  constant-set   Set of ignored values that will not be covered.                                                  
// Comments:                                                                   
//       - In order to clarify, the difference between ONE_OF and ALL_VALUES_WITH_IGNORE is:
//           - ONE_OF is implemented as a cover property and covers the case where the expression 
//             has one of the values passed as an argument.
//           - ALL_VALUES_WITH_IGNORE is implemented as a covergroup, and the tool collecting 
//             coverage will automatically create a bin for each possible non-ignored value. 
//             Coverage is collected per bin.
//       - For this macro, the 'name' argument is used as the base name of the condition. 
//         If the covered integral expression is of an enumerated type, each created bin will be
//         named <name>.val.auto[<enum_value>]. Otherwise, each created bin will be named 
//         <name>.val.auto[<integral_value>].                                                
// Related:
//       ONE_OF
//       ALL_VALUES
//       VALUES
//       VALUES_WITH_IGNORE
// Example:                                                                    
//       The following example separately covers values of variable imph.GfxTileTypeU267H of 
//       an enumerated type with the following possible values: TILE_LINEAR, TILE_X, TILE_Y,
//       GTT, IOBAR. All values except GTT and IOBAR are covered. A total of three bins will
//       be created, one per non-ignored value of the variable, which will be named 
//          imph_gfx_tile_type_hit_gtlb.val.auto[TILE_LINEAR], 
//          imph_gfx_tile_type_hit_gtlb.val.auto[TILE_X], 
//       and so on.
// 
// Code sample:
//      `ip2211ringpll_COVERG_ALL_VALUES_WITH_IGNORE(
//          imph_gfx_tile_type_hit_gtlb,
//          imph.GfxTileTypeU267H,
//          { GTT, IOBAR },
//          posedge imph.Uclk,
//          imph.mpcohtrk.NCRadecspwrgoodU002H);
//                                           
// ------------------------------------------------------------------------------------------ //


`define ip2211ringpll_COVERG_ALL_VALUES_WITH_IGNORE(name, int_expr, ignored_values, clk, rst, DESC) \
    `ifndef INTC_SVA_LIB_COVERG_ENABLE                                               \
        typedef bit t_``name                                                    \
    `else                                                                       \
        (* cover_lib_macro = "COVERG_ALL_VALUES_WITH_IGNORE" *)                 \
        covergroup cg``name @(clk);                                                 \
            option.comment = DESC;                                              \
            name: coverpoint (int_expr) iff (!(rst))                            \
            {                                                                   \
                ignore_bins ignored = ignored_values;                           \
            }                                                                   \
        endgroup                                                                \
        cg``name name = new                                                     \
    `endif


// ****************************************************************************************** //



// --- --- ---       



// ****************************************************************************************** //
// Name:   values                                                             
// Category: CoverGroups                                                     
// Description:                                                                
//       Separately covers values of an integral expression. Each given value of the 
//       expression results with a separate bin.
// Arguments:   
//       - int_exp  expression       The Combinational expression of which are covered.  
//       - values   constant-set     Set of values that will be covered.
// Comments:                                                                   
//       - In order to clarify, the difference between ONE_OF and VALUES is as follows:
//           - ONE_OF is implemented as a cover property and covers the case where the expression 
//             has one of the values passed as an argument.
//           - VALUES is implemented as a covergroup, and the tool collecting coverage will 
//             create a bin for each given value. Coverage is collected per bin.
//             Using VALUES will result in detailed coverage per bin while using ONE_OF results
//             in total coverage result.
//       - For this macro, the 'name' argument is used as the base name of the condition. 
//         If the covered integral expression is of an enumerated type, each created bin will be
//         named <name>.val.auto[<enum_value>]. Otherwise, each created bin will be named 
//         <name>.val.auto[<integral_value>].
// Related:
//       ONE_OF
//       ALL_VALUES
//       ALL_VALUES_WITH_IGNORE
//       VALUES_WITH_IGNORE
// Example:                                                                    
//       The following example separately covers values TILE_X and TILE_Y of variable 
//       imph.GfxTileTypeU267H of an enumerated type with the following possible values: 
//       TILE_LINEAR, TILE_X, TILE_Y, GTT, IOBAR. A total of two bins will be created,
//       one per each covered value, which will be named
//            imph_gfx_tile_type_hit_gtlb.val[0], 
//            imph_gfx_tile_type_hit_gtlb.val[1].
// 
// Code sample:
//       `ip2211ringpll_COVERG_VALUES(
//           imph_gfx_tile_type_hit_gtlb,
//           imph.GfxTileTypeU267H,
//           { TILE_X, TILE_Y },
//           posedge imph.Uclk,
//           imph.mpcohtrk.NCRadecspwrgoodU002H);
//                                     
// ------------------------------------------------------------------------------------------ //



`define ip2211ringpll_COVERG_VALUES(name, int_expr, values, clk, rst, DESC)               \
    `ifndef INTC_SVA_LIB_COVERG_ENABLE                                               \
        typedef bit t_``name                                                    \
    `else                                                                       \
        (* cover_lib_macro = "COVERG_VALUES" *)                                 \
        covergroup cg``name @(clk);                                                 \
            option.comment = DESC;                                              \
            name: coverpoint (int_expr) iff (!(rst))                            \
            {                                                                   \
                bins val[] = values;                                            \
            }                                                                   \
        endgroup                                                                \
        cg``name name = new                                                     \
    `endif


// ****************************************************************************************** //



// --- --- ---  



// ****************************************************************************************** //
// Name:   values_with_ignore                                                             
// Category: CoverGroups                                                     
// Description:                                                                
//       Separately covers the given values of an integral expression, with the exception of 
//       some explicitly specified ignored values. Each given non-ignored value of the 
//       expression results with a separate bin.
// Arguments:   
//       - int_exp         expression     Combinational expression values of which are covered.                                                             
//       - values          constant-set   Set of values that will be covered.
//       - ignored_values  constant-set   Set of values that will be ignored.
// Comments:                                                                   
//       - In order to clarify, the difference between ONE_OF and ALL_VALUES_WITH_IGNORE is:
//           - ONE_OF is implemented as a cover property and covers the case where the expression 
//             has one of the values passed as an argument.
//           - ALL_VALUES_WITH_IGNORE is implemented as a covergroup, and the tool collecting 
//             coverage will automatically create a bin for each possible non-ignored value. 
//             Coverage is collected per bin.
//       - For this macro, the 'name' argument is used as the base name of the condition. 
//         If the covered integral expression is of an enumerated type, each created bin will be
//         named <name>.val.auto[<enum_value>]. Otherwise, each created bin will be named 
//         <name>.val.auto[<integral_value>].                                                
// Related:
//       ONE_OF
//       ALL_VALUES
//       ALL_VALUES_WITH_IGNORE
//       VALUES
// Example:   
//       The following example separately covers all values of variable my_var in the range [0:63],
//       except those that are a power of two. A total of 58 bins will be created, one per covered 
//       value, which will be named
//           my_var.val[0]
//           my_var.val[1] 
//       and so on up to my_var.val[57].
// 
// Code sample:
//       `ip2211ringpll_COVERG_VALUES_WITH_IGNORE(
//            not_power_of_two,
//            my_var,
//            { [0:63] },
//            { 0, 2, 4, 8, 16, 32 },
//            posedge clk,
//            ~pwrgood);                                                      
//                                                                
// ------------------------------------------------------------------------------------------ //


`define ip2211ringpll_COVERG_VALUES_WITH_IGNORE(name, int_expr, values, ignored_values, clk, rst, DESC) \
    `ifndef INTC_SVA_LIB_COVERG_ENABLE                                               \
        typedef bit t_``name                                                    \
    `else                                                                       \
        (* cover_lib_macro = "COVERG_VALUES_WITH_IGNORE" *)                     \
        covergroup cg``name @(clk);                                                 \
            option.comment = DESC;                                              \
            name: coverpoint (int_expr) iff (!(rst))                            \
            {                                                                   \
                bins val[] = values;                                            \
                ignore_bins ignored = ignored_values;                           \
            }                                                                   \
        endgroup                                                                \
        cg``name name = new                                                     \
    `endif



// ****************************************************************************************** //
`endif	// `ifdef ip2211ringpll_INTEL_CHECKERS_COVERG_EXT_VS

`ifndef ip2211ringpll_RINGPLL_MACROS_SV
`define ip2211ringpll_RINGPLL_MACROS_SV

//`ifndef VCSSIM_OR_EMU
//   `ifdef INTC_EMULATION
//      `define VCSSIM_OR_EMU
//   `endif
//`endif
//
//`ifndef VCSSIM_OR_EMU
//   `ifdef VCSSIM
//      `define VCSSIM_OR_EMU
//   `endif
//`endif

//`include "soc_macros.sv"
`ifndef ip2211ringpll_SVA_OFF
//`include "intel_checkers.sv"
`endif

`ifndef ip2211ringpll_MACRO_XDEFAULT
    `define ip2211ringpll_MACRO_XDEFAULT
    `define ip2211ringpll_XDefault(var)                                   \
        `ifndef ip2211ringpll_NO_VCSSIM                                       \
            default : var = {$bits(var){1'bx}};             \
        `endif
`endif

`ifndef INTC_NO_VCSSIM_OR_EMU

`ifndef ip2211ringpll_NHM_DUALEDGEMSFF_MODULE
`define ip2211ringpll_NHM_DUALEDGEMSFF_MODULE
module ip2211ringpll_nhm_dualedgemsff #(
   parameter DWIDTH = 1
) 
( 
   output logic [DWIDTH-1:0] qout,
   input  logic [DWIDTH-1:0] din,
   input  logic              clk
);

  // 0in set_clock clk -default
  logic clk_inv;
  logic [DWIDTH-1:0] pos_d , neg_d;
  assign clk_inv = ~clk;
  `ifndef INTC_NO_VCSSIM_OR_EMU
    `ip2211ringpll_MSFF(pos_d,din,clk) // novas s-21013 
    `ip2211ringpll_MSFF(neg_d,din,clk_inv) // novas s-51508, s-21013
    always_comb
     `ifdef INTEL_EMULATION
       qout <=  clk ? pos_d : neg_d; 
     `else 
       qout <= #1 clk ? pos_d : neg_d;  /* novas s-50523,s-23089,s-23016 */
     `endif
  `endif

endmodule
`endif
`endif

`define ip2211ringpll_DUAL_EDGE_MSFF(q,i,clock)                                                               \
`ifndef INTC_NO_VCSSIM_OR_EMU                                                                               \
  `ifdef ip2211ringpll_MACRO_ATTRIBUTE                                                                        \
    (* macro_attribute = `"DUAL_EDGE_MSFF(q``,i``,clock``)`" *)                                 \
  `endif                                                                                        \
  ip2211ringpll_nhm_dualedgemsff #(.DWIDTH($bits(q))) \demsff_``q (.qout(q),.din(i),.clk(clock));             \
`else                                                                                           \
   always_comb                                                                                  \
     $display("Error: ip2211ringpll_DUAL_EDGE_MSFF unsupported for implementation.  Please move to INST_ON"); \
`endif

///=====================================================================================================================
/// The ip2211ringpll_INST_ARG macro allows instrumentation-only signals to be used as predicate valid bits.
///=====================================================================================================================
`define ip2211ringpll_INST_ARG(valid)                                      \
`ifndef INTC_NO_VCSSIM_OR_EMU                                         \
   valid                                                     \
`else                                                        \
   1'b0                                                      \
`endif

// The ip2211ringpll_SX macro is used to SIGN-EXTEND packed data to a desired size.
`define ip2211ringpll_SX(in,sz) {{sz-$bits(in){in[$bits(in)-1]}},in}

// The ip2211ringpll_ZX macro is used to ZERO-EXTEND packed data to a desired size.  This macro is generally not needed.
// Standard verilog will zero-extend data.  However, it is included here for completeness.
`define ip2211ringpll_ZX(in,sz) {{sz-$bits(in){1'b0}},in}

// The ip2211ringpll_OX macro is used to ONES-EXTEND packed data to a desired size.
`define ip2211ringpll_OX(in,sz) {{sz-$bits(in){1'b1}},in}

///=====================================================================================================================
///
/// NON-BLOCKING ASSIGNMENT MACRO:  This macro assigns the input to the output with a non-blocking assignment.
///
///=====================================================================================================================
`ifdef INTEL_EMULATION
 `define ip2211ringpll_NB_ASSIGN(out, in)         \
    always_ff @(posedge `EMULATION_FAST_CLK)  \
         out <= in;       
 `else              
   `define ip2211ringpll_NB_ASSIGN(out, in)         \
      always_comb begin                                         \
      out <= #1 in; /* novas s-60029 */       \
       end             
   `endif                 

//=======================================================================================
// No X injection: Randomized 0 or 1 when X on signal
//  The following macro implements randomness only during a valid window. 
//  Outside the window, "in" is simply passed to "out" and Xs will propagate. 
//  The window should fully encompass the duration of Xs on "in" to avoid 
//  unnecessary glitches on "out".
//
// NOTE: Primarily meant for clocks, but can be used for data too (not recommended)
//=======================================================================================

`define ip2211ringpll_RANDOM_VAL_WHEN_X(out,in,window)                                \
   `ifndef ip2211ringpll_NO_VCSSIM                                                        \
         localparam width_``out = $bits(out);                           \
         localparam width_``in  = $bits(in);                            \
                                                                        \
         integer RANDOM_VAL_SEED_``out;                       \
         bit  [width_``out-1:0] RANDOM_VAL_``out;                       \
         always @(window) begin                                                 \
            if (window !== 1'bx) begin                                  \
               RANDOM_VAL_SEED_``out = $get_initial_random_seed;   \
               for (int j_``out=0; j_``out<width_``out; ++j_``out) begin                     \
                  RANDOM_VAL_``out[j_``out] = $dist_uniform(RANDOM_VAL_SEED_``out, 0, 1); \
               end                                                         \
            end                                                         \
         end                                                            \
                                                                        \
         bit  [width_``out-1:0] bit_``out;                              \
         logic [width_``in-1:0]  packed_``in;                           \
                                                                        \
         assign packed_``in = in;                                       \
                                                                        \
         generate begin : i_``out                                       \
            genvar i_``out;                                             \
            for(i_``out=0; i_``out<=width_``out-1; i_``out++) begin     \
               assign bit_``out[i_``out] = (packed_``in[i_``out] === 1'bX) ? RANDOM_VAL_``out[i_``out] : packed_``in[i_``out]; \
            end                                                         \
         end : i_``out                                                  \
         endgenerate                                                    \
                                                                        \
         assign out = (window)? bit_``out : in;                         \
         `else \
         assign out = in;  \
         `endif

///=====================================================================================================================
///
/// ip2211ringpll_XDefault Macros for partial case. Both Macros support Packed elements (var, exp)
/// ip2211ringpll_XDefault_Part - Drive instrumental 'X to solve 'X propagation issues in Partial Case w/o default and check for 2-value violation 
///                 uniqueness and fullness of the case
/// ip2211ringpll_XDefault_Part_Def - Drive instrumental 'X to solve 'X propagation issues in Partial Case with 2-value default. The 
///                     Macro is replacing the 2-value default

`ifndef ip2211ringpll_MACRO_XDEFAULT_PART
    `define ip2211ringpll_MACRO_XDEFAULT_PART
    `define ip2211ringpll_XDefault_Part(var,exp)                          \
        `ifndef ip2211ringpll_NO_VCSSIM                                       \
            default:  begin : \Default_``var                \
            `ifndef ip2211ringpll_SVA_OFF                                 \
            `ip2211ringpll_ASSERTC_FORBIDDEN(Illegal_Case_select,(!(^(exp) === 1'bX)),0,  \
                 `ip2211ringpll_ERR_MSG("Illegal case selector: exp = %h", exp)); \
            `endif                                          \
                           var = {$bits(var){1'bx}};        \
                      end                                   \
        `elsif INTC_LINT_ON                                      \
            default:                                        \
            (* macro_attribute = `"XDefault_Part(var``,exp``)`" *) \
            if (&exp) begin /* novas s-2050 */                                \
               {>>{var}} = {>>{{$bits(var){1'b0}}}};        \
            end                                             \
            else begin                                      \
               {>>{var}} = {>>{{$bits(var){1'b0}}}};        \
            end                                             \
         `endif
`endif

`ifndef ip2211ringpll_MACRO_XDEFAULT_PART_NAME
    `define ip2211ringpll_MACRO_XDEFAULT_PART_NAME
    `define ip2211ringpll_XDefault_Part_Name(var,exp,name)                \
        `ifndef ip2211ringpll_NO_VCSSIM                                       \
            default:  begin : \Default_``name               \
            `ifndef ip2211ringpll_SVA_OFF                                 \
            `ip2211ringpll_ASSERTC_FORBIDDEN(Illegal_Case_select,(!(^(exp) === 1'bX)),0,  \
                 `ip2211ringpll_ERR_MSG("Illegal case selector: exp = %h", exp)); \
            `endif                                          \
                           {>>{var}} = {>>{{$bits(var){1'bX}}}};  \
                      end                                   \
        `elsif INTC_LINT_ON                                      \
            default:                                        \
            (* macro_attribute = `"XDefault_Part_Name(var``,exp``,name``)`" *) \
            if (&exp) /* novas s-2050 */                                      \
               {>>{var}} = {>>{{$bits(var){1'b0}}}};        \
            else                                            \
               {>>{var}} = {>>{{$bits(var){1'b0}}}};        \
         `endif
`endif

`ifndef ip2211ringpll_MACRO_XDEFAULT_PART_DEF
    `define ip2211ringpll_MACRO_XDEFAULT_PART_DEF
    `define ip2211ringpll_XDefault_Part_Def(var,def,exp)                  \
        `ifdef INTC_LINT_ON                                      \
            default: begin                                  \
            (* macro_attribute = `"XDefault_Part_Def(var``,def``,exp``)`" *) \
            if (&exp) /* novas s-2050 */                                      \
               var = def;                                  \
            else                                            \
               var = def;                                  \
          `else                                             \
            default:  begin : \Default_``var                \
                        var = def;                          \
        `ifndef ip2211ringpll_NO_VCSSIM                                       \
                        if (^(exp) === 1'bX)                \
                                 var = {$bits(var){1'bX}};  \
        `endif                                              \
        `endif                                              \
            end
`endif

`ifndef ip2211ringpll_MACRO_XDEFAULT_PART_DEF_NAME
    `define ip2211ringpll_MACRO_XDEFAULT_PART_DEF_NAME
    `define ip2211ringpll_XDefault_Part_Def_Name(var,def,exp,name)        \
        `ifdef INTC_LINT_ON                                      \
            default: begin                                  \
            (* macro_attribute = `"XDefault_Part_Def_Name(var``,def``,exp``,name``)`" *) \
            if (&exp) /* novas s-2050 */                                      \
               var = def;                                  \
            else                                            \
                var = def;                                 \
        `else                                               \
            default:  begin : \Default_``name               \
                        var = def;                          \
        `ifndef ip2211ringpll_NO_VCSSIM                                       \
                        if (^(exp) === 1'bX)                \
                           {>>{var}} = {>>{{$bits(var){1'bX}}}};  \
        `endif                                              \
        `endif                                              \
            end
`endif
 
`ifndef ip2211ringpll_MACRO_XDEFAULT_PART_DEF_LATCH
    `define ip2211ringpll_MACRO_XDEFAULT_PART_DEF_LATCH
    `define ip2211ringpll_XDefault_Part_Def_Latch(var,def,exp,name)       \
        `ifdef INTC_LINT_ON                                      \
            default: begin                                  \
            (* macro_attribute = `"XDefault_Part_Def_Latch(var``,def``,exp``,name``)`" *) \
            if (&exp) /* novas s-2050 */                                      \
               var <= def;                                  \
            else                                            \
               var <= def;                                  \
         `else                                              \
            default:  begin                                 \
                        var <= def;                         \
        `ifndef ip2211ringpll_NO_VCSSIM                                       \
                        if (^(exp) === 1'bX)                \
                           {>>{var}} <= {>>{{$bits(var){1'bX}}}};  \
        `endif                                              \
        `endif                                              \
            end
`endif


 `define ip2211ringpll_XDefault_ENDCASE(var,exp)                               \
        endcase                                                  \
        `ifndef ip2211ringpll_NO_VCSSIM                                       \
           if (^({exp}) === 1'bX)                                \
              var = {$bits(var){1'bX}};                          \
        `elsif INTC_LINT_ON                                           \
           (* macro_attribute = `"XDefault_ENDCASE(var``,exp``)`" *) \
            if (&exp) /* novas s-60043 s-2050 */            \
               {>>{var}} = {>>{{$bits(var){1'b0}}}};        \
        `endif


 `define ip2211ringpll_XDefault_ENDIF(var,exp)                                 \
        `ifndef ip2211ringpll_NO_VCSSIM                                       \
           if (^({exp}) === 1'bX)                                \
              var = {$bits(var){1'bX}};                          \
        `elsif INTC_LINT_ON                                           \
           (* macro_attribute = `"XDefault_ENDIF(var``,exp``)`" *) \
            if (&exp) /* novas s-60043 s-2050 */            \
               {>>{var}} = {>>{{$bits(var){1'b0}}}};        \
        `endif

`endif // ip2211ringpll_RINGPLL_MACROS_SV

`ifndef ip2211ringpll_LJPLL_DFX_VH
`define ip2211ringpll_LJPLL_DFX_VH

typedef struct packed { 
      logic        base0;
      logic        base1;
      logic        val0;
      logic        val1;
} t_odcs_state ;

typedef struct packed {
  logic                  odcsenable;           // ODCS :: ODCS enable
  logic                  dualtrigswap;         // ODCS :: Swap dual trigger functions
  logic                  dualtrigen;           // ODCS :: Enable dual triggering mode
  logic                  stayinbase1;          // ODCS :: Configure FSM to stay in B1
  logic [3:0]            riseoncnt;            // ODCS :: ON counter initial value
  logic [3:0]            riseoffcnt;           // ODCS :: OFF counter initial value
  logic [4:0]            risebase0;            // ODCS :: Base0 delay code
  logic [4:0]            risebase1;            // ODCS :: Base1 delay code
  logic [4:0]            riseval0;             // ODCS :: Val0 delay code
  logic [4:0]            riseval1;             // ODCS :: Val1 delay code
  logic [3:0]            falloncnt;            // ODCS :: ON counter initial value
  logic [3:0]            falloffcnt;           // ODCS :: OFF counter initial value
  logic [4:0]            fallbase0;            // ODCS :: Base0 delay code
  logic [4:0]            fallbase1;            // ODCS :: Base1 delay code
  logic [4:0]            fallval0;             // ODCS :: Val0 delay code
  logic [4:0]            fallval1;             // ODCS :: Val0 delay code
} t_odcs_config;

typedef struct packed {
  logic                  usetaptrig;           // OPSP :: Trigger using Tap instead of ubp
  logic                  trigger;              // OPSP :: Opsp tap based trigger
  logic                  opspen;               // OPSP :: Feature enable
  logic                  finedelsel;           // OPSP :: Add 40ps
  logic [1:0]            coursedelsel;         // OPSP :: 1|2|3|4 phase selection
  logic                  drvedgesel;           // OPSP :: Select falling edge driver
} t_opsp_config;

typedef struct packed {
  logic                  odcsfalltrig;         // ODCS :: FallTrigStatus
  logic                  odcsrisetrig;         // ODCS :: RiseTrigStatus
  logic                  stmtrig;              // STM :: StmTrigSeen
  logic [4:0]            dummydldelay;         // DUMMYDL :: DLDelaySetting
  logic                  opspfallsamp;         // OPSP :: OpspFallSamp
  logic                  opsprisesamp;         // OPSP :: OpspRiseSamp
} t_odcs_status;

typedef struct packed {
  logic                  stmwren;              // STM :: Disable clock modulation; can be used to stop mod...
  logic                  usetaptrigger;        // STM :: Trigger from ClkModStart instead of ubkpoint (not...
  logic                  clkmodstop;           // STM :: Stop clock modulation
  logic                  clkmodstart;          // STM :: Start clock modulation if UseTapTrigger=1 (not en...
  logic [27:0]           modcount;             // STM :: Period of modulation in PLL output clock cycles
  logic [1:0]            modesel;              // STM :: Mode select
  logic                  stoplevel;            // STM :: Level at which clock stops
} t_stm_config;

typedef struct packed {
  logic                  usedlclk;             // reg[8]     DUMMYDL :: Use DL clk in pll FB div
  logic [4:0]            dldelayovrd;          // reg[7:3]   DUMMYDL :: Delay line override encoding
  logic                  dldelayovrden;        // reg[2]     DUMMYDL :: Select delay override setting
  logic                  dlrun;                // reg[1]     DUMMYDL :: Enable delay locking loop
  logic                  dlylineen;            // reg[0]     DUMMYDL :: Enable delay line clock only
} t_dummydl_config;

typedef struct packed {
   logic [1:0]  view_dig_out;
} t_ljpll_view_out_ifc;

typedef struct packed {
//   logic [9:0]              misc_cfg;            // SPARES! -- these are spare fuse bits routed to the HIP
   logic                    disable_run_upd;     // Disable SSC/ratio runtime updates. When this bit is set, all SSC reg writes are rejected after PLL lock.
   logic                    tight_loop;          // Tight Loop Select Bit (optional as a fuse for tight loop only PLLs) // fz_tight_loopb
   //logic                    tie_lockrst_zero;    // Force the lock reset to 0 until after sticky lock asserts // fz_lockforce
   logic                    fz_lockforce;    // Force the lock reset to 0 until after sticky lock asserts // fz_lockforce
   logic [3:0]              startup_rdac;        // Startup RDAC setting
   logic [2:0]              pfd_chop_val;        // ip2211ringpll_PFD chop value
   logic [2:0]              pfd_residual_pw;     // ip2211ringpll_PFD residual pulse width - maps to fz_pfd_pw
// logic [2:0]              fz_pfd_pw;	         // NEW - maps to pfd_residual_pw  ^^^
   logic [4:0]              cp1_trim;            // Charge pump 1 trim 	// fz_cp1trim
   logic [4:0]              cp2_trim;            // Charge pump 2 trim	// fz_cp2trim
   logic [4:0]              skadj_ctrl;          // Skew Adjust Control // fz_skadj
   logic [2:0]              fz_lockcnt;             // lock count before lock assert // fz_lockcnt
   logic [2:0]              startcnt;            // iref ramp time counter
   logic [3:0]              lockthresh;          // lock threshold setting to AIP // fz_lockthresh
   logic		    lockstickyb;         //NEW fuse: Lock detect sticky enable bar Fusedefault value = 0 // fz_lockstickyb
   logic [2:0]              iref_ctune;          // IREF course tune bits
   logic [3:0]              iref_ftune;          // IREF fine tune bits
   logic                    mash_order_plus_one; // MASH modulator order control
   logic                    lp_cp_en;            // Low power charge pump mode chicken bit
   logic [1:0]              lpf_itrim;           // SR-LPF (internal to AIP) current trim
   logic [3:0]              ro_freq_sel;         // Ring oscillator frequency control
   logic [2:0]              iref_mode;           // IREF operating mode
   logic [2:0]              cp_mode;             // CP operating mode
   logic [1:0]              sr_lpf_mode;         // SR LPF Mode
   logic [1:0]              dca_cb;              // Static DCA capacitor bank control // fz_dca_cb
   logic                    start_mode;          // 2 different start modes 0=parallel iref/vctl pulldn, 1=serial iref 1st, vctl 2nd
   logic [3:0]              vco_trim_pg;         // PG trim
   logic [2:0]              vco_trim_cb;         // CB trim
//   logic [1:0]              pvd_mode;            // PVD mode (/1, /2, /4, /8)
   logic                    tllm_en;             // tight loop lock mode enable
   logic                    tllm_prchg_mode;     // gate clock distribution during tight loop lock
   logic [1:0]              tllm_sw_latency;     // wait some cycles after distribution ungated before switching to long loop
   logic [5:0]              dca_ctrl;            // Static DCA control bits // fz_dca_ctrl
   logic                    fz_vcosel ;            //NEW fuse: ip2211ringpll_VCO select (0=low freq., 1=high freq range)
   logic                          fz_ldo_faststart;       //NEW PIN: Enables LDO fast startup mode
   logic                          fz_ldo_bypass;          //NEW PIN: Enables LDO bypass
   logic [1:0]                    fz_ldo_vinvoltsel;           //NEW PIN: set to 1 if using 1.24v ldo input
   logic                          fz_ldo_extrefsel;       //NEW PIN: Selects external voltage ref (ldo_vref)
   logic [3:0]                    fz_ldo_fbtrim;          //NEW PIN: Adjust LDO feedback divider
   logic [3:0]                    fz_ldo_reftrim;         //NEW PIN: Adjust LDO internal voltage ref
   logic [1:0]                   fz_cpnbias;        //NEW fuse: CP nbias tuning
   logic [4:0]                   fz_irefgen;    //NEW fuse: Iref current
   logic                         fz_nopfdpwrgate;   //NEW fuse: Disable ip2211ringpll_PFD power gating
   logic                         fz_lpfclksel;      //NEW fuse: LPF clock selection
   logic [1:0]                   fz_pfddly;         //NEW fuse: ip2211ringpll_PFD power gating delay section
   logic [4:0]                   fz_spare;          //NEW fuse: spare bits
   logic [5:0]                   fz_startup;    //NEW fuse: PLL startup circuit tuning
  logic [10:0]                  fz_vcotrim;        //NEW fuse: ip2211ringpll_VCO trim
} t_ljpll_fuse_ifc;

typedef struct packed {
   logic                    ovrd_enable_sel;
   logic                    ovrd_enable_val;
   logic                    ovrd_powergood_sel;
   logic                    ovrd_powergood_val;
   logic                    ovrd_bypass_sel;
   logic                    ovrd_bypass_val;
   logic                    ovrd_ratio_sel;
   logic [9:0]              ovrd_ratio_val;
   logic                    ovrd_frac_sel;
   logic [23:0]             ovrd_frac_val;
   logic                    openloop;
   logic                    adc_start;
   logic [1:0]              adc_start_cnt;
   logic [1:0]              adc_clkdiv;
   logic                    adc_freeze;
   logic                    adc_chop_en;
   logic                    adc_use_vref;
   logic [2:0]              adc_sel_in;
   logic [1:0]              view_en;
   logic [1:0]              view_ana_en;
   logic [1:0][4:0]         view_sel;
   logic                    ssc_mod_dfx_en;
   logic                    ssc_mod_dfx_trigger;
   logic [1:0]              ssc_mod_dfx_steps;
   logic [1:0]              ssc_mod_dfx_clkdiv;

   logic                    tap_fuseoverride;	 // 1= enabled, 0=disbled
//   logic [9:0]              ovrd_misc_cfg;            // SPARES! -- these are spare fuse bits routed to the HIP
//   logic                    ovrd_disable_run_upd;     // Disable SSC/ratio runtime updates. When this bit is set, all SSC reg writes are rejected after PLL lock.
   logic                    ovrd_tight_loop;          // Tight Loop Select Bit (optional as a fuse for tight loop only PLLs)
   //logic                    ovrd_tie_lockrst_zero;    // Force the lock reset to 0 until after sticky lock asserts
   logic                    ovrd_fz_lockforce;    // Force the lock reset to 0 until after sticky lock asserts
//   logic [3:0]              ovrd_startup_rdac;        // Startup RDAC setting
//   logic [2:0]              ovrd_pfd_chop_val;        // ip2211ringpll_PFD chop value
   logic [2:0]              ovrd_pfd_residual_pw;     // ip2211ringpll_PFD residual pulse width
   logic [4:0]              ovrd_cp1_trim;            // Charge pump 1 trim
   logic [4:0]              ovrd_cp2_trim;            // Charge pump 2 trim
   logic [4:0]              ovrd_skadj_ctrl;          // Skew Adjust Control
   logic [2:0]              ovrd_fz_lockcnt;             // lock count before lock assert
//   logic [2:0]              ovrd_startcnt;            // iref ramp time counter
   logic [3:0]              ovrd_lockthresh;          // lock threshold setting to AIP
   logic                    ovrd_lockstickyb;         //NEW fuse: Lock detect sticky enable bar Fusedefault value = 0
//   logic [2:0]              ovrd_iref_ctune;          // IREF course tune bits
//   logic [3:0]              ovrd_iref_ftune;          // IREF fine tune bits
   logic                    ovrd_mash_order_plus_one; // MASH modulator order control
//   logic                    ovrd_lp_cp_en;            // Low power charge pump mode chicken bit
//   logic [1:0]              ovrd_lpf_itrim;           // SR-LPF (internal to AIP) current trim
//   logic [3:0]              ovrd_ro_freq_sel;         // Ring oscillator frequency control
//   logic [2:0]              ovrd_iref_mode;           // IREF operating mode
//   logic [2:0]              ovrd_cp_mode;             // CP operating mode
//   logic [1:0]              ovrd_sr_lpf_mode;         // SR LPF Mode
   logic [1:0]              ovrd_dca_cb;              // Static DCA capacitor bank control
//   logic                    ovrd_start_mode;          // 2 different start modes 0=parallel iref/vctl pulldn, 1=serial iref 1st, vctl 2nd
//   logic [3:0]              ovrd_vco_trim_pg;         // PG trim
//   logic [2:0]              ovrd_vco_trim_cb;         // CB trim
//   logic [1:0]              ovrd_pvd_mode;            // PVD mode (/1, /2, /4, /8)
   logic                    ovrd_tllm_en;             // tight loop lock mode enable
//   logic                    ovrd_tllm_prchg_mode;     // gate clock distribution during tight loop lock
//   logic [1:0]              ovrd_tllm_sw_latency;     // wait some cycles after distribution ungated before switching to long loop
   logic [5:0]              ovrd_dca_ctrl;            // Static DCA control bits

   // Brought in to over write via TAP
   //
   logic [1:0]                   ovrd_fz_cpnbias;        //NEW fuse: CP nbias tuning
   logic [4:0]                   ovrd_fz_irefgen;    //NEW fuse: Iref current
   logic                         ovrd_fz_nopfdpwrgate;   //NEW fuse: Disable ip2211ringpll_PFD power gating
   logic [2:0]                   ovrd_fz_pfd_pw;	    // NEW
   logic                         ovrd_fz_lpfclksel;      //NEW fuse: LPF clock selection
   logic [1:0]                   ovrd_fz_pfddly;         //NEW fuse: ip2211ringpll_PFD power gating delay section
   logic [4:0]                   ovrd_fz_spare;          //NEW fuse: spare bits
   logic [5:0]                   ovrd_fz_startup;    //NEW fuse: PLL startup circuit tuning
   logic                         ovrd_fz_vcosel;    //NEW fuse: ip2211ringpll_VCO sel 
   logic [10:0]                  ovrd_fz_vcotrim;        //NEW fuse: ip2211ringpll_VCO trim

   logic                         ovrd_ldo_enable;             //new -nd
   logic [1:0]                   ovrd_fz_ldo_vinvoltsel;      //new -nd
   logic                         ovrd_fz_ldo_bypass;          //new -nd
   logic                         ovrd_fz_ldo_extrefsel;       //new -nd
   logic                         ovrd_fz_ldo_faststart;       //new -nd
   logic [3:0]                   ovrd_fz_ldo_fbtrim;          //new -nd
   logic [3:0]                   ovrd_fz_ldo_reftrim;         //new -nd
   logic [5:0]                   ovrd_mdiv_ratio;             //new -nd
   logic [1:0]                   ovrd_vcodiv_ratio;           //new -nd
   logic [9:0]                   ovrd_zdiv0_ratio;            //new -nd
   logic                         ovrd_zdiv0_ratio_p5;         //new -nd
   logic [9:0]                   ovrd_zdiv1_ratio;            //new -nd
   logic                         ovrd_zdiv1_ratio_p5;         //new -nd
   logic			 start_measurement;	      //new -nd

   logic                         ta_ldo_hiz_debug;            //new -nd
   logic                         ta_ldo_idq_debug;            //new -nd
   logic [4:0]                   ta_spare;                    //NEW TAP: spare bits

   logic			 ta_openloop2;                 //new -nd
   logic [3:0]                   ta_vctlrdac;                  //new -nd


   // IDV interface
 //  logic                         ovrd_idvdisable_bi;          // new -nd
 //  logic                         ovrd_idvfreqai;              // new -nd
 //  logic                         ovrd_idvfreqbi;              // new -nd
 //  logic                         ovrd_idvpulsei;              // new -nd
 //  logic                         ovrd_idvvtclki;              // new -nd
 //  logic                         ovrd_idvvtctrli;             // new -nd
 //  logic                         ovrd_idvtdi;                 // new -nd
 //  logic                         ovrd_idvtresi;               // new -nd
 //  logic                         ovrd_clkidvih;               // new -nd
 //  logic                         ovrd_pllen;                  // new -nd

   //t_stm_config             stm_config;
   //t_odcs_config            odcs_dig_config;
   //t_dummydl_config         odcs_dll_config;
   //t_opsp_config            opsp_config;
   //logic [1:0]              odcs_tuner_cb;
} t_ljpll_tap_in_ifc;

typedef struct packed {
   logic [7:0]   ssc_ratio_step;
   logic [23:0]  ssc_frac_step;
   logic         ssc_en;              // SSC enable bit
   logic [1:0]   ssc_mode;            // SSC spread mode (upspread/downspread/centerspread)
   logic [8:0]   ssccyctopeakm1;     
} t_ljpll_reg_ifc;

typedef struct packed {
   logic idvtclki;
   logic idvtdi;
   logic idvtresi;
   logic idvtctrli;
   logic idvdisable_bi;
   logic idvfreqai;
   logic idvfreqbi;
   logic idvpulsei;
} t_ljpll_idv_in_ifc;

typedef struct packed {
   logic idvtclko;
   logic idvtdo;
   logic idvtreso;
   logic idvtctrlo;
   logic idvdisable_bo;
   logic idvfreqao;
   logic idvfreqbo;
   logic idvpulseo;
} t_ljpll_idv_out_ifc;

typedef struct packed {
   logic OdcsActTrigM736H;
   logic AnalogActTrigM736H;
} t_ljpll_odcs_trig_ifc;

typedef struct packed {
   logic         pll_enable;
   logic         dist_pwr_good;
   logic         iref_done;
   logic         pfd_en;
   logic [1:0]   unlock_count;
   logic [11:0]  lock_time;
   logic [9:0]   pll_ratio;
   logic         pll_half_int;
   logic         lock;
   logic         raw_lock;
   logic [9:0]   adc_dig_out;
   logic         adc_start;
   logic         adc_done;
   logic         ssc_mod_dfx_run;
   logic         ssc_mod_dfx_trig;
   logic [1:0]   tctrlfsmstate;
   logic [14:0]  view_freq_count;
   //t_odcs_status odcs;
} t_ljpll_tap_out_ifc;

typedef struct packed {
   t_ljpll_fuse_ifc    fuse;
   t_ljpll_reg_ifc     register;
   t_ljpll_tap_in_ifc  tap;
   t_ljpll_idv_in_ifc  idv; // Is directly used
   t_ljpll_odcs_trig_ifc odcs;
   logic                 ip2211ringpll_global_align;
   logic                 ssc_prof_update_req;
   logic                 ratio_update_req;
} t_ljpll_dfx_in_ifc;

typedef struct packed {
   t_ljpll_view_out_ifc view;
//   t_ljpll_tap_out_ifc  tap;
   t_ljpll_idv_out_ifc  idv; //Is directly used
   logic                ssc_prof_update_ack;
   logic                ratio_update_ack;
} t_ljpll_dfx_out_ifc;

`endif	// `ifdef ip2211ringpll_LJPLL_DFX_VH

`ifndef ip2211ringpll_TCU_TPSB_STAP_DATA_REG_SV 
`define ip2211ringpll_TCU_TPSB_STAP_DATA_REG_SV 

module ip2211ringpll_tcu_tpsb_stap_data_reg
   #(
   parameter DATA_REG_STAP_SIZE_OF_EACH_TEST_DATA_REGISTER           = 1,
   parameter DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS       = 0
   )
   (
   input  logic                                                         sync_reset,
   input  logic                                                         ftap_tck,
   input  logic                                                         ftap_tdi,
   input  logic                                                         reset_b,
   input  logic                                                         stap_irdecoder_drselect,
   input  logic                                                         stap_fsm_capture_dr,
   input  logic                                                         stap_fsm_shift_dr,
   input  logic                                                         stap_fsm_update_dr,
   input  logic [(DATA_REG_STAP_SIZE_OF_EACH_TEST_DATA_REGISTER - 1):0] tdr_data_in,
   output logic                                                         data_reg_tdo,
   output logic [(DATA_REG_STAP_SIZE_OF_EACH_TEST_DATA_REGISTER - 1):0] tdr_data_out
   );

   // *********************************************************************
   // Localparameters
   // *********************************************************************
   localparam HIGH = 1'b1;
   localparam LOW  = 1'b0;

   // *********************************************************************
   // Internal Signals
   // *********************************************************************
   logic [(DATA_REG_STAP_SIZE_OF_EACH_TEST_DATA_REGISTER - 1):0] shift_register;

   // *********************************************************************
   // shift register implementation - the value of tdi pin will come to this
   // reg during shift_DR state. Implementation support single bit register
   // *********************************************************************
   generate
      if (DATA_REG_STAP_SIZE_OF_EACH_TEST_DATA_REGISTER > 1)
      begin:generate_tdr_shift_capture
         always_ff @(posedge ftap_tck or negedge reset_b)
         begin
            if (!reset_b)
            begin
               shift_register <= DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS;
            end
            else if (sync_reset)
            begin
               shift_register <= DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS;
            end
            else if (stap_fsm_capture_dr & stap_irdecoder_drselect)
            begin
               shift_register <= tdr_data_in;
            end
            else if (stap_fsm_shift_dr & stap_irdecoder_drselect)
            begin
               shift_register <= {ftap_tdi, shift_register[(DATA_REG_STAP_SIZE_OF_EACH_TEST_DATA_REGISTER - 1):1]};
            end
         end
      end
      else
      begin:generate_tdr_shift_capture
         always_ff @(posedge ftap_tck or negedge reset_b)
         begin
            if (!reset_b)
            begin
               shift_register <= DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS;
            end
            else if (sync_reset)
            begin
               shift_register <= DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS;
            end
            else if (stap_fsm_capture_dr & stap_irdecoder_drselect)
            begin
               shift_register <= tdr_data_in;
            end
            else if (stap_fsm_shift_dr & stap_irdecoder_drselect)
            begin
               shift_register <= ftap_tdi;
            end
         end
      end
   endgenerate

   // *********************************************************************
   // Bit0 is assigned to data_reg_tdo and this is going to the TDOmux FUB.
   // *********************************************************************
   assign data_reg_tdo = shift_register[0];

   // *********************************************************************
   // parallel register implementation - the value will be updated to parallel
   // reg during update_DR state and negedge of tck
   // *********************************************************************


logic tup_treg;
logic ftap_tck_gated;
assign tup_treg = stap_irdecoder_drselect & stap_fsm_update_dr ; 
 
//ctech_dlat clk_gate_tdr_data_out_reg_latch_sh   ( .clkout(ftap_tck_gated),  .clk(ftap_tck), .en(tup_treg), .te(1'b0)); 
`ip2211ringpll_CLKGATE_TE(ftap_tck_gated, ftap_tck, tup_treg, 1'b0)
   always_ff @(negedge ftap_tck or negedge reset_b)
   begin
      if (!reset_b)
      begin
         tdr_data_out[103:0] <= DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS ;
      end
      else if (sync_reset)
      begin
         tdr_data_out[103:0]  <= DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS ;
      end
      else if (stap_fsm_update_dr & stap_irdecoder_drselect)
      begin
         tdr_data_out[103:0]  <= shift_register [103:0];
      end
   end
always_ff @(negedge ftap_tck_gated or negedge reset_b)
   begin
      if (!reset_b)
      begin
         tdr_data_out[104] <= DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS ;
      end
      else if (sync_reset)
      begin
         tdr_data_out[104]  <= DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS ;
      end
      else if (stap_fsm_update_dr & stap_irdecoder_drselect)
      begin
         tdr_data_out[104]  <= shift_register [104];
      end
   end
always_ff @(negedge ftap_tck or negedge reset_b)
   begin
      if (!reset_b)
      begin
         tdr_data_out[126:105] <= DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS ;
      end
      else if (sync_reset)
      begin
         tdr_data_out[126:105]  <= DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS ;
      end
      else if (stap_fsm_update_dr & stap_irdecoder_drselect)
      begin
         tdr_data_out[126:105]  <= shift_register [126:105];
      end
   end
always_ff @(negedge ftap_tck_gated or negedge reset_b)
   begin
      if (!reset_b)
      begin
         tdr_data_out[129:127] <= DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS ;
      end
      else if (sync_reset)
      begin
         tdr_data_out[129:127]  <= DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS ;
      end
      else if (stap_fsm_update_dr & stap_irdecoder_drselect)
      begin
         tdr_data_out[129:127]  <= shift_register [129:127];
      end
   end
always_ff @(negedge ftap_tck or negedge reset_b)
   begin
      if (!reset_b)
      begin
         tdr_data_out[268:130] <= DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS ;
      end
      else if (sync_reset)
      begin
         tdr_data_out[268:130]  <= DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS ;
      end
      else if (stap_fsm_update_dr & stap_irdecoder_drselect)
      begin
         tdr_data_out[268:130]  <= shift_register [268:130];
      end
   end


// Assertions and coverage
`ifndef INTC_DFX_FPV_ENABLE
   `ifdef INTEL_SIMONLY     //  Pragma no longer supported /   /synopsys translate_off
`else
   //\\`ifdef INTEL_SIMONLY     //  Pragma no longer supported /   /synopsys translate_off /  / synopsys translate_off  note:1
`endif

   // Assertions and coverage
 //  //`include "tcu_tpsb_stap_data_reg_include.sv"

`ifndef INTC_DFX_FPV_ENABLE
   `endif     //  Pragma no longer supported /   / synopsys translate_on
`else
   //\\`ifdef INTEL_SIMONLY     //  Pragma no longer supported / / synopsys translate_on
`endif

endmodule
`endif
	// `ifdef ip2211ringpll_tcu_tpsb_stap_data_reg


//`define ip2211ringpll_SVA_LIB_SVA2005
//`define ip2211ringpll_UPF

`ifndef ip2211ringpll_cpaclkphdelana_SV
`define ip2211ringpll_cpaclkphdelana_SV

//`ifndef VCSSIM_OR_EMU
//   `ifdef INTC_EMULATION
//      `define VCSSIM_OR_EMU
//   `endif
//`endif
//
//`ifndef VCSSIM_OR_EMU
//   `ifdef VCSSIM
//      `define VCSSIM_OR_EMU
//   `endif
//`endif

`ifndef INTC_NO_VCSSIM_OR_EMU
   //`include "soc_macros.sv"
`endif

module ip2211ringpll_cpaclkphdelana (
  //  vccxx is a powerpin   input  wire  vccxx,
   input  logic rst,
   input  logic cueh,
   input  logic clkin,
   output logic clkoutb
);


`ifndef INTC_NO_VCSSIM_OR_EMU
   // NOTE: MH_b = clkout high phase (!clkoutb)
   //
   logic ClkInMH;
   logic ClkInMH_b;
   logic UseInvClkMH_b;
   logic EnInvClkMH_b;
   logic EnInvClkMH, EnClkML;
   logic overlap_pulse;
   // This implementation more closely represents the hardware
   //
   `ip2211ringpll_ASYNC_RST_MSFF(UseInvClkMH_b, !UseInvClkMH_b, cueh, rst)

   // This implementation is timeable since cueh is generated on negedge
   // clkoutb (posedge clkout).
   //
   //`ip2211ringpll_ASYNC_RST_MSFF_P(UseInvClkMH_b, (CuehEdgeMH_b ^ UseInvClkMH_b), clkoutb, rst)

   // In the worst case, there is a phase path between clkoutb and clkin
   // (both flops have a phase path) so the circuit can be timed with the
   // above flop stamped on both clocks.
   //
   // This circuit
   // ensures that the enables for clk and ip2211ringpll_clkinv are staged such that
   // there is guaranteed to be a phase overlap in order to insert a phase
   // during clock switching.
   //
   `ip2211ringpll_ASYNC_RST_MSFF_P(EnClkML,       UseInvClkMH_b, clkin, rst)
   `ip2211ringpll_ASYNC_RST_MSFF  (EnInvClkMH_b,  UseInvClkMH_b, clkin, rst)
   assign EnInvClkMH = !EnInvClkMH_b;
assign overlap_pulse = EnClkML & EnInvClkMH; 
   // Gating clock and ip2211ringpll_clkinv
   //   Clk and ClkInv enables are always guaranteed to be opposite except
   //   during switching (when both are enabled for 1 phase)
   //
   assign ClkInMH   = clkin && EnClkML;
   assign ClkInMH_b = !clkin && EnInvClkMH;


   // OR clkin gated and clkin_b gated
   //
   assign clkoutb = ClkInMH | ClkInMH_b | overlap_pulse;
`endif


endmodule

`endif


`ifndef ip2211ringpll_IP22_ip2211ringpll_cpafdivcore_SV
`define ip2211ringpll_IP22_ip2211ringpll_cpafdivcore_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
`ifndef ip2211ringpll_SVA_OFF
   //`include "intel_checkers.sv"
`endif

module ip2211ringpll_ip2211ringpll_cpafdivcore 
//#( parameter     RATIO_BITS = 10)
(
   //input  logic [8:0]   ratio2x,
   input  logic [10:0]   ratio2x,
   input  logic         clkinb,
   output logic         clkout,
   output logic         cueh,
   output logic         rstd,
   input  logic         rst
);

///========================================================================================================
/// Reset Generation
///========================================================================================================

   logic RstCntMH;

   // Rename reset
   //
   always_comb RstCntMH = rst;


   // Reset to ip2211ringpll_cpaclkphdelana
   //
   always_comb rstd = rst;


///========================================================================================================
/// Reload Logic
///========================================================================================================

   logic [6:0] CountMH;
   logic Clk0MH;
   logic ReloadMH;
   logic CountToZeroMH;
   logic RatioOddMH;
   logic Zero61MH;
   logic Zero63MH;
   logic HiPhaseMH; // indicates whether divider is currently outputing clkout=1

   // More readable name for Odd ratio
   //
   always_comb RatioOddMH = ratio2x[1];

   // Compute the segmented zero values to execute a reload
   //
   always_comb begin : ZERO_CALCULATION
      Zero61MH = (CountMH[6:1] == 6'd0);
      Zero63MH = (CountMH[6:3] == 4'd0);
   end : ZERO_CALCULATION

   always_comb begin : RELOAD
      // Determine whether or not to count to zero on a reload
      //   Changes between 0/1 every cycle when the ratio is odd.
      //
      CountToZeroMH = (!HiPhaseMH && RatioOddMH);

      // Reload the counter based on the count to zero flag.
      //   If counting to zero, wait until counter matches zero,
      //   else reload at one.
      //
      ReloadMH = (CountToZeroMH) ? (CountMH == 7'd0) :
                                   (CountMH <= 7'd1) ;

   end : RELOAD

///========================================================================================================
/// Segmented 1+2+4 Reloadable Counter
///========================================================================================================

   logic [1:0] CountM1Nxt21MH;
   logic [3:0] CountM1Nxt63MH;
   logic [6:0] CountStartMH;
   logic [6:0] RatioD2MH;
   logic [6:0] CountNxtMH;
   logic       Clk21MH, Clk63MH;
   logic       EnClk21MH, EnClk63MH;
   logic       EnClk21ML, EnClk63ML;

   `ip2211ringpll_CLK_NOR(Clk0MH, clkinb, 1'b0)


   // Segmented counter declaration
   //
   `ip2211ringpll_RST_MSFF(CountMH[0],   CountNxtMH[0],   Clk0MH,  RstCntMH)
   `ip2211ringpll_RST_MSFF(CountMH[2:1], CountNxtMH[2:1], Clk21MH, RstCntMH)
   `ip2211ringpll_RST_MSFF(CountMH[6:3], CountNxtMH[6:3], Clk63MH, RstCntMH)

   always_comb EnClk21MH = (~( CountMH[0]  ) || ReloadMH);
   always_comb EnClk63MH = (~(|CountMH[2:0]) || ReloadMH);

   // Count Clock Generation
   //
   `ip2211ringpll_LATCH(EnClk21ML, EnClk21MH, clkinb)
   `ip2211ringpll_LATCH(EnClk63ML, EnClk63MH, clkinb)

   `ip2211ringpll_CLK_NOR(Clk21MH, clkinb, ~EnClk21ML)
   `ip2211ringpll_CLK_NOR(Clk63MH, clkinb, ~EnClk63ML)

   // Count start is ratio / 2
   //
   //always_comb CountStartMH    = ratio2x[8:2];
   always_comb CountStartMH    = ratio2x[8:2];

   always_comb begin : COUNT_NXT

      CountM1Nxt21MH = (CountMH[2:1] - 2'b01);
      CountM1Nxt63MH = (CountMH[6:3] - 4'b0001);

      CountNxtMH[0]   = (ReloadMH) ? CountStartMH [0]  :
                                     ~CountMH[0]       ;

      CountNxtMH[2:1] = (Zero61MH) ? CountStartMH [2:1] :
                                     CountM1Nxt21MH     ;

      CountNxtMH[6:3] = (Zero63MH) ? CountStartMH [6:3] :
                                     CountM1Nxt63MH     ;

   end : COUNT_NXT


///========================================================================================================
/// Output Clock
///========================================================================================================

   logic PhaseStretchML;

   // Every reload changes the output state of the divider clkout
   //  Since the counter uses /2 ratio value, this serves as a toggle flop
   //  for the state of the output clock.
   //
   `ip2211ringpll_EN_RST_MSFF(HiPhaseMH, ~HiPhaseMH, Clk0MH, ReloadMH, RstCntMH)

   // For odd ratios, we need to phase stretch
   //
   `ip2211ringpll_LATCH_P(PhaseStretchML, HiPhaseMH, Clk0MH)

   always_comb begin : CLKOUT
      clkout = (PhaseStretchML & RatioOddMH) || HiPhaseMH;
   end : CLKOUT

///========================================================================================================
/// Pulse extention logic
///========================================================================================================

   logic ForceSwStateLowMH;

   // For powerup, force a low state until everything factoring into the
   //   cueh signal is stable.
   //
   `ip2211ringpll_ASYNC_SET_LATCH(ForceSwStateLowMH, 1'b0, HiPhaseMH, rst)

   // Switch the clock state (clkinb) when we are in half int mode and
   //   clkout is 0 (switch every cycle)
   //
   always_comb begin : CLKIN_STATE_SELECT
      cueh = ForceSwStateLowMH ? 1'b0                    :
                                 ratio2x[0] & ~HiPhaseMH ;
   end : CLKIN_STATE_SELECT


///========================================================================================================
/// Assertions
///========================================================================================================

   `ifndef ip2211ringpll_SVA_OFF
	// IP22: It is ok for have div value 0 or 1 so commenting out. -
      //`ip2211ringpll_ASSUMEC_MUST(A_ratio_gte_2,
      //              //(ratio2x[8:1] >= 8'd2),
      //              (ratio2x[10:1] >= 10'd2),
      //              (rst!==1'b0),
      //              `ip2211ringpll_ERR_MSG("[PLL-AIP] F-divider ratio must be set >=2"));

      `ip2211ringpll_ASSERTC_FORBIDDEN(R_fdiv_core_reload_only_when_count_lte_1,
                         (ReloadMH & (CountMH > 7'd1)),
                         (rst!==1'b0),
                         `ip2211ringpll_ERR_MSG("[PLL-AIP] F-divider reloaded its internal counter unexpectedly. The counter should only reload when Count<=1"));
   `endif

endmodule

`endif

`ifndef ip2211ringpll_IP22_CPAFDIVTOP_SV
`define ip2211ringpll_IP22_CPAFDIVTOP_SV

//`include "ip2211ringpll_cpaclkphdelana.sv"
//`include "ip2211ringpll_cpafdivcore.sv"
//`include "soc_macros.sv"

//module ip2211ringpll_ip2211cpafdivtop 
//#( parameter     RATIO_BITS = 10)
// to match postdividers module w,r,t netlist 
module ip2211ringpll_ip2211cpafdivtop 
//#( parameter     ratio_bits = 10)
(
   input  logic         clkin,
   input  logic         rst,
   input  logic [10:0]   ratio2x,
//
 input logic 		enb,
    
  
   output logic         clkout,
  //added by  
   output logic 	divbygt1

 
);


   logic cueh;
   logic clkinb;
   logic rstd;
 logic clkdiv;
logic divby0or1;
logic n1;
logic n2;
logic enbi;
logic en;
logic endivclk;
logic divby1;
logic clktodiv;
logic reset_sync;
logic reset_sync_b;
logic zdiv_sync_rst;
assign en = ~enb ;
assign enbi = ~en ;
assign endivclk = en & divbygt1 ; 
assign divbygt1 = ~divby0or1 ;
assign divby0or1 = ~ (enbi | n1 | n2 | (ratio2x[10]) ) ;
assign n1 = (ratio2x[9]) |  (ratio2x[8]) |  (ratio2x[7]) |  (ratio2x[6])  ;
assign n2 = (ratio2x[5]) |  (ratio2x[4]) |  (ratio2x[3]) |  (ratio2x[2])  ;

assign clktodiv = endivclk & clkin ; 
 assign clkout = divby1 ? clkin : clkdiv ;
assign divby1 = (ratio2x[1]) & divby0or1;  



   // Phase delay insertion for half integer ratios
   //
   ip2211ringpll_cpaclkphdelana phdel_core (
      //.vccxx   ( 1'b1    ),
      .rst     ( rstd    ),
      .cueh    ( cueh    ),
      .clkin   ( clktodiv   ),
      .clkoutb ( clkinb  )
   );
   
   // F-divider counter cores for integer logic
   //
   ip2211ringpll_cpafdivcore    fdiv_core ( .clkout(clkdiv),
                                            .rst(zdiv_sync_rst),
				.*); 

   //ip2211ringpll_ip2211ringpll_cpafdivcore    fdiv_core (.*);

     `ip2211ringpll_ASYNC_SET_2MSFF_META(zdiv_sync_rst,1'b0,clkin,rst )

endmodule

//added to match refclkdiv heirarchy to netlist 

module ip2211ringpll_ip2211cpafdivtop_refclk 
(
input logic clkin ,
input logic fz_tight_loopb,
input  logic         rst,
input  logic [5:0] mdiv_ratio ,

output logic         clkout
);

logic clktodiv_1;
logic clkin_1 ;
logic selnot ;
logic tightloopnor ;
logic divbygt1;

assign clktodiv_1 = selnot ? clkin :clkin_1 ;
assign clkin_1 = clkin & tightloopnor ;
assign tightloopnor = ~ (fz_tight_loopb | divbygt1) ;
assign selnot = ~ tightloopnor ;     

 logic cueh;
   logic clkinb;
   logic rstd;
 logic clkdiv;
logic divby0or1;
logic n1;
logic n2;
logic enbi;
logic enb;
logic en;
logic endivclk;
logic divby1;
logic clktodiv;
logic reset_sync;
logic reset_sync_b;
logic [10:0]   ratio2x;
logic ratio2x_1;
assign enb = 1'b0 ;
assign en = ~enb ;
assign enbi = ~en ;
assign endivclk = en & divbygt1 ; 
assign divbygt1 = ~divby0or1 ;
assign divby0or1 = ~ (enbi | n1 | n2 | (ratio2x[10]) ) ;
assign n1 = (ratio2x[9]) |  (ratio2x[8]) |  (ratio2x[7]) |  (ratio2x[6])  ;
assign n2 = (ratio2x[5]) |  (ratio2x[4]) |  (ratio2x[3]) |  (ratio2x[2])  ;

assign clktodiv = endivclk & clktodiv_1 ; 
assign clkout = divby1 ? clktodiv_1 : clkdiv ;
assign divby1 = (ratio2x[1]) & divby0or1;

 

assign ratio2x_1 = (~ divbygt1) | (mdiv_ratio[0]) ;
assign ratio2x = ({1'b0,1'b0,1'b0,1'b0,mdiv_ratio[5],mdiv_ratio[4],mdiv_ratio[3],mdiv_ratio[2],mdiv_ratio[1],ratio2x_1,1'b0 }) ;




// Phase delay insertion for half integer ratios
   //
   ip2211ringpll_cpaclkphdelana phdel_core (
      //.vccxx   ( 1'b1    ),
      .rst     ( rstd    ),
      .cueh    ( cueh    ),
      .clkin   ( clktodiv   ),
      .clkoutb ( clkinb  )
   );
   
   // F-divider counter cores for integer logic
   //
   ip2211ringpll_cpafdivcore    fdiv_core ( .clkout(clkdiv),
				.*); 

   //ip2211ringpll_ip2211ringpll_cpafdivcore    fdiv_core (.*);


endmodule

`endif



`ifndef ip2211ringpll_CLKGEN_SV
`define ip2211ringpll_CLKGEN_SV
module ip2211ringpll_clkgen 
//#(parameter RATIO_BITS = 10)
(
   input  logic clk_ref,
   input  logic enable,
   input  logic [9:0] ratio,
   input  logic                     half_int,
   output bit clk_out
);

int T1, T2, ref_period;
logic en_calc;

always @(enable) begin : ENABLE_BLOCK
   if (enable === 1'b1) begin
      T1 = $realtime;
      en_calc <= 1'b1;
   end
   else begin
      en_calc <= 1'b0;
   end
end : ENABLE_BLOCK

always @(posedge clk_ref) begin
   if (en_calc) begin
      T2 = $realtime;
      ref_period = (T2 - T1);
      T1 = T2;
      gen_clk(ref_period, ratio, half_int);
   end else begin
      clk_out = 1'b0;
   end
end


task gen_clk;
   // Input variables are ref period and ratio
   input int ref_period_samp;
   input logic [9:0] ratio_samp;
   input logic half_int_samp;

   // Local variables
   //
   int toggle_repeat;
   int sum_until_now;
   int phase_number;
   int effective_ref_period;
   int clk_out_phase;
      
   toggle_repeat = (ratio_samp << (1-half_int_samp)) - 1;
   effective_ref_period = (ref_period_samp << half_int_samp);
   sum_until_now = 0;
   phase_number = 1;
  
   // Generate initial edge
   //
   clk_out = ~clk_out;
   
   repeat (toggle_repeat) begin : CLKGEN
      clk_out_phase = phase_number * effective_ref_period / (2 * ratio_samp) - sum_until_now;
      sum_until_now = sum_until_now + clk_out_phase;
      if (~enable)
         return;
      #(clk_out_phase) clk_out = ~clk_out;
      phase_number = phase_number + 1;
   end : CLKGEN

endtask

endmodule
`endif


`ifndef ip2211ringpll_VIEWMUXANA_SV
`define ip2211ringpll_VIEWMUXANA_SV

module ip2211ringpll_viewmuxana (
    `ifndef ip2211ringpll_INTC_NO_PWR_PINS
        input wire     vccvdd2,
        input wire     vccpll,
    `endif
    input  logic [1:0] viewanaen,
    input  logic       adc_in,	// from adc_in mux
    input  logic       anadft_ldo,
    output logic [1:0] viewanabus
    );//Module begin

    // Analog view mux drive the outputs tristate when not enabled
    // When viewanaen[1] = 1, ViewPinNH[1] = iref_view; When viewanaen[1] = 0,  ViewPinNH[1] = ldo output
    `ifndef ip2211ringpll_LJPLL_MSV
    `ifndef INTC_NO_VCSSIM_OR_EMU
        logic [1:0] ViewPinNH;
        always_comb begin : VIEW
            ViewPinNH[0] = viewanaen[0] ? adc_in : 1'bz;
            ViewPinNH[1] = viewanaen[1] ? 1'b1 : anadft_ldo;
        end : VIEW
        assign viewanabus = ViewPinNH;
    `endif
    `endif
endmodule //Module end
`endif

`ifndef ip2211ringpll_pllljtopana_SV
`define ip2211ringpll_pllljtopana_SV

//`ifndef VCSSIM_OR_EMU
//   `ifdef INTC_EMULATION
//      `define VCSSIM_OR_EMU
//   `endif
//`endif
//
//`ifndef VCSSIM_OR_EMU
//   `ifdef VCSSIM
//      `define VCSSIM_OR_EMU
//   `endif
//`endif

`ifndef INTC_NO_VCSSIM_OR_EMU
   //`include "soc_macros.sv"
   //`include "ringpll_macros.sv"
`endif
//`ifndef ip2211ringpll_SVA_OFF
   //`include "intel_checkers.vs"
//`endif

`ifndef ip2211ringpll_NO_VCSSIM
   //`include "PLL_AIP.sv"
   //`include "clkgen.sv"
`endif

//`include "viewmuxana.sv"
// added and commented few pins at the interface of pll_core by taking netlist and lib as referance
module ip2211ringpll_pllljtopana
//`ifndef ip2211ringpll_LJPLL_MSV
//`ifndef ip2211ringpll_NO_VCSSIM
//#(parameter bit INTC_USE_DETAILED_AIP_MODEL = 0,
//  parameter     RATIO_BITS = 10)
//`endif
//`endif
(
   `ifndef ip2211ringpll_LJPLL_MSV
   `ifndef INTC_NO_VCSSIM_OR_EMU
      // The PLL clock generator needs to be aware of the ratio in
      // instrumentation mode. In analog, all of this is done through phase
      // detection and frequency multiplication
      //
      //input logic [7:0] ratio,
      input logic [9:0] ratio,
      input logic       half_int,

      // Whenever the ip2211ringpll_pll_inst_align halts the clock, we should reset the lock
      // detector
      //
      input logic                      pllfbgen__haltclk_inst,
  
   `endif
   `ifndef ip2211ringpll_SVA_OFF
      // Feedback clock should be driven when EarlyLock asserts
      input logic                      EarlyLockXXH,
      
      // Lock is used to reset feedback clock alignment SVAs
      input logic                      LockXXL,
      
   `endif
   `endif
  
   `ifndef ip2211ringpll_INTC_NO_PWR_PINS
      input wire                       vccpll,
      input wire                       vccref,
      input wire                       vccvdd2,
   `endif

   // RDAC interface
   //
   input  logic [3:0]                vctlrdac,
   
   // PLL Startup Controls
   //
   input  logic                      vctlrdacen,
   input  logic                      rdactovctlen,
   input  logic                      pfden,
 // input  logic                      cmpen,
 // input  logic                      vctl_pullup,
 // input  logic                      vctl_pulldn,
   

   // Charge Pump Controls
   //
//   input  logic                      lpcpen,
//   input  logic                      cpdisfbampsamp,
//   input  logic                      cpenfbamp,
//   input  logic                      cpselfbamp,
//   input  logic                      cpirefaltmode,
//   input  logic                      pfd_chop_en, 
//   input  logic [2:0]                pfd_chop_val, 
   input  logic [2:0]                pfd_residual_pw,
   input  logic [4:0]                cp1_trim,
   input  logic [4:0]                cp2_trim,
   input  logic [4:0]                skadj_ctrl,
`ifdef INTC_NO_VCSSIM_OR_EMU
   input logic [10:0]  fz_vcotrim,
   input logic [1:0] fz_cpnbias,
   input logic [1:0] fz_pfddly,
   input logic [4:0] fz_irefgen,
   input logic [5:0] fz_startup,
   input logic fz_nopfdpwrgate,
`endif
   // IREF
   //
`ifndef INTC_NO_VCSSIM_OR_EMU
   input  logic                      clk_iref,
`endif
   input  logic                      irefvcoclksel,
//   input  logic                      irefbypassamp_mode, // IREF amplifier disable
//   input  logic                      irefrmodeen,
//   input  logic                      en_vcodiv16toiref,
//   input  logic                      en_vcodiv32toiref,
//   input  logic                      irefhighcurr_en,
   
//   input  logic [2:0]                iref_ctune,
//   input  logic [3:0]                iref_ftune,
   

   // LPF
   //
//   input  logic                      lpf_pg_en,
//   input  logic [1:0]                lpf_itrim,


//   input  logic [1:0]                pvd_mode, 
   input  logic [1:0]                pdivrat, 
   input  logic [3:0]                lockthresh,
  `ifndef INTC_NO_VCSSIM_OR_EMU
   input  logic [3:0]                vco_trim_pg,
   input  logic [2:0]                vco_trim_cb,
   input  logic [3:0]                viewsel0 ,
   input  logic [3:0]                viewsel1 ,
  `endif  
   input  logic [1:0]                viewanaen,


   input  logic                      clkref,
   input  logic                      clkfb,
   input  logic                      reset_b,
         
   output wire                       adc_in,
   input  wire  [2:0]                adc_sel_in,	 
  
   // LDO outputs 
   input  logic			     anadft_ldovfb,
   input  logic			     anadft_ldovref,
   input  logic			     anadft_ldo,
   
   // PLL core DFX outputs
   `ifdef INTC_NO_VCSSIM_OR_EMU
    output logic                      cp1clk,
    output logic                      cp1aclk,
    output logic                      cp2clk,
    output logic                      cp2aclk,
   `endif
   output tri   [1:0]                viewanabus,
   output logic                      pfdlockrst,
  // output logic                      compout,
   output logic                      clkpll
);

   logic                      cp1clk;
   logic                      cp1aclk;
   logic                      cp2clk;
   logic                      cp2aclk;


//parameter bit INTC_USE_DETAILED_AIP_MODEL = 0;

`ifndef INTC_NO_VCSSIM_OR_EMU

`ifndef ip2211ringpll_LJPLL_MSV
   logic ResetBXXnnnH;
   logic ClkFbDelayMXH;
   logic [1:0] FbEdgeVecNnnnH;
   logic FbEdgeNnnnH;
   logic FbTickXXnnnH;
   logic FbIsTickingXXnnnH;
   //logic [7:0] ratio_samp;
   logic [9:0] ratio_samp;
   logic half_int_samp;
   //logic [8:0] vco_ratio;
   logic [9:0] vco_ratio;
   logic [9:0] vco_divider;
// These clocks are not used in ip22 ringpll anymore.
assign cp1clk = 1'b0;
assign cp1aclk = 1'b0;
assign cp2clk = 1'b0;
assign cp2aclk = 1'b0;

//   logic CmpReset;
  // logic CmpChangeGo;
//   logic StartupCmpInitNH;
//  `ifndef ip2211ringpll_NO_VCSSIM
//     always @(posedge reset_b) begin
//        StartupCmpInitNH <= $dist_uniform($get_initial_random_seed, 0, 1);
//     end
//  `else
//     assign StartupCmpInitNH = 1'b0;
//  `endif

//   always_comb CmpReset = ~reset_b /*| ~cmpen*/;
//   always_comb CmpChangeGo = StartupCmpInitNH ? vctl_pullup
//                                              : vctl_pulldn  ;

  // logic [2:0] StartupDoneNnnnH;

 //  always_comb StartupDoneNnnnH[0] = 1'b1;
//   `ip2211ringpll_EN_ASYNC_RST_MSFF(StartupDoneNnnnH[2:1], StartupDoneNnnnH[1:0], clkref, CmpChangeGo, CmpReset)

   // Initial conditions
   //    compout = 1 means startup should pull down
   //    compout = 0 means startup should pull up
   //
//   always_comb begin 
  //    compout = StartupCmpInitNH ? ~StartupDoneNnnnH[2]
 //                                :  StartupDoneNnnnH[2]  ;
   //   compout = compout & cmpen;
//   end

   `ip2211ringpll_ASYNC_RST_MSFF(ResetBXXnnnH, 1'b1, clkref, ~reset_b)
  
   `ip2211ringpll_LATCH_P(ratio_samp, ratio, reset_b)
   `ip2211ringpll_LATCH_P(half_int_samp, half_int, reset_b)

   assign vco_ratio = half_int_samp ? {ratio_samp,1'b1} : {1'b0,ratio_samp};


   `ifndef ip2211ringpll_NO_VCSSIM
      //if (INTC_USE_DETAILED_AIP_MODEL) begin : AIP_DETAILED_MODEL
     `ifdef INTC_USE_DETAILED_AIP_MODEL  //AIP_DETAILED_MODEL
      ip2211ringpll_PLL_AIP #(
                     // ip2211ringpll_PFD Parameters
                     .PFD_SIGN       ( -1 ),  // if ip2211ringpll_VCO frequency is inversely proportional to Vctrl, put PFD_SIGN = -1, otherwise put it 1

                     // Charge Pump Parameters
                     .I_INTEGRAL     ( 0.000002 ),        // Amp
                     .I_PROPORTIONAL ( 0.0000357 ),    // Amp
                     
                     // SC Loop Filter Parameters
                     .C1_VALUE       ( 0.000000000001 ),    // Farad
                     .C2_VALUE       ( 0.000000000090 ),    // Farad

                     .VCTRL_INITIAL  ( 0.5 ),          // Volt
                     .VINT_INITIAL   ( 0.5 ),          // Volt
                     .VPROP_INITIAL  ( 0 ),            // Volt

                     // ip2211ringpll_VCO Parameters:
                     .F0_VALUE       ( 7966 ),         // MHz
                     .KVCO_VALUE     ( -12936.666 )
               )                  vco (.CLK_REF     ( clkref   ),
                                       .CLK_FED     ( clkfb    ),
                                       .pvdmode     ( pdivrat  ),
                                       .VCO_RESET   ( reset_b  ),
                                       .RESET       ( pfden    ),
                                       .CLK_VCO     ( clkpll   ));
      //`end : AIP_DETAILED_MODEL
      `else  //AIP_DETAILED_MODEL
      //else begin : SIMPLE_MODEL
      // Clock Generator for RTL Simulation
      //
      ip2211ringpll_clkgen 
		//#(.RATIO_BITS(RATIO_BITS))    
				vco (.clk_ref(clkref),
                                       .enable(ResetBXXnnnH),
                                       .ratio(vco_ratio),
                                       .half_int(half_int_samp),
                                       .clk_out(clkpll));
      //end : SIMPLE_MODEL
      `endif //AIP_DETAILED_MODEL
      
      //if (INTC_USE_DETAILED_AIP_MODEL) begin : PHASE_ERROR_MODEL
      `ifdef INTC_USE_DETAILED_AIP_MODEL  //PHASE_ERROR_MODEL
         time clkref_period;
         time clkref_start;
         time clkfb_start;
         time ph_error;
         time true_ph_error;
         time lock_threshold_time;

         always_comb begin : LOCKTHRESH
            unique casez (lockthresh)
               4'b0000 : lock_threshold_time = 29ps;
               4'b0001 : lock_threshold_time = 68ps;
               4'b0010 : lock_threshold_time = 94ps;
               4'b0011 : lock_threshold_time = 132ps;
               4'b0100 : lock_threshold_time = 158ps;
               4'b0101 : lock_threshold_time = 196ps;
               4'b0110 : lock_threshold_time = 224ps;
               4'b0111 : lock_threshold_time = 263ps;
               4'b1000 : lock_threshold_time = 484ps;
               4'b1001 : lock_threshold_time = 522ps;
               4'b1010 : lock_threshold_time = 743ps;
               4'b1011 : lock_threshold_time = 782ps;
               4'b1100 : lock_threshold_time = 1002ps;
               4'b1101 : lock_threshold_time = 1041ps;
               4'b1110 : lock_threshold_time = 1262ps;
               4'b1111 : lock_threshold_time = 1300ps;
               default : lock_threshold_time = 1ps;
            endcase
         end : LOCKTHRESH
         
         always @(posedge clkref) begin
            clkref_period <= ($realtime() - clkref_start);
            clkref_start <= $realtime();
         end

         always @(posedge clkfb)
            clkfb_start <= $realtime();

         always_ff @(posedge clkref)
            ph_error <= ABS(clkref_start - clkfb_start);

         assign true_ph_error = MIN(ph_error, ABS(ph_error-clkref_period));

         assign pfdlockrst = (true_ph_error > lock_threshold_time);
	
	 // =============================================================== //
   	 // adc_in:  							    //
   	 // 0 - vss							    //
   	 // 1 - cp bias						     	    //
  	 // 2 - vctl							    //
   	 // 3 - vro							    //
   	 // 4 - vccpll						      	    //
    	 // 5 - vss							    //
   	 // 6 - ldo vfb						            //
   	 // 7 - ldo vref					 	    //
   	 // viewanabus[0] = adc_in					    //
   	 // viewanabus[1] = iref_view (= vccpll on voltmeter)		    //
   	 // viewanabus[1] is shared with LDO and debug		     	    //
   	 // =============================================================== //
   	 logic to_adc;

   	 always_comb begin
	   	case (adc_sel_in)
		   3'd0 : to_adc = 1'b0;
		   3'd1 : to_adc = realZ;
		   3'd2 : to_adc = vco.SC_LPF_i1.Vctrl;
		   3'd3 : to_adc = realZ;
		   3'd4 : to_adc = vccpll;
		   3'd5 : to_adc = 1'b0;
		   3'd6 : to_adc = anadft_ldovfb;
		   3'd7 : to_adc = anadft_ldovref;
		   default : to_adc = 1'b0;
	   	endcase
   	 end

   	 assign adc_in = to_adc;

      //end : PHASE_ERROR_MODEL
      //else begin : SIMPLE_FBTICK_MODEL
	`else //SIMPLE_FBTICK_MODEL
      `ip2211ringpll_NB_ASSIGN(ClkFbDelayMXH, clkfb)


      always_comb begin : FB_EDGE_DETECT
         FbEdgeVecNnnnH = {ClkFbDelayMXH, clkfb};
         FbEdgeNnnnH    = (FbEdgeVecNnnnH == 2'b01) || (FbEdgeVecNnnnH == 2'b10);
      end : FB_EDGE_DETECT

      `ip2211ringpll_ASYNC_SET_MSFF(FbTickXXnnnH, 1'b0, clkref, FbEdgeNnnnH)
      `ip2211ringpll_ASYNC_RST_MSFF(FbIsTickingXXnnnH, FbTickXXnnnH, clkref, ~reset_b)
   
      assign pfdlockrst   = ~FbIsTickingXXnnnH | pllfbgen__haltclk_inst ;
      logic to_adc;

   	 always_comb begin
	   	case (adc_sel_in)
		   3'd0 : to_adc = 1'b0;
		   3'd1 : to_adc = 1'bz;
		   3'd2 : to_adc = 1'bz;
		   3'd3 : to_adc = 1'bz;
		   3'd4 : to_adc = anadft_ldo;
		   3'd5 : to_adc = 1'b0;
		   3'd6 : to_adc = anadft_ldovfb;
		   3'd7 : to_adc = anadft_ldovref;
		   default : to_adc = 1'b0;
	   	endcase
   	 end

   	 assign adc_in = to_adc;
               
      //end : SIMPLE_FBTICK_MODEL
	`endif //SIMPLE_FBTICK_MODEL

   `else //ip2211ringpll_NO_VCSSIM
     `ifdef INTEL_EMULATION 

	bit [15:0] vco_ratio_zero_ext, vco_divide_zero_ext;

	
	 assign vco_divider = half_int_samp ? 2 : 1;
      assign vco_ratio_zero_ext  = {{$bits(vco_ratio_zero_ext)-$bits(vco_ratio){1'b0}}, vco_ratio};
      assign vco_divide_zero_ext = {{$bits(vco_ratio_zero_ext)-$bits(vco_ratio){1'b0}}, vco_divider};

      // VCO clock generator delayed reset
      //    EMU clock generator samples reference clock frequency only when
      //    reset is asserted. Delaying reset de-assertion provides more
      //    time for the PLL's reference clock frequency to stabilize in emulation.
      //
      bit vco_delayed_reset;
      bit [7:0] vco_reset_timer;
      bit [7:0] vco_reset_timer_init;

      assign vco_reset_timer_init = 8'd30;

      always @(posedge clkref) begin
        if(~ResetBXXnnnH) begin
            vco_reset_timer = vco_reset_timer_init;

        end
        else begin
            if(vco_reset_timer) begin
                vco_reset_timer = vco_reset_timer - 1;
            end
        end
      end
      assign vco_delayed_reset = ~ResetBXXnnnH || (vco_reset_timer!=0);

		emu_clk_pll emu_ringpll_vco (
               .enable             (!vco_delayed_reset),               // active high enable for the clk_out
               .numerator          (vco_ratio_zero_ext),          // numerator, can be changed on the fly
               .denominator        (vco_divide_zero_ext),         // denominator, can be changed on the fly
               .lock_delay         (0),                           // num of ref clks from enable to lock ?? can this be calculated
               .ref_clk            (clkref),                      // optional used if edge alignment is need
               .outclk_alignment   (0),                           // align out clock to refclk  (0 = pos edge , 1 neg )
               .lock_alignment     (0),                           // align lock enable to refclk (0)pos/(1)neg egdge
               .lock               (),                           
               .clk_out            (clkpll)                       // output clock
          );

      `ip2211ringpll_NB_ASSIGN(ClkFbDelayMXH, clkfb)


      always_comb begin : FB_EDGE_DETECT
         FbEdgeVecNnnnH = {ClkFbDelayMXH, clkfb};
         FbEdgeNnnnH    = (FbEdgeVecNnnnH == 2'b01) || (FbEdgeVecNnnnH == 2'b10);
      end : FB_EDGE_DETECT

      `ip2211ringpll_ASYNC_SET_MSFF(FbTickXXnnnH, 1'b0, clkref, FbEdgeNnnnH)
      `ip2211ringpll_ASYNC_RST_MSFF(FbIsTickingXXnnnH, FbTickXXnnnH, clkref, ~reset_b)
   
      assign pfdlockrst   = ~FbIsTickingXXnnnH | pllfbgen__haltclk_inst ;
     `else 

      assign pfdlockrst   = pllfbgen__haltclk_inst ;
      assign adc_in = 'z;
      `endif
   `endif

 
`endif
`endif
    
   // Analog view mux
   ip2211ringpll_viewmuxana viewana(
    `ifndef ip2211ringpll_INTC_NO_PWR_PINS
           .vccvdd2 (vccvdd2),
           .vccpll  (vccpll),
    `endif
		.*);
`ifndef ip2211ringpll_SVA_OFF

///========================================================================================================
/// Assertions
///========================================================================================================

//   `ip2211ringpll_ASSERTS_KNOWN_DRIVEN(R_pllljtopana_X_inputs,
//   {vctlrdac, vctlrdacen, rdactovctlen, pfden,
//   /*cmpen, vctl_pullup, vctl_pulldn,*/ lpcpen, cpdisfbampsamp,
//   cpenfbamp, cpselfbamp, cpirefaltmode, pfd_chop_en,
//   pfd_chop_val, pfd_residual_pw, cp1_trim, cp2_trim,
//   clk_iref, irefvcoclksel, irefbypassamp_mode, irefrmodeen,
//   en_vcodiv16toiref, en_vcodiv32toiref, irefhighcurr_en,
//   iref_ctune, iref_ftune, lpf_pg_en, lpf_itrim, pdivrat,
//   lockthresh, vco_trim_pg, vco_trim_cb, viewsel0, viewsel1,
//   viewanaen, clkref, reset_b, adc_sel_in},
//   clkref, ~(reset_b===1'b1),
//   `ip2211ringpll_ERR_MSG("[LJPLL] X inputs to ip2211ringpll_pllljtopana after powerup"));
   

   `ip2211ringpll_ASSERTS_KNOWN_DRIVEN(R_pllljtopana_X_inputs,
   {vctlrdac, vctlrdacen, rdactovctlen, pfden,
   pfd_residual_pw, cp1_trim, cp2_trim,
   clk_iref, irefvcoclksel, 
   lockthresh, vco_trim_pg, vco_trim_cb, viewsel0, viewsel1,
   viewanaen, clkref, reset_b, adc_sel_in},
   clkref, ~(reset_b===1'b1),
   `ip2211ringpll_ERR_MSG("[LJPLL] X inputs to ip2211ringpll_pllljtopana after powerup"));


   `ip2211ringpll_ASSERTS_KNOWN_DRIVEN(R_pllljtopana_X_clkfb, clkfb,
            clkref, (~(reset_b===1'b1) | (pfden===1'b0)),
   `ip2211ringpll_ERR_MSG("[LJPLL] X inputs to ip2211ringpll_pllljtopana after powerup"));

`ifndef ip2211ringpll_LJPLL_MSV
   `ip2211ringpll_ASSERTC_SAME(R_pllljtopana_fb_align, (clkref && !$sampled(clkref) && !$sampled(clkfb)), (clkfb  && !$sampled(clkfb)  && !$sampled(clkref)), (~(reset_b===1'b1) | ~(LockXXL===1'b1)),   `ip2211ringpll_ERR_MSG("[LJPLL] Reference clock and feedback clock are not aligned after lock"));
`endif

`endif


endmodule

`ifndef ip2211ringpll_NO_VCSSIM
function int ABS (int num);
   ABS = (num <0) ? -num : num;
endfunction // ABS 

function int MIN (int num1, num2);
   MIN = (num1 < num2) ? num1 : num2;
endfunction // ABS
`endif

`endif

`ifndef ip2211ringpll_PLL_AIP_SV
`define ip2211ringpll_PLL_AIP_SV

///============================================================================================================================================================================================
/// Included Files
///============================================================================================================================================================================================

//`include "PFD.sv"
//`include "SC_LPF.sv"
//`include "VCO.sv"
//`include "SecondOrderLoopFilter.sv"

module ip2211ringpll_PLL_AIP
#(
   // ip2211ringpll_PFD Parameters
   parameter real PFD_SIGN = -1,  // if ip2211ringpll_VCO frequency is inversely proportional to Vctrl, put PFD_SIGN = -1, otherwise put it 1

   // Charge Pump Parameters
   parameter real I_INTEGRAL = 0.000002,        // Amp
   parameter real I_PROPORTIONAL = 0.0000357,    // Amp

   // SC Loop Filter Parameters
   parameter real C1_VALUE = 0.000000000001,    // Farad
   parameter real C2_VALUE = 0.000000000090,    // Farad

   parameter real VCTRL_INITIAL = 0.5,          // Volt
   parameter real VINT_INITIAL  = 0.5,          // Volt
   parameter real VPROP_INITIAL = 0,            // Volt

   // ip2211ringpll_VCO Parameters:
   parameter real F0_VALUE = 7966,         // MHz
   parameter real KVCO_VALUE = -12936.666, //MHz
   parameter real TIME_INCREASE = 0.000000000001 // increase time by 1ps
)

(CLK_VCO, CLK_REF, CLK_FED, RESET, VCO_RESET, pvdmode);

// INPUTS AND OUTPUTS
output logic CLK_VCO;
input  logic CLK_REF, RESET, VCO_RESET;
input  logic CLK_FED;
input  logic [1:0] pvdmode;

// INTERNAL SIGNALS
logic PhaseErrorSign, PhaseErrorMag;
real Vctrl;


///============================================================================================================================================================================================
/// Phase Frequency Detector
///============================================================================================================================================================================================

ip2211ringpll_PFD PFD_i1 (PhaseErrorSign, PhaseErrorMag, CLK_REF, CLK_FED, RESET, 1'b1);


///============================================================================================================================================================================================
/// Switched Capacitor Loop Filter
///============================================================================================================================================================================================

ip2211ringpll_SC_LPF #(
         .PFD_SIGN(PFD_SIGN),
         .I_INTEGRAL(I_INTEGRAL),
         .I_PROPORTIONAL(I_PROPORTIONAL),
         .C1_VALUE(C1_VALUE),
         .C2_VALUE(C2_VALUE),

         .VCTRL_INITIAL(VCTRL_INITIAL),
         .VINT_INITIAL(VINT_INITIAL),
         .VPROP_INITIAL(VPROP_INITIAL),
         .TIME_INCREASE(TIME_INCREASE)

)

SC_LPF_i1 (Vctrl, PhaseErrorMag, PhaseErrorSign, RESET);

///============================================================================================================================================================================================
/// Voltage Controlled Oscillator
///============================================================================================================================================================================================

ip2211ringpll_VCO  #(
         .F0_VALUE(F0_VALUE),
         .KVCO_VALUE(KVCO_VALUE)
)

VCO_i1  (CLK_VCO, Vctrl, pvdmode, VCO_RESET);


endmodule

`endif

`ifndef ip2211ringpll_PFD_SV
`define ip2211ringpll_PFD_SV


module ip2211ringpll_PFD (PhaseErrorSign, PhaseErrorMag, CLK_REF, CLK_FED, RESET, dco_reset);

    // INPUTS AND OUTPUTS
    output bit PhaseErrorSign, PhaseErrorMag;
    input CLK_REF, CLK_FED, dco_reset;
    input bit RESET;

    // INTERNAL SIGNALS
    bit  n1, n2, n3, n4, n5, n6, n7, n8, n9, UP;
    bit n11, DN, n13, n14, n16, n17, n18;
    bit PhaseErrorSign_neg;

    bit PhaseErrorMagGlitchy, PhaseErrorMagGlitchy_delayed;


///============================================================================================================================================================================================
/// ip2211ringpll_PFD Circuit Discription
///============================================================================================================================================================================================

    nand  #20   g1(n1, n7, !CLK_REF),
                   g2(n2, n1, n3),
                   g3(n3, n2, n13),
                   g4(n4, n13, n5),
                   g5(n5, n4, n6),
                   g6(n6, !CLK_FED, n9);

    nand  #40   u1(n7, n1, n2, n13),
                   u3(n9, n13, n5, n6);

    nand  #60   u2(n8, n2, n1, n6, n5);

    nand  #40   k1(n11, n8, RESET, dco_reset);

    ip2211ringpll_my_buffer  buff (n14, n11);

    not #10     i1(UP, n7),
                   i2(n13, n14),
                   i3(DN, n9);


    ip2211ringpll_dff_pos_nr ff (PhaseErrorSign_neg, DN, UP, RESET);


    not         i7 (PhaseErrorSign,PhaseErrorSign_neg);

    xor         z9 (PhaseErrorMagGlitchy, UP, DN);    //EVENT is an output representing the magnitude of the phase error

    // Remove Glitches if any from PhaseErrorMag
    assign #2fs PhaseErrorMagGlitchy_delayed = PhaseErrorMagGlitchy;
    assign PhaseErrorMag = PhaseErrorMagGlitchy_delayed & PhaseErrorMagGlitchy;


///============================================================================================================================================================================================
/// Measure Phase Error
///============================================================================================================================================================================================

real PhaseErrorMag_REAL_pre, PhaseErrorMag_REAL, PhaseErrorMag_RISE, PhaseErrorMag_FALL;
real sign;

always @(PhaseErrorSign) sign = (PhaseErrorSign == 1'b1)? 1 : -1;

always_ff @(posedge PhaseErrorMag) begin if (PhaseErrorMag == 1'b1) PhaseErrorMag_RISE = $realtime; end
always_ff @(negedge PhaseErrorMag) begin if (PhaseErrorMag == 1'b0) PhaseErrorMag_FALL = $realtime; end

always @(PhaseErrorMag_FALL) if (PhaseErrorMag_FALL > PhaseErrorMag_RISE) PhaseErrorMag_REAL_pre = PhaseErrorMag_FALL - PhaseErrorMag_RISE;

// PhaseErrorMag_REAL represents phase error between CLKREF and CLKFED in ps
always @(PhaseErrorMag_FALL) if (PhaseErrorMag_FALL > PhaseErrorMag_RISE) PhaseErrorMag_REAL = PhaseErrorMag_REAL_pre * sign;


///============================================================================================================================================================================================
/// Indicate Lock Based on Phase Error
///============================================================================================================================================================================================

// Assign raw_lock 1 if phase error is less than 100 ps, even for 1 ref cycle.
bit raw_lock, lock;
assign raw_lock = (~RESET)? 1'b0 : (PhaseErrorMag_REAL_pre < 100)? 1'b1 : 1'b0;  // PhaseErrorMag_REAL_pre is the absolute value

// use the raw_lock as a counter enable. the counter counts for # cycles to make sure phase error is stable and PLL is locked
bit [4:0] lock_count;
always @(negedge RESET or posedge CLK_REF) begin lock_count <= (~RESET)? 5'd0 : (lock_count == 5'd30)? 5'd30 : (raw_lock == 1'b1)? (lock_count + 1) : 5'd0; end

// Sticky Lock
assign lock = (~RESET)? 1'b0 : (lock_count == 5'd30)? 1'b1 : 1'b0;

// Check that phase error shouldn't be higher than bounded value when lock is asserted, NOTE: PhaseErrorMag_Real_pre is the absolute value for phase error
always @(PhaseErrorMag_REAL) begin
if (  (lock == 1'b1) && (PhaseErrorMag_REAL_pre > 2000)  ) $display ("[INFO]: Phase Error is higher than 2ns while PLL is locked");
end


endmodule



///============================================================================================================================================================================================
/// Buffer to delay RESET signal
///============================================================================================================================================================================================

   module ip2211ringpll_my_buffer (out, in);

    output bit out;
    input bit in;
    bit w1, w2, w3, w4, w5, w6, w7, w8, w9;

    assign #10 w1 = !in;
    assign #10 w2 = !w1;
    assign #10 w3 = !w2;
    assign #10 w4 = !w3;
    assign #10 w5 = !w4;
    assign #10 w6 = !w5;
    assign #10 w7 = !w6;
    assign #10 w8 = !w7;
    assign #10 w9 = !w8;
    assign #10 out = !w9;


   endmodule


///============================================================================================================================================================================================
/// Flip Flop to determine ip2211ringpll_PFD Output Sign
///============================================================================================================================================================================================

   module ip2211ringpll_dff_pos_nr (q, din, clk, reset);
      output q;
      input din,clk, reset;
      reg q;
      always @ (posedge clk or negedge reset)
         begin
            if (~reset) q <= 1'b0;
            else q <= din;

         end
   endmodule

`endif

`ifndef ip2211ringpll_SC_LPF_SV
`define ip2211ringpll_SC_LPF_SV

///============================================================================================================================================================================================
/// Module Inputs/Outputs
///============================================================================================================================================================================================


module ip2211ringpll_SC_LPF
#(
  parameter real PFD_SIGN = 1,                 // if ip2211ringpll_VCO frequency is inversely proportional to Vctrl, put PFD_SIGN = -1, otherwise put it 1

  parameter real I_INTEGRAL = 0.000002,        // Amp
  parameter real I_PROPORTIONAL = 0.0000357,    // Amp
  parameter real C1_VALUE = 0.000000000001,    // Farad
  parameter real C2_VALUE = 0.000000000090,    // Farad

  parameter real VCTRL_INITIAL = 0.5,          // Volt
  parameter real VINT_INITIAL  = 0.5,          // Volt
  parameter real VPROP_INITIAL = 0,            // Volt
  parameter real TIME_INCREASE =0.000000000001 // Increase time by 1ps
)

(Vctrl, PhaseErrorMag, PhaseErrorSign, RESET);

`ifdef INTEL_EMULATION
 output logic Vctrl; // Units in Volt
`else
 output real Vctrl; // Units in Volt
`endif
 input logic PhaseErrorMag, PhaseErrorSign;
 input bit RESET;

 real Vctrl_initial; // Initial value for ip2211ringpll_VCO control voltage, this determines ip2211ringpll_VCO initial frequency when PLL starts its operation
 real time_t, time_t_stored;  // real number representing time (factored in loop filter equations)

 real Vint, Vprop;  // Vint --> integral voltage generated due to integral CP current. Vprop --> proportional voltage generated due to proportioanl CP current. Vctrl = Vint + Vprop
 real Vint_initial, Vprop_initial;  // iniital values for integer and proportional voltages.

 real Ii, Ip;  // Units in Amp, integral and proportional charge pump currents
 real C1, C2;  // Units in Farad, Capacitors of Loop Filter. C1 is the cap that effectively integrates the charges to generate Vctrl for ip2211ringpll_VCO.

 real sign, sign_stored;  // phase error sign

 logic very_first_cycle;
 logic ClkSample; // Very high frequency clock to smoothly incerase time_t to emulate time. this clock toggles only in the presense of phase error for performance optimization
 bit initial_trig; // used to make sure the "always" block that includes design parameters, get accessed one time. (represents initial block).

 real ClkSample_delay_pre, ClkSample_delay;


///============================================================================================================================================================================================
/// Converting phase error logic sign into real sign
///============================================================================================================================================================================================

 always @(PhaseErrorSign) begin
   if (PhaseErrorSign == 1'b1) sign = PFD_SIGN; else sign = -PFD_SIGN;
 end

///============================================================================================================================================================================================
/// Vctrl Generation through Switched Capacitor Loop Filter
///============================================================================================================================================================================================


 always @(negedge ClkSample or posedge ClkSample or PhaseErrorMag or RESET) begin
 if (~RESET) begin Vint = 0.02; Vprop = 0.02; end  // when PFD_EN is 0, cap should discharge, Vctrl should go to ~0
 else begin

   if (PhaseErrorMag == 1'b0)  // if phase error is zero, resets everything, time should be 0, loop filter is assumed to hold its final Vctrl
    //----------------------------------------------------------------------------------------------------------------------------------------
    begin

     Vint_initial = Vint;
     Vprop_initial = Vprop;

     if (ClkSample == 1'b0) begin  // this check because it might be accessed twice if ClkSample = 1 when PhaseErrorMag = 0, as after 1ps ClkSample will be 0 and will access it again making time_t_store = 0
       time_t_stored = time_t;
       sign_stored = sign;
       time_t = 0;
     end

    end



    else // if phase error is 1, time should increase gradually to update the loop filter equations
    //----------------------------------------------------------------------------------------------------------------------------------------
    begin

      // once phase error is 1 (only instantinuous action), reset Vprop, because the charges accumulated over C2 should be gone during reset phase, Vctrl should have ~Vint value only
      if ( (time_t == 0) && (very_first_cycle == 0) ) begin Vprop = 0; Vprop_initial = 0;

         Vint = Vint  -  ( Ii/(C1+C2) ) * time_t_stored * sign_stored  +  ( Ii/(C1+ 2*C2) ) * time_t_stored * sign_stored;
         ////   ----     ---------------------------------------------    ------------------------------------------------
         Vint_initial = Vint; time_t = time_t + TIME_INCREASE;
      end

      // After Vprop gets reset, Vint and Vprop will increase gradually becuase of the integration of the CP currents over the caps, forming Vctrl
      else begin

        Vint = Vint_initial + ( Ii/(C1+C2) ) * time_t * sign;
        Vprop = Vprop_initial + ( Ip/(C1+C2) ) * time_t * sign;
        time_t = time_t + TIME_INCREASE;
        very_first_cycle = 0;

      end


    end
    //---------------------------------------------------------------------------------------------------------------------------------------

  // be careful, at begining of simulation, this statement will be valid, and Vctrl will be calculated
  // becuase at time 0, simulater considers ClkSample as negedge or posedge depending on initial value
  // in the testbench put the following, #0 Vctrl2 = 0.5; #1 Vctrl2 = 0.5 --> to guarantee right value
end  // end if (~RESET)
end  // end always

///============================================================================================================================================================================================
/// Vctrl is Vint + Vprop
///============================================================================================================================================================================================

 always @( Vint or Vprop) begin Vctrl = Vint + Vprop; end


///============================================================================================================================================================================================
/// Create ClkSample to increase/decrease Vctrl linearly and smoothly
///============================================================================================================================================================================================


  assign #(ClkSample_delay) ClkSample = (PhaseErrorMag == 1'b0)? 1'b0 : !ClkSample;  // PhaseError MUST be zero at #0 in order not to have unknown values for ClkSample(add reset signal to reset ip2211ringpll_PFD out at #0)



///============================================================================================================================================================================================
/// Always block equivalent to initial block. All ip2211ringpll_VCO related parameters are defined here
///============================================================================================================================================================================================


 always @(PhaseErrorMag)  begin  // at 0 time, reset is zero, so PhaseErrorMag in (ip2211ringpll_PFD.sv) is zero, so this always block is triggered

  // Equivalent to Initial Block for MPP Simulations that do not accept initial block

  if (initial_trig == 1'b0) begin


      time_t = 0;
      time_t_stored = 0;
      very_first_cycle = 1;

   // CP and Loop Filter Parameters
   //-------------------------------------------
      Ii = I_INTEGRAL;            // uA
      Ip = I_PROPORTIONAL;            // uA

      C1 = C1_VALUE;      // pF
      C2 = C2_VALUE;      // pf


   // Initial Voltages Values
   //-------------------------------------------
   Vctrl = VCTRL_INITIAL;
   Vint_initial = VINT_INITIAL;
   Vint = VINT_INITIAL;

   Vprop_initial = VPROP_INITIAL;
   Vprop = VPROP_INITIAL;

   ClkSample_delay_pre = TIME_INCREASE;
   ClkSample_delay =  ClkSample_delay_pre * 1000000 * 1000000;   // Convert TIME_INCREASE from seconds to ps, then this value is used to determine the pulse width of the ClkSample in ps

   initial_trig = 1'b1;  // to access this always block only one time in the beginning (as an initial block).

  end
end
 ////////////////////////////////////////////////////////////////////////////////////

endmodule

`endif

`ifndef ip2211ringpll_VCO_SV
`define ip2211ringpll_VCO_SV

///============================================================================================================================================================================================
/// Module Inputs/Outputs
///============================================================================================================================================================================================

module ip2211ringpll_VCO
#(
   parameter real F0_VALUE = 7966,         // MHz
   parameter real KVCO_VALUE = -12936.666  // MHz/Volt
)

(CLKPVD, Vctrl, pvdmode, VCO_RESET);

  input logic [1:0] pvdmode;
  input bit VCO_RESET;
`ifdef INTEL_EMULATION
  input logic Vctrl;        // Units in Volt
`else
  input real Vctrl;        // Units in Volt
`endif
  output logic CLKPVD;     // Output logic clock

  real F0;                 // Initial ip2211ringpll_VCO frequency if Vctrl = 0, Units in MHz
  real Kvco;               // Gain of ip2211ringpll_VCO, Units in MHz/Volt
  real Td, Td_pre;         // Delay of each inverter stage in ps

  logic ClkVCO, ClkVCO1, ClkVCO2;  // Output clocks of each stage of the ring osccilator.

  real VCO_Period, VCO_Freq, CLKPVD_Freq;  // real number represents the period and frequency of ip2211ringpll_VCO. You can plot VCO_Freq vs. time to see how PLL locks.

  bit initial_trig;        // used to make sure the "always" block that includes design parameters, get accessed one time. (represents initial block).

  bit ClkVCO_div_by_2, ClkVCO_div_by_4, ClkVCO_div_by_8;

///============================================================================================================================================================================================
/// Ring Oscillator (3 Inverter stages), Td is the delay of each stage
///============================================================================================================================================================================================

  always @ (ClkVCO1 or VCO_RESET)  begin #Td ClkVCO   = (~VCO_RESET)? 1'b0 : !ClkVCO1;  end  // Kill output clock if PFD_EN is 0
  always @ (ClkVCO2)  begin #Td ClkVCO1  = !ClkVCO2;  end
  always @ (ClkVCO)   begin #Td ClkVCO2  = !ClkVCO ;  end

  // NOTE: what happens here is that once ClkVCO1 changes, its always block gets activated, and the last Td is taken to calculate ClkVCO
  // The same happens with each always block above.
  // so for one ClkVCO cycle, we have total of 6 changes in Ring Oscillator internal signals.
  // So at least 6 steps for Td (6 ClkSample edges) are required for each ClkVCO cycle.
  // assume a 5GHz ClkVCO Max freq, 200 ps period. And assume we will provide 10 steps, so every step is 20 ps. ClkSample may toggle every 20 ps.
  // You can not make the step so high, because in lock, phase error is small (~20 ps), so it should be less than that, or you can make it higher, but phase error will be higher
  // smaller steps give better accuracy but higher run time.


///============================================================================================================================================================================================
/// Calculating Td (Delay of each stage in Ring Oscillator)
///============================================================================================================================================================================================

  // For a ip2211ringpll_VCO --> Fvco = F0 + Kvco * Vctrl
  // For a 3-stage Ring Oscillator --> Fro = 1/(2*3*Td) where Td is the delay of each stage
  // So, by equating above equations (Fvco = Fro), and doing some math we get the following equation
  // Td = 1 /  6(F0 +  Kvco*Vctrl)
  // NOW, we deal with this as a ip2211ringpll_VCO, with controlled parameters for F0 and Kvco.
  // Td is calculated automatically from the given F0 and Kvco parameters

  always @(Vctrl) begin
    Td_pre = 1/( 6*(F0 + (Kvco * Vctrl) ) ) * 1000_000;   // Td is in ps --> look at units, this should be multiplied by 1000_000 to get ps
    //NOTE: from the equation above, if Vctrl = 0.6157, the denominator will be 0, giving an infinite value of Td_pre.
    // Also, if Vctrl is slightly higher than 0.6157, Td_pre will be very small, maybe 1 Hz, to Period in range of seconds, not acceptable.
    // Based on that, Vctrl value has to be protected from any wrong value (the designer should give a value that lies in the F-V curve)
    // NOTE: if Vctrl = 0.608 V --> F = 100 MHz. --> ALWAYS Limit Vctrl_min to 0.608, the minimum allowed freq of the ip2211ringpll_VCO is 100 MHz
    // because this ip2211ringpll_VCO is used in LCPLL as well that has different F-V curve, DO NOT limit Vctrl, just limit Td, so that minimum F is 100 MHz

    Td = ( ( 0 < Td_pre) && (Td_pre <= 1666.6667) ) ? Td_pre : Td;  // Td has to be less than or equal to  1666.6667 ps --> Minimum allowed frequency is 100 MHz
    //Td = Td_pre;   // It is allwed that Td be less than zero to terminate simulation

    //if ( 0 > Td_pre) begin $display ("[INFO]: ip2211ringpll_VCO output period cannot be negative, fixed to last positive value, please check ip2211ringpll_VCO F-V Curve, warning time = %0t" , $time); end
    //if (Td_pre > 1666.6667) begin $display ("[INFO]: ip2211ringpll_VCO output frequency cannot be less than 100 MHz, fixed to 100 MHz, please check ip2211ringpll_VCO F-V Curve, warning time = %0t" , $time); end
  end


///============================================================================================================================================================================================
/// Generating PVD Clock
///============================================================================================================================================================================================

// ip2211ringpll_VCO Clock Divided by 2
//-----------------------
   always @(posedge ClkVCO)          begin if (pvdmode !== 2'b00)  ClkVCO_div_by_2 = !ClkVCO_div_by_2; end

// ip2211ringpll_VCO Clock Divided by 4
//-----------------------
   always @(posedge ClkVCO_div_by_2) begin if (pvdmode[1] == 1'b1) ClkVCO_div_by_4 = !ClkVCO_div_by_4; end

// ip2211ringpll_VCO Clock Divided by 8
//-----------------------
   always @(posedge ClkVCO_div_by_4) begin if (pvdmode == 2'b11)   ClkVCO_div_by_8 = !ClkVCO_div_by_8; end

// Assign CLKPVD any of the above:
//--------------------------------
   assign CLKPVD = (pvdmode == 2'b00)? ClkVCO : (pvdmode == 2'b01)? ClkVCO_div_by_2 : (pvdmode == 2'b10)? ClkVCO_div_by_4 : ClkVCO_div_by_8;


///============================================================================================================================================================================================
/// Calculating ip2211ringpll_VCO related Period and Frequency
///============================================================================================================================================================================================

  always @(Td) begin VCO_Period = Td * 6; VCO_Freq = 1 / VCO_Period * 1000000; end  // VCO_Freq to be plotted vs. time to see PLL dynamics

  always @(VCO_Freq) CLKPVD_Freq = (pvdmode == 2'b00)? VCO_Freq : (pvdmode == 2'b01)? VCO_Freq/2 : (pvdmode == 2'b10)? VCO_Freq/4 : VCO_Freq/8;

///============================================================================================================================================================================================
/// Always block equivalent to initial block. All ip2211ringpll_VCO related parameters are defined here
///============================================================================================================================================================================================

  always @(Vctrl) begin  // at 0 time, VCO_RESET is zero, so PhaseErrorMag in (ip2211ringpll_PFD.sv) is zero, so Vctrl in (ip2211ringpll_SC_LPF.sv) triggers, so this "always" block triggers

   if (initial_trig == 1'b0) begin

    // Initial Values for ClkVCO:
    //------------------------------------------------
    #0 ClkVCO = 0; ClkVCO2 = 1; ClkVCO1 = 0;
       ClkVCO_div_by_2 = 0; ClkVCO_div_by_4 = 0; ClkVCO_div_by_8 = 0;

    // Important Parameters:
    //-------------------------------------------
    F0 = F0_VALUE;   // MHz
    Kvco = KVCO_VALUE;  // MHz/Volt

    // Calculating Td (Delay of each stage in Ring Oscillator):
    //---------------------------------------------------------

    Td_pre = 1/( 6*(F0 + (Kvco * Vctrl) ) ) * 1000_000;

    //Td = (Td_pre > 0)? Td_pre : 250;   // Td has to be greater than zero. Output clock period can not be zero or negative number.
    Td = Td_pre;   // It is allwed that Td be less than zero to terminate simulation

    if (~(( 0 < Td_pre) && (Td_pre <= 1666.6667))) begin $display (" [INFO]: ip2211ringpll_VCO output Frequency can't be less than 100 MHz, Please check ip2211ringpll_VCO F-V Curve, initial Vctrl with a reasonable value"); end

    initial_trig = 1'b1;  // to access this always block only one time in the beginning (as an initial block).
   end

  end


 endmodule

`endif

`ifndef ip2211ringpll_SECONDORDERLOOPFILTER_SV
`define ip2211ringpll_SECONDORDERLOOPFILTER_SV

module ip2211ringpll_SecondOrderLoopFilter (Vctrl, PhaseErrorMag, PhaseErrorSign);
`ifdef INTEL_EMULATION
  output logic Vctrl;
`else
  output real Vctrl;
`endif
  input bit PhaseErrorMag, PhaseErrorSign;

  real Ip;                // in Ampere
  real Rp;                // in Ohm
  real C1, C2;             // in Farad
  real Vctrl_R, Vctrl_EXP, Vctrl_Linear;    // in Volt
  real sign;              // 1 or -1
  logic ClkSample;

  logic PhaseErrorSign_delayed, PhaseErrorSign_EdgeDetect;

  real A, B, C, D, E;
  real Vfinal_exp, Vinitial_exp, Vinitial_linear, Linear_Const;
  real Vctrl_initial;
  real time_t;
  logic C2_bit;

   bit initial_trig;



  //////////////////////////////   Creating Edge Detector for PhaseErrorMag   /////////////////////////////////////////////////////////////
  assign #0.001 PhaseErrorSign_delayed = PhaseErrorSign;
  assign PhaseErrorSign_EdgeDetect = PhaseErrorSign ^ PhaseErrorSign_delayed;

  //////////////////////////////   Vctrl Generation   /////////////////////////////////////////////////////////////////////////////////////
  // Convertin phase error logic sign into real sign
  always @(PhaseErrorSign) begin
    if (PhaseErrorSign == 1'b1) sign = -1; else sign =  1;
  end

  always @(negedge ClkSample or posedge ClkSample or posedge PhaseErrorSign_EdgeDetect) begin

     if (PhaseErrorSign_EdgeDetect == 1'b1)
     begin
      time_t = 24'd0;
      Vinitial_exp = Vctrl_EXP;
      Vinitial_linear = Vctrl_Linear;
     end

     else
     begin
      time_t = time_t + 10;

      if (C2 > 0) Vctrl_EXP =  Vfinal_exp * sign  +  ( Vinitial_exp   -   Vfinal_exp * sign ) * ( 2.718281828**(E * time_t / 1000000/1000000) );
    //  else        Vctrl_EXP =  Vfinal_exp * sign * PhaseErrorMag  +  ( Vinitial_exp   -   Vfinal_exp * sign * PhaseErrorMag) * ( 2.718281828**(E * time_t / 1000000/1000000) );
      Vctrl_Linear = Vinitial_linear + Linear_Const * sign * time_t / 1000000 / 1000000;

     end


   // be careful, at begining of simulation, this statement will be valid, and Vctrl will be calculated
   // becuase at time 0, simulater considers ClkSample as negedge or posedge depending on initial value
   // in the testbench put the following, #0 Vctrl2 = 0.5; #1 Vctrl2 = 0.5 --> to guarantee right value
  end

  always @(PhaseErrorMag) begin if (C2 == 0) Vctrl_EXP = Vfinal_exp * sign * PhaseErrorMag; end  //  C2 == 0 --> exponential = 0, Vfinal_exp = Ip*R
  // Calculating Final Voltage Value
  always @( Vctrl_EXP or Vctrl_Linear) begin Vctrl = Vctrl_EXP + Vctrl_Linear; end

  // Creating ClkSample to linearize Vctrl2
  assign #10 ClkSample = (PhaseErrorMag == 1'b0)? 1'b0 : !ClkSample;  // PhaseError MUST be zero at #0 in order not to have unknown values for ClkSample(add reset signal to reset ip2211ringpll_PFD out at #0)
  ////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////    Parameters Values    /////////////////////////////////
  always @(PhaseErrorMag) begin
    // Initial Values for Vctrl_R and Vctrl_Cq (to be parametrized):
    //--------------------------------------------------------------
    if (initial_trig == 1'b0) begin
     //  Vinitial_exp = 0.00000001;
     //  Vinitial_linear = 0.00000001;


       time_t = 24'd0;
    // Important Parameters (to be parametrized):
    //-------------------------------------------
       Ip = 0.000001;                  // 1 uA
       Rp = 200;                          // 3.25K Ohm
       C1 = 0.000000000500;      // 1300 pF
       C2 = 0.000000000050;

    // Second Order Loop Filter Parameters:
    //------------------------------------
    A = Ip;
    B = Rp * C1;
    C = C1 + C2;
    D = C1 * C2 * Rp;
    E = (0-C)/D;
    Vfinal_exp = A * (B*C - D) / (C**2);
    Linear_Const = A / C;

    // At the beginning of simulation (time = 0fs), Vctrl_EXP is almost equal to Vinitial_exp, and Vctrl_linear is almost equal to Vinitial_linear
    // So Vctrl will have the initial value described below
    Vctrl_initial = 0.33;
    Vctrl = Vctrl_initial;  // If initially Vctrl = 0, there will be 0 iteration limmit Error, don't know why yet

    Vinitial_exp = Vfinal_exp/3;
    Vctrl_EXP = Vinitial_exp;  // Making sure that Vctrl_EXP should be equal to Vinitial_exp in the beginning of simulation.

    // If C2 = 0, this means first order loop filter, Vinitial should be on the cap only and the resisitance should have a zero voltage value
    // Vinitial_exp represents the resistance in the first loop filter when C2 = 0;
    Vinitial_linear = (C2>0)? (Vctrl_initial - Vinitial_exp) : Vctrl_initial;
    //Vctrl_Linear = Vinitial_linear; // Making sure that Vctrl_linear is equal to Vinitial_linear in the beginning of simulation

   //#1ps
   // Vctrl_EXP = Vinitial_exp;  // Making sure that Vctrl_EXP should be equal to Vinitial_exp in the beginning of simulation.

    Vctrl_Linear = Vinitial_linear; // Making sure that Vctrl_linear is equal to Vinitial_linear in the beginning of simulation
   //Vctrl_initial = 1;
      initial_trig = 1'b1;

   end

   end
  ////////////////////////////////////////////////////////////////////////////////////

endmodule

`endif

///========================================================================================================
///                                 ip2211ringpll_pll_inst_align Defines, Structures, Interfaces
///========================================================================================================

`ifndef ip2211ringpll_PLL_INST_ALIGN_VS
`define ip2211ringpll_PLL_INST_ALIGN_VS

//`include "soc_macros.sv"
//`include "ringpll_macros.sv"

module ip2211ringpll_pll_inst_align (
         input  logic       aligndis,         // Alignment scheme enable (during PLL lock)
         input  bit         clkin,            // Non-stop instrumentation clock from PLL ip2211ringpll_VCO
         input  logic       clkfb,            // Feedback clock from Q-div being used by PLL
         input  logic       clkref,           // Reference clock being used by PLL
         input  logic       reset_b,          // Async reset to avoid initial Xs
         output logic       haltclk           // Command to clock generator whithin PLL to stop output clock
      );

///========================================================================================================
/// Internal Signal Declarations
///========================================================================================================

   logic        init_reset, align_reset;
   logic        refclk_masked, fbclk_masked;
   logic        refclk_delay, fbclk_delay;
   bit   [1:0]  refclk_samp,  fbclk_samp;
   logic        refclk_rise,  fbclk_rise;
   logic [2:0]  haltclk_delay;
   logic        haltclkin;
   logic        inhibit_correction;

///========================================================================================================
/// Main Procedure
///========================================================================================================

   // Initialize all states with the following reset to avoid Xs if the
   //  "aligndis" reset never asserts (common in lower level DUTs)
   //
   `ip2211ringpll_ASYNC_SET_MSFF(init_reset, 1'b0, clkin, ~reset_b)
   always_comb align_reset = init_reset | aligndis;


   // Randomly convert any Xs on the reference or feedback clock to known 
   //  values so the below code does not get corrupted by Xs on the inputs.
   //
   `ip2211ringpll_RANDOM_VAL_WHEN_X(refclk_masked, clkref, 1'b1)
   `ip2211ringpll_RANDOM_VAL_WHEN_X(fbclk_masked,  clkfb,  1'b1)

   // Delay the clkref and clkfb by 1 VCS tick before sampling them with
   //  clkin to avoid races in VCS when sampled and sampling clock change
   //  in the same tick.
   //
   `ip2211ringpll_NB_ASSIGN(refclk_delay, refclk_masked)
   `ip2211ringpll_NB_ASSIGN(fbclk_delay,  fbclk_masked)

   // Sample the clkref and clkfb with falling clkin and do a rising edge
   //  detect give an indication of the rising clkref and clkfb edges in
   //  the clkin domain. Mask out subsequent clkfb edges immediately after
   //  an alignment correction.
   //
   `ip2211ringpll_DUAL_EDGE_MSFF(refclk_samp, {refclk_samp[0],refclk_delay}, clkin)
   `ip2211ringpll_DUAL_EDGE_MSFF(fbclk_samp,  {fbclk_samp[0], fbclk_delay},  clkin)

   always_comb refclk_rise = (refclk_samp == 2'b01);
   always_comb fbclk_rise  = (fbclk_samp  == 2'b01) & ~inhibit_correction;


   // If enabled to correct the clkfb alignment, use the rising clkfb to 
   //  set the haltclk control (used to gate the clkfb source clock with 
   //  clkin cycle granularity) and the rising clkref to reset it.
   //
   // When clkref and clkfb are aligned, the reset condition should take
   //  priority and prevent haltclk from asserting.
   //
   always_comb haltclkin = (refclk_rise)? 1'b0 : (fbclk_rise)? 1'b1 : haltclk;
   `ip2211ringpll_ASYNC_RST_MSFF(haltclk, haltclkin, clkin, align_reset)


   // Once the haltclk control asserts we need to prevent it from asserting
   //  again for a few clkref cycles to allow things to settle. Sample
   //  haltclk with clkref to create a delayed version with which to
   //  inhibit successive assertions. Force the state high during reset to
   //  allow some time for clkfb to settle after reset de-asserts.
   //
   `ip2211ringpll_EN_ASYNC_RSTD_MSFF(haltclk_delay, {haltclk_delay[1:0],haltclk}, clkin, refclk_rise, align_reset, '1)
   always_comb inhibit_correction = |haltclk_delay;

endmodule   // module ip2211ringpll_pll_inst_align

`endif // ip2211ringpll_PLL_INST_ALIGN_VS


`ifndef ip2211ringpll_cpafdivcore_SV
`define ip2211ringpll_cpafdivcore_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
`ifndef ip2211ringpll_SVA_OFF
   //`include "intel_checkers.sv"
`endif

module ip2211ringpll_cpafdivcore 
//#( parameter     RATIO_BITS = 10)
(
   //input  logic [8:0]   ratio2x,
   input  logic [10:0]   ratio2x,
   input  logic         clkinb,
   output logic         clkout,
   output logic         cueh,
   output logic         rstd,
   input  logic         rst
);

///========================================================================================================
/// Reset Generation
///========================================================================================================

   logic RstCntMH;

   // Rename reset
   //
   always_comb RstCntMH = rst;


   // Reset to ip2211ringpll_cpaclkphdelana
   //
   always_comb rstd = rst;


///========================================================================================================
/// Reload Logic
///========================================================================================================

   logic [6:0] CountMH;
   logic Clk0MH;
   logic ReloadMH;
   logic CountToZeroMH;
   logic RatioOddMH;
   logic Zero61MH;
   logic Zero63MH;
   logic HiPhaseMH; // indicates whether divider is currently outputing clkout=1

   // More readable name for Odd ratio
   //
   always_comb RatioOddMH = ratio2x[1];

   // Compute the segmented zero values to execute a reload
   //
   always_comb begin : ZERO_CALCULATION
      Zero61MH = (CountMH[6:1] == 6'd0);
      Zero63MH = (CountMH[6:3] == 4'd0);
   end : ZERO_CALCULATION

   always_comb begin : RELOAD
      // Determine whether or not to count to zero on a reload
      //   Changes between 0/1 every cycle when the ratio is odd.
      //
      CountToZeroMH = (!HiPhaseMH && RatioOddMH);

      // Reload the counter based on the count to zero flag.
      //   If counting to zero, wait until counter matches zero,
      //   else reload at one.
      //
      ReloadMH = (CountToZeroMH) ? (CountMH == 7'd0) :
                                   (CountMH <= 7'd1) ;

   end : RELOAD

///========================================================================================================
/// Segmented 1+2+4 Reloadable Counter
///========================================================================================================

   logic [1:0] CountM1Nxt21MH;
   logic [3:0] CountM1Nxt63MH;
   logic [6:0] CountStartMH;
   logic [6:0] RatioD2MH;
   logic [6:0] CountNxtMH;
   logic       Clk21MH, Clk63MH;
   logic       EnClk21MH, EnClk63MH;
   logic       EnClk21ML, EnClk63ML;

   `ip2211ringpll_CLK_NOR(Clk0MH, clkinb, 1'b0)


   // Segmented counter declaration
   //
   //`ip2211ringpll_RST_MSFF(CountMH[0],   CountNxtMH[0],   Clk0MH,  RstCntMH)
   //`ip2211ringpll_RST_MSFF(CountMH[2:1], CountNxtMH[2:1], Clk21MH, RstCntMH)
   //`ip2211ringpll_RST_MSFF(CountMH[6:3], CountNxtMH[6:3], Clk63MH, RstCntMH)
   `ip2211ringpll_ASYNC_RST_MSFF(CountMH[0],   CountNxtMH[0],   Clk0MH,  RstCntMH)
   `ip2211ringpll_ASYNC_RST_MSFF(CountMH[2:1], CountNxtMH[2:1], Clk21MH, RstCntMH)
   `ip2211ringpll_ASYNC_RST_MSFF(CountMH[6:3], CountNxtMH[6:3], Clk63MH, RstCntMH)

   always_comb EnClk21MH = (~( CountMH[0]  ) || ReloadMH);
   always_comb EnClk63MH = (~(|CountMH[2:0]) || ReloadMH);

   // Count Clock Generation
   //
   `ip2211ringpll_LATCH(EnClk21ML, EnClk21MH, clkinb)
   `ip2211ringpll_LATCH(EnClk63ML, EnClk63MH, clkinb)

   `ip2211ringpll_CLK_NOR(Clk21MH, clkinb, ~EnClk21ML)
   `ip2211ringpll_CLK_NOR(Clk63MH, clkinb, ~EnClk63ML)

   // Count start is ratio / 2
   //
   //always_comb CountStartMH    = ratio2x[8:2];
   always_comb CountStartMH    = ratio2x[8:2];

   always_comb begin : COUNT_NXT

      CountM1Nxt21MH = (CountMH[2:1] - 2'b01);
      CountM1Nxt63MH = (CountMH[6:3] - 4'b0001);

      CountNxtMH[0]   = (ReloadMH) ? CountStartMH [0]  :
                                     ~CountMH[0]       ;

      CountNxtMH[2:1] = (Zero61MH) ? CountStartMH [2:1] :
                                     CountM1Nxt21MH     ;

      CountNxtMH[6:3] = (Zero63MH) ? CountStartMH [6:3] :
                                     CountM1Nxt63MH     ;

   end : COUNT_NXT


///========================================================================================================
/// Output Clock
///========================================================================================================

   logic PhaseStretchML;

   // Every reload changes the output state of the divider clkout
   //  Since the counter uses /2 ratio value, this serves as a toggle flop
   //  for the state of the output clock.
   //
   //`ip2211ringpll_EN_RST_MSFF(HiPhaseMH, ~HiPhaseMH, Clk0MH, ReloadMH, RstCntMH)
   `ip2211ringpll_EN_ASYNC_RST_MSFF(HiPhaseMH, ~HiPhaseMH, Clk0MH, ReloadMH, RstCntMH)

   // For odd ratios, we need to phase stretch
   //
   `ip2211ringpll_LATCH_P(PhaseStretchML, HiPhaseMH, Clk0MH)

   always_comb begin : CLKOUT
      clkout = (PhaseStretchML & RatioOddMH) || HiPhaseMH;
   end : CLKOUT

///========================================================================================================
/// Pulse extention logic
///========================================================================================================

   logic ForceSwStateLowMH;

   // For powerup, force a low state until everything factoring into the
   //   cueh signal is stable.
   //
   `ip2211ringpll_ASYNC_SET_LATCH(ForceSwStateLowMH, 1'b0, HiPhaseMH, rst)

   // Switch the clock state (clkinb) when we are in half int mode and
   //   clkout is 0 (switch every cycle)
   //
   always_comb begin : CLKIN_STATE_SELECT
      cueh = ForceSwStateLowMH ? 1'b0                    :
                                 ratio2x[0] & ~HiPhaseMH ;
   end : CLKIN_STATE_SELECT


///========================================================================================================
/// Assertions
///========================================================================================================

   `ifndef ip2211ringpll_SVA_OFF
      `ip2211ringpll_ASSUMEC_MUST(A_ratio_gte_2,
                    //(ratio2x[8:1] >= 8'd2),
                    (ratio2x[10:1] >= 10'd2),
                    (rst!==1'b0),
                    `ip2211ringpll_ERR_MSG("[PLL-AIP] F-divider ratio must be set >=2"));

      `ip2211ringpll_ASSERTC_FORBIDDEN(R_fdiv_core_reload_only_when_count_lte_1,
                         (ReloadMH & (CountMH > 7'd1)),
                         (rst!==1'b0),
                         `ip2211ringpll_ERR_MSG("[PLL-AIP] F-divider reloaded its internal counter unexpectedly. The counter should only reload when Count<=1"));
   `endif

endmodule

`endif


`ifndef ip2211ringpll_CPAFDIVTOP_SV
`define ip2211ringpll_CPAFDIVTOP_SV

//`include "ip2211ringpll_cpafdivcore.sv"
//`include "ip2211ringpll_cpaclkphdelana.sv"
//`include "soc_macros.sv"

module ip2211ringpll_cpafdivtop 
//#( parameter     RATIO_BITS = 10)
(
   input  logic         clkin,
   input  logic         rst,
   input  logic [10:0]   ratio2x,

   output logic         clkout
);

///========================================================================================================
/// Module Begin
///========================================================================================================

   logic cueh;
   logic clkinb;
   logic rstd;


   // Phase delay insertion for half integer ratios
   //
   ip2211ringpll_cpaclkphdelana phdel_core (
      // in netlist it is not tied to 1 .vccxx   ( 1'b1    ),
      .rst     ( rstd    ),
      .cueh    ( cueh    ),
      .clkin   ( clkin   ),
      .clkoutb ( clkinb  )
   );
   
   // F-divider counter cores for integer logic
   //
   ip2211ringpll_cpafdivcore    fdiv_core ( .* );

///========================================================================================================
/// Module End
///========================================================================================================

endmodule

`endif

`ifndef ip2211ringpll_cpafdivcore_SV
`define ip2211ringpll_cpafdivcore_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
`ifndef ip2211ringpll_SVA_OFF
   //`include "intel_checkers.sv"
`endif

module ip2211ringpll_cpafdivcore 
//#( parameter     RATIO_BITS = 10)
(
   //input  logic [8:0]   ratio2x,
   input  logic [10:0]   ratio2x,
   input  logic         clkinb,
   output logic         clkout,
   output logic         cueh,
   output logic         rstd,
   input  logic         rst
);

///========================================================================================================
/// Reset Generation
///========================================================================================================

   logic RstCntMH;

   // Rename reset
   //
   always_comb RstCntMH = rst;


   // Reset to ip2211ringpll_cpaclkphdelana
   //
   always_comb rstd = rst;


///========================================================================================================
/// Reload Logic
///========================================================================================================

   logic [6:0] CountMH;
   logic Clk0MH;
   logic ReloadMH;
   logic CountToZeroMH;
   logic RatioOddMH;
   logic Zero61MH;
   logic Zero63MH;
   logic HiPhaseMH; // indicates whether divider is currently outputing clkout=1

   // More readable name for Odd ratio
   //
   always_comb RatioOddMH = ratio2x[1];

   // Compute the segmented zero values to execute a reload
   //
   always_comb begin : ZERO_CALCULATION
      Zero61MH = (CountMH[6:1] == 6'd0);
      Zero63MH = (CountMH[6:3] == 4'd0);
   end : ZERO_CALCULATION

   always_comb begin : RELOAD
      // Determine whether or not to count to zero on a reload
      //   Changes between 0/1 every cycle when the ratio is odd.
      //
      CountToZeroMH = (!HiPhaseMH && RatioOddMH);

      // Reload the counter based on the count to zero flag.
      //   If counting to zero, wait until counter matches zero,
      //   else reload at one.
      //
      ReloadMH = (CountToZeroMH) ? (CountMH == 7'd0) :
                                   (CountMH <= 7'd1) ;

   end : RELOAD

///========================================================================================================
/// Segmented 1+2+4 Reloadable Counter
///========================================================================================================

   logic [1:0] CountM1Nxt21MH;
   logic [3:0] CountM1Nxt63MH;
   logic [6:0] CountStartMH;
   logic [6:0] RatioD2MH;
   logic [6:0] CountNxtMH;
   logic       Clk21MH, Clk63MH;
   logic       EnClk21MH, EnClk63MH;
   logic       EnClk21ML, EnClk63ML;

   `ip2211ringpll_CLK_NOR(Clk0MH, clkinb, 1'b0)


   // Segmented counter declaration
   //
   //`ip2211ringpll_RST_MSFF(CountMH[0],   CountNxtMH[0],   Clk0MH,  RstCntMH)
   //`ip2211ringpll_RST_MSFF(CountMH[2:1], CountNxtMH[2:1], Clk21MH, RstCntMH)
   //`ip2211ringpll_RST_MSFF(CountMH[6:3], CountNxtMH[6:3], Clk63MH, RstCntMH)
   `ip2211ringpll_ASYNC_RST_MSFF(CountMH[0],   CountNxtMH[0],   Clk0MH,  RstCntMH)
   `ip2211ringpll_ASYNC_RST_MSFF(CountMH[2:1], CountNxtMH[2:1], Clk21MH, RstCntMH)
   `ip2211ringpll_ASYNC_RST_MSFF(CountMH[6:3], CountNxtMH[6:3], Clk63MH, RstCntMH)

   always_comb EnClk21MH = (~( CountMH[0]  ) || ReloadMH);
   always_comb EnClk63MH = (~(|CountMH[2:0]) || ReloadMH);

   // Count Clock Generation
   //
   `ip2211ringpll_LATCH(EnClk21ML, EnClk21MH, clkinb)
   `ip2211ringpll_LATCH(EnClk63ML, EnClk63MH, clkinb)

   `ip2211ringpll_CLK_NOR(Clk21MH, clkinb, ~EnClk21ML)
   `ip2211ringpll_CLK_NOR(Clk63MH, clkinb, ~EnClk63ML)

   // Count start is ratio / 2
   //
   //always_comb CountStartMH    = ratio2x[8:2];
   always_comb CountStartMH    = ratio2x[10:2];

   always_comb begin : COUNT_NXT

      CountM1Nxt21MH = (CountMH[2:1] - 2'b01);
      CountM1Nxt63MH = (CountMH[6:3] - 4'b0001);

      CountNxtMH[0]   = (ReloadMH) ? CountStartMH [0]  :
                                     ~CountMH[0]       ;

      CountNxtMH[2:1] = (Zero61MH) ? CountStartMH [2:1] :
                                     CountM1Nxt21MH     ;

      CountNxtMH[6:3] = (Zero63MH) ? CountStartMH [6:3] :
                                     CountM1Nxt63MH     ;

   end : COUNT_NXT


///========================================================================================================
/// Output Clock
///========================================================================================================

   logic PhaseStretchML;

   // Every reload changes the output state of the divider clkout
   //  Since the counter uses /2 ratio value, this serves as a toggle flop
   //  for the state of the output clock.
   //
   //`ip2211ringpll_EN_RST_MSFF(HiPhaseMH, ~HiPhaseMH, Clk0MH, ReloadMH, RstCntMH)
   `ip2211ringpll_EN_ASYNC_RST_MSFF(HiPhaseMH, ~HiPhaseMH, Clk0MH, ReloadMH, RstCntMH)

   // For odd ratios, we need to phase stretch
   //
   `ip2211ringpll_LATCH_P(PhaseStretchML, HiPhaseMH, Clk0MH)

   always_comb begin : CLKOUT
      clkout = (PhaseStretchML & RatioOddMH) || HiPhaseMH;
   end : CLKOUT

///========================================================================================================
/// Pulse extention logic
///========================================================================================================

   logic ForceSwStateLowMH;

   // For powerup, force a low state until everything factoring into the
   //   cueh signal is stable.
   //
   `ip2211ringpll_ASYNC_SET_LATCH(ForceSwStateLowMH, 1'b0, HiPhaseMH, rst)

   // Switch the clock state (clkinb) when we are in half int mode and
   //   clkout is 0 (switch every cycle)
   //
   always_comb begin : CLKIN_STATE_SELECT
      cueh = ForceSwStateLowMH ? 1'b0                    :
                                 ratio2x[0] & ~HiPhaseMH ;
   end : CLKIN_STATE_SELECT


///========================================================================================================
/// Assertions
///========================================================================================================

   `ifndef ip2211ringpll_SVA_OFF
      `ip2211ringpll_ASSUMEC_MUST(A_ratio_gte_2,
                    //(ratio2x[8:1] >= 8'd2),
                    (ratio2x[10:1] >= 10'd2),
                    (rst!==1'b0),
                    `ip2211ringpll_ERR_MSG("[PLL-AIP] F-divider ratio must be set >=2"));

      `ip2211ringpll_ASSERTC_FORBIDDEN(R_fdiv_core_reload_only_when_count_lte_1,
                         (ReloadMH & (CountMH > 7'd1)),
                         (rst!==1'b0),
                         `ip2211ringpll_ERR_MSG("[PLL-AIP] F-divider reloaded its internal counter unexpectedly. The counter should only reload when Count<=1"));
   `endif

endmodule

`endif


`ifndef ip2211ringpll_LJPLL_PLLFBGEN_SV
`define ip2211ringpll_LJPLL_PLLFBGEN_SV

//`ifndef VCSSIM_OR_EMU
//   `ifdef INTC_EMULATION
//      `define VCSSIM_OR_EMU
//   `endif
//`endif
//   
//`ifndef VCSSIM_OR_EMU
//   `ifdef VCSSIM
//      `define VCSSIM_OR_EMU
//   `endif
//`endif
//
//`ifdef VCSSIM_OR_EMU
//   `ifndef ip2211ringpll_LJPLL_MSV
//      `define VCSSIM_OR_EMU_NOT_MSV
//   `endif
//`endif

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
////`include "cpafdivtop.sv"
//`include "ringpll_macros.sv"
//`ifdef VCSSIM_OR_EMU_NOT_MSV
   //`include "pll_inst_align.sv"
//`endif

module ip2211ringpll_ljpll_pllfbgen
//#(
//`ifndef ip2211ringpll_LJPLL_MSV
//`ifdef VCSSIM
//   parameter bit INTC_USE_DETAILED_AIP_MODEL = 1,
//`endif
//`endif
//   parameter RATIO_BITS =10 
//)
(

   `ifndef INTC_NO_VCSSIM_OR_EMU_NOT_MSV
      // Use reference clock to align the feedback clock in simulation
      //
      input  logic ClkRefXXH,

      // Halt clock should be used to reset the lock detector
      //
      output logic pllfbgen__haltclk_inst,
   `endif

   `ifdef ip2211ringpll_LJPLL_NO_UPF_SUPPORT
      input wire   vccpll,
   `endif

   input  logic reset_b_xxl,
   input  logic idv_gate_en,
   input  logic pll_core__clk_pll_div1,
   input  logic post_dist_mux__ClkPostDistMH,
   input  logic pfdennh,
   input  logic tight_loop,
   input  logic tlctrl_hip__TightLoopMnn0L,
   input  logic tlctrl_hip__GateGridClkMnnnL,
   input  logic                      half_int,
   input  logic [9:0] ratio,
//   output logic [9:0] pll_fbgen__RatioSampMXH,
   output logic pll_fbgen__tight_loop,
//   output logic pll_fbgen__ClkPllFdivMH,
   //output logic ClkFbMXH
   output logic clkfb,
   output logic clkfb2
);

///========================================================================================================
/// Module Begin
///========================================================================================================
  
   parameter bit INTC_USE_DETAILED_AIP_MODEL = 0;
   logic ClkPllMH;
   logic ClkPllSyncMH;
   logic QdivReset_b_MnnnH;
   logic ClkPostDistGateMH;
   logic pll_fbgen__ClkPllFdivMH;
   logic ClkFbMXH;
 
   // Squash X for syncronizer (modeling)
   //
   `ip2211ringpll_RANDOM_VAL_WHEN_X(ClkPllSyncMH, ClkPllMH, 1'b1)

   // Only deassert the reset after it has been sampled downstream by ClkPllMH
   //
   //   SPEC Assumption: This assumes that the IDV chain is not changing at
   //   all between PLL enable and ip2211ringpll_PFD Enable assertion
   //
   //   When the PLL IDV is targeted, openloop is assumed to be asserted
   //   before PLL enable is asserted.  This allows the IDV chain to toggle
   //   as it sees fit.
   //
   `ip2211ringpll_ASYNC_RST_2MSFF_META(QdivReset_b_MnnnH, (pfdennh | idv_gate_en), ClkPllSyncMH, reset_b_xxl)

   // Tight loop select - could come from tap OR tight loop lock mode
   //
   always_comb begin : TIGHT_LOOP_SELECT
      pll_fbgen__tight_loop =  tight_loop | (~ tlctrl_hip__TightLoopMnn0L) ;

   end : TIGHT_LOOP_SELECT

   // Gate grid clock from the tight loop lock mode FSM
   // 
   `ip2211ringpll_CLKAND(ClkPostDistGateMH, post_dist_mux__ClkPostDistMH, tlctrl_hip__GateGridClkMnnnL)

   // Tight Loop Mux
   //   Selects between a post distribution clock, odcs clock
   //   and the internal pll clock output as an input to
   //   the feedback divider
   //
   always_comb begin : FEEDBACK_SELECT
     
      // Feedback Clock Mux Selection Logic
      //                  
      //        tight_loop     | CLK To F-Div
      //   -------------------------------------------------------------
      //           0           | POST DIST CLOCK or  ODCS DLL Clock Out
      //           1           | PLL Div1 Clock (From ANA)
      //
      ClkPllMH = pll_fbgen__tight_loop ? pll_core__clk_pll_div1
                                       : ClkPostDistGateMH       ;

   end : FEEDBACK_SELECT


   // Ratio Sampling on FBCLK to facilitate SIP/HIP timing
   //  SIP drives the ratio on rising FBCLK and has falling REFCLK logic
   //  fan-in. Sampling in the HIP on rising FBCLK allows a safe transfer
   //  and lets partition timing analyze the path properly.
   //  To initialize the ratio before the divider is released from reset we
   //  use the raw ratio, then switch to the sampled ratio after seeing
   //  a couple of feedback clocks. Note the divider is reset by !pfden
   //  synchronized to the full speed clock.
   //
   logic [9:0] RatioSampMXH, Ratio2FbDivMXH;
   logic                  HalfIntSampMXH, HalfInt2FbDivMXH;
   logic                  SelRatioSampMXH, SampEnable;

   `ip2211ringpll_EN_MSFF({RatioSampMXH, HalfIntSampMXH}, {ratio, half_int}, ClkFbMXH, SampEnable)

   `ip2211ringpll_ASYNC_RST_2MSFF_META(SelRatioSampMXH, 1'b1, ClkFbMXH, pfdennh)

   always_comb {Ratio2FbDivMXH, HalfInt2FbDivMXH} = (SelRatioSampMXH)? {RatioSampMXH, HalfIntSampMXH} : {ratio, half_int};


   // Send the sampled ratio out to SyncGen block
   //
   //always_comb pll_fbgen__RatioSampMXH = Ratio2FbDivMXH;


   // If VCSSIM_OR_EMU, Align feedback and PLL clocks unless using the detailed model
   //
   `ifndef INTC_NO_VCSSIM_OR_EMU_NOT_MSV
      logic haltclk_inst_lat;
      logic clkfb_inst;

        `ifndef ip2211ringpll_NO_VCSSIM
      
// NOTE: Following is commented out dur to Macroprep parameter issue.
//       Later on uncomment it so AIP model can be tested. -
      if (INTC_USE_DETAILED_AIP_MODEL) begin : FBDIV_FEEDTHRU
         assign pll_fbgen__ClkPllFdivMH = ClkPllMH;
         assign SampEnable              = 1'b1;
      end : FBDIV_FEEDTHRU
      else begin : INST_ALIGN
      `endif

      always_comb clkfb_inst = ClkFbMXH;

      // Prevent the ratio from changing after sampling it from the SIP because 
      // the standard PLL behavioral model does not support SSC or frac-N
      //
 assign SampEnable      = !SelRatioSampMXH;

      ip2211ringpll_pll_inst_align ip2211ringpll_pll_inst_align (
         .aligndis   (1'b0),
         .clkin      (ClkPllMH),
         .clkfb      (clkfb_inst),
         .clkref     (ClkRefXXH),
         .reset_b    (pfdennh),
         .haltclk    (pllfbgen__haltclk_inst)
      );

      `ip2211ringpll_LATCH_P(haltclk_inst_lat, pllfbgen__haltclk_inst, ClkPllMH)
      always_comb pll_fbgen__ClkPllFdivMH = ClkPllMH & ~haltclk_inst_lat;
      `ifndef ip2211ringpll_NO_VCSSIM
      end : INST_ALIGN
      `endif
   `else   
      assign pll_fbgen__ClkPllFdivMH = ClkPllMH;
      assign SampEnable              = 1'b1;
   `endif

   // Feedback Divider Instantiation
   //
   ip2211ringpll_cpafdivtop  fdiv (
      .clkin      (pll_fbgen__ClkPllFdivMH),
      .rst        (~QdivReset_b_MnnnH),
      .ratio2x    ({Ratio2FbDivMXH, HalfInt2FbDivMXH}),
      .clkout     (ClkFbMXH)
   );

	// Output buffers
	assign clkfb = ClkFbMXH;
	assign clkfb2 = ClkFbMXH;

///========================================================================================================
/// Assertions
///========================================================================================================

/* -----\/----- EXCLUDED -----\/-----
   `ifndef ip2211ringpll_SVA_OFF
      `ip2211ringpll_ASSERTS_TRIGGER(R_sampled_and_raw_ratio_equal_at_ratio_switch,
                    $rose(SelRatioSampMXH), 
                    $past({ratio,half_int})==$past({RatioSampMXH,HalfIntSampMXH}),
                    posedge ClkFbMXH,
                    !reset_b_xxl,
                  `ip2211ringpll_ERR_MSG("[LJPLL] Sampled feedback ratio (%d) is not equal to the raw ratio (%d) at ratio mux switch",
                           {RatioSampMXH,HalfIntSampMXH}, {ratio,half_int}));
   `endif
 -----/\----- EXCLUDED -----/\----- */

///========================================================================================================
/// Module End
///========================================================================================================

endmodule

`endif


`ifndef ip2211ringpll_PLLLSVCCPLL2VCCDIST_SV
`define ip2211ringpll_PLLLSVCCPLL2VCCDIST_SV

//`include "soc_power_macros.sv"

module ip2211ringpll_plllsvccpll2vccdist (
   `ifdef ip2211ringpll_LJPLL_NO_UPF_SUPPORT
      input  wire vccpll,
      input  wire vccdist,
   `endif
  
   input  logic pll_core__clk_pll_div1,
   input  logic gate_trunk_sync__GateClkTrunkML,
   input  logic reset_b_xxl,

   output logic pll_core__clk_pll_div1_ls_dist,
   output logic gate_trunk_sync__GateClkTrunkML_ls_dist
);

`ifdef ip2211ringpll_LJPLL_NO_UPF_SUPPORT
   `ip2211ringpll_LS_WITH_AND_FW_CLK(pll_core__clk_pll_div1_ls_dist,  vccdist, pll_core__clk_pll_div1, vccpll, reset_b_xxl)
  // `ip2211ringpll_LS_WITH_AND_FW    (gate_trunk_sync__GateClkTrunkML_ls_dist,  vccdist, gate_trunk_sync__GateClkTrunkML, vccpll, reset_b_xxl)
`else
   assign pll_core__clk_pll_div1_ls_dist          = pll_core__clk_pll_div1;
  // assign gate_trunk_sync__GateClkTrunkML_ls_dist = gate_trunk_sync__GateClkTrunkML;
`endif

endmodule

`endif

`ifndef ip2211ringpll_GATE_TRUNK_SYNC_SV
`define ip2211ringpll_GATE_TRUNK_SYNC_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"

module ip2211ringpll_gate_trunk_sync (
   input  logic Reset_b_XXL,
   input  logic ClkFbMXH,
   input  logic pll_core__clk_pll_div1,
   input  logic tllm_gate_clk_trunk,
   output logic gate_trunk_sync__GateClkTrunkML
);

///========================================================================================================
/// Syncronize Clock Trunk Gating
///========================================================================================================
   
   logic GateClkTrunkRstXXL;
   logic GateClkTrunkMXH;
   logic GateClkTrunkMH;
   logic GateClkTrunkML;
   logic ClkPllMH_b;

   // Generate reset condition from PLL Enable
   //
   assign GateClkTrunkRstXXL = ~Reset_b_XXL;

   // Syncronize falling refclk aligned tllm_gate_clk_trunk to rising edge
   //   feedback and rising edge MCLK
   //
   //   Handshake:
   //    Falling Refclk -> Rising Feedback Clock -> Rising MCLK
   //
   `ip2211ringpll_ASYNC_RST_MSFF(GateClkTrunkMXH, tllm_gate_clk_trunk, ClkFbMXH,               GateClkTrunkRstXXL)
   `ip2211ringpll_ASYNC_RST_MSFF(GateClkTrunkMH,  GateClkTrunkMXH,     pll_core__clk_pll_div1, GateClkTrunkRstXXL)

   // Add a latch so that the clock gate only changes on falling edge of
   // MCLK
   //
   `ip2211ringpll_CLKINV(ClkPllMH_b, pll_core__clk_pll_div1)
   `ip2211ringpll_ASYNC_RST_LATCH(GateClkTrunkML, GateClkTrunkMH, ClkPllMH_b, GateClkTrunkRstXXL)
   
   // Always gate the clock distribution immediately whenever the clock
   //   trunk gate asserts
   //
   always_comb begin : ASYNC_DRIVE
      gate_trunk_sync__GateClkTrunkML = (tllm_gate_clk_trunk | GateClkTrunkML);
   end : ASYNC_DRIVE

endmodule

`endif

`ifndef ip2211ringpll_PLL_GLITCHLESSMUX_SV 
`define ip2211ringpll_PLL_GLITCHLESSMUX_SV 

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "ringpll_macros.sv"

module ip2211ringpll_pll_glitchlessmux 
(
   `ifndef ip2211ringpll_INTC_NO_PWR_PINS
      input wire vccpll,
      input wire vss,
   `endif

   input  logic bypass,
   input  logic bypassen,
   input  logic pllclk,
   input  logic refclk,
   input  logic rb,
   output logic muxclk
);

///========================================================================================================
/// Module Begin
///========================================================================================================
      //   State Table:
      //   | bypass | bypassen     |  muxclk
      //   -------------------------------------------
      //   |    1   |     1        |  refclk
      //   |    1   |     0        |  vss
      //   |    0   |     0        |  pllclk 
      //   |    0   |     1        |  pllclk
      //

    logic pllclki;
    logic refclki;
    logic n4;
    logic n3;
    logic n2;
    logic n1;
    logic refclkbuf;
    logic refclkb;
    logic enref;
    logic enrefb;
    logic enref2;
    logic bypassb;
    logic pllclkb;
    logic pllclkbuf;
    logic enclk;
logic bypassb_shwe ;



    //ip2211ringpll_ASYNC_RST_2MSFF_META(q,i,clkin,rst_b)
    `ip2211ringpll_ASYNC_RST_2MSFF_META(n4,n3,refclkbuf,rb)

    //ip2211ringpll_ASYNC_RST_LATCH(q,i,clock,rst)
    //`ip2211ringpll_ASYNC_RST_LATCH(enref,n4,refclkb,rb)
    //ip2211ringpll_RST_LATCH_P(q,i,clock,rst)
    //`ip2211ringpll_RST_LATCH_P(enref,n4,refclkb,rb)

    //`ASYNC_RST_LATCH_P(enref,n4,refclkb,rb)
        //`define ASYNC_RST_LATCH_P(q,i,clock,rst)      
   	always_comb begin : async_reset_latch_p       
         if      (~rb) enref <= '0; /* lintra s-30529 */ 
         else if (refclkb) enref <= n4;                
   	end : async_reset_latch_p



    `ip2211ringpll_ASYNC_RST_2MSFF_META(n2,n1,pllclkbuf,rb)
    //`ip2211ringpll_ASYNC_RST_LATCH(enclk, n2,pllclkb, rb)
    //`ip2211ringpll_RST_LATCH_P(enclk, n2,pllclkb, rb)

    //`ASYNC_RST_LATCH_P(enclk, n2,pllclkb, rb)
        //`define ASYNC_RST_LATCH_P(q,i,clock,rst)    
   	always_comb begin : async_reset_latch_p_1    
         if      (~rb) enclk <= '0; /* lintra s-30529 */ 
         else if (pllclkb) enclk <= n2;                 
   	end : async_reset_latch_p_1

    always_comb begin : MUX

 bypassb_shwe = ~bypassen | bypass ;
// REFCLK path
//
    n3 = (bypassb_shwe & ~enclk);
    refclkbuf = refclk;
    refclkb = ~refclk;

    enref2 = (bypassen && enref);
    refclki = ~(enref2 && refclk);

// PLLCLK path
//
    bypassb = ~bypass;
    enrefb = ~enref;
    n1 = (enrefb && ~bypassb_shwe);
// fix for SPG LINT 60000_a
// bypassb_shwe = ~bypassen | bypass ;
    pllclkb = ~pllclk;
    pllclkbuf = pllclk;
    pllclki = ~(enclk && pllclk);
 
// Output MUX clock
//
    muxclk = ~(pllclki & refclki); 
   end : MUX

endmodule
`endif

`ifndef ip2211ringpll_cpadcaana_SV
`define ip2211ringpll_cpadcaana_SV

`ifndef ip2211ringpll_NO_VCSSIM
//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "intel_checkers.vs"
`endif

///=====================================================================================================================
///                                  Defines, Structures, Interfaces
///=====================================================================================================================

module ip2211ringpll_cpadcaana (
      `ifndef ip2211ringpll_NO_VCSSIM 
         input   logic         sva_reset,
      `endif
         input   logic [1:0]   cb,
         input   logic          clkin,
         input   logic [5:0]    ctrl,
         input   logic          vccxx,

         output  logic          clkout
);


///=====================================================================================================================
///                                  Non-VCS simulation code
///=====================================================================================================================
`ifdef ip2211ringpll_LJPLL_PERF_SIM
assign clkout = clkin;
`else
// To disable ev injection inside VCSSIM instrumentation code
//`ifndef VCSSIM
`ifdef ip2211ringpll_NO_VCSSIM

   always_comb clkout = clkin;

`endif

///=====================================================================================================================
///                                  VCS simulation code
///
/// This code allows the TE to enable duty cycle offset injection and behavioral duty 
///  cycle adjustment.  To use this code the TE needs to pound the following controls:
///
///  1) Behavioral duty cycle model enable
///  2) Magnitude of initial duty cycle offset in VCS ticks (or ps if you prefer)
///  3) Direction of initial duty cycle offset
///
/// Note that initial offset mangnitude must be less than one ideal phase of the input 
///  clock.
/// An offset direction of 1'b1 corresponds to a postive DCO, or elongated high phase.
/// An offset direction of 1'b0 corresponds to a negative DCO, or elongated low phase.
///
///=====================================================================================================================


`ifndef ip2211ringpll_NO_VCSSIM

///=================================================================================
/// Duty Cycle Offset Injection
///
///   Assumes incoming clock is 50% duty cycle and injects programmable 
///   duty cycle distortion of offset that can be corrected by the DCC loop.
///=================================================================================

   bit  [7:0]  dco_magnitude;       // TE must pound a non-zero value
   bit         dco_direction;       // TE must pound either 1'b0 or 1'b1
   bit         clkin_delay; 
   logic        clkin_dca;

   initial begin

      dco_magnitude = '0;           // 0 = no DCO , >0 = DCO in VCS ticks
      dco_direction = '0;           // 0 = negative DCO, 1 = postitive DCO

   end//initial


   // Generate a delayed version of clkin used to inject a duty cycle offset.
   // Note that this is a blocking assignment because clocks should evaluate
   //  in the blocking queue. The delay magnitude should never be equal to
   //  or greater than one phase of clkin; that will not evaluate correctly.
   //
   always @(clkin)
      clkin_delay = #dco_magnitude clkin;


   // If the DCO magnitude is set to 0, pass clkin directly to clkout
   // To add positive DCO (elongated high phase), OR clkin with clkin_delay
   // To add negative DCO (elongated low phase), AND clkin with clkin_delay
   // 
   assign clkin_dca = (dco_magnitude == 0)? clkin : 
                     ((dco_direction)? (clkin | clkin_delay) : (clkin & clkin_delay));
   
   

///=================================================================================
/// Duty Cycle Adjustment
///
///   Behavioral modeling of DCA functionality. Converts the incoming
///   "ctrl" code into a programmable amount of duty cycle adjustment.
///=================================================================================

   bit         en_dca_model;        // TE must pound to 1'b1
   logic [2:0]  dca_step_size;       // TE can adjust the adjustement step in VCS ticks
   logic [5:0]  step_magnitude;
   logic [8:0]  delay_amount;
   bit         clkdly_dca;
   logic        clkout_dca;

   initial begin

      en_dca_model  = 1'b0;         // 0 = no behavioral adjustment modeling; 1 = yes
      dca_step_size = 3'd3;         // duty cycle adjust step size in VCS ticks

   end//initial


   // Determine the magnitude of the duty cycle adjustment by finding the
   //  difference from the mid-point setting of 0x20 (decimal 32). If the
   //  MSB of the DCA code is '1, adjustments are in the positive DCO
   //  direction and the LSBs indicate the true magnitude. If the MSB is
   //  '0, adjustments are in the negative direction and we need to
   //  subtract the LSB value from the unsigned midpoint of 0x4.
   //  the LSBs.
   //  
   always_comb step_magnitude = (ctrl[5]) ? {1'b0,ctrl[4:0]} : (9'd32 - {1'b0,ctrl[4:0]});


   // Multiply the magnitude by the step size to get the required
   //  adjustment in VCS ticks. Quality the delay with the behavioral
   //  modeling enable to avoid undesired delay events in simulation.
   //
   always_comb delay_amount = (en_dca_model)? (step_magnitude * dca_step_size) : '0;


   // Generate a delayed version of clkin_dca used to adjust the duty cycle.
   // Note that this is a blocking assignment because clocks should evaluate
   //  in the blocking queue. The delay magnitude should never be equal to
   //  or greater than one phase of clkin; that will not evaluate correctly.
   //
   always @(clkin_dca)
      clkdly_dca = #delay_amount clkin_dca;


   // Skew the outbound clock based on the calculated duty cycle offset
   //  magnitude and direction. For postitive adjustments (MSB=1), OR the
   //  incoming and delayed clocks to elongate the high phase. For negative
   //  adjustments (MSB=0), AND the incoming and delayed clocks to shorten
   //  the high phase.
   //
   always_comb clkout_dca = (ctrl[5]) ? (clkin_dca | clkdly_dca) : (clkin_dca & clkdly_dca);


   //  Modelling output as a function of vccxx "primary" domain of this AIP
   //  This should realistically inject an X on clkout in non-MPP DUTs
   //
   always_comb clkout = (vccxx)? ((en_dca_model)? clkout_dca : clkin_dca) : 1'bX;



///=================================================================================
/// Duty Cycle Monitoring
///
///   Monitors the high and low phase time percentages of the DCA output 
///   clock in order to facilitate testing in a closed loop system.
///=================================================================================

   bit      clkout_inst;
   integer  rise_time, fall_time, hi_phase, lo_phase, HI_TIME_PERCENT, LO_TIME_PERCENT;


   // Generate a gated clock so this logic does not evaluate when the
   // behavioral model is not being used
   //
   `ip2211ringpll_CLKAND(clkout_inst, clkout_dca, en_dca_model)


   // Sample the simulation time at the rising and falling edges of the
   //  output clock
   //
   always @(posedge(clkout_inst)) rise_time <= $realtime;
   always @(negedge(clkout_inst)) fall_time <= $realtime;


   // Compute delta simlation time for high and low phases of the clock
   //
   `ip2211ringpll_ASYNC_RSTD_MSFF  (hi_phase, (fall_time-rise_time), clkout_inst, ~en_dca_model, 1)
   `ip2211ringpll_ASYNC_RSTD_MSFF  (lo_phase, (rise_time-fall_time), ~clkout_inst, ~en_dca_model, 1)


   // Calculate the high and low time percentages
   //
   always_comb HI_TIME_PERCENT = (hi_phase*100)/(hi_phase+lo_phase);
   always_comb LO_TIME_PERCENT = (lo_phase*100)/(hi_phase+lo_phase);



`endif

   logic [1:0]    cb_nc;
   logic [5:0]    ctrl_nc;

   // Dummy assignments so MPP can see receivers in this hierarchy
   //
   always_comb cb_nc   = cb;
   always_comb ctrl_nc = ctrl;

///=====================================================================================================================
/// Black Box Assertions
///=====================================================================================================================

`ifndef ip2211ringpll_NO_VCSSIM 
`ifndef ip2211ringpll_SVA_OFF
   // Check for 1'b1 on vccxx when this BB outputs are ready to be consumed downstream
   //  NOTE: Disabling the assertions when in modes other than REGULATION and JITTER
   //
   `ip2211ringpll_ASSERTC_MUST(R_cpadcaana_vccxx_1, vccxx == 1'b1, sva_reset,
   `ip2211ringpll_ERR_MSG("ERROR, vccxx in ip2211ringpll_cpadcaana is not '1 !!"));

   // Check for inputs that are X when  this BB outputs are ready to be consumed downstream
   //  NOTE: Disabling the assertions when in modes other than REGULATION and JITTER
   //
   `ip2211ringpll_ASSERTC_KNOWN_DRIVEN(R_cpadcaana_X_inputs, {cb,clkin,ctrl,vccxx}, sva_reset,
   `ip2211ringpll_ERR_MSG("ERROR, Some inputs to ip2211ringpll_cpadcaana are unknown!"));

`endif //  `ifndef ip2211ringpll_SVA_OFF 
`endif //  `ifdef VCSSIM 



///=====================================================================================================================
/// Trailer Files
///=====================================================================================================================
`endif

endmodule // ip2211ringpll_cpadcaana

`endif //  `ifndef ip2211ringpll_cpadcaana_SV

`ifndef ip2211ringpll_PLLDCA_SV
`define ip2211ringpll_PLLDCA_SV

//`include "cpadcaana.sv"

module ip2211ringpll_plldca(

          
         `ifndef ip2211ringpll_NO_VCSSIM
	`ifdef INTC_SIM
// @ hip/dca level  reset_b_xxl was not present 
        input   logic         reset_b_xxl,
 	`endif
         `endif
         input   logic [5:0]   dca_ctrl,
         input   logic [1:0]   dca_cb,
         //input   logic         trunk_mux__ClkPllMH,
         input   logic         pll_core_clkm,

         output  logic         clkpllmh
);

   logic reset_b_xxl ;
   // DCA AIP
   //
   ip2211ringpll_cpadcaana dca_ana (
         `ifndef ip2211ringpll_NO_VCSSIM 
            .sva_reset   ( ~reset_b_xxl        ),
         `endif
            .vccxx       ( 1'b1                ),
            .ctrl        ( dca_ctrl            ),
            .cb          ( dca_cb              ),
            //.clkin       ( trunk_mux__ClkPllMH ),
            .clkin       ( pll_core_clkm ),

            .clkout      ( clkpllmh            )
   );

endmodule

`endif

`ifndef ip2211ringpll_VIEW_MUX_SV
`define ip2211ringpll_VIEW_MUX_SV

//`include "ringpll_macros.sv"
//`include "soc_clock_macros.sv"

module ip2211ringpll_view_mux (
   `ifdef ip2211ringpll_LJPLL_NO_UPF_SUPPORT
      input wire   vccpll,
   `endif
   
   input  logic                                       pll_core__clk_pll_div1,
   input  logic                                       ClkPostDistMH,
   input  logic                                       clkref_prediv,
   input  logic                                       VctlRdacEnNL,
   input  logic                                       ClkRefXXH,
   input  logic                                       ClkFbMXH,
   input  logic                                       Reset_b_XXL,
   input  logic                                       pfdennh,
   input  logic                                       pll_fbgen__tight_loop,
   input  logic                                       powergood,
   input  logic [1:0]                                 ViewDigEnNH,
   input  logic [4:0]                                 viewsel0,
   input  logic [4:0]                                 viewsel1,
   input  logic                                       RawLockXXL,
   input  logic                                       LockXXL,
   input  logic                                       EarlyLockXXH,
   input  logic                                       ssc_reload,
   input  logic                                       mod_clk_to_view,

   // View Signals
   //
//   input  logic                                       clk_sync,
//   input  logic                                       stm_ifdim__StmStopMnnnH,
//   input  logic                                       odcs_dll__OdcsDllAddDelayMnnnL ,
//   input  logic                                       odcs_dll__OdcsDllPhDetEarlyMnnnH ,
//   input  logic                                       odcs_dll__OdcsDllPhDetLateMnnnH ,
//   input  logic                                       odcs_dll__OdcsDllUpdateMnnnL ,
//   input  logic                                       odcs_dig__OdcsRiseBase0MnnnH ,
//   input  logic                                       odcs_dig__OdcsFallBase0MnnnH ,
//   input  logic                                       odcs_dig__OdcsRiseVal1MnnnH ,
//   input  logic                                       odcs_dig__OdcsFallVal1MnnnH ,
//   input  logic                                       vctl_pullupnh,
//   input  logic                                       vctl_pulldnnh,
//   input  logic                                       pll_core__cp1clk,
//   input  logic                                       pll_core__cp1aclk,
//   input  logic                                       pll_core__cp2clk,
//   input  logic                                       pll_core__cp2aclk,
//   input  logic                                       trunk_mux__ClkRoRH,
//   input  logic                                       cmpenxxh,

   output logic [1:0]                                 view_mux__ViewOutNnnnH
);

///========================================================================================================
/// Module Begin
///========================================================================================================
   
   ///==========================================================
   /// PLL pre- and post-distribution clock division
   ///==========================================================

      logic        GatedClkEnNnnnH;

      logic        ClkPreGatedMH, ClkPostGatedMH;
      logic        ClkRoGatedRH;
      logic  ClkPreDivMH_0 ; 
	logic ClkPostDivMH_0 ;
	logic  ClkPreDivMH_1 ;
	logic ClkPostDivMH_1 ;
logic [1:0] ClkPreDivMH , ClkPostDivMH ;
      logic        ClkModToViewDXH;
      logic        ClkPreDivMH_nf, ClkPostDivMH_nf;
      logic        ClkPreDivMH_f,  ClkPostDivMH_f;

      always_comb GatedClkEnNnnnH = (|ViewDigEnNH);

      // Gate the pre- and post-dist clocks with the enable. Note that the
      //  enable can be considered static and used without synchronization to
      //  the clock source.
      //
      `ip2211ringpll_CLKAND(ClkPostGatedMH, ClkPostDistMH,          GatedClkEnNnnnH)
      `ip2211ringpll_CLKAND(ClkPreGatedMH,  pll_core__clk_pll_div1, GatedClkEnNnnnH)

      // Gate the RO clock with the enable.
      //
      //`ip2211ringpll_CLKAND(ClkRoGatedRH,   trunk_mux__ClkRoRH,     GatedClkEnNnnnH)

      // Gate SSC DFX clock with the enable.
      //
      `ip2211ringpll_CLKAND(ClkModToViewDXH, mod_clk_to_view,       GatedClkEnNnnnH)

      // Use simple 2-bit counters to divide the clocks by 2 and 4. The
      //  timing alignment between pre- and post-dist is not important, nor is
      //  the initializtion of the counter states.
      //
      //  `ip2211ringpll_ASYNC_RST_MSFF(ClkPreDivMH,  (ClkPreDivMH  + 2'b1), ClkPreGatedMH,  ~GatedClkEnNnnnH)
      //  `ip2211ringpll_ASYNC_RST_MSFF(ClkPostDivMH, (ClkPostDivMH + 2'b1), ClkPostGatedMH, ~GatedClkEnNnnnH)
	

// to resolve view_mux issue/noneq  ,  clock and data pin assignment for flops  were different fro different bits  
logic ClkPreDivMH_0_b;
logic ClkPostDivMH_0_b; 
 
assign ClkPreDivMH_0_b = ~ ClkPreDivMH_0; 
assign ClkPostDivMH_0_b = ~ClkPostDivMH_0; 
       `ip2211ringpll_ASYNC_RST_MSFF(ClkPreDivMH_0,  ~(ClkPreDivMH_0 ), ClkPreGatedMH,  ~GatedClkEnNnnnH)
       `ip2211ringpll_ASYNC_RST_MSFF(ClkPreDivMH_1, ~ (ClkPreDivMH_1 ),  ClkPreDivMH_0_b ,  ~GatedClkEnNnnnH)

       `ip2211ringpll_ASYNC_RST_MSFF(ClkPostDivMH_0,~ (ClkPostDivMH_0 ), ClkPostGatedMH, ~GatedClkEnNnnnH)
       `ip2211ringpll_ASYNC_RST_MSFF(ClkPostDivMH_1,~ (ClkPostDivMH_1 ), ClkPostDivMH_0_b , ~GatedClkEnNnnnH)


      // Flopping to create signals one cycle apart
      //
      /* -> Redundant Logic : Not driven/driving any logic. This 2 bit reg was removed and replaced with T-FF based implementation ; see comment from  above
      assign ClkPreDivMH_nf  = ClkPreDivMH[1];
      assign ClkPostDivMH_nf = ClkPostDivMH[1];
      `ip2211ringpll_MSFF(ClkPreDivMH_f,  ClkPreDivMH[1],  ClkPreGatedMH)
      `ip2211ringpll_MSFF(ClkPostDivMH_f, ClkPostDivMH[1], ClkPostGatedMH)
      */  
   logic [1:0] ViewSigBusNnnnH;

   // TODO: need to figure out if it's possible to parameterize the view
   //       selects properly.  Perhaps through RDL?
   //
   ///==========================================================
   /// View mux signal decode
   ///==========================================================
   always_comb begin : VIEW_SIGNALS

      unique casez(viewsel0)
         5'h0  : ViewSigBusNnnnH[0] = 1'b0;
         5'h1  : ViewSigBusNnnnH[0] = 1'b1;
         5'h2  : ViewSigBusNnnnH[0] = ClkRefXXH;
         5'h3  : ViewSigBusNnnnH[0] = RawLockXXL;
         5'h4  : ViewSigBusNnnnH[0] = ClkFbMXH;
         5'h5  : ViewSigBusNnnnH[0] = LockXXL;
         5'h6  : ViewSigBusNnnnH[0] = pll_fbgen__tight_loop;
         5'h7  : ViewSigBusNnnnH[0] = Reset_b_XXL;
         5'h8  : ViewSigBusNnnnH[0] = pfdennh;
         5'h9  : ViewSigBusNnnnH[0] = ssc_reload;	
         5'hA  : ViewSigBusNnnnH[0] = powergood;
         5'hB  : ViewSigBusNnnnH[0] = EarlyLockXXH;
         5'hC  : ViewSigBusNnnnH[0] = VctlRdacEnNL;
         5'hD  : ViewSigBusNnnnH[0] = 1'b0;
         5'hE  : ViewSigBusNnnnH[0] = mod_clk_to_view;
         5'hF  : ViewSigBusNnnnH[0] = 1'b0;
         5'h10 : ViewSigBusNnnnH[0] = ClkPostGatedMH;
         5'h11 : ViewSigBusNnnnH[0] = 1'b0;
         5'h12 : ViewSigBusNnnnH[0] = ClkPreGatedMH;
         5'h13 : ViewSigBusNnnnH[0] = 1'b0;
         5'h14 : ViewSigBusNnnnH[0] =~ ClkPreDivMH_1; // plldiv4
         5'h15 : ViewSigBusNnnnH[0] = 1'b0;
         5'h16 : ViewSigBusNnnnH[0] = ~ ClkPreDivMH_0; // plldiv2
         5'h17 : ViewSigBusNnnnH[0] = 1'b0;
         5'h18 : ViewSigBusNnnnH[0] = ~ ClkPostDivMH_0; // postdiv2
         5'h19 : ViewSigBusNnnnH[0] = 1'b0;
         5'h1A : ViewSigBusNnnnH[0] =~ ClkPostDivMH_1; // postdiv4
         5'h1B : ViewSigBusNnnnH[0] = 1'b0;
         5'h1C : ViewSigBusNnnnH[0] = 1'b0;
         5'h1D : ViewSigBusNnnnH[0] = 1'b0;
         5'h1E : ViewSigBusNnnnH[0] = 1'b0;
         5'h1F : ViewSigBusNnnnH[0] = clkref_prediv;
         `ip2211ringpll_XDefault(ViewSigBusNnnnH[0])
      endcase
      
      unique casez(viewsel1)
         5'h0  : ViewSigBusNnnnH[1] = 1'b0;
         5'h1  : ViewSigBusNnnnH[1] = 1'b1;
         5'h2  : ViewSigBusNnnnH[1] = ClkRefXXH;
         5'h3  : ViewSigBusNnnnH[1] = RawLockXXL;
         5'h4  : ViewSigBusNnnnH[1] = ClkFbMXH;
         5'h5  : ViewSigBusNnnnH[1] = LockXXL;
         5'h6  : ViewSigBusNnnnH[1] = pll_fbgen__tight_loop;
         5'h7  : ViewSigBusNnnnH[1] = Reset_b_XXL;
         5'h8  : ViewSigBusNnnnH[1] = pfdennh;
         5'h9  : ViewSigBusNnnnH[1] = ssc_reload;	
         5'hA  : ViewSigBusNnnnH[1] = powergood;
         5'hB  : ViewSigBusNnnnH[1] = EarlyLockXXH;
         5'hC  : ViewSigBusNnnnH[1] = VctlRdacEnNL;
         5'hD  : ViewSigBusNnnnH[1] = 1'b0;
         5'hE  : ViewSigBusNnnnH[1] = mod_clk_to_view;
         5'hF  : ViewSigBusNnnnH[1] = 1'b0;
         5'h10 : ViewSigBusNnnnH[1] = ClkPostGatedMH;
         5'h11 : ViewSigBusNnnnH[1] = 1'b0;
         5'h12 : ViewSigBusNnnnH[1] = ClkPreGatedMH;
         5'h13 : ViewSigBusNnnnH[1] = 1'b0;
         5'h14 : ViewSigBusNnnnH[1] = ~ClkPreDivMH_1; // plldiv4
         5'h15 : ViewSigBusNnnnH[1] = 1'b0;
         5'h16 : ViewSigBusNnnnH[1] =~ ClkPreDivMH_0; // plldiv2
         5'h17 : ViewSigBusNnnnH[1] = 1'b0;
         5'h18 : ViewSigBusNnnnH[1] =~ ClkPostDivMH_0; // postdiv2
         5'h19 : ViewSigBusNnnnH[1] = 1'b0;
         5'h1A : ViewSigBusNnnnH[1] =~ ClkPostDivMH_1; // postdiv4
         5'h1B : ViewSigBusNnnnH[1] = 1'b0;
         5'h1C : ViewSigBusNnnnH[1] = 1'b0;
         5'h1D : ViewSigBusNnnnH[1] = 1'b0;
         5'h1E : ViewSigBusNnnnH[1] = 1'b0;
         5'h1F : ViewSigBusNnnnH[1] = clkref_prediv;
         `ip2211ringpll_XDefault(ViewSigBusNnnnH[1])
      endcase

   end : VIEW_SIGNALS


   ///==========================================================
   /// View Mux select internal/external signal
   ///==========================================================
   logic [1:0] ViewOutNnnnH;

   always_comb begin : VIEW_MUX
  
      unique casez (ViewDigEnNH)
         2'b00   : ViewOutNnnnH = 2'b00;
         2'b01   : ViewOutNnnnH = {1'b0,ViewSigBusNnnnH[0]};
         2'b10   : ViewOutNnnnH = {ViewSigBusNnnnH[1],1'b0};
         2'b11   : ViewOutNnnnH = ViewSigBusNnnnH;
         `ip2211ringpll_XDefault(ViewOutNnnnH)
      endcase
   
   end : VIEW_MUX

   assign view_mux__ViewOutNnnnH = ViewOutNnnnH;

endmodule

`endif


`ifndef ip2211ringpll_TSADCSDMOD10ANA_SV
`define ip2211ringpll_TSADCSDMOD10ANA_SV 

//`include "soc_macros.sv"     // Project generic macros.
`ifndef ip2211ringpll_SVA_OFF
//`include "intel_checkers.sv"
//`include "ringpll_macros.sv"
`endif

module ip2211ringpll_tsadcsdmod10ana (
`ifndef ip2211ringpll_LJPLL_ADC_MSV
`ifndef ip2211ringpll_SVA_OFF
input logic     ADCen_inst,
`endif
`endif

//Reference Voltage selects
input logic     selvsense_b,
input logic     selvccthm_b,
input logic     selvccio_b,
//Reference voltage selects
`ifndef INTEL_EMULATION
input tri      vref_a,
`else 
input logic     vref_a,
`endif
input logic     vccthmxx,
input logic     vccioxx,
//ADC inputs
`ifdef INTEL_EMULATION
input logic    vangin_a,
`else
input tri      vangin_a,
`endif
//Clocks
input logic     ckph1,
input logic     ckph2,
output logic    ckph1dfb,
output logic    ckph2dfb,
//Other inputs
input logic     en_b,         //Turns off current source in the circuit (Disables circuit)
input logic     fdbkin,       //Digital Feedback loop input
input logic     adj,          //PRBS noise source
input logic     chop,         //ADC ChopEn TapCfg bit
output logic    sdout
);

`ifndef ip2211ringpll_NO_VCSSIM
   logic       ckfben;
   logic       ckinpen;

  `ifndef ip2211ringpll_NO_VCSSIM
   logic [9:0] Vref_inst;   //This is the inst declaration for the reference voltage (VCCIO,VCCTHM or external vref)
   logic [9:0] VGnd_inst;   //This is the inst declaration for the SDinNeg value
   logic [9:0] VinPos_inst; //This is the inst declaration for SDinPos value
   logic [9:0] VinNeg_inst; //This is the inst declaration for the actual VNeg. It could either be 0 or SDinNeg
   logic       sdouteval;

   real SDFeedback;        //SigmaDelta Feedback value
   real SDIntegrateOutL;   //SigmaDelta Integrated value
   real SDIntegrateInL;    //SigmaDelta Evaluated but Pre-Integrated value
   real SDInputNormalized; //Normalized SDInput value

//TE can pound these logics to simulate the usage in different voltage values
(* vcs_ignore_drive *)
initial begin
 Vref_inst = 10'h3ff;
 VinPos_inst = 10'h0ff;
 VGnd_inst = 10'h00f;
 SDIntegrateInL = 0; 
end

//Modelling chopped non-overlap clocks (moved inside AIP for BDW)
assign ckinpen =  chop ? ckph2 : ckph1;
assign ckfben  = chop ? ckph1 : ckph2;

//Vin Negative is the remote ground value in differential mode, else it's 0
//BDW: Diff mode removed
assign VinNeg_inst = 10'h0 ; 

//Final Normalized SD input
assign SDInputNormalized = (VinPos_inst - VinNeg_inst)/(1.0 * Vref_inst);

//SD feedback
assign SDFeedback = chop ? (fdbkin - SDInputNormalized) : (SDInputNormalized - fdbkin);

//ADC is evaluated in Phase 2 ADC clk 
`ip2211ringpll_MSFF(SDIntegrateInL, SDIntegrateOutL, ckph2)
assign SDIntegrateOutL = SDIntegrateInL + SDFeedback;

//1-bit quantizer
assign sdouteval = (SDIntegrateOutL > 0);

//Output of SigmaDelta ADC
assign sdout = ( (!vccioxx & !selvccio_b) | (!vccthmxx & !selvccthm_b) | (!vref_a & !selvsense_b) ) ? 1'bx : (~en_b ? sdouteval : 1'b1);  

`endif //ip2211ringpll_NO_VCSSIM



//=====================================================================================================================
//Output feedback clock (to generate non-overlapping clocks)
//=====================================================================================================================
assign ckph1dfb = ckph1;
assign ckph2dfb = ckph2;


`endif   //ip2211ringpll_NO_VCSSIM



endmodule 
`endif

`ifndef ip2211ringpll_TSADCSDMOD10TOP_SV
`define ip2211ringpll_TSADCSDMOD10TOP_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "tsadcsdmod10ana.sv"
//`include "ringpll_macros.sv"
`ifndef ip2211ringpll_SVA_OFF
//`include "intel_checkers.sv"
`endif
module ip2211ringpll_tsadcsdmod10top (
//   input    logic         VCCIOxx,  		// Removed to match SCH -
//   input    logic         ADCEnDizzX1nnnH_b,  // Removed to match SCH -
//   input    logic         ADCContModeX1nnnH,  // Removed to match SCH -
//   input    logic  [1:0]  SDVrefSelX1nnnH,	// Removed to match SCH -
//   input    logic         BGTrimMode,		// Removed to match SCH -
   input    logic         VCCxx,
   input    logic         ClkInXH,
   input    logic         ADCEnX1nnnH,
   input    logic         ADCRstX1nnnH_b,
   input    logic         ADCFreezeX1nnnH,
   input    logic         ADCChopEnX1nnnH,
   input    logic  [1:0]  ADCClkDivX1nnnH,
`ifdef INTEL_EMULATION
   input    logic         SDinPos_a, 
   input    logic         Vref_a,
`else 
   input    tri           SDinPos_a, 
   input    tri           Vref_a,
`endif
   output   logic         ADCDoneX1nnnH,  
   output   logic  [9:0]  ADCDigOutX1nnnH,
   output   logic         CkDigOutValU2N00 
);

//logic declarations
logic [1:0] ADCClkDivX1nnnH_DC;

// Tied to a specific value as these signals are not used in SCH. -
logic  [1:0]  SDVrefSelX1nnnH;	// Removed to match SCH -
assign SDVrefSelX1nnnH = 2'b01; // Tied to => 2b’01 (choose VREF_A as a reference) -
logic         BGTrimMode;		// Removed to match SCH -
assign BGTrimMode = 1'b0;		
logic         ADCEnDizzX1nnnH_b;  // Removed to match SCH -
assign ADCEnDizzX1nnnH_b = 1'b1;
logic         ADCContModeX1nnnH;
assign ADCContModeX1nnnH = 1'b1;


//ADC Clock logics
logic Clk25MhzX1H, Clk50MhzX1H, Clk12p5MhzX1H, Clk6p25MhzX1H; //Divided input clock
logic ClkDivOutAngX1H;  //Selected Divided clock
logic ClkSigmaDeltaX1H; //Divided clock gated with ADCFreeze
logic ClkADCCounterX1H;    //Counter divided clock, will be gated after 1024 cycles if not in Continuous mode
logic ADCCountClkEnX1nnnL; //ADC counter clk enable

//Selects for voltage reference to sigma delta 
logic SelVSenseX1nnnH, SelVccioX1nnnH, SelVccthmX1nnnH;  

//Sigma Delta ADC output and flopped version
logic SDModOut_AngX1nnnH, SDModOutX1nnnH;   
logic SDModOut_Ang_ModX1nnnH;   

//Flop repeated signals
logic  ADCEnSyncX1nnnH, ADCChopEnX1nnnH_mcp;
logic  FreezeSyncX1nnnH_b, FreezeSyncLatOutX1nnnL_b;

//counter related logics
logic PrimCntr_WrapX1nnnH;
logic [9:0] Prim_CountX1nnnH;
logic [9:0] Next_Sec_CountX1nnnH, Sec_CountX1nnnH;

//ADC Done Bit, non flopped version
logic         ADCDoneX1nn0H;

//ADC Data ip2211ringpll_MSFF Output
logic [9:0]   ADCDigOutX1nnnH_b;

//Non-overlap clocks to be sent to AIP
logic         ClkSDinX1H;
logic         ClkSDinX1L;

//Delayed clock from AIP
logic         ClkSDinX1H_d, ClkSDinX1L_d;

// PRBS related Signals
logic         PrbsXnn0H, PrbsXnn1H, PrbsXnn2H, PrbsXnn3H, PrbsXnn4H, PrbsXnn5H, PrbsXnn6H, RstLFSRXnnnH_b;

/////////////////////////////////////////////////////////////////////////////
//ADC DFT clock divider

//`ASYNC_RST_MSFF_CLK(Clk50MhzX1H,   ~Clk50MhzX1H,   ClkInXH,       ~ADCRstX1nnnH_b)   
//`ASYNC_RST_MSFF_CLK(Clk25MhzX1H,   ~Clk25MhzX1H,   Clk50MhzX1H,   ~ADCRstX1nnnH_b)
//`ASYNC_RST_MSFF_CLK(Clk12p5MhzX1H, ~Clk12p5MhzX1H, Clk25MhzX1H,   ~ADCRstX1nnnH_b)
//`ASYNC_RST_MSFF_CLK(Clk6p25MhzX1H, ~Clk6p25MhzX1H, Clk12p5MhzX1H, ~ADCRstX1nnnH_b)
   logic ClkDiv2XXH;
   logic ClkDiv2NbXXH;
   logic ClkDiv4XXH;
   logic ClkDiv4NbXXH;
   logic ClkDiv8XXH;
   logic ClkDiv8NbXXH;
   logic ClkDiv16XXH;
   logic ClkDiv16NbXXH;

   `ip2211ringpll_NB_ASSIGN(ClkDiv2NbXXH, ClkDiv2XXH)
   `ip2211ringpll_MAKE_CLK_DIV2_RESET(ClkDiv2XXH,  ~ClkDiv2NbXXH,  ClkInXH,    ADCRstX1nnnH_b)
   `ip2211ringpll_NB_ASSIGN(ClkDiv4NbXXH, ClkDiv4XXH)
   `ip2211ringpll_MAKE_CLK_DIV2_RESET(ClkDiv4XXH,  ~ClkDiv4NbXXH,  ClkDiv2XXH, ADCRstX1nnnH_b)
   `ip2211ringpll_NB_ASSIGN(ClkDiv8NbXXH, ClkDiv8XXH)
   `ip2211ringpll_MAKE_CLK_DIV2_RESET(ClkDiv8XXH,  ~ClkDiv8NbXXH,  ClkDiv4XXH, ADCRstX1nnnH_b)
   `ip2211ringpll_NB_ASSIGN(ClkDiv16NbXXH, ClkDiv16XXH)
   `ip2211ringpll_MAKE_CLK_DIV2_RESET(ClkDiv16XXH, ~ClkDiv16NbXXH, ClkDiv8XXH, ADCRstX1nnnH_b)

   assign Clk50MhzX1H  = ClkDiv2XXH;
   assign Clk25MhzX1H  = ClkDiv4XXH;
   assign Clk12p5MhzX1H = ClkDiv8XXH;
   assign Clk6p25MhzX1H = ClkDiv16XXH;

//In DTS we sync to local clock, in some other places its not sync'd to local clock.
//Also the clock divider override in BE creates funky pessimistic hold checks.
//`CUTDC(ADCClkDivX1nnnH_DC, ADCClkDivX1nnnH, ~ADCEnX1nnnH)
assign ADCClkDivX1nnnH_DC = ADCClkDivX1nnnH;

always_comb begin: ADCClk_div
     unique casez (ADCClkDivX1nnnH_DC)
         2'b00   : ClkDivOutAngX1H = Clk25MhzX1H;
         2'b01   : ClkDivOutAngX1H = Clk12p5MhzX1H;
         2'b10   : ClkDivOutAngX1H = Clk50MhzX1H;
         2'b11   : ClkDivOutAngX1H = Clk6p25MhzX1H;
         `ip2211ringpll_XDefault(ClkDivOutAngX1H)
     endcase
end


//Sending the non-overlap clocks to ADC blackbox
//Feedback causes HW loop in emulation
//`ifndef INTC_EMULATION  
`ifndef ip2211ringpll_NO_VCSSIM 
assign ClkSDinX1H =   ClkDivOutAngX1H & ~ClkSDinX1L_d;
assign ClkSDinX1L =  ~ClkDivOutAngX1H & ~ClkSDinX1H_d;
`else
assign ClkSDinX1H =   ClkDivOutAngX1H;
assign ClkSDinX1L =  ~ClkDivOutAngX1H;
`endif

//Flops replaced with Meta which will be used by the Counters as reset 
//`METAFLOP_2(ADCEnSyncX1nnnH, ADCEnX1nnnH, ClkSDinX1H)
logic AdcEnX1nn1H;
`ip2211ringpll_MSFF(AdcEnX1nn1H, ADCEnX1nnnH, ClkSDinX1H)
`ip2211ringpll_MSFF(ADCEnSyncX1nnnH, AdcEnX1nn1H, ClkSDinX1H)


////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//Sigma Delta Analog Block 

//Decoder to obtain the Vref to be used for Sigma Delta Analog block
assign SelVccthmX1nnnH  = (SDVrefSelX1nnnH == 2'b00) ;
assign SelVccioX1nnnH   = (SDVrefSelX1nnnH == 2'b01) ;
assign SelVSenseX1nnnH  = (SDVrefSelX1nnnH == 2'b10) ;

// PRBS for HW Dithering: Reset only is we are stuck at 0000001, otherwise we are fine.
assign RstLFSRXnnnH_b = ~PrbsXnn0H | PrbsXnn1H | PrbsXnn2H | PrbsXnn3H | PrbsXnn4H | PrbsXnn5H | PrbsXnn6H;

// LFSR chain
`ip2211ringpll_ASYNC_RST_MSFF(PrbsXnn0H, ~(PrbsXnn5H ^ PrbsXnn6H), ClkSDinX1H, (ADCEnDizzX1nnnH_b | ~RstLFSRXnnnH_b))
`ip2211ringpll_MSFF(PrbsXnn1H, ~PrbsXnn0H, ClkSDinX1H)
`ip2211ringpll_MSFF(PrbsXnn2H,  PrbsXnn1H, ClkSDinX1H)
`ip2211ringpll_MSFF(PrbsXnn3H,  PrbsXnn2H, ClkSDinX1H)
`ip2211ringpll_MSFF(PrbsXnn4H,  PrbsXnn3H, ClkSDinX1H)
`ip2211ringpll_MSFF(PrbsXnn5H,  PrbsXnn4H, ClkSDinX1H)
`ip2211ringpll_MSFF(PrbsXnn6H,  PrbsXnn5H, ClkSDinX1H)

// You reset only when stuck at 0000001. Even if it inadvertently resets becuase of
// a glitch its not a fatal/functional problem, as its on dither generation block.
//`ip2211ringpll_ASSERTS_GRAY_CODE(GLITCH_PrbsRst, {PrbsXnn0H, `GWAIVE(PrbsXnn1H), `GWAIVE(PrbsXnn2H), `GWAIVE(PrbsXnn3H), `GWAIVE(PrbsXnn4H), `GWAIVE(PrbsXnn5H), `GWAIVE(PrbsXnn6H), ADCEnDizzX1nnnH_b}, ClkSDinX1H, 1'b0,`ip2211ringpll_ERR_MSG("PrbsRst glitch detected."));

//The ADCChopEnX1nnnH is from tap/fuse endpoint. Even if it cause X to be captured in 
//SDModOutX1nnnH flop, it'll get resolved the next cycle. That X is harmless (possible
//bad ADC value the first time its enabled. If its written before ADCen & ADCRst then
//we don't run into that risk either.
//`CUTMCP_HP1(ADCChopEnX1nnnH_mcp, ADCChopEnX1nnnH, 1'b0, ClkInXH, ClkInXH, 3, '0, '1)
assign ADCChopEnX1nnnH_mcp = ADCChopEnX1nnnH;

ip2211ringpll_tsadcsdmod10ana ip2211ringpll_tsadcsdmod10ana (
//Inputs
   .en_b                   (~ADCRstX1nnnH_b),
   .fdbkin                 (SDModOutX1nnnH),
   .vangin_a               (SDinPos_a),
   .selvsense_b            (~SelVSenseX1nnnH),
   .selvccthm_b            (~SelVccthmX1nnnH),
   .selvccio_b             (~SelVccioX1nnnH),
   .ckph1                  (ClkSDinX1H),
   .ckph2                  (ClkSDinX1L),
   .ckph1dfb               (ClkSDinX1H_d),
   .ckph2dfb               (ClkSDinX1L_d),

   //.vccioxx                (VCCIOxx),
   .vccioxx                (1'b1),

   .vccthmxx               (VCCxx),
   .vref_a                 (Vref_a),
   .adj                    (PrbsXnn0H),
   .chop                   (ADCChopEnX1nnnH_mcp),
`ifndef ip2211ringpll_LJPLL_ADC_MSV
`ifndef ip2211ringpll_SVA_OFF
   .ADCen_inst             (ADCEnX1nnnH),
`endif
`endif
//Outputs
   .sdout                  (SDModOut_AngX1nnnH)
);

//Output of Sigma Delta Converter is flopped once before it's sent to the
//secondary counter to sample the number of 1s in the bitstream
//
// if chop=1, then flip SDMod bit
//
assign SDModOut_Ang_ModX1nnnH = ADCChopEnX1nnnH_mcp ? ~SDModOut_AngX1nnnH : SDModOut_AngX1nnnH;
`ip2211ringpll_MSFF(SDModOutX1nnnH, SDModOut_Ang_ModX1nnnH, ClkSDinX1H)

 //Freeze Logic for DFT
 //In continuous mode, the ADC clock will only be gated if freeze config bit is asserted. 
//`METAFLOP_2(FreezeSyncX1nnnH_b,       ~ADCFreezeX1nnnH,     ClkSDinX1H)
logic AdcFreezeX1nn1H_b;
`ip2211ringpll_MSFF(AdcFreezeX1nn1H_b, ~ADCFreezeX1nnnH,     ClkSDinX1H)
`ip2211ringpll_MSFF(FreezeSyncX1nnnH_b, AdcFreezeX1nn1H_b,   ClkSDinX1H)
`ip2211ringpll_LATCH_P(FreezeSyncLatOutX1nnnL_b,    FreezeSyncX1nnnH_b,   ClkSDinX1H)

assign ClkSigmaDeltaX1H = FreezeSyncLatOutX1nnnL_b & ClkSDinX1H;

//Gate the clocks to the counters
//Counters Clock will be gated after 1024 cycles ClkSDinX1H if we are
//in non-continuous mode. In continuous mode, the ADC clock will only be
//gated if freeze config bit is asserted. 
`ip2211ringpll_LATCH_P(ADCCountClkEnX1nnnL , ADCContModeX1nnnH | ~ADCDoneX1nn0H, ClkSigmaDeltaX1H)
`ip2211ringpll_CLKAND(ClkADCCounterX1H, ClkSigmaDeltaX1H, ADCCountClkEnX1nnnL)

/////////////////////////////////////////////////////////////////////////////////////////////////////
//Primary Counter to generate 1024 sync
/////////////////////////////////////////////////////////////////////////////////////////////////////
`ip2211ringpll_RST_MSFF(Prim_CountX1nnnH, Prim_CountX1nnnH + 10'd1, ClkADCCounterX1H, ~ADCEnSyncX1nnnH )

assign PrimCntr_WrapX1nnnH = BGTrimMode ? (Prim_CountX1nnnH[5:0] == 6'b111111) :
                                          (Prim_CountX1nnnH == 10'b1111111111) ;

//Secondary Counter to calculate number of 1s in the 1024 bitstream
always_comb begin : Secondary_Counter
      unique casez ({BGTrimMode,SDModOutX1nnnH, PrimCntr_WrapX1nnnH})
        3'b?00   : Next_Sec_CountX1nnnH = Sec_CountX1nnnH;
        3'b?01   : Next_Sec_CountX1nnnH = {9'd0, 1'b0};    //New cycle with output of 0 from ADC
        3'b?10   : Next_Sec_CountX1nnnH = Sec_CountX1nnnH + 10'd1;
        3'b011   : Next_Sec_CountX1nnnH = {9'd0, 1'b0};    //New cycle with output of 1 from ADC (rst to 0 to prevent wrap around)
	3'b111   : Next_Sec_CountX1nnnH = {9'd0, 1'b1};    //New cycle with output of 1 from ADC (preset to 1 for BGTrim Mode)
        `ip2211ringpll_XDefault(Next_Sec_CountX1nnnH)
      endcase
end
`ip2211ringpll_RST_MSFF(Sec_CountX1nnnH, Next_Sec_CountX1nnnH, ClkADCCounterX1H, ~ADCEnSyncX1nnnH)

//In non continuous mode, final counter values will stay stuck and will be
//sent to the Tap statu shadow register for update.
//In continuous mode, final counter values will be updated every 1024 cycles. 
//Together with the ADC done valid bit, the tap status shadow register will be updated
assign CkDigOutValU2N00 = (~ClkSigmaDeltaX1H & PrimCntr_WrapX1nnnH & FreezeSyncX1nnnH_b);
`ip2211ringpll_ASYNC_SET_MSFF(ADCDigOutX1nnnH_b, ~Sec_CountX1nnnH, CkDigOutValU2N00, ~ADCEnX1nnnH)
assign ADCDigOutX1nnnH = ~ADCDigOutX1nnnH_b;

//HoldMCP for the above flop on ADCEnX1nnnH (as it bypasses the Metaflop)
//When ADCEN transitions first time, the clock doesn't toggle. When the clock starts to toggle, we know ADCEN wont toggle.
//`HOLDMCP2(ADCEnX1nnnH, 1'b1, CkDigOutValU2N00, ClkInXH, 2, ~ADCRstX1nnnH_b, holdmcp_adcen)

//ADC done valid bit after 1024 cycles of sampling. 
//In non-continuous mode, this will stay stuck on after 1024 cycles.
//In continuous mode, this will turn on every 1024 cycles to update the
//status register shadow registers with the new values.
assign ADCDoneX1nn0H   = PrimCntr_WrapX1nnnH & ADCEnSyncX1nnnH;
`ip2211ringpll_MSFF(ADCDoneX1nnnH, ADCDoneX1nn0H, ClkSigmaDeltaX1H)

//===================================================================
//Assertions
//===================================================================

`ifndef ip2211ringpll_SVA_OFF
`ip2211ringpll_ASSERTC_FORBIDDEN(ADC_VrefSel_Forbids, SDVrefSelX1nnnH == 2'b11, 1'b0, `ip2211ringpll_ERR_MSG("Reference voltage selections cannot be 11"));
`endif

endmodule
`endif



`ifndef ip2211ringpll_pllljviewadc_VS
`define ip2211ringpll_pllljviewadc_VS

//`include "soc_macros.sv"
//`include "tsadcsdmod10top.sv"

module ip2211ringpll_pllljviewadc (
   
         `ifndef ip2211ringpll_INTC_NO_PWR_PINS
            input wire   vccpll,
         `endif
            input logic   vccref,

         input  logic       ClkRefXXH,
         input  logic       adc_Reset_bXXL,
         input  logic       adc_StartXXH,
         input  logic [1:0] adc_clkdiv,
         input  logic       adc_freeze,
         input  logic       adc_chop_en,
         // input  logic       adc_use_vref,
         input  logic       pll_core__adc_in,

         output logic  [9:0] adc_dig_out,
         output logic        adc_done  

);


///========================================================================================================
/// Main Procedure
///========================================================================================================

ip2211ringpll_tsadcsdmod10top hvmadc  (
   `ifndef ip2211ringpll_INTC_NO_PWR_PINS
//      .VCCIOxx          ( vccpll               ),
      .VCCxx            ( vccpll               ),
      .Vref_a           ( vccref               ),
   `else
//      .VCCIOxx          ( 1'b1                 ),
      .VCCxx            ( 1'b1                 ),
      .Vref_a           ( 1'b1                 ),
   `endif
   
   .ClkInXH             ( ClkRefXXH            ),
   .ADCEnX1nnnH         ( adc_StartXXH         ),
   .ADCRstX1nnnH_b      ( adc_Reset_bXXL       ),
//   .ADCEnDizzX1nnnH_b   ( 1'b1                 ),
   .ADCFreezeX1nnnH     ( adc_freeze           ),
   .ADCChopEnX1nnnH     ( adc_chop_en          ),
//   .ADCContModeX1nnnH   ( 1'b0                 ),
   .ADCClkDivX1nnnH     ( adc_clkdiv           ),
//   .SDVrefSelX1nnnH     ( {adc_use_vref,1'b0}  ),
//   .BGTrimMode          ( 1'b0                 ),
   .SDinPos_a           ( pll_core__adc_in     ), 
   .ADCDoneX1nnnH       ( adc_done             ),  
   .ADCDigOutX1nnnH     ( adc_dig_out          ),
   .CkDigOutValU2N00    (                      )

);                     


endmodule // ip2211ringpll_pllljviewadc

`endif

`ifndef ip2211ringpll_LJPLL_IDV_GATE_SV
`define ip2211ringpll_LJPLL_IDV_GATE_SV

//`include "soc_clock_macros.sv"
//`include "ringpll_macros.sv"

module ip2211ringpll_ljpll_idv_gate (
   `ifdef ip2211ringpll_LJPLL_NO_UPF_SUPPORT
      input wire                     vccpll,
   `endif

   input  logic                      ClkFbMXH,
   input  logic                      idv_gate_en,
   output logic                      clkidvih
);

///========================================================================================================
/// Module Begin
///========================================================================================================

   logic ClkIdvIntIH;
   logic ClkIdvNbIH;

   // Only pass the IDV clock in openloop
   //
   `ip2211ringpll_CLKAND(ClkIdvIntIH, ClkFbMXH, idv_gate_en)

   // Add a toggle flop on the clock output in order to make the
   // duty cycle 50%
   //
   `ip2211ringpll_NB_ASSIGN(ClkIdvNbIH, clkidvih)
   `ip2211ringpll_MAKE_CLK_DIV2_RESET(clkidvih, ~ClkIdvNbIH, ClkIdvIntIH, idv_gate_en)

///========================================================================================================
/// Module End
///========================================================================================================

endmodule

`endif

`ifndef ip2211ringpll_TLCTRL_HIP_VS
`define ip2211ringpll_TLCTRL_HIP_VS

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "ringpll_macros.sv"
`ifndef ip2211ringpll_SVA_OFF
   //`include "intel_checkers.vs"
`endif
// tlctrl module is changed completely to match netlist
//module ip2211ringpll_tlctrl_hip
module ip2211ringpll_tlctrl_hip
(
 input  logic pll_core__clk_pll_div1,
 input  logic Reset_b_XXL,
 input  logic post_dist_mux__ClkPostDistMH,
 input  logic tllm_force_tight_loop,
 input logic fz_tightloop,

 output logic tlctrl_hip__TightLoopMnn0L,
 output logic tlctrl_hip__GateGridClkMnnnL
 );



///========================================================================================================
/// Module Begin
///========================================================================================================

///========================================================================================================
/// TL -> LL transition control (input to feedback divider) 
///========================================================================================================
  
   logic ClkPllMH;
   logic ClkPllMH_b;
   logic ClkPostDistNonXMH;
   logic TightLoopBMnn0L, TightLoopBMnn0H, TightLoopBMnn1L;
   logic TightLoopMnn0L;
   logic ClkSampLeadMH;
   logic GridLeadsTlMnn0H, GridLeadsTlMnn1H;
   logic ResetXXL;
   logic gridleads ;
   logic ClkPostMH_b;

   always_comb begin : RESET_GEN
      ResetXXL = ~Reset_b_XXL;
   end : RESET_GEN

 // Set post-dist clock to random value to sample at phase detector to
   // prevent faulty x-injection
  //
  //`ip2211ringpll_RANDOM_VAL_WHEN_X(ClkPostDistNonXMH, post_dist_mux__ClkPostDistMH, 1'b1)

   // Assign PLL clock to a standard name
   //
 // assign ClkPllMH = pll_core__clk_pll_div1;

   // Stage TightLoop Indicator for gating ClkGridMH
   //
   //`ip2211ringpll_CLKINV(ClkPllMH_b, pll_core__clk_pll_div1)

   ` ip2211ringpll_CLK_NAND (ClkPllMH_b, pll_core__clk_pll_div1 ,fz_tightloop)
   `ip2211ringpll_ASYNC_RST_2MSFF_META(TightLoopBMnn0L, tllm_force_tight_loop, ClkPllMH_b, Reset_b_XXL) //  SET flops were made RST flops  

  // `ip2211ringpll_ASYNC_SET_LATCH(TightLoopBMnn0H, TightLoopBMnn0L, ClkPllMH,   ResetXXL) // cmt
  // `ip2211ringpll_ASYNC_SET_LATCH(TightLoopBMnn1L, TightLoopBMnn0H, ClkPllMH_b, ResetXXL) // cmt

`ifndef ip2211ringpll_SVA_OFF
  // Custom async_drv to allow post metaflop, pre gate drive clock to be
   //  used.
   //
  //do we need to cmt this ? `ip2211ringpll_ASSERTS_GRAY_CODE(tight_loop_lock_fsm_async_drv_clksamp, {TightLoopBMnn0L, tllm_force_tight_loop}, ClkPllMH_b, ~Reset_b_XXL, `ip2211ringpll_ERR_MSG("Glitch on set or reset in tight loop lock async_drv"));
`endif

  // Create switch to disable sampling Grid with Alt FB clock & to switch
   //  feedback divider input clock
   //
 
always_comb tlctrl_hip__TightLoopMnn0L = ~ (tllm_force_tight_loop | TightLoopBMnn0L); //
  
//`ip2211ringpll_CLKAND(ClkSampLeadMH, pll_core__clk_pll_div1, TightLoopMnn0L)

   // Sample Grid clock with altfb clock to see if grid leads altfb clock
  // NOTE: GridLeadsT1Mnn0H needs to be generated using a custom phase detector cell as in BDW
 // 
  // `ip2211ringpll_MSFF(GridLeadsTlMnn0H, ClkPostDistNonXMH, pll_core__clk_pll_div1) // cmt
  // `ip2211ringpll_MSFF(GridLeadsTlMnn1H, GridLeadsTlMnn0H, ClkSampLeadMH) // cmt


 ` ip2211ringpll_CLK_NAND (ClkPostMH_b, post_dist_mux__ClkPostDistMH ,fz_tightloop)

   `ip2211ringpll_ASYNC_RST_2MSFF_META(GridLeadsTlMnn0H,TightLoopBMnn0L , ClkPostMH_b, Reset_b_XXL) //  SET flop was changed  to RST     
  assign tlctrl_hip__GateGridClkMnnnL = ~GridLeadsTlMnn0H ; //



endmodule // module tlctrl


`endif // TLCTRL_VS

`ifndef ip2211ringpll_pll_dist_lsbank_sv 
`define ip2211ringpll_pll_dist_lsbank_sv

module ip2211ringpll_pll_dist_lsbank 
(
   input  logic reset_b_xxl,
   input  logic clkpll_pre,
//   input  logic clkplldiv0_pre,
//   input  logic clkplldiv1_pre,

   output logic clkpllmh
//   output logic clkplldiv0,
//   output logic clkplldiv1
);
logic clkpllmh_3 ;
//pll_clk_ls  csb01_3 ( .out0(clkpllmh_3), .clk(clkpll_pre), .en(reset_b_xxl), .vcc_in(), .vcc_out(), .vssx());
//assign clkpllmh = ~clkpllmh_3 ;


`ifndef ip2211ringpll_INTC_NO_PWR_PINS
assign clkpllmh = clkpll_pre  ;

//pll_clk_ls  csb01_3 ( .out0(clkpllmh_3), .clk(clkpll_pre), .en(reset_b_xxl), .vcc_in(), .vcc_out(), .vssx());
//assign clkpllmh = ~clkpllmh_3 ;
 
//assign clkplldiv0 = clkplldiv0_pre & reset_b_xxl;
//assign clkplldiv1 = clkplldiv1_pre & reset_b_xxl;
`else // !`ifndef ip2211ringpll_INTC_NO_PWR_PINS
assign clkpllmh = clkpll_pre & reset_b_xxl;
//assign clkplldiv0 = clkplldiv0_pre;
//assign clkplldiv1 = clkplldiv1_pre;
`endif   

   
endmodule
`endif


`ifndef ip2211ringpll_pll_dig_lsbank_sv 
`define ip2211ringpll_pll_dig_lsbank_sv

module ip2211ringpll_pll_dig_lsbank 
(
   input  logic reset_b_xxl,
   input  logic lockrst,
   input  logic clkidv_pre,
   input  logic clkfb2,
   input  logic [9:0] adc_dig_out_pre,
   input  logic adc_done_pre,
   input  logic [1:0] viewout_pre,

   output logic pfdlockrstnh,
   output logic clkidvih,
   output logic clkfbmxh,
   output logic [9:0] adc_dig_out,
   output logic adc_done,
   output logic [1:0] viewoutnh
);
logic viewoutnh_1;
logic viewoutnh_0;
`ifndef ip2211ringpll_INTC_NO_PWR_PINS

assign pfdlockrstnh = lockrst;
assign clkidvih = clkidv_pre;
assign clkfbmxh = clkfb2;
assign adc_dig_out = adc_dig_out_pre;
assign adc_done = adc_done_pre;
assign viewoutnh = viewout_pre;

//pll_clk_ls  csb01_1 ( .out0(viewoutnh_1), .clk(viewout_pre[1]), .en(reset_b_xxl), .vcc_in(), .vcc_out(), .vssx());
//pll_clk_ls  csb01_0 ( .out0(viewoutnh_0), .clk(viewout_pre[0]), .en(reset_b_xxl), .vcc_in(), .vcc_out(), .vssx());
//assign viewoutnh = ({~viewoutnh_1,~viewoutnh_0}) ;

`else // !`ifndef ip2211ringpll_INTC_NO_PWR_PINS

assign pfdlockrstnh = lockrst & reset_b_xxl ;
assign clkidvih = clkidv_pre & reset_b_xxl;
assign clkfbmxh = clkfb2 & reset_b_xxl;
assign adc_dig_out = adc_dig_out_pre & {10{reset_b_xxl}};
assign adc_done = adc_done_pre & reset_b_xxl;
assign viewoutnh = viewout_pre & {2{ reset_b_xxl }};

//pll_clk_ls  csb01_1 ( .out0(viewoutnh_1), .clk(viewout_pre[1]), .en(reset_b_xxl), .vcc_in(), .vcc_out(), .vssx());
//pll_clk_ls  csb01_0 ( .out0(viewoutnh_0), .clk(viewout_pre[0]), .en(reset_b_xxl), .vcc_in(), .vcc_out(), .vssx());
//assign viewoutnh = ({~viewoutnh_1,~viewoutnh_0}) ;


`endif   
   
endmodule
`endif


module pll_rstdly (
output logic dlyout ,
input logic dlyin 
//input logic vccdig ,
//input logic vssx
);
assign dlyout = dlyin ;
endmodule

module pll_clk_ls ( 
output logic out0 ,
input logic clk ,
input logic en,
input logic vcc_in,
input logic vssx,
output logic vcc_out
); 
assign out0 = !(en & clk) ;
endmodule

`ifndef ip2211ringpll_IP22_RINGPLL_HIP_SV
`define ip2211ringpll_IP22_RINGPLL_HIP_SV 

//`ifndef VCSSIM_OR_EMU
//   `ifdef INTC_EMULATION
//      `define VCSSIM_OR_EMU
//   `endif
//`endif
//
//`ifndef VCSSIM_OR_EMU
//   `ifdef VCSSIM
//      `define VCSSIM_OR_EMU
//   `endif
//`endif

//`include "ljpll_dfx.vh"
//`include "soc_power_macros.sv"

//`include "ljpll_idv_gate.sv"
//`include "pllljtopana.sv"
//`include "pllljviewadc.sv"
//`include "ljpll_pllfbgen.sv"
//`include "gate_trunk_sync.sv"
////`include "trunk_mux.sv"
//`include "post_dist_mux.sv"
//`include "view_mux.sv"
//`include "pll_dist_lsbank.sv"
//`include "pll_dig_lsbank.sv" 
//`include "plllsvccpll2vccdist.sv"
//`include "tlctrl_hip.sv"
////`include "sync_gen.sv"
//`include "plldca.sv"
//`include "cpafdivtop.sv"
//`include "pll_glitchlessmux.sv"
//`include "ip2211cpafdivtop.sv"


//module cpfljfulla
module ip2211ringpll_hip
//`ifndef ip2211ringpll_LJPLL_MSV
//`ifndef ip2211ringpll_NO_VCSSIM
//#(parameter bit INTC_USE_DETAILED_AIP_MODEL = 0,
// parameter     RATIO_BITS = 10)
//`endif
//`endif
(
   `ifndef ip2211ringpll_INTC_NO_PWR_PINS
      input  wire                       vccdig,
      input  wire                       vccpll,
      input  wire                       vccdist,
      input  wire                       vccvdd2,
      input  wire                       vss,
   `endif
      input  logic                       vccref,
   input  logic                      clkrefxxh,
//   input  logic                      clkirefxih,
   input  logic                      clkpostdistmh,
   input  logic                      reset_b_xxl,
   input  logic                      bypassenxxl,
   input  logic                      bypassxxl,
   input  logic                      powergood,
   input  logic [9:0]   	     ratio,
   input  logic                      ratio_halfint,
//   input  logic                      half_int,

   input  logic [9:0]   	     ratiozdiv0,
   input  logic                      zdiv0ratiop5,
   input  logic [9:0]                ratiozdiv1,
   input  logic                      zdiv1ratiop5,

//   input  logic                      tight_loop,
   input  logic                      adc_startxxh,
   input  logic                      adc_reset_bxxl,
   input  logic [1:0]                adc_clkdiv,
   input  logic                      adc_freeze,
   input  logic                      adc_chop_en,
   input  logic                      adc_use_vref,
   input  logic [2:0]                adc_sel_in,
   
   output logic                      clkfbmxh,
   
 
   // To view pins
   //
   input  logic                      rawlockxxl,
   input  logic                      lockxxl,
   input  logic                      earlylockxxh,

   // PLL core specific DFX inputs
   //
   //input  logic                      lpcpenxxl,
   //input  logic                      cp_dis_fb_amp_samp,
   //input  logic                      cp_en_fb_amp,
   //input  logic                      cp_sel_fb_amp,
   //input  logic                      cp_iref_alt_mode,
   //input  logic                      iref_amp_disable,
   //input  logic                      iref_high_current_en,
   //input  logic                      pfd_chop_en, 
   //input  logic [2:0]                pfd_chop_val, 
   //input  logic [1:0]                pvd_mode, 
   //input  logic [2:0]                pfd_residual_pw,
   //input  logic [4:0]                cp1_trim,
   //input  logic [4:0]                cp2_trim,
   //input  logic [4:0]                skadj_ctrl,
   //input  logic [1:0]                lpf_itrim,
   //input  logic                      lpf_pg_en,
   //input  logic                      en_vco_div_16_to_iref,
   //input  logic                      en_vco_div_32_to_iref,
   //input  logic                      vco_ref_sel,
   //input  logic [3:0]                lockthresh,
   //input  logic [2:0]                iref_ctune,
   //input  logic [3:0]                iref_ftune,
   //input  logic [3:0]                vco_trim_pg,
   //input  logic [1:0]                vco_trim_cb,
   //input  logic [9:0]                misc_cfg,

   // New pins
   input  logic				fz_lpfclksel,
   input  logic				fz_nopfdpwrgate,
   input  logic				fz_tight_loopb,
   input  logic			        fz_vcosel,
   input  logic [4:0]			fz_cp1trim,
   input  logic [4:0]			fz_cp2trim,
   input  logic [1:0]			fz_cpnbias,
   input  logic [1:0]			fz_dca_cb,
   input  logic [5:0]			fz_dca_ctrl,
   input  logic [4:0]			fz_irefgen,
   input  logic [3:0]			fz_lockthresh,
   input  logic [2:0]			fz_pfd_pw,
   input  logic [1:0]			fz_pfddly,
   input  logic [4:0]			fz_skadj,
   input  logic [4:0]			fz_spare,
   input  logic [5:0]			fz_startup,
   input  logic [10:0]			fz_vcotrim,

   // LDO analog dft pins
   input  logic                 	anadft_ldovref,
   input  logic                 	anadft_ldo,
   input  logic                 	anadft_ldovfb,
  
   // Duty Cycle Adjustor Inputs
   //
   //input  logic [5:0]                dca_ctrl,
   //input  logic [1:0]                dca_cb,

   // SSC to view
   //
   input  logic                      ssc_reload,

   // SSC DFX to view
   //
   input  logic                      mod_clk_to_view,

   //input  logic [3:0]                ro_freq_sel,

   // PLL RDAC control
   //
   input  logic [3:0]                vctlrdacctlnh,

   // PLL Startup Controls
   //
   //input  logic                      irefrmodenh,
   input  logic                      vctlrdacennl,
   input  logic                      rdactovctlennh,
   input  logic                      pfdennh,
  // input  logic                      cmpenxxh,
  // input  logic                      vctl_pullupnh,
  // input  logic                      vctl_pulldnnh,
  // output logic                      compoutnh,

   // View pin settings
   //
   input  logic [1:0]                viewdigennh,
   input  logic [1:0]                viewanaennh,
   input  logic [4:0]                viewsel0 ,
   input  logic [4:0]                viewsel1 ,
   output logic [1:0]                viewoutnh,
   //output tri   [1:0]                viewanabusnh,
   output logic   [1:0]                viewanabusnh,
 
   // Tight Loop Lock Mode Inputs
   //
   input  logic                      tllm_force_tight_loop,
   input  logic                      tllm_gate_clk_trunk,

   // IDV/PLL Core Interface
   //
   input  logic                      idv_gate_en,
   output logic                      clkidvih,
   
   // SYNC Generator
   //
   //input  logic                      sync_en,
   //input  logic [4:0]                sync_pipe,
   //output logic                      sync_out,
   //output logic                      clk_sync,

   // ODCS config
   //
//   input    logic [59:0]             odcs_dig_config,
//   input    logic [34:0]             stm_config,
//   input    logic [8:0]              odcs_dll_config,
//   input    logic [1:0]              odcs_tuner_config,
//   input    logic [6:0]              opsp_config,
   
   // ODCS status 
   //
//   output   logic [4:0]              odcs_dll_delay,
//   output   logic [1:0]              odcs_trig,
//   output   logic                    stm_trig,
//   output   logic                    opsp_rise_samp,
//   output   logic                    opsp_fall_samp,

   // ODCS triggers
   //
//   input    logic                    odcsacttrig ,
//   input    logic                    analogacttrig ,

	// NEW Pins
   input logic [4:0]			ta_spare,	// some spare tap bits to the custom block
   input logic [1:0]			vcodiv_ratio,	// post vco divider setting to analog block;  was a fuse in bxt, regular input for us
   input logic [5:0]			mdiv_ratio,	// for refclk divider ratio


   // ODCS to GT
   //
//   output   logic                    odcs_kill_obsv ,


   // ADC specific DFX outputs
   //
   output logic [9:0]                adc_dig_out,
   output logic                      adc_done,
   
   output logic                      pfdlockrstnh,
   output logic                      clkplldiv0,
   output logic                      clkplldiv1,
   output logic                      clkpllmh
);

//###adding inst for RST_dleay 

logic reset_b_dly;

pll_rstdly  irstdly ( .dlyout(reset_b_dly), .dlyin(reset_b_xxl));


// `ifdef INTEL_EMULATION
// // For Emulation model only
//   assign viewoutnh[1:0] = 2'b00;
//   assign viewanabusnh[1:0] = 2'b00;
//   assign adc_dig_out[9:0] = 10'b0000000000;
//   assign adc_done = 1'b0;
//   assign pfdlockrstnh = 1'b1;

//   assign clkidvih = 1'b0; //IDV signal,  not needed for LKF
  
//   // clkpllmh = (ratio X clkref/mdivratio)
//   // clkplldiv0 = clkpllmh / ratiozdiv0
//   // clkplldiv1 = clkpllmh / ratiozdiv1

// bit [31:0] num1;
// bit [31:0] num2;
// bit [31:0] num3;

// assign num1 = (ratiozdiv0 == 4) && ( ratiozdiv1 == 125) ? 'd3072 :
//                 (ratiozdiv0 == 6) && ( ratiozdiv1 == 0) ? 'd2400 :
//                                                           32'h77359400;

// assign num2 = (ratiozdiv0 == 4) && ( ratiozdiv1 == 125) ? 'd768 :
//                 (ratiozdiv0 == 6) && ( ratiozdiv1 == 0) ? 32'h17d78400 :
//                                                           32'h1dcd6500;

// //assign num3 = (ratiozdiv0 == 4) && ( ratiozdiv1 == 125) ? 32'h24.576 :
// assign num3 = (ratiozdiv0 == 4) && ( ratiozdiv1 == 125) ? 'd25 :
//                 (ratiozdiv0 == 6) && ( ratiozdiv1 == 0) ? 32'h0:
//                                                           32'h0;
//   emu_clk_osc emu_ip22_ringpll_1 (
//         .enable(reset_b_xxl),
//         .numerator(num1), //Need to fill in this from the clk_ref, ratio and half_int
//         .denominator(1'b1), //Need to fill in this from the clk_ref, ratio and half_int
//         .clk_out(clkpllmh));

//   emu_clk_osc emu_ip22_ringpll_2 (
//         .enable(reset_b_xxl),
//         .numerator(num2), //Need to fill in this from the clk_ref, ratio and half_int
//         .denominator(1'b1), //Need to fill in this from the clk_ref, ratio and half_int
//         .clk_out(clkplldiv0));

//   emu_clk_osc emu_ip22_ringpll_3 (
//         .enable(reset_b_xxl),
//         .numerator(num3), //Need to fill in this from the clk_ref, ratio and half_int
//         .denominator(1'b1), //Need to fill in this from the clk_ref, ratio and half_int
//         .clk_out(clkplldiv1));

// `else  // NOT in EMULATION

   // Lowercase to uppercase assignments due to schematic limitation
   //
   logic                      ClkRefXXH;
   //logic                      ClkFbMXH;
   logic                      clkfb;
   logic                      clkfb2;
   logic                      ClkPostDistMH;
   logic                      Reset_b_XXL;
   logic                      VctlRdacEnNL;
   logic [1:0]                ViewDigEnNH;
   logic [1:0]                view_mux__ViewOutNnnnH;
   logic                      RawLockXXL;
   logic                      LockXXL;
   logic                      EarlyLockXXH;
   logic                      adc_StartXXH;
   logic                      adc_Reset_bXXL;
   logic 		      half_int;
   logic		      tight_loop;

   logic                      cmpenxxh;
//   logic                      vctl_pullupnh;
//   logic                      vctl_pulldnnh;
 //  logic                      compoutnh;
   // Duty Cycle Adjustor Inputs
   logic [5:0]                dca_ctrl;
   logic [1:0]                dca_cb;


//----------------------------------------------------
       logic clkrefdiv;

       // ip2211ringpll_cpafdivtop: Divider with0.5 support
        // REFCLK DIVIDER
        // if mdiv_ratio is set to 0 or 1 then bypass and use refclk only.
        //
// module definition for refclkdiv is cahnged and thus teh instantiation 
//reclkdiv        ip2211ringpll_ip2211cpafdivtop                                      refclkdiv       (
//reclkdiv                                                                       // .clkin (clkrefxxh),
//reclkdiv                                                                        .//rst (~reset_b_xxl),
//reclkdiv                                                                        // .ratio2x ({4'b0,mdiv_ratio,1'b0}),
//reclkdiv								 	// .ratio2x ({4'b0,mdiv_ratio[5],(mdiv_ratio[4]),(mdiv_ratio[3]),(mdiv_ratio[2]),(mdiv_ratio[1]) ,(ratio2x[1])}) ,
//reclkdiv                                                                        //.clkout (clkrefdiv)
//reclkdiv									 //);
// new inst for refclkdiv 
ip2211ringpll_ip2211cpafdivtop_refclk                                      refclkdiv       (
                                                                        .clkin (clkrefxxh),
                                                                        //.rst (~reset_b_xxl),
                                                                        .rst(~reset_b_dly),
									.clkout (clkrefdiv),
									 .* );


        logic refclkbypass;
        logic clkrefmux;

        always_comb begin : REFCLKDIVIDE
        // if the refclk divide mdiv_ratio is 0 or 1 then pass refclk as is.
        // For any value > 1 provide divided refclk to pllcore.
        //
        //refclkbypass = ((mdiv_ratio == 6'd0) || (mdiv_ratio == 6'd1));
        //clkrefmux = (refclkbypass) ? clkrefxxh :
      //                               clkrefdiv ;
        clkrefmux = clkrefdiv;     

        end : REFCLKDIVIDE
//----------------------------------------------------

       logic clkref_prediv;
       assign clkref_prediv = clkrefxxh;

   //assign ClkRefXXH           = clkrefxxh;
   assign ClkRefXXH           = clkrefmux;

   assign tight_loop		= ~fz_tight_loopb;
   assign dca_ctrl		= fz_dca_ctrl;
   assign dca_cb		= fz_dca_cb;
   assign half_int	      = ratio_halfint;
   assign ClkPostDistMH       = clkpostdistmh;
   assign Reset_b_XXL         = reset_b_xxl;
   assign ViewDigEnNH         = viewdigennh;
   assign RawLockXXL          = rawlockxxl;
   assign LockXXL             = lockxxl;
   assign EarlyLockXXH        = earlylockxxh;
   assign adc_StartXXH        = adc_startxxh;
   assign adc_Reset_bXXL      = adc_reset_bxxl;
   assign VctlRdacEnNL        = vctlrdacennl;

   //assign clkfbmxh            = ClkFbMXH;
   //assign clkfbmxh            = clkfb2;

   //=============================================================================
   // Internal Wire Declaration
   //
   //    Declare wires for internal connectivity grouped by driver
   //=============================================================================

   // Post Dist Mux
   //
   logic             post_dist_mux__ClkPostDistMH;

   // ODCS Dig
   //
//   logic   [4:0]     odcs_dig__OdcsRiseCodeMnn0L;
//   logic   [4:0]     odcs_dig__OdcsFallCodeMnn1H;
//   logic             odcs_dig__OdcsKillRiseMnn0L;
//   logic             odcs_dig__OdcsKillFallMnn1H;
//   logic             odcs_dig__OdcsModeEnNH;
//   logic             odcs_dig__CguBrkAnalogActM759H;
//   logic             odcs_dig__CkOdcsStmM1N22 ;
//   logic             odcs_dig__OdcsRiseBase0MnnnH ;
//   logic             odcs_dig__OdcsFallBase0MnnnH ;
//   logic             odcs_dig__OdcsRiseVal1MnnnH ;
//   logic             odcs_dig__OdcsFallVal1MnnnH ;

   // STM/IFDIM block
   //
//   logic             stm_ifdim__StmEnableNnnnH;
//   logic             stm_ifdim__StmStopHiNnnnH;
//   logic             stm_ifdim__StmStopMnnnH;

   // Gate Trunk Sync
   //
   logic gate_trunk_sync__GateClkTrunkML;

   // Trunk Mux
   //
   logic trunk_mux__ClkTrunkMH;
   logic trunk_mux__DistPwrGoodRL;
   logic trunk_mux__ClkRoRH;
   logic trunk_mux__ClkPllMH;

   // ODCS DLL
   //
//   logic odcs_dll__ClkOdcsDllOutMH;
//   logic odcs_dll__CguBrkActOdcsM756H ;
//   logic odcs_dll__CguBrkAnalogActM756H ;
//   logic odcs_dll__AnalogActTrigM738H ;
//   logic odcs_dll__OdcsDllAddDelayMnnnL ;
//   logic odcs_dll__OdcsDllPhDetEarlyMnnnH ;
//   logic odcs_dll__OdcsDllPhDetLateMnnnH ;
//   logic odcs_dll__OdcsDllUpdateMnnnL ;
//   logic odcs_dll__ForceUseDllNH ;
//   logic odcs_dll__ClkDlGatedMH ;

   // ODCS Tuner
   //
//   logic odcs_tuner__ClkTuneMH;

   // PLL Core
   //
   logic pll_core__clk_pll_div1;
   wire  pll_core__adc_in;
   logic pll_core__cp1clk;
   logic pll_core__cp1aclk;
   logic pll_core__cp2clk;
   logic pll_core__cp2aclk;

   // LS -> DIST
   //
   logic pll_core__clk_pll_div1_ls_dist;
   logic gate_trunk_sync__GateClkTrunkML_ls_dist;

   // PLL feedback generator
   //
   logic pll_fbgen__tight_loop;
//   logic pll_fbgen__ClkPllFdivMH;
   //logic [7:0] pll_fbgen__RatioSampMXH;
//   logic [9:0] pll_fbgen__RatioSampMXH;

   // Tight Loop Lock Mode
   //
   logic    tlctrl_hip__TightLoopMnn0L;
   logic    tlctrl_hip__GateGridClkMnnnL;
                
   //`ifdef VCSSIM_OR_EMU
   `ifndef INTC_NO_VCSSIM_OR_EMU
   logic pllfbgen__haltclk_inst;
   `endif


   // pllclk divider0 and divider1
	logic pll_core_clkd;
	logic pll_core_clkm;
        logic clkplldiv0gated;
        logic clkplldiv1gated;
        logic clkplldiv0bypass;
        logic clkplldiv1bypass;
        logic clkplldiv0mux;
        logic clkplldiv1mux;
   	logic clkplldiv0_pre;
   	logic clkplldiv1_pre;

   // Output level shifters
	logic lockrst;
 	logic clkidv_pre;
   	logic [9:0] adc_dig_out_pre;
   	logic       adc_done_pre;
   	logic [1:0] viewout_pre;

   assign viewout_pre         = view_mux__ViewOutNnnnH;

   //=============================================================================
   // Submodule Declarations
   //
   //   Declare the top level SIP hierarchy of LJPLL
   //
   //   The top level hierarchy is as follows:
   //    -hip
   //    --ljpll_core
   //    --pllfbgen
   //    --trunk_mux
   //    --tlctrl
   //=============================================================================
    
      // LJPLL Core
      //   LJPLL Analog components (e.g. ip2211ringpll_PFD, CP, ip2211ringpll_VCO, etc.)
      //
      ip2211ringpll_pllljtopana
         //`ifndef ip2211ringpll_LJPLL_MSV
         //`ifndef ip2211ringpll_NO_VCSSIM
         //   #(.INTC_USE_DETAILED_AIP_MODEL(INTC_USE_DETAILED_AIP_MODEL),
         //     .RATIO_BITS(RATIO_BITS))
         //`endif
         //`endif
// pin names are changed by taking SCh as reference 
pll_core   (
            //`ifdef ip2211ringpll_LJPLL_MSV
             `ifndef ip2211ringpll_INTC_NO_PWR_PINS
               .vccpll          (vccpll),
               .vccref          (vccdig),
               .vccvdd2         (vccvdd2),
             `endif
            //.clkfb              (     ClkFbMXH                ),
            .clkfb                (     clkfb                   ),
            .clkref               (     clkrefmux               ),
            .cp1_trim            (    fz_cp1trim              ),
            .cp2_trim             (           fz_cp2trim              ),
            .vctlrdac             (     vctlrdacctlnh           ),
            .vctlrdacen           (     vctlrdacennl            ),
            .rdactovctlen         (     rdactovctlennh          ),
            .pfden                (     pfdennh                 ),
           `ifndef INTC_NO_VCSSIM_OR_EMU
              .clk_iref             (    clkrefmux               ),
           `endif
            .irefvcoclksel        (         fz_vcosel               ),
            .pfd_residual_pw      (   fz_pfd_pw               ),
            .skadj_ctrl           (       fz_skadj                ),
          `ifdef INTC_NO_VCSSIM_OR_EMU
            .fz_vcotrim           ( fz_vcotrim), 
	    .fz_cpnbias    (~fz_cpnbias),
            .fz_pfddly      ({fz_pfddly[1],!fz_pfddly[0]}),
	    .fz_irefgen (fz_irefgen),
	    .fz_startup (fz_startup),
	    .fz_nopfdpwrgate (fz_nopfdpwrgate),
          `endif
            .lockthresh           (          fz_lockthresh           ),
          `ifndef INTC_NO_VCSSIM_OR_EMU
            .vco_trim_pg          (   fz_vcotrim[9:6]         ),
            .vco_trim_cb          (   fz_vcotrim[2:0]         ),
            .viewsel0             (           viewsel0[3:0]           ),
            .viewsel1             (           viewsel1[3:0]           ),
          `endif
            .viewanaen            (     viewanaennh             ),
            // .reset_b              (     reset_b_xxl             ),
            .reset_b              (     reset_b_dly             ),
            .adc_sel_in           (     adc_sel_in              ),
            `ifdef INTC_NO_VCSSIM_OR_EMU
             .cp1clk               (           pll_core__cp1clk        ),
             .cp1aclk              (           pll_core__cp1aclk       ),
             .cp2clk               (           pll_core__cp2clk        ),
             .cp2aclk              (           pll_core__cp2aclk       ),
            `endif
            .pfdlockrst           (        lockrst                 ),
            .viewanabus           (     viewanabusnh            ),
            .adc_in               (     pll_core__adc_in        ),
            .pdivrat              (     vcodiv_ratio            ),
            .anadft_ldovfb        (     anadft_ldovfb           ),      // LDO DFT pins
            .anadft_ldovref       (     anadft_ldovref          ),
            .anadft_ldo           (     anadft_ldo              ),
            //.lpf_itrim            ( 2'b00   ),
            //.pfd_chop_en          ( 1'b0  ),
            //.pfd_chop_val         (3'b000   ),
            //.pvd_mode             ( 2'b00  ),
            //.irefrmodeen          (1'b0  ),
            //.en_vcodiv16toiref    (1'b0  ),
            //.en_vcodiv32toiref    (1'b0  ),
            //.irefhighcurr_en      (1'b0   ),
            //.lpcpen               (1'b0   ),
            //.cpdisfbampsamp       (1'b0   ),
            //.cpenfbamp            ( 1'b0  ),
            //.cpselfbamp           (1'b0   ),
            //.cpirefaltmode        (1'b0   ),
            //.iref_ctune           (3'b000   ),
            //.iref_ftune           (4'b0000   ),
            //.irefbypassamp_mode   (1'b0  ),
            //.lpf_pg_en            (1'b0  ),
            .clkpll               (   pll_core__clk_pll_div1   )
                       `ifndef ip2211ringpll_LJPLL_MSV
            , .*
            `endif
      );


      // PLL Post Distribution MUX
      //   This mux selects the post distribution clock feedback path to
      //   the F-Divider and the tight loop lock mode HIP.  The DLL is
      //   expected to operate as a distribution replica.
      //
      //ip2211ringpll_post_dist_mux                           ip2211ringpll_post_dist_mux ( .* );
	assign	post_dist_mux__ClkPostDistMH = ClkPostDistMH;


      // PLL Feedback Generator
      //   Generates the feedback clock to the PLL
      //
      ip2211ringpll_ljpll_pllfbgen   
	 //#(
         //`ifndef ip2211ringpll_LJPLL_MSV
         //`ifndef ip2211ringpll_NO_VCSSIM
         //   .INTC_USE_DETAILED_AIP_MODEL(1)
         //`endif
         //`endif
	//)
         //   .RATIO_BITS(10))                   pll_fbgen  ( .* );
                                                 pll_fbgen  (
								.reset_b_xxl(reset_b_dly),
								 .half_int(ratio_halfint),
								 .* );

      // Level shifter PLL->DIST
      //   Include level shifters for tools that dont support ip2211ringpll_UPF
      //
      //ip2211ringpll_plllsvccpll2vccdist                      lspll2dist ( .* );

      // Trunk Gate Syncronizer
      //   Allows for TLLM to deterministically enable the clock
      //   distribution (no chopping) and also allows for deterministic
      //   global alignment points for HVM debug
      //
      //ip2211ringpll_gate_trunk_sync                          ip2211ringpll_gate_trunk_sync ( 
		//			.Reset_b_XXL			(Reset_b_XXL),
		//			.ClkFbMXH			(clkfb),
		//			.pll_core__clk_pll_div1		(pll_core__clk_pll_div1),
		//			//.tllm_gate_clk_trunk		(tllm_gate_clk_trunk),
		//			.tllm_gate_clk_trunk		(1'b0),  // TBD: Connect it if we use it for long loop in the future.
		//			.gate_trunk_sync__GateClkTrunkML	(gate_trunk_sync__GateClkTrunkML)
 		//				);

      // Trunk Mux
      //   Chooses the correct trunk based on PLL mode and power/reset
      //   state.
      //
      //
      //trunk_mux      #(.HAS_RO(0))             trunk_mux  ( 
      //							.ro_freq_sel (4'b0000),
      //							.* );

      // GMUX
      // Glichless mux between refclk and pllclk
      // This is used in place of Trunk Mux.
      //
      ip2211ringpll_pll_glitchlessmux		ip2211ringpll_pll_glitchlessmux (
		  `ifndef ip2211ringpll_INTC_NO_PWR_PINS
      		.vccpll		(vccpll),
      		.vss		(vss),
   		`endif

   		.bypass		(bypassxxl),
   		// in netlist bypassen was not usedat hip interface ,  where as rst pin was connected to bypassen pin of gmux ,  .bypassen	(bypassenxxl),
		.bypassen	(reset_b_xxl),

   		.pllclk		(pll_core_clkm),
   		.refclk		(clkrefxxh),
   	//	.rb		(reset_b_xxl),
		.rb		(reset_b_dly),
   		//.rb		(bypassenxxl),

   		.muxclk		(pll_core_clkd)
	);

      // PLL DCA
      //   Static duty cycle corrector used to correct duty cycle offset
      //   introduced in the forward clock path
      //
     ip2211ringpll_plldca                                   dca       ( 
		`ifndef ip2211ringpll_NO_VCSSIM
		`ifdef INTC_SIM
		 .reset_b_xxl		(reset_b_xxl),
		`endif
		`endif
		.dca_ctrl		(dca_ctrl),
		.dca_cb			(dca_cb),
		.pll_core_clkm		(pll_core__clk_pll_div1),
		.clkpllmh		(pll_core_clkm)
			);

      // ODCS DIG
      //   This block sits on VCCDIST and acts as the control logic for the
      //   tuner.  It receives a microbreakpoint from the salmon ladder and
      //   feeds delay codes to the tuner to shape the clock to the
      //   distribution.
      //
//      pllodcsdig                               odcs_dig  ( .* );

      // ODCS IFDIM/STM
      //   This block contains the IFDIM/STM logic that extend the ODCS
      //   architecture to provide additional debug capability
      //
//      pllodcsstm                               stm_ifdim ( .* );

      // ODCS DLL
      //   This delay line should be calibrated with the RO from the trunk
      //   mux to match the distribution delay.  When enabled, the delay
      //   of the delay line should approximate that of the distribution.
      //
//      pllodcsdll                               odcs_dll   ( .* );

      // ODCS Tuner
      //   This block sits in the forward clock path and acts as a rise
      //   delay / fall delay tuner when ODCS is disabled.  It otherwise
      //   acts as a buffer feeding the clock distribution
      //
//      odcs_tuner                               odcs_tuner ( .* );

      // OPSP
      //    On purpose speedpath allows ODCS to be tested by forcing
      //    a speedpath to occur when shmooing ref clock then using ODCS to
      //    correct the speedpath.
      //
//      pllopsp                                  odcs_opsp  ( .* );

      // SYNC Generator
      //    This block generates the sync signal used for deterministic
      //    clock crossing schemes on chip.
      //
      //sync_gen                                 sync_gen   ( .* );
      //sync_gen                                 sync_gen #(.RATIO_BITS(RATIO_BITS))  ( .* );

      // View Mux
      //   Visibility muxes for output of signals onto the DFX view pins
      //
      //ip2211ringpll_view_mux                                 ip2211ringpll_view_mux   ( .* );
      ip2211ringpll_view_mux                                 ip2211ringpll_view_mux   ( 
					`ifdef ip2211ringpll_LJPLL_NO_UPF_SUPPORT
						.vccpll		(vccpll),
					`endif
					.pll_core__clk_pll_div1	(pll_core__clk_pll_div1),
					.ClkPostDistMH		(ClkPostDistMH),
					.clkref_prediv		(clkref_prediv),
					.VctlRdacEnNL		(VctlRdacEnNL),
					.ClkRefXXH		(ClkRefXXH),
					//.ClkFbMXH		(ClkFbMXH),
					.ClkFbMXH		(clkfb),
					//.Reset_b_XXL		(Reset_b_XXL),
					.Reset_b_XXL		(reset_b_dly),
					.pfdennh		(pfdennh),
					.pll_fbgen__tight_loop	(pll_fbgen__tight_loop),
					.powergood		(powergood),
					.ViewDigEnNH		(ViewDigEnNH),
					.viewsel0		(viewsel0),
					.viewsel1		(viewsel1),
					.RawLockXXL		(RawLockXXL),
					.LockXXL		(LockXXL),
					.EarlyLockXXH		(EarlyLockXXH),
					.ssc_reload		(ssc_reload),
					.mod_clk_to_view	(mod_clk_to_view),
					.view_mux__ViewOutNnnnH	(view_mux__ViewOutNnnnH)
					);
// View adc pin names are changed to match netlist , pins are case sensitive 
      // View ADC
      //   Used for DFT debug of analog signals. This ADC is capable of
      //   sending analog voltages in the form of a digital code to the TAP
      //
      //ip2211ringpll_pllljviewadc                             view_adc   ( .* );
        ip2211ringpll_pllljviewadc                             view_adc   ( 
                                        `ifndef ip2211ringpll_INTC_NO_PWR_PINS
                                                .vccpll             (1'b1),
                                        `endif
                                                .vccref                (1'b1),

                                        .ClkRefXXH              (clkref_prediv),
                                        .adc_Reset_bXXL         (adc_Reset_bXXL),
                                        .adc_StartXXH            (adc_StartXXH),
                                        .adc_clkdiv             (adc_clkdiv),
                                        .adc_freeze             (adc_freeze),
                                        .adc_chop_en            (adc_chop_en),
                                        //.adc_use_vref          (adc_use_vref),
                                        .pll_core__adc_in        (pll_core__adc_in),
                                        .adc_dig_out            (adc_dig_out_pre),
                                        .adc_done               (adc_done_pre)
                                        );

      
      // IDV Gate
      //   Gate IDV clock during normal PLL operation (openloop=0)
      //
      ip2211ringpll_ljpll_idv_gate                           idv_gate   ( 
					`ifdef ip2211ringpll_LJPLL_NO_UPF_SUPPORT
					.vccpll		(vccpll),
					`endif

					.ClkFbMXH	(clkfb2),
					.idv_gate_en	(idv_gate_en),
					.clkidvih	(clkidv_pre)
					);

      // IDV GateTight loop lock control
      //   Tight loop lock mode logic on high freq clock
      //
      ip2211ringpll_tlctrl_hip                               ip2211ringpll_tlctrl_hip ( .fz_tightloop(fz_tight_loopb), 
                                                                                        .Reset_b_XXL(reset_b_dly), 
											.* );

logic zdiv1_sync_rst,zdiv0_sync_rst;

      // ip2211ringpll_cpafdivtop: Divider with0.5 support
      // ZDIV0


    // synchronizing the reset from clkref domain to vco clock domain
     //`ip2211ringpll_ASYNC_SET_2MSFF_META(zdiv0_sync_rst,1'b0,clkpllmh ,EarlyLockXXH )
//     `ip2211ringpll_ASYNC_SET_2MSFF_META(zdiv0_sync_rst,1'b0,clkpllmh , reset_b_dly)
      //
      //ip2211ringpll_cpafdivtop	#(.RATIO_BITS(RATIO_BITS))		vcozdiv0   ( 
      //ip2211ringpll_cpafdivtop			vcozdiv0   ( 
      ip2211ringpll_ip2211cpafdivtop			vcozdiv0   ( 
											.clkin (clkpllmh),
											//.rst (~reset_b_xxl),
											.rst (reset_b_dly),
										//	.rst (~EarlyLockXXH),
											.ratio2x ({ratiozdiv0,zdiv0ratiop5}),
											// .clkout (clkplldiv0mux) ,
											.clkout(clkplldiv0) ,
                                                                                        .enb(1'b0),
											.divbygt1() 
										);

      // ip2211ringpll_cpafdivtop: Divider with0.5 support
      // ZDIV1
      //
    // synchronizing the reset from clkref domain to vco clock domain
     //`ip2211ringpll_ASYNC_SET_2MSFF_META(zdiv1_sync_rst,1'b0,clkpllmh,EarlyLockXXH )
//     `ip2211ringpll_ASYNC_SET_2MSFF_META(zdiv1_sync_rst,1'b0,clkpllmh,reset_b_dly )
      //ip2211ringpll_cpafdivtop	#(.RATIO_BITS(RATIO_BITS))		vcozdiv1   ( 
      //ip2211ringpll_cpafdivtop			vcozdiv1   ( 
      ip2211ringpll_ip2211cpafdivtop			vcozdiv1   ( 
											.clkin (clkpllmh),
											//.rst (~reset_b_xxl),
											.rst (reset_b_dly ),
											//.rst (~EarlyLockXXH),
											.ratio2x ({ratiozdiv1,zdiv1ratiop5}),
											// .clkout (clkplldiv1mux),
                                                                                        .enb(1'b0),
											.clkout(clkplldiv1),
                                                                                        .divbygt1()
										);


        always_comb begin : CLKPLLDIV0DIVIDE 
        // if the refclk divide ratiozdiv0 is 0 or 1 then pass clkpllmh as is.
        // For any value > 1 provide divided refclk to pllcore.
        //
        clkplldiv0gated = (ratiozdiv0 == 10'd0);

        //clkplldiv0bypass = ((ratiozdiv0 == 10'd0) || (ratiozdiv0 == 10'd1));
        clkplldiv0bypass = (ratiozdiv0 == 10'd1);

        // defined inside module definition clkplldiv0 = (clkplldiv0gated) ? 1'b0 : (clkplldiv0bypass) ? clkpllmh : clkplldiv0mux ;

        end : CLKPLLDIV0DIVIDE


        always_comb begin : CLKPLLDIV1DIVIDE 
        // if the refclk divide ratiozdiv1 is 0 or 1 then pass clkpllmh as is.
        // For any value > 1 provide divided refclk to pllcore.
        //
        clkplldiv1gated = (ratiozdiv1 == 10'd0);

        //clkplldiv1bypass = ((ratiozdiv1 == 10'd0) || (ratiozdiv1 == 10'd1));
        clkplldiv1bypass = (ratiozdiv1 == 10'd1);

        // defined inside module def  clkplldiv1 = clkplldiv1gated ? 1'b0 : (clkplldiv1bypass) ? clkpllmh : clkplldiv1mux ;

        end : CLKPLLDIV1DIVIDE

///========================================================================================================
// OUTPUT Level shifters
// ip2211ringpll_LS_WITH_AND_FW(o, pro, a, vcc_in, en)
//
logic clkpll_pre;
assign clkpll_pre = pll_core_clkd;


ip2211ringpll_pll_dist_lsbank ipll_dist_lsbank 
(
 .reset_b_xxl(reset_b_dly),
 .clkpll_pre,
// .clkplldiv0_pre,
// .clkplldiv1_pre,

 .clkpllmh
// .clkplldiv0,
// .clkplldiv1
);

ip2211ringpll_pll_dig_lsbank ipll_dig_lsbank
(
   .reset_b_xxl,
   .lockrst,
   .clkidv_pre,
   .clkfb2,
   .adc_dig_out_pre,
   .adc_done_pre,
   .viewout_pre,

   .pfdlockrstnh,
   .clkidvih,
   .clkfbmxh,
   .adc_dig_out,
   .adc_done,
   .viewoutnh
);

   
`ifndef ip2211ringpll_INTC_NO_PWR_PINS
//`ip2211ringpll_LS_WITH_AND_FW(clkpllmh, vccdist, clkpll_pre, vccpll, reset_b_xxl)
//`ip2211ringpll_LS_WITH_AND_FW(clkplldiv0, vccdist, clkplldiv0_pre, vccpll, reset_b_xxl)
//`ip2211ringpll_LS_WITH_AND_FW(clkplldiv1, vccdist, clkplldiv1_pre, vccpll, reset_b_xxl)

//`ip2211ringpll_LS_WITH_AND_FW(pfdlockrstnh, vccdist, lockrst, vccdig, reset_b_xxl)
//`ip2211ringpll_LS_WITH_AND_FW(clkidvih, vccdist, clkidv_pre, vccdig, reset_b_xxl)
//`ip2211ringpll_LS_WITH_AND_FW(clkfbmxh, vccdist, clkfb2, vccdig, reset_b_xxl)
//`ip2211ringpll_LS_WITH_AND_FW(adc_dig_out, vccdist, adc_dig_out_pre, vccdig, reset_b_xxl)
//`ip2211ringpll_LS_WITH_AND_FW(adc_done, vccdist, adc_done_pre, vccdig, reset_b_xxl)
//`ip2211ringpll_LS_WITH_AND_FW(viewoutnh, vccdist, viewout_pre, vccdig, reset_b_xxl)
`else // !`ifndef ip2211ringpll_INTC_NO_PWR_PINS
//assign clkpllmh = clkpll_pre;
//assign clkplldiv0 = clkplldiv0_pre;
//assign clkplldiv1 = clkplldiv1_pre;

//assign pfdlockrstnh = lockrst & reset_b_xxl;
//assign clkidvih = clkidv_pre & reset_b_xxl;
//assign clkfbmxh = clkfb2 & reset_b_xxl;
//assign adc_dig_out = adc_dig_out_pre & reset_b_xxl;
//assign adc_done = adc_done_pre & reset_b_xxl;
//assign viewoutnh = viewout_pre & reset_b_xxl;

`endif   

endmodule

`endif

`ifndef ip2211ringpll_POST_DIST_MUX_SV
`define ip2211ringpll_POST_DIST_MUX_SV

module ip2211ringpll_post_dist_mux (
   input  logic clkpostdistmh,
//   input  logic odcs_dll__ClkOdcsDllOutMH,
//   input  logic odcs_dll__ForceUseDllNH,
//   input  logic odcs_dig__OdcsModeEnNH,
   output logic post_dist_mux__ClkPostDistMH
);


   // When ODCS mode is enabled or when usedl is selected, select the delay
   // line for the feedback path
   //
   always_comb begin : POST_DIST_MUX
//      post_dist_mux__ClkPostDistMH = (odcs_dll__ForceUseDllNH | odcs_dig__OdcsModeEnNH) ? odcs_dll__ClkOdcsDllOutMH
//                                                                                        : clkpostdistmh               ;
	post_dist_mux__ClkPostDistMH = clkpostdistmh;

   end : POST_DIST_MUX


endmodule

`endif


//`celldefine
//
// LDO model created for P1222. -
//
`ifndef ip2211ringpll_ldopgd_sv
`define ip2211ringpll_ldopgd_sv

//`include "soc_macros.sv"

module ip2211ringpll_ldopgd
(   
//`ifdef PWRPINS
`ifndef ip2211ringpll_INTC_NO_PWR_PINS
    `ifdef SFE_BMOD_PWR_USE_REAL
        input  real vnnaon_nom,
        input  real vccdig,		//vcc_main,
        input  real vccldo,		//vcc_hv,
        input  real vssx,
        output real vccpll,
    `else
        input  logic vnnaon_nom,
        input  logic vccdig,		//vcc_main,
        input  logic vccldo,		//vcc_hv,
        input  logic vssx,
        output logic vccpll,
    `endif
`endif

// Analog Signals
`ifdef SFE_BMOD_ANA_USE_REAL
    input real  ldo_vref,
`else
    input logic ldo_vref,
`endif


    input logic		powergood_vnn,
    input logic [1:0] 	fz_ldo_vinvoltsel,	//d_ldo_en_1p24v,
    input logic 	fz_ldo_faststart,	//d_fast_start_i,
    input logic 	clkref,			//d_refclk_i,
    input logic 	fz_ldo_bypass,		//d_ldo_bypass_i,
    input logic 	fz_ldo_extrefsel,	//d_ldo_extrefsel_i,
    input logic [3:0] 	fz_ldo_fbtrim,		//d_ldo_fbtrim,
    input logic [3:0] 	fz_ldo_reftrim,		//d_ldo_reftrim,
    input logic 	ldo_enable,		//d_ldo_pon_i,
    input logic 	ta_ldo_hiz_debug,
    input logic 	ta_ldo_idq_debug,

    input logic         powergood_vccdig,
    input logic         fz_spare_4_strong_ladder_en,

    //inout tri   viewana,
    output tri          viewana,
    // LDO analog dft pins
    output logic        anadft_ldovref,
    output logic        anadft_ldovfb
);


`ifdef SFE_BMOD_ANA_USE_REAL
// Parameter declaration
parameter real vnnaon_nom_min  = 0.675;   // Typ voltage 0.77V
parameter real vnnaon_nom_max  = 0.825;
parameter real vccdig_min      = 0.675;   // Typ voltage 0.77V
parameter real vccdig_max      = 0.825;
parameter real vccldo_min      = 1.15;   // Typ voltage 1.25V
parameter real vccldo_max      = 1.32;
parameter real vssx_min        = -0.05;   // Typ voltage 0V
parameter real vssx_max        = 0.05;
parameter real vref_min        = 0.985; // ideal val=1.0V
parameter real vref_max        = 1.015; 
parameter real R_resunit       = 1.649e03;
parameter real ldo_vref_K1     = 36;
parameter real ldo_vref_K2     = 54;
parameter real vccldo_K1       = 48;
parameter real vccldo_K2       = 42;
parameter real maxreftrimval   = 15;
`endif

// ELS - HSD 16013510558
parameter real OUTDELAY_RISE   = 4;  // in us
parameter real OUTDELAY_FALL   = 0.1;  // in us
//`endif

// Internal variables
logic ldo_vref_ok, vnnaon_nom_ok, vccdig_ok, vccldo_ok, vssx_ok, supply_ok;
logic pwr_vccdig_ok, pwr_vnn_ok;
logic d_ldo_bypass_i_delay, d_ldo_bypass_i_int, ldo_enabled;
logic d_ldo_pon_i_delay, d_ldo_pon_i_int;
logic debugen;
//TODO : need to check the type
//logic analog_debug_out_o;
wire analog_debug_out_o;

`ifdef SFE_BMOD_ANA_USE_REAL
real vref_int, vccpll_real;
real ldo_vref_is, vccldo_is;
real del;
`else
logic vref_int;
`endif

//real del;

`ifdef SFE_BMOD_ANA_USE_REAL
  real vccpll_int;
`else
  logic vccpll_int;
`endif


// Supply range checks
`ifndef ip2211ringpll_INTC_NO_PWR_PINS
  `ifdef SFE_BMOD_PWR_USE_REAL // Full AMS Mode
	assign vnnaon_nom_ok = ((vnnaon_nom >= vnnaon_nom_min) & (vnnaon_nom <= vnnaon_nom_max)) ? 1'b1 : 1'b0 ;
	assign vccdig_ok = ((vccdig >= vccdig_min) & (vccdig <= vccdig_max)) ? 1'b1 : 1'b0 ;
	assign vccldo_ok = ((vccldo >= vccldo_min) & (vccldo <= vccldo_max)) ? 1'b1 : 1'b0 ;
	assign vssx_ok   = ((vssx   >= vssx_min)   & (vssx   <= vssx_max))   ? 1'b1 : 1'b0 ;

	assign supply_ok = vnnaon_nom_ok & vccdig_ok & vccldo_ok & vssx_ok ;

  `else // Digital Functional Mode
	assign supply_ok = vnnaon_nom & vccdig & vccldo & ~vssx ;
  `endif
`else // UPF Mode
	assign supply_ok = 1'b1 ;
`endif // end of `ifndef ip2211ringpll_INTC_NO_PWR_PINS


// ldo_vref range check
`ifdef SFE_BMOD_ANA_USE_REAL
    assign ldo_vref_ok = ( (ldo_vref >= vref_min) & (ldo_vref <= vref_max) ) ? 1'b1 : 1'b0 ;
`else
    assign ldo_vref_ok = ldo_vref ;
`endif


// powergood enables
assign pwr_vccdig_ok = supply_ok ? powergood_vccdig : 1'b0 ;
assign pwr_vnn_ok    = supply_ok ? powergood_vnn : 1'b0 ;


// vref selection
`ifndef ip2211ringpll_INTC_NO_PWR_PINS
 `ifdef SFE_BMOD_ANA_USE_REAL
    assign vref_int = fz_ldo_extrefsel ? ldo_vref_is : vccldo_is ;
 `else
    assign vref_int = fz_ldo_extrefsel ? ldo_vref : vccldo ;
 `endif
 `else
    assign vref_int = (ldo_enabled & pwr_vnn_ok) ? 1'b1 : 1'b0;
 `endif

// vref calculation  // if reftrim = 0000 => interbal setting to code 9
`ifdef SFE_BMOD_ANA_USE_REAL
    assign ldo_vref_is = ((ldo_vref_K2 + fz_ldo_reftrim) / (ldo_vref_K2 + ldo_vref_K1 + maxreftrimval)) * ldo_vref ;
// vccldo_is calc: reftrim = vccldo=1.2V => reftrim= 9
    assign vccldo_is   = ((vccldo_K2 + fz_ldo_reftrim) / (vccldo_K2 + vccldo_K1 + maxreftrimval)) * vccldo ;
`endif

`ifdef SFE_BMOD_ANA_USE_REAL
// fbtrim
always @ (fz_ldo_fbtrim or fz_ldo_reftrim)
begin
    casex (fz_ldo_fbtrim)
	4'b0000:    vccpll_real = 0.855 ; 
	4'b0001:    vccpll_real = 0.735 ; 
	4'b0010:    vccpll_real = 0.749 ; 
	4'b0011:    vccpll_real = 0.762 ; 
	4'b0100:    vccpll_real = 0.776 ; 
	4'b0101:    vccpll_real = 0.791 ; 
	4'b0110:    vccpll_real = 0.806 ; 
	4'b0111:    vccpll_real = 0.822 ;
	4'b1000:    vccpll_real = 0.838 ; 
	4'b1001:    vccpll_real = 0.855 ; 
	4'b1010:    vccpll_real = 0.873 ; 
	4'b1011:    vccpll_real = 0.891 ; 
	4'b1100:    vccpll_real = 0.910 ; 
	4'b1101:    vccpll_real = 0.930 ; 
	4'b1110:    vccpll_real = 0.951 ; 
	4'b1111:    vccpll_real = 0.973 ; 
	default:    vccpll_real = 0.855 ; // same as 4'b0000 and 4'b1001
    endcase

    casex (fz_ldo_reftrim)
	4'b0000:    vccpll_real = 0.855 ; 
	4'b0001:    vccpll_real = 0.722 ; 
	4'b0010:    vccpll_real = 0.739 ; 
	4'b0011:    vccpll_real = 0.755 ; 
	4'b0100:    vccpll_real = 0.772 ; 
	4'b0101:    vccpll_real = 0.789 ; 
	4'b0110:    vccpll_real = 0.805 ; 
	4'b0111:    vccpll_real = 0.822 ;
	4'b1000:    vccpll_real = 0.838 ; 
	4'b1001:    vccpll_real = 0.855 ; 
	4'b1010:    vccpll_real = 0.872 ; 
	4'b1011:    vccpll_real = 0.888 ; 
	4'b1100:    vccpll_real = 0.905 ; 
	4'b1101:    vccpll_real = 0.921 ; 
	4'b1110:    vccpll_real = 0.938 ; 
	4'b1111:    vccpll_real = 0.954 ; 
	default:    vccpll_real = 0.855 ; // same as 4'b0000 and 4'b1001
    endcase

end  // end of always 
`endif

   `ifdef INTEL_EMULATION
      assign d_ldo_bypass_i_delay = fz_ldo_bypass;
      assign d_ldo_pon_i_delay    = ldo_enable;
   `else
      assign #50ps  d_ldo_bypass_i_delay = fz_ldo_bypass;
      assign #500ps d_ldo_pon_i_delay    = ldo_enable;
   `endif


   assign d_ldo_pon_i_int = d_ldo_pon_i_delay & ldo_enable & pwr_vnn_ok & pwr_vccdig_ok;
   assign d_ldo_bypass_i_int = d_ldo_bypass_i_delay & fz_ldo_bypass & pwr_vccdig_ok;

   assign ldo_enabled = d_ldo_pon_i_int | d_ldo_bypass_i_int;

// ============================================================================================================================================== //
// vfb generated by triming ldo_out vccpll by signal fb_trim[3:0], just refer to SPEC, if enable signal ta_ldo_hiz_debug = 1, got anadft_ldovfb.  //
// When fz_ldo_extrefsel = 1, vref came from ldo_vref, then enable signal ta_ldo_hiz_debug = 1, got anadft_ldovref; When fz_ldo_extrefsel = 0,    //
// vref came from vref_int which generated by triming vccldo by signal ref_trim[3:0], just refer to SPEC, if enable signal ta_ldo_hiz_debug = 1,  // 
// got anadft_ldovfb.															     //
// ============================================================================================================================================== //
// DFT feature
   assign debugen = pwr_vnn_ok ? ta_ldo_hiz_debug : 1'b0;
   assign anadft_ldovfb = ldo_enabled ? (debugen ? 1'b1 : 1'b0) : 1'b0;
   assign anadft_ldovref = debugen ? vref_int : 1'b0;
//`ifndef ip2211ringpll_INTC_NO_PWR_PINS
//   assign analog_debug_out_o = ta_ldo_hiz_debug ? (ta_ldo_idp_debug == 0 ? vccpll :  : 1'bz;
   assign analog_debug_out_o = ta_ldo_hiz_debug ? (ta_ldo_idq_debug == 0 ? anadft_ldovfb : (ldo_enabled & powergood_vnn)) : 1'bz;
   assign viewana = analog_debug_out_o;


// Output assignment
`ifndef ip2211ringpll_INTC_NO_PWR_PINS
    `ifdef SFE_BMOD_ANA_USE_REAL
	assign vccpll_int = ldo_enabled ? (ldo_vref_ok ? vccpll_real : 0.0) : 0.0 ;

    `else
	assign vccpll_int = ldo_enabled ? ldo_vref_ok : 1'b0 ;


    `endif  // end of `ifdef SFE_BMOD_PWR_USE_REAL

`endif  // end of `ifndef ip2211ringpll_INTC_NO_PWR_PINS


`ifdef INTEL_SIMONLY
`ifndef ip2211ringpll_INTC_NO_PWR_PINS 
  `ifdef SFE_BMOD_ANA_USE_REAL
	always @ (vccpll_int)
    	begin
    	    if(vccpll_int == 0)
    	        assign del =  OUTDELAY_FALL;
    	    else
    	        assign del =  OUTDELAY_RISE;
    	end

	always_comb  vccpll <= #(del*1us) (supply_ok == 1'b1) ? vccpll_int : `wrealZState ;

  `else
	always @ (vccpll_int)
    	begin
    	    if(vccpll_int == 1'b0)
    	        #(OUTDELAY_FALL*1us) vccpll = supply_ok ? vccpll_int : 1'bz ;
    	    else
    	        #(OUTDELAY_RISE*1us) vccpll = supply_ok ? vccpll_int : 1'bz ;
    	end

	//if (vccpll_int != 1'b0) #(OUTDELAY_RISE*1us) vccpll = supply_ok ? vccpll_int : 1'bz ;
        //else                    #(OUTDELAY_FALL*1us) vccpll = supply_ok ? vccpll_int : 1'bz ;
  `endif
  `endif

`else  // emulation mode

    //if (vccpll_int != 1'b0) vccpll = supply_ok ? vccpll_int : 1'bz ;
    //else                    vccpll = supply_ok ? vccpll_int : 1'bz ;

	assign vccpll = supply_ok ? vccpll_int : 1'bz ;

`endif


endmodule // ip2211ringpll_ldopgd

`endif //  `ifndef ip2211ringpll_ldopgd_sv
//`endcelldefine




/*

//`ifndef PWRPINS
//supply1  vccdig,
//         vccldo;
//supply0  vss;
//`endif

   logic d_ldo_pon_i_delay;
   logic d_ldo_bypass_i_delay;

   logic d_ldo_pon_i_int;
   logic d_ldo_bypass_i_int;

   logic ldo_enabled;
   
   logic debugen;
   logic vref;
   logic vref_int;
   logic en_1p24;
   logic analog_debug_out_o;
//   assign anadft_ldovref = 1'b0;
//   assign anadft_ldovfb = 1'b0;
   assign debugen = powergood_vnn ? ta_ldo_hiz_debug : 1'b0;
   assign vref    = fz_ldo_extrefsel ? ldo_vref : vref_int;
   assign en_1p24 = powergood_vnn ? ~fz_ldo_vinvoltsel[0] : 1'b0;

   `ifdef INTEL_EMULATION
   assign d_ldo_pon_i_delay = ldo_enable;
   `else 
   assign #500ps  d_ldo_pon_i_delay = ldo_enable;
   `endif 

   //assign d_ldo_pon_i_int = d_ldo_pon_i_delay & ldo_enable;
   assign d_ldo_pon_i_int = d_ldo_pon_i_delay & ldo_enable & powergood_vnn;

   `ifdef INTEL_EMULATION
      assign  d_ldo_bypass_i_delay = fz_ldo_bypass;
   `else
      assign #50ps  d_ldo_bypass_i_delay = fz_ldo_bypass;
   `endif

   assign d_ldo_bypass_i_int = d_ldo_bypass_i_delay & fz_ldo_bypass;

   assign ldo_enabled = d_ldo_pon_i_int | d_ldo_bypass_i_int;
  
   assign vref_int = (ldo_enabled & en_1p24) ? 1'b1 : 1'b0;
   // ============================================================================================================================================== //
   // vfb generated by triming ldo_out vccpll by signal fb_trim[3:0], just refer to SPEC, if enable signal ta_ldo_hiz_debug = 1, got anadft_ldovfb.  //
   // When fz_ldo_extrefsel = 1, vref came from ldo_vref, then enable signal ta_ldo_hiz_debug = 1, got anadft_ldovref; When fz_ldo_extrefsel = 0,    //
   // vref came from vref_int which generated by triming vccldo by signal ref_trim[3:0], just refer to SPEC, if enable signal ta_ldo_hiz_debug = 1,  // 
   // got anadft_ldovfb.															     //
   // ============================================================================================================================================== //
   assign anadft_ldovfb = ldo_enabled ? (debugen ? 1'b1 : 1'b0) : 1'b0;
   assign anadft_ldovref = debugen ? vref : 1'b0;
//`ifndef ip2211ringpll_INTC_NO_PWR_PINS
//   assign analog_debug_out_o = ta_ldo_hiz_debug ? (ta_ldo_idp_debug == 0 ? vccpll :  : 1'bz;
   assign analog_debug_out_o = ta_ldo_hiz_debug ? (ta_ldo_idq_debug == 0 ? anadft_ldovfb : (ldo_enabled & powergood_vnn)) : 1'bz;
   assign viewana = analog_debug_out_o;

/// -----\/----- EXCLUDED -----\/-----
//
//   bit sampleclk;
//   longint sampleclk_period;
//
//   initial begin
//      sampleclk_period = 1000;//1GHz   
//      sampleclk = 1;
//      forever begin
//	 #(sampleclk_period/2) sampleclk = ~sampleclk;
//	 #(sampleclk_period-(sampleclk_period/2)) sampleclk = ~sampleclk;
//      end
//   end
//
//    real  VoltageIn, Ires, VoltageOut;
//   
//   always @(posedge sampleclk or ldo_enable) begin
//       if (ldo_enable == 1'b0) begin 
//	  VoltageIn = 0;
//       end
//       else begin
//	  VoltageIn = 1.0;
//       end
//   end
//  
//   always @(posedge sampleclk or ldo_enable) begin
//       if (ldo_enable == 1'b0) begin 
//	  Ires = 0;
//       end
//       else begin
//	  Ires = (VoltageIn - VoltageOut) / 1e3;
//       end
//   end
//
//   always @(posedge sampleclk or ldo_enable) begin
//       if (ldo_enable == 1'b0) begin 
//	  VoltageOut = 0;
//       end
//       else begin
//	  VoltageOut = VoltageOut + Ires / 1e-6;      
//       end
//   end
// -----/\----- EXCLUDED -----/\----- */
//
//endmodule // ip2211ringpll_ldopgd
//
//`endif //  `ifndef ip2211ringpll_ldopgd_sv
//`endcelldefine
//
//*/
//`endcelldefine


`ifdef INTC_SYNTHESIS
`define ip2211ringpll_SVA_OFF 
`define ip2211ringpll_SVA_LIB_SVA2005 
`define ip2211ringpll_NO_VCSSIM
`endif


`ifndef ip2211ringpll_LOCK_DETECTOR_SV
`define ip2211ringpll_LOCK_DETECTOR_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "ringpll_macros.sv"
//`include "ljpll_dfx.vh"

module ip2211ringpll_lock_detector (

   // DFX settings
   //
   //input  t_ljpll_dfx_in_ifc dfx_in,
   input logic 				fz_lockforce,
   input logic [2:0]                    fz_lockcnt,

   // functional inputs
   //
   input  logic ClkRefXXH,
   input  logic dfx__openloop,
   input  logic dfx__GlobalAlignXXL,
   input  logic pll_core__PfdLockRstNnnnH,
   input  logic reset_sync__Reset_b_XXnnnL,
   input  logic reset_sync__BypassXXnnnL,
   input  logic reset_sync__BypassEnXXnnnL,
   input  logic startup_gen__PfdEnXXH,
   input  logic tlctrl_sip__LockRstXXnnnH,
   output logic lock_detector__RawLockXXnnnL,
   output logic lock_detector__EarlyLockXXnnnH,
   output logic LockXXnnnL,

   input   logic                         idfx_fscan_rstbypen,
   input   logic                         idfx_fscan_clkungate,
   input   logic                         idfx_fscan_byprstb


);

///========================================================================================================
/// Module Begin
///========================================================================================================

   //=============================================================================
   // Lock Counter
   //
   //  The lock counter acts as a digital filter for the PLL lock indicator. The 
   //  counter gets reset by the ip2211ringpll_PFD while the PLL acquires phase/frequency
   //  alignment. Once the phase error is stable within a specified threshold, 
   //  the counter is allowed to count. When the counter saturates we declare
   //  the PLL locked by asserting the "lock" signal. The counter also provides
   //  an early indication that the phase error is stable called "EarlyLockXXnnnH".
   //
   //               Lock Clock Divider and Counter Saturation Values
   //
   //                      lockcnt  |    Lock   | Early Lock
   //                       [2:0]   |  (cntclk) |  (cntclk)  
   //                    ------------------------------------
   //                        000    |     16    |     8
   //                        001    |     24    |     8
   //                        010    |     32    |     8
   //                        011    |     40    |     8
   //                        100    |     48    |     8
   //                        101    |     56    |     8
   //                        110    |     60    |     8
   //                        111    |     63    |     8
   //
   //=============================================================================
 
   logic       ResetXXnnnL;
//   logic       ResetXXnnnL_pre;
  
   logic       PfdLockRstNH;

   logic       ClkRefXXH_b;
   logic       ClkLockCntXXH;
   logic [5:0] LockCntValXXnnnH;

   logic       RawLockNnnnL;
   logic       LockCntRstNnnnH;
   logic       LockCntRstNnnnH_pre;
   logic       StkyLockCntRstNnnnH;
   logic       StkyLockCntRstNnnnH_pre;
   logic       LockCntTripXXnnnH;

   logic       PllLockXXnnnL;
   logic       PllEarlyLockXXnnnH;
  
   // Create inverted clock for use downstream
   //
   `ip2211ringpll_CLKINV(ClkRefXXH_b, ClkRefXXH)

   // Create a positive polarity reset
   //
   always_comb begin : RESET_GEN

      ResetXXnnnL = ~reset_sync__Reset_b_XXnnnL;

   end : RESET_GEN

   always_comb begin : LOCK_TRIP_AND_RESET

      // Determine when to trip the Lock Done indicator based on the
      //  lock count configuration control
      //
      unique casez (fz_lockcnt)
         3'b000 : LockCntTripXXnnnH =   LockCntValXXnnnH[4];                        // Count = 16
         3'b001 : LockCntTripXXnnnH =  &LockCntValXXnnnH[4:3];                      // Count = 24
         3'b010 : LockCntTripXXnnnH =   LockCntValXXnnnH[5];                        // Count = 32
         3'b011 : LockCntTripXXnnnH =  &{LockCntValXXnnnH[5],LockCntValXXnnnH[3]};  // Count = 40
         3'b100 : LockCntTripXXnnnH =  &LockCntValXXnnnH[5:4];                      // Count = 48
         3'b101 : LockCntTripXXnnnH =  &LockCntValXXnnnH[5:3];                      // Count = 56
         3'b110 : LockCntTripXXnnnH =  &LockCntValXXnnnH[5:2];                      // Count = 60
         3'b111 : LockCntTripXXnnnH =  &LockCntValXXnnnH[5:0];                      // Count = 63
         `ip2211ringpll_XDefault(LockCntTripXXnnnH)
      endcase
 
      // Force the lock reset to 0 until sticky lock asserts when tie
      //    lockrst zero asserts.
      //
      //PfdLockRstNH = (dfx_in.fuse.tie_lockrst_zero & !LockXXnnnL) ? 1'b0
      PfdLockRstNH = (fz_lockforce & !LockXXnnnL) ? 1'b0
                                                                  : pll_core__PfdLockRstNnnnH ;

      // Lock Reset Logic
      //  Reset the lock counter during startup, openloop mode, a yank
      //  condition, or when the PLL is disabled. Also reset the lock
      //  counter if the phase error between the reference and feedback
      //  clocks exceeds the specified threshold (given by 
      //  "pfdlockrst".) Finally, provide an external reset input
      //  that could be used to reset the lock counter under other
      //  conditions, like during a ratio change for example.
      //
      LockCntRstNnnnH_pre = ResetXXnnnL | dfx__openloop | PfdLockRstNH | ~startup_gen__PfdEnXXH | tlctrl_sip__LockRstXXnnnH;

      StkyLockCntRstNnnnH_pre = ResetXXnnnL | tlctrl_sip__LockRstXXnnnH;

   end : LOCK_TRIP_AND_RESET

   // Counter state is ASYNC reset so that short reset pulses from the ip2211ringpll_PFD
   //  can reset the state
   //
   `ip2211ringpll_ASYNC_RST_MSFF(LockCntValXXnnnH, (LockCntValXXnnnH + 6'h1), ClkLockCntXXH, LockCntRstNnnnH)
 //Changes done for scan 
assign LockCntRstNnnnH =  idfx_fscan_rstbypen ? ~idfx_fscan_byprstb : LockCntRstNnnnH_pre;


 
   // Latch the count trip condition to use as the count done indicator and
   //  the counter clock enable
   //
   `ip2211ringpll_LATCH_P(RawLockNnnnL, LockCntTripXXnnnH, ClkRefXXH)

   // Note that this gate is controlled by lock which is OK only if
   //  LockCntTrip does not use LockCntValXXnnnH[0] since the counter will
   //  count 1 extra cycle in order to assert the sticky lock bit
   //
//idfx_fscan_clkungate change added for scan
   `ip2211ringpll_CLKAND(ClkLockCntXXH, ClkRefXXH, (~RawLockNnnnL || idfx_fscan_clkungate))

   // Metaflop rawlock so that it is not metastable if the ip2211ringpll_PFD lock reset
   //  asserts
   //
   `ip2211ringpll_ASYNC_RST_2MSFF_META(lock_detector__RawLockXXnnnL, RawLockNnnnL, ClkRefXXH_b, reset_sync__Reset_b_XXnnnL)

   // Generate a sticky lock indicator when the counter trips
   //
   `ip2211ringpll_ASYNC_RST_MSFF_P(PllLockXXnnnL, (~dfx__GlobalAlignXXL & (lock_detector__RawLockXXnnnL || PllLockXXnnnL)), ClkRefXXH, ResetXXnnnL)

//assign ResetXXnnnL =  idfx_fscan_rstbypen ? ~idfx_fscan_byprstb : ResetXXnnnL_pre;


   // Generate a sticky early-lock indicator when the lock counter hits 0x8
   //
   `ip2211ringpll_ASYNC_RST_MSFF(PllEarlyLockXXnnnH, (LockCntValXXnnnH[3] || PllEarlyLockXXnnnH), ClkLockCntXXH, StkyLockCntRstNnnnH)
  
 //Changes done for scan 
assign StkyLockCntRstNnnnH =  idfx_fscan_rstbypen ? ~idfx_fscan_byprstb : StkyLockCntRstNnnnH_pre;
 
   // Override the lock in bypass mode
   //   The lock signal is based on bypass enable when in bypass mode
   //   Else, lock is based on the actual PLL lock
   //
   always_comb begin : LOCK_GEN
      LockXXnnnL =      (reset_sync__BypassXXnnnL) ? reset_sync__BypassEnXXnnnL
                                                   : PllLockXXnnnL                       ;
      lock_detector__EarlyLockXXnnnH = (reset_sync__BypassXXnnnL) ? reset_sync__BypassEnXXnnnL
                                                                  : (PllEarlyLockXXnnnH) ;
   end : LOCK_GEN

///========================================================================================================
/// Module End
///========================================================================================================

endmodule

`endif

`ifndef ip2211ringpll_LOCK_TIMER_SV
`define ip2211ringpll_LOCK_TIMER_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "ringpll_macros.sv"

module ip2211ringpll_lock_timer #(parameter LOCKCNT_WIDTH = 12) (
   input  logic ClkRefXXH,
   input  logic reset_sync__Reset_b_XXnnnL,
   input  logic LockXXnnnL,
   output logic [LOCKCNT_WIDTH - 1 : 0] lock_timer__LockTimeCntXXnnnH,
   input   logic                         idfx_fscan_clkungate
//   input   logic                         idfx_fscan_rstbypen,
//   input   logic                         idfx_fscan_byprstb
);

///========================================================================================================
/// Module Begin
///========================================================================================================

   logic ClkLockCntXXH;
   logic CountSatXXnnnH;
   logic CountSatXXnnnL;
   logic ResetXXnnnL;
//   logic ResetXXnnnL_pre;
   
   // Create a positive polarity reset
   //
   always_comb begin : RESET_GEN

      ResetXXnnnL = ~reset_sync__Reset_b_XXnnnL;

   end : RESET_GEN

   // Lock counter flops
   //   Counts up until lock is asserted.  Counter is reset by inverted
   //   global reset_b
   //
   `ip2211ringpll_ASYNC_RST_MSFF(lock_timer__LockTimeCntXXnnnH, (lock_timer__LockTimeCntXXnnnH + `ip2211ringpll_ZX(1'b1,LOCKCNT_WIDTH)), ClkLockCntXXH, ResetXXnnnL)

//assign ResetXXnnnL = idfx_fscan_rstbypen ? ~idfx_fscan_byprstb : ResetXXnnnL_pre;

   // Counter Saturation Logic
   //
   always_comb begin: COUNT_SAT
      CountSatXXnnnH = (lock_timer__LockTimeCntXXnnnH == '1);
   end : COUNT_SAT

   // Counter sat latch for clock gate
   //
   `ip2211ringpll_LATCH_P(CountSatXXnnnL, CountSatXXnnnH, ClkRefXXH)

   // Lock signal will come in on low phase of ClkRefXXH
   //   The lock signal is sticky so does not need to be syncronized
   //
//idfx_fscan_clkungate change added for scan
   `ip2211ringpll_CLKAND(ClkLockCntXXH, ClkRefXXH, ((~LockXXnnnL & reset_sync__Reset_b_XXnnnL & ~CountSatXXnnnL) || idfx_fscan_clkungate))


endmodule

`endif

`ifndef ip2211ringpll_UNLOCK_COUNTER_SV
`define ip2211ringpll_UNLOCK_COUNTER_SV

`ifndef ip2211ringpll_SVA_OFF
//`include "intel_checkers.vs"
`endif
//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "ringpll_macros.sv"

module ip2211ringpll_unlock_counter #(parameter UNLOCK_COUNT_BITS = 2) (
   input  logic                            ClkRefXXH,
   input  logic                            reset_sync__Reset_b_XXnnnL,

   input  logic                            LockXXnnnL,
   input  logic                            lock_detector__RawLockXXnnnL,
   input  logic                            idfx_fscan_clkungate,

   output logic [UNLOCK_COUNT_BITS - 1 :0] unlock_counter__UnlockCountXXnnnH
);


   logic UnlockXXnn0L, UnlockXXnn1L;

   logic CounterSatXXnnnH;
   logic CounterSatXXnnnL;

   logic UnlockClkEnXXnnnL;
   logic ClkUnlockXXH;

   logic ResetXXnnnL;

   always_comb begin : RESET_GEN

      ResetXXnnnL = ~reset_sync__Reset_b_XXnnnL;

   end : RESET_GEN

   // Unlock detector circuit
   //   Edge detect an unlock to enable the counter
   //   An unlock is defined as sticky lock asserted and rawlock deasserted
   //
   `ip2211ringpll_ASYNC_RST_MSFF_P(UnlockXXnn0L, (LockXXnnnL & ~lock_detector__RawLockXXnnnL), ClkRefXXH, ResetXXnnnL)
   `ip2211ringpll_ASYNC_RST_MSFF_P(UnlockXXnn1L,                     UnlockXXnn0L, ClkRefXXH, ResetXXnnnL)

   // Detect Unlock signal assertion
   //
   always_comb begin : UNLOCK_ASSERTION_DETECT

      UnlockClkEnXXnnnL = UnlockXXnn0L & ~UnlockXXnn1L;

   end : UNLOCK_ASSERTION_DETECT

   // Unlock Counter Flops
   //  Counts up when an unlock is detected and the counter is not saturated
   //
   `ip2211ringpll_ASYNC_RST_MSFF(unlock_counter__UnlockCountXXnnnH, (unlock_counter__UnlockCountXXnnnH + `ip2211ringpll_ZX(1'b1, UNLOCK_COUNT_BITS)), ClkUnlockXXH, ResetXXnnnL)

   // Detect Counter Saturation
   //
   always_comb begin : COUNTER_SAT

      CounterSatXXnnnH = (unlock_counter__UnlockCountXXnnnH == '1);

   end : COUNTER_SAT

   // Latch saturation signal to low phase
   //
   `ip2211ringpll_LATCH_P(CounterSatXXnnnL, CounterSatXXnnnH, ClkRefXXH)

   // Lock signal and rawlock signal are both low phase signals
   //
//idfx_fscan_clkungate change added for scan
   `ip2211ringpll_CLKAND(ClkUnlockXXH, ClkRefXXH, ((UnlockClkEnXXnnnL & ~CounterSatXXnnnL) || idfx_fscan_clkungate) )

///========================================================================================================
/// Assertions
///========================================================================================================

   `ifndef ip2211ringpll_SVA_OFF
      `ip2211ringpll_ASSERTC_FORBIDDEN(R_unlock_counter_nonzero, (|unlock_counter__UnlockCountXXnnnH), ResetXXnnnL, `ip2211ringpll_ERR_MSG("[LJPLL] Unlock counter is >0 which means the PLL has unlocked!"));
   `endif

endmodule

`endif

`ifndef ip2211ringpll_LJPLL_DFX_SV
`define ip2211ringpll_LJPLL_DFX_SV

//`include "ljpll_dfx.vh"
//`include "ringpll_macros.sv"

module ip2211ringpll_ljpll_dfx 
//#(parameter RATIO_BITS = 10, parameter FRAC_BITS = 24, parameter FMOD_BITS = 9) 
(
   // Fuse/View Input
   //
   //input  t_ljpll_dfx_in_ifc         dfx_in,
   
   // View Output
   //
   output t_ljpll_dfx_out_ifc        dfx_out,

   // Accommodate RTDR - dfx - to SIP programming for TAP bits.
   input  t_ljpll_tap_in_ifc       tap_in,
   output t_ljpll_tap_out_ifc      tap_out,

  
   // Non-Override Values (LJPLL Inputs)
   //
   input  logic                      Reset_b_NnnnH,
   input  logic                      PllDistPwrGoodNnnnH,
   input  logic                      BypassNnnnH,
   input  logic [9:0] 		     RatioNnnnH,
   input  logic [23:0] 		     FractionNnnnH,
   
   input  logic [1:0]                unlock_counter__UnlockCountXXnnnH,
   input  logic [11:0]               lock_timer__LockTimeCntXXnnnH,
   input  logic                      lock_detector__RawLockXXnnnL,
   input  logic [1:0]                tlctrl_sip__StateXXnnnH,                                                            
   input  logic [9:0]                view_adc__dig_out,
   input  logic                      adc_ctl__StartXXH,
   input  logic                      view_adc__done,

   // ODCS signals from HIP
   //
   //input  logic                        odcs_dig__odcsrisetrig,
   //input  logic                        odcs_dig__odcsfalltrig,
   //input  logic [4:0]                  odcs_dll__DlyLineSettingNH,
   //input  logic                        stm_ifdim__StmTrigStatusNH,
   //input  logic                        odcs_opsp__RiseSampNH,
   //input  logic                        odcs_opsp__FallSampNH,

   // Lock signal for low power charge pump enable and status
   //
   input  logic                        LockXXnnnL,

   input  logic [9:0]   		mash__RatioMXH,
   input  logic                        mash__HalfIntMXH,
   
   input  logic                        ssc_mod_dfx__TriggerRegXDH,
   input  logic                        ssc_mod_dfx__ModulatorEnNH,

   input  logic                        iref_ctrl__IrefDoneXXH,
   input  logic                        startup_gen__PfdEnXXH,

   input  logic [14:0]                 view_freq_count,

   // Enable signal for tap out encode
   //
   input  logic                        reset_sync__Reset_b_XXnnnL,

   // Tap in decode
   //
   output logic                                     dfx__openloop,
   output logic [1:0]                               dfx__ViewDigEnNnnnH,
   output logic [1:0]                               dfx__ViewAnaEnNnnnH,
   output logic [1:0] [4:0]                         dfx__ViewSelNnnnH,
   output logic [1:0]                               dfx__adc_clkdiv,
   output logic					    dfx__adc_start,
   output logic [1:0]				    dfx__adc_start_cnt,
   output logic                                     dfx__adc_freeze,
   output logic                                     dfx__adc_chop_en,
   output logic                                     dfx__adc_use_vref,
   output logic [2:0]                               dfx__adc_sel_in,
   //output t_opsp_config                             dfx__opsp_config,
   //output logic [1:0]                               dfx__odcs_tuner_cb,
   output logic                                     dfx__GlobalAlignXXL,
  
   // IDV encode/decode
   //
   input  t_ljpll_idv_out_ifc                       idv_fub__idv_out,

   // Fuse decode to SIP
   //
   output logic                                     dfx__disable_run_upd,
   output logic                                     dfx__mash_order_plus_one,
   output logic                                     dfx__ssc_en,
//   output logic [1:0]                               dfx__ssc_mode,
//   output logic [2:0]                               dfx__cp_mode,
//   output logic                                     dfx__lp_cp_en,
//   output logic [1:0]                               dfx__lpf_itrim,
//   output logic [1:0]                               dfx__sr_lpf_mode,
//   output logic [3:0]                               dfx__startup_rdac,
   //output logic [3:0]                               dfx__vco_trim_pg,
   //output logic [2:0]                               dfx__vco_trim_cb,
//   output logic [2:0]                               dfx__iref_mode,
//   output logic [2:0]                               dfx__startcnt,
   output logic                                     dfx__SscModTrigNH,
   output logic  [1:0]                              dfx__SscModStepsNH,
   output logic                                     dfx__SscDfxEnNH,
   output logic  [1:0]                              dfx__SscModClkDivNH,
//   output logic                                     dfx__start_mode,

   // Fuse decode to HIP
   //
   output logic                                     dfx__tight_loop,
//   output logic                                     dfx__pfd_chop_en, 
//   output logic [2:0]                               dfx__pfd_chop_val, 
//   output logic [1:0]                               dfx__pvd_mode, 
   output logic [2:0]                               dfx__pfd_residual_pw,
   output logic [4:0]                               dfx__cp1_trim,
   output logic [4:0]                               dfx__cp2_trim,
   output logic [4:0]                               dfx__skadj_ctrl,
   output logic [3:0]                               dfx__lockthresh,
   output logic                                     dfx__lockstickyb,
//   output logic [2:0]                               dfx__iref_ctune,
//   output logic [3:0]                               dfx__iref_ftune,
//   output logic [3:0]                               dfx__ro_freq_sel,
   output logic [5:0]                               dfx__dca_ctrl,
   output logic [1:0]                               dfx__dca_cb,
   output logic                                     dfx__tllm_en,   // new -nd Using fz_spare[3]
  
   // Register decode to ip2211ringpll_ssc_mod
   //
   //output logic [9:0]                    dfx__RatioStepNH,
   output logic [23:0]                     dfx__FracStepNH,
   output logic [8:0]                     dfx__ssc_cyc_to_peak_m1,

   // Req/Ack to/from Ratio sync
   //
   output logic                                    dfx__ratio_update_req,
   input  logic                                    reg_req_ack__RatioUpdAckMXH,

   // Req/Ack to/from SSC modulator
   //
   output logic                                     dfx__ssc_prof_update_req,
   input  logic                                     reg_req_ack__SscProfUpdAckMXH,

   // View Pins In
   //
   input  logic [1:0]                               view_mux__ViewOutNnnnH,
   
//--------------------------------------------------------------------------
   // Brought these in for over writing via TAP
   //
input  logic [4:0]                     fz_cp1trim,             // Part of DFX_IN bus
input  logic [4:0]                     fz_cp2trim,             // Part of DFX_IN bus
input  logic [1:0]                     fz_cpnbias,        //NEW fuse: CP nbias tuning				// part of dfx_in
input  logic [1:0]                     fz_dca_cb,              // Part of DFX_IN bus
input  logic [5:0]                     fz_dca_ctrl,            // Part of DFX_IN bus
input  logic [4:0]                     fz_irefgen,    //NEW fuse: Iref current				// part of dfx_in
input  logic [2:0]                     fz_lockcnt,           // Part of DFX_IN bus
input  logic                           fz_lockforce,         // Part of DFX_IN bus
input  logic                           fz_lockstickyb,         // Part of DFX_IN bus
input  logic [3:0]                     fz_lockthresh,          // Part of DFX_IN bus
input  logic                           fz_lpfclksel,      //NEW fuse: LPF clock selection				// part of dfx_in
input  logic                           fz_nopfdpwrgate,   //NEW fuse: Disable ip2211ringpll_PFD power gating				// part of dfx_in
input  logic [2:0]                     fz_pfd_pw,              // Part of DFX_IN bus
input  logic [1:0]                     fz_pfddly,         //NEW fuse: ip2211ringpll_PFD power gating delay section				// part of dfx_in
input  logic [4:0]                     fz_skadj,               // Part of DFX_IN bus
input  logic [4:0]                     fz_spare,          //NEW fuse: spare bits				// part of dfx_in
input  logic [5:0]                     fz_startup,    //NEW fuse: PLL startup circuit tuning				// part of dfx_in
input  logic                           fz_tight_loopb,         // Part of DFX_IN bus
input  logic			       fz_vcosel,
input  logic [10:0]                    fz_vcotrim,        //NEW fuse: ip2211ringpll_VCO trim				// part of dfx_in
input  logic [1:0]                   fz_ldo_vinvoltsel,      //new -nd				// part of dfx_in
input  logic                         fz_ldo_bypass,          //new -nd				// part of dfx_in
input  logic                         fz_ldo_extrefsel,       //new -nd				// part of dfx_in
input  logic                         fz_ldo_faststart,       //new -nd				// part of dfx_in
input  logic [3:0]                   fz_ldo_fbtrim,          //new -nd				// part of dfx_in
input  logic [3:0]                   fz_ldo_reftrim,         //new -nd				// part of dfx_in
 input  logic                           mash_order_plus_one,    // Part of DFX_IN bus
 input  logic [8:0]                     ssc_cyc_to_peak_m1,         // Part of DFX_IN bus
 input  logic                           ssc_en,                 // Part of DFX_IN bus
 input  logic [23:0]                    ssc_frac_step,          // Part of DFX_IN bus


   input  logic                         ldo_enable,             //new -nd
   input  logic [5:0]                   mdiv_ratio,             //new -nd
   input  logic [1:0]                   vcodiv_ratio,           //new -nd
   input  logic [9:0]                   zdiv0_ratio,            //new -nd
   input  logic                         zdiv0_ratio_p5,         //new -nd
   input  logic [9:0]                   zdiv1_ratio,            //new -nd
   input  logic                         zdiv1_ratio_p5,         //new -nd
          // IDV interface
//   input  logic                         idvdisable_bi,          // new -nd
//   input  logic                         idvfreqai,              // new -nd
//   input  logic                         idvfreqbi,              // new -nd
//   input  logic                         idvpulsei,              // new -nd
//   input  logic                         idvvtclki,              // new -nd
//   input  logic                         idvvtctrli,             // new -nd
//   input  logic                         idvtdi,                 // new -nd
//   input  logic                         idvtresi,               // new -nd
//   input  logic                         clkidvih,               // new -nd
//   input  logic                         pllen,                  // new -nd  // same as Reset_b_NnnnH

   output logic                         dfx__ldo_enable_a,           // new -nd
   output logic                         dfx__ta_ldo_hiz_debug,       // new -nd
   output logic                         dfx__ta_ldo_idq_debug,       // new -nd
   output logic [4:0]                   dfx__ta_spare,       	     // new -nd
   output logic [3:0]			dfx__ta_vctlrdac,	     // new -nd
   output logic				dfx__ta_openloop2,	     // new -nd
   output logic [1:0]                   dfx__fz_ldo_vinvoltsel_a,    // new -nd
   output logic                         dfx__fz_ldo_bypass_a,        // new -nd
   output logic                         dfx__fz_ldo_extrefsel_a,     // new -nd
   output logic                         dfx__fz_ldo_faststart_a,     // new -nd
   output logic [3:0]                   dfx__fz_ldo_fbtrim_a,        // new -nd
   output logic [3:0]                   dfx__fz_ldo_reftrim_a,       // new -nd
   output logic [5:0]                   dfx__mdiv_ratio_a,           // new -nd
   output logic [1:0]                   dfx__vcodiv_ratio_a,         // new -nd
   output logic [9:0]                   dfx__zdiv0_ratio_a,          //new -nd
   output logic                         dfx__zdiv0_ratio_p5_a,       //new -nd
   output logic [9:0]                   dfx__zdiv1_ratio_a,          //new -nd
   output logic                         dfx__zdiv1_ratio_p5_a,       //new -nd
   output logic [1:0]                   dfx__cpnbias,           //new -nd
   output logic [4:0]                   dfx__fz_irefgen_a,           //new -nd
   output  logic                        dfx__fz_lpfclksel_a,         //new -nd
   output  logic                        dfx__fz_nopfdpwrgate_a,      //new -nd
   output  logic [2:0]                  dfx__fz_pfd_pw_a,            //new -nd
   output  logic [1:0]                  dfx__fz_pfddly_a,            //new -nd
   output  logic [4:0]                  dfx__fz_spare_a,             //new -nd
   output  logic [5:0]                  dfx__fz_startup_a,           //new -nd
   output  logic                        dfx__fz_vcosel_a,            //new -nd
   output  logic                        dfx__fz_lockforce_a,         //new -nd
   output  logic [2:0]                  dfx__fz_lockcnt_a,           //new -nd
   output  logic [10:0]                 dfx__fz_vcotrim_a,           //new -nd
   output  logic			dfx__start_measurement,	     //new -nd
//--------------------------------------------------------------------------

   // Post-Mux Outputs
   //
   output logic                         dfx__reset_b,
   output logic                         dfx__powergood,
   output logic                         dfx__bypass,
   output logic [9:0]                   dfx__ratio,
   output logic [23:0]                  dfx__fraction
);

///========================================================================================================
/// Module Begin
///========================================================================================================
   logic 		    dfx__fuseoverride;
//   logic [9:0]              ovrd_misc_cfg;            // SPARES! -- these are spare fuse bits routed to the HIP
//   logic                    ovrd_disable_run_upd;     // Disable SSC/ratio runtime updates. When this bit is set, all SSC reg writes are rejected after PLL lock.
   logic                    ovrd_tight_loop;          // Tight Loop Select Bit (optional as a fuse for tight loop only PLLs)
//   logic                    ovrd_tie_lockrst_zero;    // Force the lock reset to 0 until after sticky lock asserts
   logic                    ovrd_lockstickyb;         // 
//   logic [3:0]              ovrd_startup_rdac;        // Startup RDAC setting
//   logic [2:0]              ovrd_pfd_chop_val;        // ip2211ringpll_PFD chop value
   logic [2:0]              ovrd_pfd_residual_pw;     // ip2211ringpll_PFD residual pulse width
   logic [4:0]              ovrd_cp1_trim;            // Charge pump 1 trim
   logic [4:0]              ovrd_cp2_trim;            // Charge pump 2 trim
   logic [4:0]              ovrd_skadj_ctrl;          // Skew Adjust Control
//   logic [2:0]              ovrd_lockcnt;             // lock count before lock assert
//   logic [2:0]              ovrd_startcnt;            // iref ramp time counter
   logic [3:0]              ovrd_lockthresh;          // lock threshold setting to AIP
//   logic [2:0]              ovrd_iref_ctune;          // IREF course tune bits
//   logic [3:0]              ovrd_iref_ftune;          // IREF fine tune bits
   logic                    ovrd_mash_order_plus_one; // MASH modulator order control
//   logic                    ovrd_lp_cp_en;            // Low power charge pump mode chicken bit
//   logic [1:0]              ovrd_lpf_itrim;           // SR-LPF (internal to AIP) current trim
//   logic [3:0]              ovrd_ro_freq_sel;         // Ring oscillator frequency control
//   logic [2:0]              ovrd_iref_mode;           // IREF operating mode
//   logic [2:0]              ovrd_cp_mode;             // CP operating mode
//   logic [1:0]              ovrd_sr_lpf_mode;         // SR LPF Mode
   logic [1:0]              ovrd_dca_cb;              // Static DCA capacitor bank control
//   logic                    ovrd_start_mode;          // 2 different start modes 0=parallel iref/vctl pulldn, 1=serial iref 1st, vctl 2nd
//   logic [3:0]              ovrd_vco_trim_pg;         // PG trim
//   logic [2:0]              ovrd_vco_trim_cb;         // CB trim
//   logic [1:0]              ovrd_pvd_mode;            // PVD mode (/1, /2, /4, /8)
   logic                    ovrd_tllm_en;             // tight loop lock mode enable
//   logic                    ovrd_tllm_prchg_mode;     // gate clock distribution during tight loop lock
//   logic [1:0]              ovrd_tllm_sw_latency;     // wait some cycles after distribution ungated before switching to long loop
   logic [5:0]              ovrd_dca_ctrl;            // Static DCA control bits

   // Brought in for overwriting via TAP
   //
   logic [1:0]                   ovrd_fz_cpnbias;        //NEW fuse: CP nbias tuning
   logic [4:0]                   ovrd_fz_irefgen;    //NEW fuse: Iref current
   logic                         ovrd_fz_nopfdpwrgate;   //NEW fuse: Disable ip2211ringpll_PFD power gating
   logic [2:0]			 ovrd_fz_pfd_pw;         // NEW
   logic                         ovrd_fz_lpfclksel;      //NEW fuse: LPF clock selection
   logic [1:0]                   ovrd_fz_pfddly;         //NEW fuse: ip2211ringpll_PFD power gating delay section
   logic [4:0]                   ovrd_fz_spare;          //NEW fuse: spare bits
   logic [5:0]                   ovrd_fz_startup;    //NEW fuse: PLL startup circuit tuning
   logic                         ovrd_fz_vcosel;     // NEW fuse: ip2211ringpll_VCO select
   logic [10:0]                  ovrd_fz_vcotrim;        //NEW fuse: ip2211ringpll_VCO trim

   logic			 ovrd_fz_lockforce;
   logic [2:0]			 ovrd_fz_lockcnt;    // lock count before lock assert

   logic                         ovrd_ldo_enable;             //new -nd
   logic [1:0]                   ovrd_fz_ldo_vinvoltsel;      //new -nd
   logic                         ovrd_fz_ldo_bypass;          //new -nd
   logic                         ovrd_fz_ldo_extrefsel;       //new -nd
   logic                         ovrd_fz_ldo_faststart;       //new -nd
   logic [3:0]                   ovrd_fz_ldo_fbtrim;          //new -nd
   logic [3:0]                   ovrd_fz_ldo_reftrim;         //new -nd
   logic [5:0]                   ovrd_mdiv_ratio;             //new -nd
   logic [1:0]                   ovrd_vcodiv_ratio;           //new -nd
   logic [9:0]                   ovrd_zdiv0_ratio;            //new -nd
   logic                         ovrd_zdiv0_ratio_p5;         //new -nd
   logic [9:0]                   ovrd_zdiv1_ratio;            //new -nd
   logic                         ovrd_zdiv1_ratio_p5;         //new -nd
   // IDV interface
//   logic                         ovrd_idvdisable_bi;          // new -nd
//   logic                         ovrd_idvfreqai;              // new -nd
//   logic                         ovrd_idvfreqbi;              // new -nd
//   logic                         ovrd_idvpulsei;              // new -nd
//   logic                         ovrd_idvvtclki;              // new -nd
//   logic                         ovrd_idvvtctrli;             // new -nd
//   logic                         ovrd_idvtdi;                 // new -nd
//   logic                         ovrd_idvtresi;               // new -nd
//   logic                         ovrd_clkidvih;               // new -nd
//   logic                         ovrd_pllen;                  // new -nd

     logic			dfx__ldo_enable_a_int;        // Internal befor ORing with PLLen
     logic			dfx__fz_ldo_faststart_a_pre;

   logic                    tllm_en;             // tight loop lock mode enable
   assign  tllm_en = fz_spare[3]; // Using a spare fuse as TLLM enable.

   // Register decode to SSC
   //
   //assign dfx__RatioStepNH         = ssc_ratio_step;
   assign dfx__FracStepNH          = ssc_frac_step;
   assign dfx__ssc_cyc_to_peak_m1  = ssc_cyc_to_peak_m1;
   assign dfx__ssc_en              = ssc_en;
   //assign dfx__ssc_mode            = ssc_mode;
  
   // Tap decode to SIP
   //
   assign dfx__fuseoverride        = tap_in.tap_fuseoverride;
   assign dfx__SscDfxEnNH          = tap_in.ssc_mod_dfx_en;
   assign dfx__SscModTrigNH        = tap_in.ssc_mod_dfx_trigger;
   assign dfx__SscModStepsNH       = tap_in.ssc_mod_dfx_steps;
   assign dfx__SscModClkDivNH      = tap_in.ssc_mod_dfx_clkdiv;
   assign dfx__start_measurement   = tap_in.start_measurement;

   // Tap decode to HIP
   //
   assign dfx__openloop            = tap_in.openloop;
   assign dfx__ViewDigEnNnnnH      = tap_in.view_en & ~tap_in.view_ana_en;
   assign dfx__ViewAnaEnNnnnH      = tap_in.view_en &  tap_in.view_ana_en;
   assign dfx__ViewSelNnnnH        = tap_in.view_sel;
   assign dfx__adc_start           = tap_in.adc_start;
   assign dfx__adc_start_cnt       = tap_in.adc_start_cnt; 
   assign dfx__adc_clkdiv          = tap_in.adc_clkdiv;
   assign dfx__adc_freeze          = tap_in.adc_freeze;
   assign dfx__adc_chop_en         = tap_in.adc_chop_en;
   assign dfx__adc_use_vref        = tap_in.adc_use_vref;
   assign dfx__adc_sel_in          = tap_in.adc_sel_in;
   assign dfx__ta_ldo_hiz_debug	   = tap_in.ta_ldo_hiz_debug;
   assign dfx__ta_ldo_idq_debug	   = tap_in.ta_ldo_idq_debug;
   assign dfx__ta_spare		   = tap_in.ta_spare;

   assign dfx__ta_openloop2	   = tap_in.ta_openloop2;
   assign dfx__ta_vctlrdac	   = tap_in.ta_vctlrdac;


   //assign dfx__opsp_config         = dfx_in.tap.opsp_config;
   //assign dfx__odcs_tuner_cb       = dfx_in.tap.odcs_tuner_cb;


//   	assign 	ovrd_misc_cfg 		= tap_in.ovrd_misc_cfg;
//	assign  ovrd_disable_run_upd 	= tap_in.ovrd_disable_run_upd;
	assign	ovrd_tight_loop		= tap_in.ovrd_tight_loop;
//	assign  ovrd_tie_lockrst_zero	= tap_in.ovrd_tie_lockrst_zero;
//	assign 	ovrd_startup_rdac	= tap_in.ovrd_startup_rdac;
//	assign 	ovrd_pfd_chop_val	= tap_in.ovrd_pfd_chop_val;
	assign 	ovrd_pfd_residual_pw	= tap_in.ovrd_pfd_residual_pw;
	assign 	ovrd_cp1_trim		= tap_in.ovrd_cp1_trim;
	assign	ovrd_cp2_trim		= tap_in.ovrd_cp2_trim;
	assign	ovrd_skadj_ctrl		= tap_in.ovrd_skadj_ctrl;
//	assign	ovrd_lockcnt		= tap_in.ovrd_lockcnt;
//	assign	ovrd_startcnt		= tap_in.ovrd_startcnt;
	assign	ovrd_lockthresh		= tap_in.ovrd_lockthresh;
        assign  ovrd_lockstickyb        = tap_in.ovrd_lockstickyb;
//	assign	ovrd_iref_ctune		= tap_in.ovrd_iref_ctune;
//	assign	ovrd_iref_ftune		= tap_in.ovrd_iref_ftune;
	assign	ovrd_mash_order_plus_one = tap_in.ovrd_mash_order_plus_one;
//	assign	ovrd_lp_cp_en		= tap_in.ovrd_lp_cp_en;
//	assign 	ovrd_lpf_itrim		= tap_in.ovrd_lpf_itrim;
//	assign	ovrd_ro_freq_sel	= tap_in.ovrd_ro_freq_sel;
//	assign	ovrd_iref_mode		= tap_in.ovrd_iref_mode;
//	assign	ovrd_cp_mode		= tap_in.ovrd_cp_mode;
//	assign	ovrd_sr_lpf_mode	= tap_in.ovrd_sr_lpf_mode;
	assign	ovrd_dca_cb		= tap_in.ovrd_dca_cb;
//	assign	ovrd_start_mode		= tap_in.ovrd_start_mode;
//	assign	ovrd_vco_trim_pg	= tap_in.ovrd_vco_trim_pg;
//	assign	ovrd_vco_trim_cb	= tap_in.ovrd_vco_trim_cb;
//	assign	ovrd_pvd_mode		= tap_in.ovrd_pvd_mode;
	assign	ovrd_tllm_en		= tap_in.ovrd_tllm_en;
//	assign	ovrd_tllm_prchg_mode	= tap_in.ovrd_tllm_prchg_mode;
//	assign	ovrd_tllm_sw_latency	= tap_in.ovrd_tllm_sw_latency;
	assign	ovrd_dca_ctrl		= tap_in.ovrd_dca_ctrl;
	
	// Brought in here for TAP over write.
	//
	assign  ovrd_fz_lockforce       = tap_in.ovrd_fz_lockforce;
	assign  ovrd_fz_lockcnt		= tap_in.ovrd_fz_lockcnt;

        assign  ovrd_fz_cpnbias		= tap_in.ovrd_fz_cpnbias;        //NEW fuse: CP nbias tuning
        assign  ovrd_fz_irefgen		= tap_in.ovrd_fz_irefgen;    //NEW fuse: Iref current
        assign  ovrd_fz_nopfdpwrgate	= tap_in.ovrd_fz_nopfdpwrgate;   //NEW fuse: Disable ip2211ringpll_PFD power gating
        assign  ovrd_fz_pfd_pw		= tap_in.ovrd_fz_pfd_pw;   //NEW fuse: Disable ip2211ringpll_PFD power gating
        assign  ovrd_fz_lpfclksel	= tap_in.ovrd_fz_lpfclksel;      //NEW fuse: LPF clock selection
        assign  ovrd_fz_pfddly		= tap_in.ovrd_fz_pfddly;         //NEW fuse: ip2211ringpll_PFD power gating delay section
        assign  ovrd_fz_spare		= tap_in.ovrd_fz_spare;          //NEW fuse: spare bits
        assign  ovrd_fz_startup		= tap_in.ovrd_fz_startup;    //NEW fuse: PLL startup circuit tuning
        assign  ovrd_fz_vcosel		= tap_in.ovrd_fz_vcosel;    //NEW fuse: ip2211ringpll_VCO select 
        assign  ovrd_fz_vcotrim		= tap_in.ovrd_fz_vcotrim;        //NEW fuse: ip2211ringpll_VCO trim

        assign  ovrd_ldo_enable		= tap_in.ovrd_ldo_enable;             //new -nd
        assign  ovrd_fz_ldo_vinvoltsel  = tap_in.ovrd_fz_ldo_vinvoltsel;      //new -nd [1:0]
        assign  ovrd_fz_ldo_bypass	= tap_in.ovrd_fz_ldo_bypass;          //new -nd
        assign  ovrd_fz_ldo_extrefsel   = tap_in.ovrd_fz_ldo_extrefsel;       //new -nd
        assign  ovrd_fz_ldo_faststart   = tap_in.ovrd_fz_ldo_faststart;       //new -nd
        assign  ovrd_fz_ldo_fbtrim	= tap_in.ovrd_fz_ldo_fbtrim;          //new -nd [3:0]
        assign  ovrd_fz_ldo_reftrim	= tap_in.ovrd_fz_ldo_reftrim;         //new -nd [3:0]
        assign  ovrd_mdiv_ratio		= tap_in.ovrd_mdiv_ratio;             //new -nd [5:0]
        assign  ovrd_vcodiv_ratio	= tap_in.ovrd_vcodiv_ratio;           //new -nd [1:0]
        assign  ovrd_zdiv0_ratio	= tap_in.ovrd_zdiv0_ratio;            //new -nd [9:0]
        assign  ovrd_zdiv0_ratio_p5	= tap_in.ovrd_zdiv0_ratio_p5;         //new -nd
        assign  ovrd_zdiv1_ratio	= tap_in.ovrd_zdiv1_ratio;            //new -nd [9:0]
        assign  ovrd_zdiv1_ratio_p5	= tap_in.ovrd_zdiv1_ratio_p5;         //new -nd
   		// IDV interface
//        assign  ovrd_idvdisable_bi	= tap_in.ovrd_idvdisable_bi;          // new -nd
//        assign  ovrd_idvfreqai		= tap_in.ovrd_idvfreqai;              // new -nd
//        assign  ovrd_idvfreqbi		= tap_in.ovrd_idvfreqbi;              // new -nd
//        assign  ovrd_idvpulsei		= tap_in.ovrd_idvpulsei;              // new -nd
//        assign  ovrd_idvvtclki		= tap_in.ovrd_idvvtclki;              // new -nd
//        assign  ovrd_idvvtctrli		= tap_in.ovrd_idvvtctrli;             // new -nd
//        assign  ovrd_idvtdi		= tap_in.ovrd_idvtdi;                 // new -nd
//        assign  ovrd_idvtresi		= tap_in.ovrd_idvtresi;               // new -nd
//        assign  ovrd_clkidvih		= tap_in.ovrd_clkidvih;               // new -nd
//        assign  ovrd_pllen		= tap_in.ovrd_pllen;                  // new -nd


   // Global Alignment
   //
   //assign dfx__GlobalAlignXXL      = dfx_in.ip2211ringpll_global_align;
   assign dfx__GlobalAlignXXL      = 1'b0;
   
   // Fuse decode to SIP
   //
   always_comb begin : OVRD_MUX_FUSE_SIP
//
//   dfx__cp_mode             = (dfx__fuseoverride) ? ovrd_cp_mode : dfx_in.fuse.cp_mode;
//   dfx__lp_cp_en            = (dfx__fuseoverride) ? ovrd_lp_cp_en : dfx_in.fuse.lp_cp_en;
//   dfx__lpf_itrim           = (dfx__fuseoverride) ? ovrd_lpf_itrim : dfx_in.fuse.lpf_itrim;
//   dfx__sr_lpf_mode         = (dfx__fuseoverride) ? ovrd_sr_lpf_mode : dfx_in.fuse.sr_lpf_mode;
//   dfx__startup_rdac        = (dfx__fuseoverride) ? ovrd_startup_rdac : dfx_in.fuse.startup_rdac;
//   dfx__vco_trim_cb         = (dfx__fuseoverride) ? ovrd_vco_trim_cb : dfx_in.fuse.vco_trim_cb;
//   dfx__vco_trim_pg         = (dfx__fuseoverride) ? ovrd_vco_trim_pg : dfx_in.fuse.vco_trim_pg;
//   dfx__iref_mode           = (dfx__fuseoverride) ? ovrd_iref_mode : dfx_in.fuse.iref_mode;

//   dfx__disable_run_upd     = (dfx__fuseoverride) ? ovrd_disable_run_upd : dfx_in.fuse.disable_run_upd;
   dfx__disable_run_upd     = 1'b0; 
//   dfx__startcnt            = (dfx__fuseoverride) ? ovrd_startcnt : dfx_in.fuse.startcnt;
//   dfx__start_mode          = (dfx__fuseoverride) ? ovrd_start_mode : dfx_in.fuse.start_mode;
//
   end : OVRD_MUX_FUSE_SIP

   // Fuse decode to HIP
   //
   always_comb begin : OVRD_MUX_FUSE_HIP

   dfx__tight_loop          = (dfx__fuseoverride) ? ovrd_tight_loop : fz_tight_loopb;
   dfx__lockthresh          = (dfx__fuseoverride) ? ovrd_lockthresh : fz_lockthresh;
   dfx__lockstickyb         = (dfx__fuseoverride) ? ovrd_lockstickyb : fz_lockstickyb;
//   dfx__iref_ctune          = (dfx__fuseoverride) ? ovrd_iref_ctune : dfx_in.fuse.iref_ctune;
//   dfx__iref_ftune          = (dfx__fuseoverride) ? ovrd_iref_ftune : dfx_in.fuse.iref_ftune;
//   dfx__pfd_chop_en         = (dfx__fuseoverride) ? |(ovrd_pfd_chop_val) : |(dfx_in.fuse.pfd_chop_val);
//   dfx__pfd_chop_val        = (dfx__fuseoverride) ? ovrd_pfd_chop_val : dfx_in.fuse.pfd_chop_val;
//   dfx__pvd_mode            = (dfx__fuseoverride) ? ovrd_pvd_mode : dfx_in.fuse.pvd_mode;
//   dfx__ro_freq_sel         = (dfx__fuseoverride) ? ovrd_ro_freq_sel : dfx_in.fuse.ro_freq_sel;
   dfx__pfd_residual_pw     = (dfx__fuseoverride) ? ovrd_pfd_residual_pw : fz_pfd_pw;
   dfx__cp1_trim            = (dfx__fuseoverride) ? ovrd_cp1_trim : fz_cp1trim;
   dfx__cp2_trim            = (dfx__fuseoverride) ? ovrd_cp2_trim : fz_cp2trim;
   dfx__skadj_ctrl          = (dfx__fuseoverride) ? ovrd_skadj_ctrl : fz_skadj;
   dfx__dca_ctrl            = (dfx__fuseoverride) ? ovrd_dca_ctrl : fz_dca_ctrl;
   dfx__dca_cb              = (dfx__fuseoverride) ? ovrd_dca_cb : fz_dca_cb;
   dfx__tllm_en              = (dfx__fuseoverride) ? ovrd_tllm_en : tllm_en;

   end : OVRD_MUX_FUSE_HIP

   // TAP opverride other pins here
   always_comb begin : OVRD_MUX_OTHER_HIP

   dfx__mash_order_plus_one 		= 	(dfx__fuseoverride) ? ovrd_mash_order_plus_one : mash_order_plus_one;
   dfx__ldo_enable_a_int		=	(dfx__fuseoverride) ? ovrd_ldo_enable : ldo_enable ;    // new -nd
   dfx__fz_ldo_vinvoltsel_a 		= 	(dfx__fuseoverride) ? ovrd_fz_ldo_vinvoltsel : fz_ldo_vinvoltsel;    // new -nd
   dfx__fz_ldo_bypass_a			=	(dfx__fuseoverride) ? ovrd_fz_ldo_bypass : fz_ldo_bypass;        // new -nd
   dfx__fz_ldo_extrefsel_a		=	(dfx__fuseoverride) ? ovrd_fz_ldo_extrefsel : fz_ldo_extrefsel;     // new -nd
   dfx__fz_ldo_faststart_a_pre		=	(dfx__fuseoverride) ? ovrd_fz_ldo_faststart : fz_ldo_faststart;     // new -nd
   dfx__fz_ldo_fbtrim_a			=	(dfx__fuseoverride) ? ovrd_fz_ldo_fbtrim : fz_ldo_fbtrim;        // new -nd
   dfx__fz_ldo_reftrim_a		=	(dfx__fuseoverride) ? ovrd_fz_ldo_reftrim : fz_ldo_reftrim;       // new -nd
   dfx__cpnbias		    		= 	(dfx__fuseoverride) ? ovrd_fz_cpnbias : fz_cpnbias;           //new -nd
   dfx__mdiv_ratio_a			=	(dfx__fuseoverride) ? ovrd_mdiv_ratio : mdiv_ratio;           // new -nd
   dfx__vcodiv_ratio_a			=	(dfx__fuseoverride) ? ovrd_vcodiv_ratio : vcodiv_ratio;         // new -nd
   dfx__zdiv0_ratio_a			=	(dfx__fuseoverride) ? ovrd_zdiv0_ratio : zdiv0_ratio;          //new -nd
   dfx__zdiv0_ratio_p5_a		=	(dfx__fuseoverride) ? ovrd_zdiv0_ratio_p5 : zdiv0_ratio_p5;       //new -nd
   dfx__zdiv1_ratio_a			=	(dfx__fuseoverride) ? ovrd_zdiv1_ratio : zdiv1_ratio;          //new -nd
   dfx__zdiv1_ratio_p5_a		=	(dfx__fuseoverride) ? ovrd_zdiv1_ratio_p5 : zdiv1_ratio_p5;       //new -nd
   dfx__fz_irefgen_a			=	(dfx__fuseoverride) ? ovrd_fz_irefgen : fz_irefgen;           //new -nd
   dfx__fz_lpfclksel_a			=	(dfx__fuseoverride) ? ovrd_fz_lpfclksel : fz_lpfclksel;         //new -nd
   dfx__fz_nopfdpwrgate_a		=	(dfx__fuseoverride) ? ovrd_fz_nopfdpwrgate : fz_nopfdpwrgate;      //new -nd
   dfx__fz_pfd_pw_a			=	(dfx__fuseoverride) ? ovrd_fz_pfd_pw : fz_pfd_pw;            //new -nd
   dfx__fz_pfddly_a			=	(dfx__fuseoverride) ? ovrd_fz_pfddly : fz_pfddly;            //new -nd
   dfx__fz_spare_a			=	(dfx__fuseoverride) ? ovrd_fz_spare : fz_spare;             //new -nd
   dfx__fz_startup_a			=	(dfx__fuseoverride) ? ovrd_fz_startup : fz_startup;           //new -nd
   dfx__fz_vcosel_a			=	(dfx__fuseoverride) ? ovrd_fz_vcosel : fz_vcosel;            //new -nd
   dfx__fz_vcotrim_a			=	(dfx__fuseoverride) ? ovrd_fz_vcotrim : fz_vcotrim;           //new -nd
   dfx__fz_lockcnt_a			= 	(dfx__fuseoverride) ? ovrd_fz_lockcnt : fz_lockcnt;
   dfx__fz_lockforce_a			= 	(dfx__fuseoverride) ? ovrd_fz_lockforce : fz_lockforce;

   end : OVRD_MUX_OTHER_HIP

   //logic [4:0] OdcsDlyLineSettingNH;

   // Tap Output
   //   Encode tap output bits to struct
   //
   assign tap_out.pll_enable        = reset_sync__Reset_b_XXnnnL;
   assign tap_out.dist_pwr_good     = dfx__powergood;
   assign tap_out.unlock_count      = unlock_counter__UnlockCountXXnnnH;
   assign tap_out.lock_time         = lock_timer__LockTimeCntXXnnnH;
   assign tap_out.raw_lock          = lock_detector__RawLockXXnnnL;
   assign tap_out.lock              = LockXXnnnL;
   assign tap_out.pll_ratio         = mash__RatioMXH;
   assign tap_out.pll_half_int      = mash__HalfIntMXH;
   assign tap_out.adc_dig_out       = view_adc__dig_out;
   assign tap_out.adc_start         = adc_ctl__StartXXH;
   assign tap_out.adc_done          = view_adc__done;
   assign tap_out.tctrlfsmstate     = tlctrl_sip__StateXXnnnH;
   //assign dfx_out.tap.odcs.odcsfalltrig = odcs_dig__odcsfalltrig;
   //assign dfx_out.tap.odcs.odcsrisetrig = odcs_dig__odcsrisetrig;
   //assign dfx_out.tap.odcs.dummydldelay = OdcsDlyLineSettingNH;
   //assign dfx_out.tap.odcs.stmtrig      = stm_ifdim__StmTrigStatusNH;
   //assign dfx_out.tap.odcs.opsprisesamp = odcs_opsp__RiseSampNH;
   //assign dfx_out.tap.odcs.opspfallsamp = odcs_opsp__FallSampNH;
   assign tap_out.ssc_mod_dfx_run   = ssc_mod_dfx__ModulatorEnNH;
   assign tap_out.ssc_mod_dfx_trig  = ssc_mod_dfx__TriggerRegXDH;
   assign tap_out.iref_done         = iref_ctrl__IrefDoneXXH;
   assign tap_out.pfd_en            = startup_gen__PfdEnXXH;
   assign tap_out.view_freq_count   = view_freq_count;

   //`ip2211ringpll_RANDOM_VAL_WHEN_X(OdcsDlyLineSettingNH, odcs_dll__DlyLineSettingNH, dfx__tight_loop)

   // IDV in/out
   //
   assign dfx_out.idv                  = idv_fub__idv_out;

   // Req/Ack to/from Ratio sync
   //
   //assign dfx__ratio_update_req        = dfx_in.ratio_update_req;
   assign dfx__ratio_update_req        = 1'b0; 
   assign dfx_out.ratio_update_ack     = reg_req_ack__RatioUpdAckMXH;

   // Req/Ack to/from SSC modulator
   //
   //assign dfx__ssc_prof_update_req     = dfx_in.ssc_prof_update_req;
   assign dfx__ssc_prof_update_req     = 1'b0;
   assign dfx_out.ssc_prof_update_ack  = reg_req_ack__SscProfUpdAckMXH;

   // View Output
   //
   assign dfx_out.view.view_dig_out        = view_mux__ViewOutNnnnH;


   // ldo_enable_a is OR of PLLen and Ldoenable  after TAP override
   //
	assign dfx__ldo_enable_a = (dfx__reset_b || dfx__ldo_enable_a_int);
	assign dfx__fz_ldo_faststart_a = ~(dfx__fz_ldo_faststart_a_pre || reset_sync__Reset_b_XXnnnL); 

   // Override mux
   //   Drives DFX override values when the DFX override is selected
   //
   always_comb begin : OVRD_MUX
      
      dfx__reset_b   = (tap_in.ovrd_enable_sel)    ? tap_in.ovrd_enable_val    : Reset_b_NnnnH;
      dfx__powergood = (tap_in.ovrd_powergood_sel) ? tap_in.ovrd_powergood_val : PllDistPwrGoodNnnnH;
      dfx__bypass    = (tap_in.ovrd_bypass_sel)    ? tap_in.ovrd_bypass_val    : BypassNnnnH;
      dfx__ratio     = (tap_in.ovrd_ratio_sel)     ? tap_in.ovrd_ratio_val     : RatioNnnnH;
      dfx__fraction  = (tap_in.ovrd_frac_sel)      ? tap_in.ovrd_frac_val      : FractionNnnnH;

   end : OVRD_MUX
   


endmodule

`endif

`ifndef ip2211ringpll_LJPLL_RESET_SYNC_SV
`define ip2211ringpll_LJPLL_RESET_SYNC_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "ringpll_macros.sv"

module ip2211ringpll_ljpll_reset_sync (
   input  logic ClkRefXXH,

   input  logic dfx__reset_b,		// Pllen after TAP override in ip2211ringpll_ljpll_dfx
   input  logic dfx__bypass,
   input  logic dfx__ldo_enable_a,      // This triggers TIMER before letting PLL Enable go to PLL
   input  logic [1:0] ldo_timer,

   output logic reset_sync__BypassXXnnnL,
   output logic reset_sync__Reset_b_XXnnnL,
   output logic reset_sync__BypassEnXXnnnL,
//Scan controls
   input   logic                         idfx_fscan_rstbypen,
   input   logic                         idfx_fscan_byprstb
);


   logic BypassXXnnnL;
   logic ResetSync_b_XXnnnL;
   logic ClkRefXXH_b;
   logic ResetNH;
   logic dfx__reset_b_postscan;
   logic ResetSyncResetBNH;
   logic ResetSyncResetBNH_pre;
   logic sync_dfx__ldo_enable_a;

   assign ResetNH = ~dfx__reset_b_postscan;
   assign ResetSyncResetBNH_pre = ((reset_sync__BypassXXnnnL==BypassXXnnnL) & dfx__reset_b_postscan);
//Changes done for scan
  assign dfx__reset_b_postscan =  idfx_fscan_rstbypen ? idfx_fscan_byprstb : dfx__reset_b;
  assign ResetSyncResetBNH =  idfx_fscan_rstbypen ? idfx_fscan_byprstb : ResetSyncResetBNH_pre;


   // Clock inverter for negedge flops
   //
   `ip2211ringpll_CLKINV(ClkRefXXH_b, ClkRefXXH)

   // Syncronize reset into the reference clock domain
   //
   `ip2211ringpll_ASYNC_RST_2MSFF_META(BypassXXnnnL, dfx__bypass, ClkRefXXH_b, dfx__reset_b_postscan)
   `ip2211ringpll_ASYNC_RST_MSFF(reset_sync__BypassXXnnnL, BypassXXnnnL, ClkRefXXH_b, ResetNH)
   `ip2211ringpll_ASYNC_RST_2MSFF_META(ResetSync_b_XXnnnL, 1'b1, ClkRefXXH_b, ResetSyncResetBNH)

    // Synchronize ldo_enable_a into reference clock domain.
   `ip2211ringpll_ASYNC_RST_2MSFF_META(sync_dfx__ldo_enable_a, dfx__ldo_enable_a, ClkRefXXH_b, dfx__reset_b_postscan)

   // Bypass Enable = syncronized reset_b
   //
   assign reset_sync__BypassEnXXnnnL = ResetSync_b_XXnnnL;


   // TIMER: 
   // Trigger when dfx__ldo_enable_a is asserted.
   // fz_spare[1:0] are used to determine number of refclk to be counted before asserting 
   // reset_sync__Reset_b_XXnnnL.
   //
   // fz_spare[1:0] 
   //   00 = 32 (default)
   //   01 = 48
   //   10 = 72
   //   11 = 180
   //
   logic [7:0] ldocountval;
//     logic [7:0] count;
//   logic enable_pll;
   logic ResetSync_b_XXnnnL_premux;

     always_comb begin
      unique casez (ldo_timer[1:0])
         2'b00: ldocountval = 8'b00100000; 	// d32
         2'b01: ldocountval = 8'b00110000; 	// d48 
         2'b10: ldocountval = 8'b01001000;	// d72
         2'b11: ldocountval = 8'b10110100;     	// d180
         `ip2211ringpll_XDefault(ldocountval)
      endcase // casez (ldo_timer[1:0])
     end

//	// Counter
//	always @(posedge (ClkRefXXH))
//	begin
//		if (sync_dfx__ldo_enable_a == 1'b0)
//			count <= ldocountval;   // Default
//		else
//			if (count > 8'b0)
//				count <= (count - 1);	// Decrement by 1 each Refclk
//			else
//				count <= 0;
//
//
//		if ((sync_dfx__ldo_enable_a == 1'b1) & (count == 8'b0))
//			enable_pll <= 1'b1;		// Trigger PLL enable
//		else
//			enable_pll <= 1'b0;		// Gating PLL enable till timer expires
//	end

   logic ldodly_cnt_rst, ldodly_cnt_done, ldodly_cnt_done_sticky;   
   logic [7:0] ldodly_cnt, ldodly_cnt_next;
   logic  ldodly_cnt_rst_pre;
   assign ldodly_cnt_rst_pre = ~sync_dfx__ldo_enable_a & ~ResetSync_b_XXnnnL;
  
//Changes done for scan
assign ldodly_cnt_rst = idfx_fscan_rstbypen ? ~idfx_fscan_byprstb : ldodly_cnt_rst_pre;
 
   `ip2211ringpll_ASYNC_RST_MSFF(ldodly_cnt[7:0], ldodly_cnt_next[7:0], ClkRefXXH_b, ldodly_cnt_rst) 
   assign  ldodly_cnt_next = ldodly_cnt_done_sticky ? 8'b00000000 : (ldodly_cnt + 8'b00000001);
   assign ldodly_cnt_done = (ldodly_cnt == ldocountval);
   
   `ip2211ringpll_ASYNC_RST_MSFF(ldodly_cnt_done_sticky, (ldodly_cnt_done_sticky | ldodly_cnt_done), ClkRefXXH_b, ldodly_cnt_rst) 
   
   
   // Make sure reset_b is always low when bypass = 1
   //
   always_comb begin : RESET_B_LOGIC
//SSG	ResetSync_b_XXnnnL_premux = (ResetSync_b_XXnnnL & enable_pll);
	ResetSync_b_XXnnnL_premux = (ResetSync_b_XXnnnL & ldodly_cnt_done_sticky);
      //reset_sync__Reset_b_XXnnnL = reset_sync__BypassXXnnnL ? 1'b0 : ResetSync_b_XXnnnL;

      //reset_sync__Reset_b_XXnnnL = reset_sync__BypassXXnnnL ? 1'b0 : ResetSync_b_XXnnnL_premux;

	// NOTE: For pll bypass to work (bypass=1, and we should then see refclk on clk outputs),        //  so need to take the bypass term out of the reset going to the hip.
      reset_sync__Reset_b_XXnnnL = ResetSync_b_XXnnnL_premux;

   end : RESET_B_LOGIC


endmodule

`endif

`ifndef ip2211ringpll_STARTUP_GEN_SV
`define ip2211ringpll_STARTUP_GEN_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "ringpll_macros.sv"
//`include "ljpll_dfx.vh"

module ip2211ringpll_startup_gen (
   input  logic                            ClkRefXXH,
   input  logic                            reset_sync__Reset_b_XXnnnL,
//   input  logic                            dfx__openloop,
//   input  logic                            dfx__start_mode,
//   input  logic                            iref_ctrl__IrefDoneXXH,
//   input  logic                            vctl_trim_fsm__TrimDoneXXH,

   output logic                            startup_gen__ForcePullUpXXH,
   output logic                            startup_gen__VctlTrimEnXXH,
   output logic                            startup_gen__VctlRdacEnXXH,
   output logic                            startup_gen__PfdEnXXH
);

// EVERYTHING BELOW is commented out
/*
///=====================================================================================================================
/// Reset Generation
///=====================================================================================================================
   logic ResetXXL;

   always_comb begin : RESET_GEN
      ResetXXL = ~reset_sync__Reset_b_XXnnnL;
   end : RESET_GEN

///=====================================================================================================================
/// Mode Decoding
///=====================================================================================================================
   
   logic SerialModeNH;

   // Only use serial mode if we are not in openloop
   //
   always_comb begin : SERIAL_MODE
      SerialModeNH = (~dfx__openloop) & dfx__start_mode;
   end : SERIAL_MODE

///=====================================================================================================================
/// PLL Startup FSM
///=====================================================================================================================

   // LJPLL Start FSM
   //
   enum logic [3:0] {
      START_IREF         = 4'b0100,
      START_TRIM         = 4'b1010,
      START_LOCKING      = 4'b0001
   } FsmStateXXH, FsmStateNxtXXH;
   logic TrimDonePosedgeXXH;

   always_comb begin : STARTUP_FSM

      // One-hot encoded to prevent glitching on the output
      //   Each state has a bit for the output. For more information see
      //   the default statement of the unique case below
      //
      unique case (FsmStateXXH)

         START_IREF : begin
            FsmStateNxtXXH              = (~SerialModeNH | iref_ctrl__IrefDoneXXH) ? START_TRIM : FsmStateXXH ;
         end
         
         START_TRIM : begin
            FsmStateNxtXXH              = TrimDonePosedgeXXH   ? START_LOCKING  :
                                                                 FsmStateXXH    ;
         end
         
         START_LOCKING : begin
            FsmStateNxtXXH              = FsmStateXXH ;
         end

         default : begin
            `ifndef ip2211ringpll_SVA_OFF
                 `ip2211ringpll_ASSERTC_FORBIDDEN(Illegal_Case_select, !($isunknown(FsmStateXXH)), 0, `ip2211ringpll_ERR_MSG("Illegal case selector: 'FsmStateXXH' = %h", FsmStateXXH));
            `endif
         `ifndef ip2211ringpll_NO_VCSSIM
         if (^(FsmStateXXH) === 1'bX) begin
            FsmStateNxtXXH              = 'x ;
         end else begin
         `endif
            FsmStateNxtXXH              = START_IREF ;
         `ifdef ip2211ringpll_NO_VCSSIM
         end
         `endif
         end

      endcase

   end : STARTUP_FSM

   logic VctlTrimEnPrevXXH;
   logic TrimDonePrevXXH;

   `ip2211ringpll_ASYNC_RST_MSFF(VctlTrimEnPrevXXH, FsmStateXXH[3], ClkRefXXH, ResetXXL)
   `ip2211ringpll_ASYNC_SET_MSFF(TrimDonePrevXXH, vctl_trim_fsm__TrimDoneXXH, ClkRefXXH, ResetXXL)
   `ip2211ringpll_ASYNC_RSTD_MSFF(FsmStateXXH, FsmStateNxtXXH, ClkRefXXH, ResetXXL, START_IREF)

   always_comb begin : TRIM_DONE_POSEDGE
      TrimDonePosedgeXXH = vctl_trim_fsm__TrimDoneXXH & ~TrimDonePrevXXH;
   end : TRIM_DONE_POSEDGE

//   always_comb begin : GLITCH_FREE_DECODE
//         startup_gen__VctlTrimEnXXH  = FsmStateXXH[3] & ~VctlTrimEnPrevXXH;
//         startup_gen__ForcePullUpXXH = FsmStateXXH[2];  // Glitch Protect
//         startup_gen__VctlRdacEnXXH  = FsmStateXXH[1];  // Glitch Protect
//         startup_gen__PfdEnXXH       = FsmStateXXH[0];  // Glitch Protect
//   end : GLITCH_FREE_DECODE
*/

 assign startup_gen__VctlTrimEnXXH = 1'b0;
 assign startup_gen__ForcePullUpXXH = 1'b0;
 assign startup_gen__VctlRdacEnXXH = 1'b0;

logic pfden_1;
logic pfden_2;
// assign startup_gen__PfdEnXXH = reset_sync__Reset_b_XXnnnL;
   `ip2211ringpll_ASYNC_RST_MSFF(pfden_1, 1'b1, ClkRefXXH, ~reset_sync__Reset_b_XXnnnL)
   `ip2211ringpll_ASYNC_RST_MSFF(pfden_2, pfden_1, ClkRefXXH, ~reset_sync__Reset_b_XXnnnL)
 assign startup_gen__PfdEnXXH = pfden_2;

endmodule

`endif

`ifndef ip2211ringpll_IDV_FUBLET_SV
`define ip2211ringpll_IDV_FUBLET_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "ringpll_macros.sv"
//`include "ljpll_dfx.vh"

module ip2211ringpll_idv_fublet 
//#(parameter IDV_ADDR_BITS = 10) 
(
//   input  t_ljpll_idv_in_ifc        

   input  logic                         idvdisable_bi,          // new -nd
   input  logic                         idvfreqai,              // new -nd
   input  logic                         idvfreqbi,              // new -nd
   input  logic                         idvpulsei,              // new -nd
   input  logic                         idvtclki,              // new -nd
   input  logic                         idvtctrli,             // new -nd
   input  logic                         idvtdi,                 // new -nd
   input  logic                         idvtresi,               // new -nd
//   input  logic                         clkidvih,               // new -nd

//   output t_ljpll_idv_out_ifc       
   output logic                         idvdisable_bo,  // part of dfx_out
   output logic                         idvfreqao,              // part of dfx_out
   output logic                         idvfreqbo,              // part of dfx_out
   output logic                         idvpulseo,              // part of dfx_out
   output logic                         idvtclko,               // part of dfx_out
   output logic                         idvtctrlo,              // part of dfx_out
   output logic                         idvtdo,         // part of dfx_out
   output logic                         idvtreso,               // part of dfx_out



   input  logic                     ClkIdvIH,

   output logic                     idv_fub__IdvGateEnNH,
   output logic                     idv_fub__IdvDisableTH,
   //output logic [IDV_ADDR_BITS-1:0] idv_fub__IdvAddrTH
   output logic [9:0] idv_fub__IdvAddrTH
);

   localparam IDV_ADDR_BITS = 10;
   localparam FUBLET_ADDR_BITS = IDV_ADDR_BITS;
   localparam NUM_FUBLETS = IDV_ADDR_BITS / FUBLET_ADDR_BITS;

   logic [NUM_FUBLETS-1:0] [FUBLET_ADDR_BITS-1 : 0] IdvFubletAddrTH, IdvFubletAddrNxtTH;
   logic ClkTH_b;
   logic [NUM_FUBLETS-1:0] IdvAddr0NxtTH;
   logic [NUM_FUBLETS-1:0] FubletEnTH;
   logic [NUM_FUBLETS-1:0] TdoTH;
   logic [NUM_FUBLETS-1:0] TdoTL;
   logic [NUM_FUBLETS-1:0] TctrlTL;
   genvar g_fublet;

   // Create an inverted tclk signal for low phase drivers
   //
   `ip2211ringpll_CLKINV(ClkTH_b, idvtclki)
   // adding generate block to resolve LEC issue where this module gets
   // HSD : 16014566973
   generate
   for (g_fublet=0; g_fublet<NUM_FUBLETS; g_fublet++) begin : FUBLET
      logic [FUBLET_ADDR_BITS-1:0] IdvFubletAddrTmpTH;
      logic FubletEnTmpTH_b;
      logic TdiTH;
      logic TdiTH_b;

      // If fublet is the first fublet, use TDI from the IDV chain
      // 
      // Else use the previous fublet's TDO as TDI
      //
      if (g_fublet == 0)
         assign TdiTH = idvtdi;
      else
         assign TdiTH = TdoTH[g_fublet-1];

      // TDO has 3 potential paths:
      //    TCTRL = 1    : Fublet Enable Bit (output from flop)
      //    FubletEn = 0 : TDI
      //    FubletEn = 1 : IDV Address MSB
      //
      always_comb begin : TDO
         unique casez ({idvtctrli, FubletEnTH[g_fublet]})
            2'b1? : TdoTH[g_fublet] = FubletEnTH[g_fublet];
            2'b00 : TdoTH[g_fublet] = TdiTH;
            2'b01 : TdoTH[g_fublet] = IdvFubletAddrTH[g_fublet][FUBLET_ADDR_BITS-1];
            `ip2211ringpll_XDefault(TdoTH[g_fublet])
         endcase
      end : TDO
      
      // Fublet Enable Flop
      //   Reads an enable bit from TDI whenever tctrl is asserted
      //
      always_comb begin : TDI_INV
         TdiTH_b = ~TdiTH;
      end : TDI_INV
      `ip2211ringpll_EN_ASYNC_RST_MSFF(FubletEnTmpTH_b, TdiTH_b, idvtclki, idvtctrli, idvtresi)
      assign FubletEnTH[g_fublet] = ~FubletEnTmpTH_b;

      // IDV Address Flops
      //   Decode IDV address from TDI clocked by TCLK.
      //   These flops are only enabled if the fublet is enabled and TCTRL is
      //    deselected (i.e. IDV shift mode)
      //
      `ip2211ringpll_EN_ASYNC_RST_MSFF(IdvFubletAddrTmpTH, IdvFubletAddrNxtTH[g_fublet], idvtclki, (FubletEnTH[g_fublet] & ~idvtctrli), idvtresi)
      assign IdvFubletAddrTH[g_fublet] = IdvFubletAddrTmpTH;

      // IDV Addresses are shifted from TDI except in the pulse case.
      //   When pulse is asserted, the next bit(0) is always tied to 0
      //
      always_comb begin : IDV_ADDR_NXT
         IdvAddr0NxtTH[g_fublet]      = idvpulsei ? 1'b0 : TdiTH;
         IdvFubletAddrNxtTH[g_fublet] = {IdvFubletAddrTH[g_fublet][FUBLET_ADDR_BITS-2:0], IdvAddr0NxtTH[g_fublet]};
      end : IDV_ADDR_NXT
 
      // Assign fublet address to IDV address bits
      //
      assign idv_fub__IdvAddrTH[(FUBLET_ADDR_BITS * (g_fublet+1)) - 1 : FUBLET_ADDR_BITS * g_fublet] = IdvFubletAddrTH;

   end : FUBLET

   endgenerate

   logic TdoRstTH;

   always_comb begin : TDO_RST
      TdoRstTH = idvtresi | ~(idvdisable_bi); 
   end : TDO_RST

   // Latch TDO to low phase for output
   //
   `ip2211ringpll_ASYNC_RST_LATCH(TdoTL, TdoTH[NUM_FUBLETS-1], ClkTH_b, TdoRstTH)

   // Latch TCTRL to low phase for output
   //
   `ip2211ringpll_ASYNC_RST_LATCH(TctrlTL, idvtctrli, ClkTH_b, idvtresi)

   // IDV creates the following feedthroughs:
   //   tclk
   //   tdo   (Low Phase TCLK)
   //   trst
   //   disable_b
   //   tctrl (Low Phase TCLK)
   //   pulse out
   //
   `ip2211ringpll_CLKBF(idvtclko, idvtclki)
   assign   idvtdo        = TdoTL;
   assign   idvtreso      = idvtresi;
   assign   idvdisable_bo = idvdisable_bi;
   assign   idvtctrlo     = TctrlTL;
   assign   idvpulseo     = idvpulsei;

   // Calculate a bypass to use for passing input clock to output. Also pass
   //   bypass IDV code to analog when IDV is bypassed.
   //
   //   IDV does not output a clock in the following cases:
   //     PULSE    =  1
   //     IdvAddr  = '0
   //     -- IdvAddr  = '1 note, this was beacon before, but it has been reclaimed
   //     FubletEn = 0
   //
   always_comb begin : IDV_BYPASS
     
      // rename this to something else like idv enabled
      //   IDV OSC is disabled under any of the following conditions:
      //     * IDV enable (disable_b) is 0
      //     * Fublet is disabled
      //     * IDV Pulse is asserted
      //     * IDV address is 0
      //
      //idv_fub__IdvDisableTH = ~(idvdisable_bi) | ~(&FubletEnTH) | idvpulsei | (idv_fub__IdvAddrTH == `ip2211ringpll_ZX(1'b0, IDV_ADDR_BITS));
      idv_fub__IdvDisableTH = ~(idvdisable_bi) | ~(&FubletEnTH) | idvpulsei | (idv_fub__IdvAddrTH == `ip2211ringpll_ZX(1'b0, 10));

   end : IDV_BYPASS

   // Enable the IDV clock whenever IDV is not bypassed.
   // IDV is only enabled when the PLL is in openloop and not bypassed.
   //  
   //  ClkIdvIH = idv_fub__IdvGateEnNH && ClkPll
   //
   //  openloop = tap control
   //    when openloop = 0, we ignore idv
   //
   always_comb begin : IDV_EN
      idv_fub__IdvGateEnNH = ~idv_fub__IdvDisableTH;
   end : IDV_EN

   // Generate output frequency on channel A, always pass channel B
   //
 
   logic ClkIdvFreqAIH;
   logic ClkIdvFreqAIH_b;
   logic ClkIdvIH_b;
   logic ClkStg2aIH;
   logic ClkStg2bIH;
   logic ClkIdvFreqAOH;
   logic ClkIdvFreqBIH;
   logic ClkIdvFreqBOH;

   // XNOR Channel A
   //  --> pass ClkIdvIH when freqA parked at 1
   //  --> pass not(freqA) when ClkIdvIH parked at 0
   //
   assign ClkIdvFreqAIH = idvfreqai;
   `ip2211ringpll_CLKINV(ClkIdvFreqAIH_b, ClkIdvFreqAIH)
   `ip2211ringpll_CLKINV(ClkIdvIH_b, ClkIdvIH)
   `ip2211ringpll_CLK_NAND(ClkStg2aIH, ClkIdvFreqAIH, ClkIdvIH)
   `ip2211ringpll_CLK_NAND(ClkStg2bIH, ClkIdvFreqAIH_b,       ClkIdvIH_b)
   `ip2211ringpll_CLK_NAND(ClkIdvFreqAOH, ClkStg2aIH, ClkStg2bIH)
   assign idvfreqao = ClkIdvFreqAOH;

   // Invert Channel B
   //
   assign ClkIdvFreqBIH = idvfreqbi;
   `ip2211ringpll_CLKINV(ClkIdvFreqBOH, ClkIdvFreqBIH)
   assign idvfreqbo = ClkIdvFreqBOH;


endmodule

`endif

`ifndef ip2211ringpll_LJPLL_IDV_SV
`define ip2211ringpll_LJPLL_IDV_SV

module ip2211ringpll_ljpll_idv (
   input  logic         dfx__openloop,
//   input  logic [3:0]   dfx__startup_rdac, // Not needed anymore in ip22 ringpll
   input  logic [3:0]   dfx__vco_trim_pg,
   input  logic [2:0]   dfx__vco_trim_cb,
   input  logic [9:0]   idv_fub__IdvAddrTH,
   input  logic         idv_fub__IdvDisableTH,

   output logic [3:0]   idv__RdacCtlTH,
   output logic [2:0]   idv__CbCtlTH,
   output logic [3:0]   idv__PgCtlTH
);


///========================================================================================================
/// IDV is enabled only in openloop
///========================================================================================================
   
   logic IdvEnabledTH;

   always_comb begin : IDV_EN
      IdvEnabledTH = ~idv_fub__IdvDisableTH & dfx__openloop;
   end : IDV_EN

///========================================================================================================
/// Address Decoding -- PLL specific decoding (not from IDV spec)
///========================================================================================================
  
   logic [3:0]   RdacCtlTH;
   logic [2:0]   CbCtlTH;
   logic [3:0]   PgCtlTH;
   
   // Decode the address into tuning knobs
   //
   always_comb begin : IDV_DECODE
      RdacCtlTH =  idv_fub__IdvAddrTH[9:6];
      CbCtlTH   =  {~idv_fub__IdvAddrTH[5:4], 1'b0};
      PgCtlTH   =  idv_fub__IdvAddrTH[3:0];
   end : IDV_DECODE

   always_comb begin : IDV_OVERRIDE_FUSES
      //idv__RdacCtlTH = IdvEnabledTH ? RdacCtlTH : dfx__startup_rdac;
      idv__RdacCtlTH = IdvEnabledTH ? RdacCtlTH : 4'b0;
      idv__CbCtlTH   = IdvEnabledTH ? CbCtlTH   : dfx__vco_trim_cb;
      idv__PgCtlTH   = IdvEnabledTH ? PgCtlTH   : dfx__vco_trim_pg;
   end : IDV_OVERRIDE_FUSES


endmodule

`endif

`ifndef ip2211ringpll_VCTL_TRIM_FSM_SV
`define ip2211ringpll_VCTL_TRIM_FSM_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
`ifndef ip2211ringpll_SVA_OFF
   //`include "intel_checkers.vs"
`endif

typedef enum logic [1:0] {
   VCTL_TRIM_COMP_OFF = 2'b00,
   VCTL_TRIM_PULL_UP  = 2'b10,
   VCTL_TRIM_PULL_DN  = 2'b01,
   VCTL_TRIM_COMP_ON  = 2'b11
} t_VctlTrimFSM;

module ip2211ringpll_vctl_trim_fsm (
   input  logic ClkRefXXH,
   input  logic reset_sync__Reset_b_XXnnnL,
   input  logic dfx__openloop,
   input  logic startup_gen__VctlTrimEnXXH,
   input  logic startup_gen__ForcePullUpXXH,
   input  logic iref_ctrl__IrefDoneXXH,
   input  logic pll_core__CompOutNnnnH,

   output logic vctl_trim_fsm__VctlRdacShortXXH,
   output logic vctl_trim_fsm__TrimDoneXXH,
   output logic vctl_trim_fsm__CmpEnXXH,
   output logic vctl_trim_fsm__PullUpNnnnH,
   output logic vctl_trim_fsm__PullDnNnnnH,
   input logic idfx_fscan_rstbypen,
   input logic idfx_fscan_byprstb 
);


   logic ResetXXL;

   // Reset generation for downstream logic
   //
   assign ResetXXL = ~reset_sync__Reset_b_XXnnnL;

   ///==========================================================================
   /// VCTL Trim FSM
   ///   The FSM starts up with the comparator disabled and is enabled when the
   ///   vctl pump is triggered.  The TrimDone bit starts at 1 so that gray
   ///   code transitions between the off and on state are not required.
   ///
   ///==========================================================================
   
   t_VctlTrimFSM TrimFsmStateXXH, TrimFsmNxtStateXXH;
   logic TrimDoneXXH;
   logic TrimDoneNH_b;
   logic PullUpModeXXH;
   logic PullDnModeXXH;
   logic ForceDoneSetXXH;
   logic TrimDoneRstXXH;
            
            //   syncronize comp out?
            //   This should be covered by making it so that any state
            //   transition will force pulldone to be 1 eventually (in
            //   a short period of time)
            //
   
   always_comb begin : VCTL_TRIM_FSM

      case (TrimFsmStateXXH)

         VCTL_TRIM_COMP_OFF : begin
            TrimFsmNxtStateXXH         = (startup_gen__VctlTrimEnXXH) ? VCTL_TRIM_COMP_ON : TrimFsmStateXXH;
            PullUpModeXXH              = 1'b0;
            PullDnModeXXH              = 1'b0;
            ForceDoneSetXXH            = 1'b1;
            TrimDoneRstXXH             = 1'b0;
            vctl_trim_fsm__CmpEnXXH    = 1'b0;
         end
         
         VCTL_TRIM_COMP_ON  : begin
            TrimFsmNxtStateXXH         = (TrimDoneXXH) ? TrimFsmStateXXH : ((pll_core__CompOutNnnnH) ? VCTL_TRIM_PULL_UP : VCTL_TRIM_PULL_DN);
            PullUpModeXXH              = 1'b0;
            PullDnModeXXH              = 1'b0;
            ForceDoneSetXXH            = 1'b0;
            TrimDoneRstXXH             = 1'b1;
            vctl_trim_fsm__CmpEnXXH    = 1'b1;
         end
         
         VCTL_TRIM_PULL_DN  : begin
            TrimFsmNxtStateXXH         = (vctl_trim_fsm__TrimDoneXXH) ? VCTL_TRIM_COMP_OFF : TrimFsmStateXXH;
            PullUpModeXXH              = 1'b0;
            PullDnModeXXH              = 1'b1;
            ForceDoneSetXXH            = 1'b0;
            TrimDoneRstXXH             = 1'b0;
            vctl_trim_fsm__CmpEnXXH    = 1'b1;
         end
         
         VCTL_TRIM_PULL_UP  : begin
            TrimFsmNxtStateXXH         = (vctl_trim_fsm__TrimDoneXXH) ? VCTL_TRIM_COMP_OFF : TrimFsmStateXXH;
            PullUpModeXXH              = 1'b1;
            PullDnModeXXH              = 1'b0;
            ForceDoneSetXXH            = 1'b0;
            TrimDoneRstXXH             = 1'b0;
            vctl_trim_fsm__CmpEnXXH    = 1'b1;
         end

      endcase

   end : VCTL_TRIM_FSM

   `ip2211ringpll_ASYNC_RSTD_MSFF(TrimFsmStateXXH, TrimFsmNxtStateXXH, ClkRefXXH, ResetXXL, VCTL_TRIM_COMP_OFF)

   ///==========================================================================
   /// Pull Done tracking
   ///   The pull up and pull down tracks the comparator output and stops the
   ///   pullup/pulldown when the comparator trips.
   ///
   ///==========================================================================
  
   logic TrimDoneSetNH;
   logic TrimDoneSetNH_pre;
   logic TrimDoneXXH_b;
   logic IrefDoneXXL_b;
   logic ForceDoneSetFlopXXH;
   logic PullUpModeFlopXXH;
   logic PullDnModeFlopXXH;

   // Flop Signals that are glitch sensitive
   //
   `ip2211ringpll_ASYNC_SET_MSFF(ForceDoneSetFlopXXH, ForceDoneSetXXH, ClkRefXXH, ResetXXL)
   `ip2211ringpll_ASYNC_RST_MSFF(PullUpModeFlopXXH, PullUpModeXXH, ClkRefXXH, ResetXXL)
   `ip2211ringpll_ASYNC_RST_MSFF(PullDnModeFlopXXH, PullDnModeXXH, ClkRefXXH, ResetXXL)
 //Changes done for scan   
assign TrimDoneSetNH = idfx_fscan_rstbypen ? ~idfx_fscan_byprstb : TrimDoneSetNH_pre;
 
   // Set Pull Done whenever the comparator trips
   //
   always_comb TrimDoneSetNH_pre =  ResetXXL                                      |
                                ForceDoneSetFlopXXH                           |
                                (PullUpModeFlopXXH & ~pll_core__CompOutNnnnH) |
                                (PullDnModeFlopXXH &  pll_core__CompOutNnnnH) ;

   // Allow the FSM to reset TrimDone (when the comparator switches on)
   //
   `ip2211ringpll_EN_ASYNC_RST_MSFF(TrimDoneNH_b, 1'b1, ClkRefXXH, TrimDoneRstXXH, TrimDoneSetNH)

   // Syncronize the TrimDone signal to the FSM clock domain
   //
   `ip2211ringpll_ASYNC_RST_2MSFF_META(TrimDoneXXH_b, (TrimDoneNH_b | TrimDoneRstXXH), ClkRefXXH, reset_sync__Reset_b_XXnnnL)
   assign TrimDoneXXH                     = ~TrimDoneXXH_b;
   assign vctl_trim_fsm__TrimDoneXXH      =  ~dfx__openloop & iref_ctrl__IrefDoneXXH & TrimDoneXXH;

   logic ClkRefXXH_b;

   `ip2211ringpll_CLKINV(ClkRefXXH_b, ClkRefXXH)

   `ip2211ringpll_ASYNC_SET_MSFF(IrefDoneXXL_b, ~iref_ctrl__IrefDoneXXH, ClkRefXXH_b, ResetXXL)

   // This should be glitch protected
   //   -- IrefDoneXXL must come from a flop
   //   -- TrimDoneXXH must come from a flop
   //
   //   Note that RDAC short is expected to deassert before the TrimDone is
   //   registered by the downstream FSM.
   //
   //   i.e. VctlRdacShort is low at least 1 phase before vctlrdacen is
   //   deasserted
   //
   assign vctl_trim_fsm__VctlRdacShortXXH = (dfx__openloop | IrefDoneXXL_b) & TrimDoneXXH & (PullUpModeFlopXXH | PullDnModeFlopXXH);

   // Generate pull up and pull down signals based on the comparator initial
   // reading and whether the comparator has tripped
   //
   always_comb begin : PULLUP_PULLDOWN_GEN

      vctl_trim_fsm__PullUpNnnnH = (PullUpModeFlopXXH & TrimDoneNH_b) | startup_gen__ForcePullUpXXH;
      vctl_trim_fsm__PullDnNnnnH =  PullDnModeFlopXXH & TrimDoneNH_b;

   end : PULLUP_PULLDOWN_GEN

///========================================================================================================
/// Assertions
///========================================================================================================

`ifndef ip2211ringpll_SVA_OFF
   `ip2211ringpll_ASSERTC_FORBIDDEN(R_vctl_trim_fsm_pullup_and_pulldn_both_on, vctl_trim_fsm__PullUpNnnnH & vctl_trim_fsm__PullDnNnnnH, 1'b0, `ip2211ringpll_ERR_MSG("[LJPLL] VCTL pull-up and pull-dn are both asserted at the same time. Electrical contention."));
`endif


endmodule

`endif

`ifndef ip2211ringpll_ADC_CTL_SV 
`define ip2211ringpll_ADC_CTL_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "ringpll_macros.sv"
//`include "ljpll_dfx.vh"

module ip2211ringpll_adc_ctl (
         input  logic               ClkRefXXH,
//         input  logic               reset_sync__Reset_b_XXnnnL,
         //input  t_ljpll_dfx_in_ifc  dfx_in,
         //input  t_ljpll_tap_in_ifc  tap_in,
   	input logic                 dfx__adc_start,
   	input logic [1:0]           dfx__adc_start_cnt,

         output logic               adc_ctl__StartXXH,
         output logic               adc_ctl__Reset_bXXL,

  //Scan controls
   input   logic                         idfx_fscan_rstbypen,
   input   logic                         idfx_fscan_clkungate,
   input   logic                         idfx_fscan_byprstb
   

);

///========================================================================================================
/// Module Begin
///========================================================================================================
   
   logic ClkRefXXH_b;
   logic ClkAdcCountXXH;
   logic dfx__adc_start_postscan;

   // Clock inverter for negedge flops
   //
   `ip2211ringpll_CLKINV(ClkRefXXH_b, ClkRefXXH)

   logic DfxAdcStartXXL;

   // Syncronize ADC Start
   //
   //`ip2211ringpll_ASYNC_RST_2MSFF_META(DfxAdcStartXXL, 1'b1, ClkRefXXH_b, dfx_in.tap.adc_start) 
   //`ip2211ringpll_ASYNC_RST_2MSFF_META(DfxAdcStartXXL, 1'b1, ClkRefXXH_b, tap_in.adc_start) 
   `ip2211ringpll_ASYNC_RST_2MSFF_META(DfxAdcStartXXL, 1'b1, ClkRefXXH_b, dfx__adc_start_postscan) 

//Changes done  for scan
assign dfx__adc_start_postscan = idfx_fscan_rstbypen ? idfx_fscan_byprstb : dfx__adc_start;


   logic ResetXXL;
   logic ResetXXL_pre;

   // Generate a reset from the RESET_B
   //
   always_comb begin : RESET_GEN
      ResetXXL_pre = ~DfxAdcStartXXL;
   end : RESET_GEN


//Changes done  for scan
assign ResetXXL = idfx_fscan_rstbypen ? ~idfx_fscan_byprstb : ResetXXL_pre;

   logic [7:0] AdcCountXXH;

   // Counter Flops
   //
   `ip2211ringpll_ASYNC_RST_MSFF(AdcCountXXH, (AdcCountXXH + `ip2211ringpll_ZX(1'b1,$bits(AdcCountXXH))), ClkAdcCountXXH, ResetXXL)
  
   
   logic AdcStartXXL;

   /// Programmable sticky assert ADC delay of ~1us after ADC startcount, 
   /// Based on the count of 64/96/128/160 ClkRefXXH.
   //
   always_comb begin
      //unique casez (dfx_in.tap.adc_start_cnt)
      //unique casez (tap_in.adc_start_cnt)
      unique casez (dfx__adc_start_cnt)
         2'b00 : adc_ctl__StartXXH = AdcCountXXH[6];
         2'b01 : adc_ctl__StartXXH = &AdcCountXXH[6:5];
         2'b10 : adc_ctl__StartXXH = AdcCountXXH[7];
         2'b11 : adc_ctl__StartXXH = &{AdcCountXXH[7],AdcCountXXH[5]};
         `ip2211ringpll_XDefault(adc_ctl__StartXXH)
      endcase
   end

   `ip2211ringpll_LATCH_P(AdcStartXXL, adc_ctl__StartXXH, ClkRefXXH)


   logic AdcCountClkEnXXL;
   always_comb AdcCountClkEnXXL = DfxAdcStartXXL & ~AdcStartXXL;

//idfx_fscan_clkungate Changes done  for scan
   `ip2211ringpll_CLKAND(ClkAdcCountXXH, ClkRefXXH, (AdcCountClkEnXXL || idfx_fscan_clkungate))

   always_comb adc_ctl__Reset_bXXL = DfxAdcStartXXL; 


endmodule

`endif

`ifndef ip2211ringpll_REG_REQ_ACK_SV
`define ip2211ringpll_REG_REQ_ACK_SV

//`include "soc_macros.sv"

module ip2211ringpll_reg_req_ack (
   input  logic   ssc_mod_dfx__ClkModMXH,
   input  logic   LockXXnnnL,
   input  logic   dfx__disable_run_upd,
   input  logic   dfx__ratio_update_req,
   input  logic   dfx__ssc_prof_update_req,
   input  logic   ssc__ProfUpdateMXH,
   input  logic   ssc__RatioUpdateMXH,

   output logic   reg_req_ack__SscProfUpdReqMXH,
   output logic   reg_req_ack__SscProfUpdAckMXH,
   output logic   reg_req_ack__RatioUpdReqMXH,
   output logic   reg_req_ack__RatioUpdAckMXH,
   output logic   reg_req_ack__MashStateResetMXH
);

///========================================================================================================
/// Module Begin
///========================================================================================================
   
///=====================================================================================================================
/// Reset Generation
///=====================================================================================================================
   logic ResetXXL;

   always_comb begin : RESET_GEN
      ResetXXL = ~LockXXnnnL;
   end : RESET_GEN

///=====================================================================================================================
/// Ratio Req Syncronizer
///=====================================================================================================================
   
   logic RatioUpdReqMXH;

   // Syncronize the Ratio Update Bit
   //
   `ip2211ringpll_ASYNC_RST_2MSFF_META(RatioUpdReqMXH, dfx__ratio_update_req, ssc_mod_dfx__ClkModMXH, LockXXnnnL)

   always_comb begin : RATIO_REQ_IGNORE
      reg_req_ack__RatioUpdReqMXH = RatioUpdReqMXH & ~dfx__disable_run_upd;
   end : RATIO_REQ_IGNORE

   // Track profile update done which remains sticky (acts as ack) until
   //   request deasserts. Update is done when req & profile update OK is
   //   asserted
   //
   `ip2211ringpll_ASYNC_RST_MSFF(reg_req_ack__RatioUpdAckMXH, RatioUpdReqMXH & ((ssc__RatioUpdateMXH | dfx__disable_run_upd) | reg_req_ack__RatioUpdAckMXH), ssc_mod_dfx__ClkModMXH, ResetXXL)
   
///=====================================================================================================================
/// SSC Profile Update Req Syncronizer
///=====================================================================================================================

   logic SscProfUpdReqMXH;

   // Syncronize the Profile Update Bit
   //
   `ip2211ringpll_ASYNC_RST_2MSFF_META(SscProfUpdReqMXH, dfx__ssc_prof_update_req, ssc_mod_dfx__ClkModMXH, LockXXnnnL)

   always_comb begin : PROFILE_REQ_IGNORE
      reg_req_ack__SscProfUpdReqMXH = SscProfUpdReqMXH & ~dfx__disable_run_upd;
   end : PROFILE_REQ_IGNORE

   // Track profile update done which remains sticky (acts as ack) until
   //   request deasserts.
   //
   `ip2211ringpll_ASYNC_RST_MSFF(reg_req_ack__SscProfUpdAckMXH, SscProfUpdReqMXH & ((ssc__ProfUpdateMXH | dfx__disable_run_upd) | reg_req_ack__SscProfUpdAckMXH), ssc_mod_dfx__ClkModMXH, ResetXXL)

///=====================================================================================================================
/// MASH modulator reset
///=====================================================================================================================

   // Reset MASH modulator when SSC profile is updating or ratio is
   // updating
   //
   always_comb reg_req_ack__MashStateResetMXH = (ssc__ProfUpdateMXH | ssc__RatioUpdateMXH);

// assumes prof update never asserts when disable_run_upd is 1
//   reason: disable_run_upd causes req to never assert -- the profile
//   shouldn't be updated unless req asserts (exception is reset)
endmodule

`endif

`ifndef ip2211ringpll_SYNC_RESET_CLKGEN_SV
`define ip2211ringpll_SYNC_RESET_CLKGEN_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"

module ip2211ringpll_sync_reset_clkgen (
   input  logic                    ClkRefXXH,
   input  logic                    pll_fbgen__ClkFbMXH,
   input  logic                    reset_sync__BypassEnXXnnnL,
   input  logic                    EarlyLockXXnnnH,
   input  logic                    LockXXnnnL,

   output logic                    sync_reset_clkgen__ClkFbGateMXH,

  input logic  idfx_fscan_rstbypen,
  input logic  idfx_fscan_clkungate,
  input logic  idfx_fscan_byprstb

);

///========================================================================================================
/// Module Begin
///========================================================================================================
      
///=====================================================================================================================
/// Clock Gate
///=====================================================================================================================

   logic ClkRefXXL;
   logic LockXXnn1L;
   logic LockXXnn1L_pre;
   logic EarlyLockXXnn1H;
   logic EarlyLockXXnn1H_pre;
   logic ResetXXL;
   logic ResetXXL_pre;
   logic SscMashClkEnMXL;
   logic PulseEn1MXL;
   logic PulseRiseEdgeMXL;
   logic EarlyLockMXL;
   logic ClkFbMXL;

   `ip2211ringpll_CLKINV(ClkFbMXL, pll_fbgen__ClkFbMXH)
   `ip2211ringpll_CLKINV(ClkRefXXL, ClkRefXXH)

   always_comb begin : RESET
      ResetXXL_pre = ~reset_sync__BypassEnXXnnnL;
   end : RESET

//Changes done for scan 
assign ResetXXL = idfx_fscan_rstbypen ? ~idfx_fscan_byprstb : ResetXXL_pre;
assign EarlyLockXXnn1H = idfx_fscan_rstbypen ? idfx_fscan_byprstb : EarlyLockXXnn1H_pre;
assign LockXXnn1L = idfx_fscan_rstbypen ? idfx_fscan_byprstb : LockXXnn1L_pre;


   // Flop earlylock just in case there's combo glitches upstream
   //
   `ip2211ringpll_ASYNC_RST_MSFF(EarlyLockXXnn1H_pre, EarlyLockXXnnnH, ClkRefXXH, ResetXXL)

   // cross early lock for enabling 1 cycle on earlylock assertion
   //
   `ip2211ringpll_ASYNC_RST_2MSFF_META(EarlyLockMXL, 1'b1, ClkFbMXL, EarlyLockXXnn1H)
   `ip2211ringpll_MSFF(PulseEn1MXL, EarlyLockMXL, ClkFbMXL)

   always_comb begin : RISE_EDGE_DETECT
      PulseRiseEdgeMXL = ~PulseEn1MXL & EarlyLockMXL;
   end : RISE_EDGE_DETECT
   
   // Flop lock just in case there's combo glitches upstream
   //
   `ip2211ringpll_ASYNC_RST_MSFF(LockXXnn1L_pre, LockXXnnnL, ClkRefXXL, ResetXXL)

   // phase path crossing before modulator enable
   //
   `ip2211ringpll_ASYNC_RST_2MSFF_META(SscMashClkEnMXL, 1'b1, ClkFbMXL, LockXXnn1L)

   // Add a clock gate to shut down feedback clock to ssc/mash before lock
   //
   `ip2211ringpll_CLKAND(sync_reset_clkgen__ClkFbGateMXH, pll_fbgen__ClkFbMXH, (SscMashClkEnMXL | PulseRiseEdgeMXL))

///========================================================================================================
/// Module End
///========================================================================================================

endmodule
`endif

`ifndef ip2211ringpll_SSC_MOD_SV
`define ip2211ringpll_SSC_MOD_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
`ifndef ip2211ringpll_SVA_OFF
//`include "intel_checkers.vs"
`endif
//`include "ringpll_macros.sv"

module ip2211ringpll_ssc_mod 
//#(parameter RATIO_BITS=10, parameter FRAC_BITS=24, parameter FMOD_BITS=9) 
(
   input  logic                    ssc_mod_dfx__ClkModMXH,
   input  logic                    LockXXnnnL,
  
   input  logic [9:0]   dfx__RatioStepNH,
   input  logic [23:0]    dfx__FracStepNH,
   input  logic                    dfx__ssc_en,
   input  logic [1:0]              dfx__ssc_mode,
   input  logic [8:0]    dfx__ssc_cyc_to_peak_m1,
   input  logic                    reg_req_ack__SscProfUpdReqMXH,
   input  logic                    reg_req_ack__SscProfUpdAckMXH,
   input  logic                    reg_req_ack__RatioUpdReqMXH,
   input  logic                    reg_req_ack__RatioUpdAckMXH,


   input  logic [9:0]   dfx__ratio,
   input  logic [23:0]    dfx__fraction,
   output logic [9:0]   ssc__RatioMXH,
   output logic [23:0]    ssc__FractionMXH,
   output logic                    ssc__DirectionMXH,
   output logic                    ssc__ProfUpdateMXH,
   output logic                    ssc__RatioUpdateMXH
);

///========================================================================================================
/// Module Begin
///========================================================================================================

///=====================================================================================================================
/// Reset Generation
///=====================================================================================================================
   logic ResetXXL;

   always_comb begin : RESET_GEN
      ResetXXL = ~LockXXnnnL;
   end : RESET_GEN

///=====================================================================================================================
/// Modulation period tracking - used to keep track of modulation period
///=====================================================================================================================
   
   logic CntUpToProfGenMXH;
   logic [8:0] CountToPeakMXH;
   logic [8:0] CountToPeakCntNxtMXH;
   logic [8:0] CountToPeakNxtMXH;
   logic [8:0] CountToPeakRstValNH;
   logic [8:0] CountToPeakSetXXL;
   logic [8:0] CountToPeakRstXXL;
   logic [1:0]           SscModeMXH;
   logic                 ReloadMXH;
   logic [8:0] CycToPeakm1MXH;
   
   logic                 SscEnMXH;


   // Generate an async set rst to load the counter prior to enable
   //
   always_comb begin : CNT_TO_PEAK_RST
      // If center spread, start at halfway to the peak
      //
      CountToPeakRstValNH = dfx__ssc_mode[1] ? {1'b0, dfx__ssc_cyc_to_peak_m1[8:1]} : dfx__ssc_cyc_to_peak_m1;
   end : CNT_TO_PEAK_RST

   // Create a counter that counts cycles_to_peak times before reloading
   //
   `ip2211ringpll_EN_MSFF(CountToPeakMXH, CountToPeakNxtMXH, ssc_mod_dfx__ClkModMXH, (SscEnMXH | ResetXXL | ssc__ProfUpdateMXH))
   
   // Whenever CountToPeak is 0, reload counter
   //
   always_comb begin : RELOAD
      ReloadMXH = (CountToPeakMXH == 9'b0);
   end : RELOAD

   always_comb begin : CNT_TO_PEAK_NXT
      CountToPeakCntNxtMXH = (ReloadMXH)   ? CycToPeakm1MXH                               :
                                                  CountToPeakMXH - {{8{1'b0}}, 1'b1} ;
      CountToPeakNxtMXH    = (ResetXXL | ssc__ProfUpdateMXH) ? CountToPeakRstValNH                          :
                                                             CountToPeakCntNxtMXH                         ;

   end : CNT_TO_PEAK_NXT
  
   // Enable flop - whenever we reach the peak or 0, change direction
   //
   `ip2211ringpll_EN_ASYNC_RST_MSFF(ssc__DirectionMXH, ssc__ProfUpdateMXH ? 1'b0 : ~ssc__DirectionMXH, ssc_mod_dfx__ClkModMXH, (ssc__ProfUpdateMXH | ReloadMXH), ResetXXL) 

   // Generate Count Up Signal Based on Mode
   //
   always_comb begin : MODE_DECODE
      CntUpToProfGenMXH = SscModeMXH[0] ? ~ssc__DirectionMXH : // Downspread / center, start @ down
                                           ssc__DirectionMXH ; // Upspread / center, start @ up

   end : MODE_DECODE

///=====================================================================================================================
/// Output Ratio/Fraction generation
///=====================================================================================================================

   logic [9:0]  RatioNxtMXH;
   logic [23:0]   FracNxtMXH;
   logic [9:0]  RatioStepMXH;
   logic [23:0]   FracStepMXH;
   logic                   DeltaEnMXH;
   logic                   RatioLoadMXH;
   logic                   ProfileUpdateOkMXH;

   // TODO: set to numcycle like hold value for n cycles
   //    if numcycle is a power of 2 then we can use
   //    CountToPeakMXH[log2(numcycle)-1:0]=='0 to be the delta enable
   //
   assign DeltaEnMXH = 1'b1;
   
   always_comb ssc__RatioUpdateMXH = (ProfileUpdateOkMXH & reg_req_ack__RatioUpdReqMXH & ~reg_req_ack__RatioUpdAckMXH);

   always_comb begin : RATIOFRAC_NXT
      RatioLoadMXH = (ResetXXL | ssc__RatioUpdateMXH);
      unique casez ({RatioLoadMXH, DeltaEnMXH, CntUpToProfGenMXH})
         3'b1?? : begin {RatioNxtMXH,FracNxtMXH} = {dfx__ratio,    dfx__fraction};                                end
         3'b00? : begin {RatioNxtMXH,FracNxtMXH} = {ssc__RatioMXH, ssc__FractionMXH};                             end
         3'b011 : begin {RatioNxtMXH,FracNxtMXH} = {ssc__RatioMXH,ssc__FractionMXH} + {RatioStepMXH,FracStepMXH}; end
         3'b010 : begin {RatioNxtMXH,FracNxtMXH} = {ssc__RatioMXH,ssc__FractionMXH} - {RatioStepMXH,FracStepMXH}; end
         `ip2211ringpll_XDefault_Part_Def_Name({RatioNxtMXH,FracNxtMXH},
                                 {ssc__RatioMXH, ssc__FractionMXH},
                                 {RatioLoadMXH,
                                 DeltaEnMXH,
                                 CntUpToProfGenMXH},
                                 ratiofrac_nxt)
      endcase
   end : RATIOFRAC_NXT

   `ip2211ringpll_EN_MSFF(ssc__RatioMXH, RatioNxtMXH, ssc_mod_dfx__ClkModMXH,   (RatioLoadMXH | SscEnMXH))
   `ip2211ringpll_EN_MSFF(ssc__FractionMXH, FracNxtMXH, ssc_mod_dfx__ClkModMXH, (RatioLoadMXH | SscEnMXH))

///=====================================================================================================================
/// Profile Update Syncronization
///=====================================================================================================================
   
   logic [8:0] CountToPeakRstValMXH;

   // When doing a dynamic update - only refresh the profile if the next
   //   cycle is the starting point. The starting point is derived by
   //   computing if:
   //   --The next cycles to peak count will be the reset val
   //   --The current direction is opposite from the start value (except in
   //      the case of centerspread for an odd # of cyc to peak
   //      (cyc_to_peak_m1 + 1) )
   //
   always_comb begin : PROFILE_UPDATE
      ProfileUpdateOkMXH = ~SscEnMXH | ((CountToPeakCntNxtMXH == CountToPeakRstValMXH) & (ssc__DirectionMXH ^ (SscModeMXH[1] & ~CycToPeakm1MXH[0])) );
      ssc__ProfUpdateMXH = ProfileUpdateOkMXH & reg_req_ack__SscProfUpdReqMXH & ~reg_req_ack__SscProfUpdAckMXH;
   end : PROFILE_UPDATE

   `ip2211ringpll_EN_MSFF(RatioStepMXH,   dfx__RatioStepNH,        ssc_mod_dfx__ClkModMXH, (ResetXXL | ssc__ProfUpdateMXH))
   `ip2211ringpll_EN_MSFF(FracStepMXH,    dfx__FracStepNH,         ssc_mod_dfx__ClkModMXH, (ResetXXL | ssc__ProfUpdateMXH))
   `ip2211ringpll_EN_MSFF(SscEnMXH,       dfx__ssc_en,             ssc_mod_dfx__ClkModMXH, (ResetXXL | ssc__ProfUpdateMXH))
   `ip2211ringpll_EN_MSFF(SscModeMXH,     dfx__ssc_mode,           ssc_mod_dfx__ClkModMXH, (ResetXXL | ssc__ProfUpdateMXH))
   `ip2211ringpll_EN_MSFF(CycToPeakm1MXH, dfx__ssc_cyc_to_peak_m1, ssc_mod_dfx__ClkModMXH, (ResetXXL | ssc__ProfUpdateMXH))

   always_comb CountToPeakRstValMXH = SscModeMXH[1] ? {1'b0, CycToPeakm1MXH[8:1]} : CycToPeakm1MXH;

///========================================================================================================
/// Assertions
///========================================================================================================

   `ifndef ip2211ringpll_SVA_OFF

   `ifndef ip2211ringpll_NO_VCSSIM
   logic [9:0]   RatioCapture_inst;
   logic [23:0]    FractionCapture_inst;

   `ip2211ringpll_EN_MSFF(RatioCapture_inst,   dfx__ratio,        ssc_mod_dfx__ClkModMXH, (ResetXXL | ssc__ProfUpdateMXH))
   `ip2211ringpll_EN_MSFF(FractionCapture_inst,    dfx__fraction,         ssc_mod_dfx__ClkModMXH, (ResetXXL | ssc__ProfUpdateMXH))

   `ip2211ringpll_ASSERTS_FORBIDDEN(R_ssc_mod_downspread_above_ratio_in,
                        {ssc__RatioMXH, ssc__FractionMXH} > {RatioCapture_inst, FractionCapture_inst},
                        posedge ssc_mod_dfx__ClkModMXH,
                        ResetXXL | (SscModeMXH!==2'b00),
                     `ip2211ringpll_ERR_MSG("[LJPLL] SSC caused the ratio to go above the programmed ratio in downspread mode"));
   
   `ip2211ringpll_ASSERTS_FORBIDDEN(R_ssc_mod_upspread_below_ratio_in,
                        {ssc__RatioMXH, ssc__FractionMXH} < {RatioCapture_inst, FractionCapture_inst},
                        posedge ssc_mod_dfx__ClkModMXH,
                        ResetXXL | (SscModeMXH!==2'b01),
                     `ip2211ringpll_ERR_MSG("[LJPLL] SSC caused the ratio to go below  the programmed ratio in upspread mode"));
   `endif


   `ip2211ringpll_ASSERTS_FORBIDDEN(R_ssc_profile_update_at_wrong_ratiofrac,
                      SscEnMXH & ssc__ProfUpdateMXH & ({RatioNxtMXH,FracNxtMXH} != {dfx__ratio, dfx__fraction}),
                      posedge ssc_mod_dfx__ClkModMXH,
                      ResetXXL,
                     `ip2211ringpll_ERR_MSG("[LJPLL] SSC profile update on wrong ratio and/or fraction"));

 
   `endif

endmodule

`endif

`ifndef ip2211ringpll_RATIO_ASYNC_MUX_SV
`define ip2211ringpll_RATIO_ASYNC_MUX_SV

module ip2211ringpll_ratio_async_mux 
//#(parameter RATIO_BITS=10, parameter FRAC_BITS=24) 
(
   input  logic                    reset_sync__BypassXXnnnL,
   input  logic                    LockXXnnnL,
   input  logic  [9:0]  dfx__ratio,
   input  logic  [9:0]  ssc__RatioMXH,
   input  logic  [23:0]   dfx__fraction,
   input  logic  [23:0]   ssc__FractionMXH,
   input logic [5:0]     mdiv_ratio, 
   output logic  [9:0]  ratio_async_mux__RatioMXH,
   output logic  [23:0]   ratio_async_mux__FractionMXH
);

logic ref_divider_active;

///========================================================================================================
/// Module Begin
///========================================================================================================
   
   // Reset changes many ref / fb clock cycles after the flops are
   //    syncronously loaded. The clock is disabled at the time of reset
   //    change (for at least 1.5 cycles of ref period)
   //
   //    1.5 cycle MCO of ref to these flop receivers
   //
   always_comb  begin : RATIOFRAC_MUX
// if refclk divider is used, then don\BFt look at ssc_ratio, as both modes are not allowed simultaneously 
      ref_divider_active = |(mdiv_ratio[5:1]);

      ratio_async_mux__RatioMXH    = (reset_sync__BypassXXnnnL | ~LockXXnnnL | ref_divider_active) ? dfx__ratio    :
                                                                                ssc__RatioMXH ;
 
      ratio_async_mux__FractionMXH = (reset_sync__BypassXXnnnL | ~LockXXnnnL | ref_divider_active) ? dfx__fraction    :
                                                                                ssc__FractionMXH ;

   end : RATIOFRAC_MUX
      
///========================================================================================================
/// Module End
///========================================================================================================

endmodule

`endif

`ifndef ip2211ringpll_SSC_MOD_DFX_SV
`define ip2211ringpll_SSC_MOD_DFX_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "ringpll_macros.sv"

module ip2211ringpll_ssc_mod_dfx (
   input  logic                    sync_reset_clkgen__ClkFbGateMXH,
//   input  logic                    reset_sync__Reset_b_XXnnnL,
   input  logic                    LockXXnnnL,
   input  logic                    dfx__SscModTrigNH,
   input  logic  [1:0]             dfx__SscModStepsNH,
   input  logic                    dfx__SscDfxEnNH,
   input  logic  [1:0]             dfx__SscModClkDivNH,
   output logic                    ssc_mod_dfx__TriggerRegXDH,
   output logic                    ssc_mod_dfx__ModulatorEnNH,
   output logic                    ssc_mod_dfx__ClkModMXH
);

///========================================================================================================
/// Module Begin
///========================================================================================================

///=====================================================================================================================
/// Clock Dividers
///=====================================================================================================================

   logic [2:0] DivCntMXL;
   logic [2:0] DivCntNxtMXL;
   logic ClkFbMXH_b;
   logic ClkDiv2MXH;
   logic ClkDiv4MXH;
   logic ClkDiv8MXH;
   logic ClkModDfx0XDH;
   logic ClkModDfx1XDH;
   logic DivEnXXL;
   logic DivEnBXXL;

   logic Div2EnMXL;
   logic Div4EnMXL;
   logic Div8EnMXL;

   // The clock dividers are enabled whenever the SSC DFX module is
   // enabled and the PLL is enabled
   //
   always_comb begin : DIV_EN
      DivEnXXL = LockXXnnnL & dfx__SscDfxEnNH; 
      // ALTERNATE: explore (& ~dfx__openloop) for cross clock justification
      DivEnBXXL = ~DivEnXXL;
   end : DIV_EN

   // Clock Div Counter
   //
   `ip2211ringpll_CLKINV(ClkFbMXH_b, sync_reset_clkgen__ClkFbGateMXH)
   always_comb begin : DIV_CNT_NXT_VAL
      DivCntNxtMXL = (DivCntMXL - 3'd1);
   end : DIV_CNT_NXT_VAL
   `ip2211ringpll_ASYNC_SET_MSFF(DivCntMXL, DivCntNxtMXL, ClkFbMXH_b, DivEnBXXL)

   always_comb begin : CLK_DIV_EN
      Div2EnMXL = (DivCntMXL[0]   == 1'b0);
      Div4EnMXL = (DivCntMXL[1:0] == 2'b00);
      Div8EnMXL = (DivCntMXL[2:0] == 3'b000);
   end : CLK_DIV_EN

   `ip2211ringpll_CLKAND(ClkDiv2MXH, sync_reset_clkgen__ClkFbGateMXH, Div2EnMXL)
   `ip2211ringpll_CLKAND(ClkDiv4MXH, sync_reset_clkgen__ClkFbGateMXH, Div4EnMXL)
   `ip2211ringpll_CLKAND(ClkDiv8MXH, sync_reset_clkgen__ClkFbGateMXH, Div8EnMXL)

   logic [1:0] SscModClkDivQualNH;
   logic ClkModDfxXDH;

   always_comb begin : SSC_MOD_CLKDIV_QUAL
      SscModClkDivQualNH = DivEnXXL ? dfx__SscModClkDivNH
                                    : 2'b00                ;
   end : SSC_MOD_CLKDIV_QUAL

   // Select the internal DFX clock to be used by the step and stop
   // counter system
   //
   //     SscModClkDiv | CLK_TO_COUNTER
   //   ---------------------------------
   //          00      |  Fb / 1
   //          01      |  Fb / 2
   //          10      |  Fb / 4
   //          11      |  Fb / 8
   //
   `ip2211ringpll_MAKE_CLK_2TO1MUX(ClkModDfx0XDH, sync_reset_clkgen__ClkFbGateMXH,         ClkDiv2MXH,    SscModClkDivQualNH[0])
   `ip2211ringpll_MAKE_CLK_2TO1MUX(ClkModDfx1XDH, ClkDiv4MXH,           ClkDiv8MXH,    SscModClkDivQualNH[0])
   `ip2211ringpll_MAKE_CLK_2TO1MUX(ClkModDfxXDH,  ClkModDfx0XDH,        ClkModDfx1XDH, SscModClkDivQualNH[1])

///=====================================================================================================================
/// Trigger Syncronization
///=====================================================================================================================

   logic TapTriggerXD0H;
   logic TapTriggerXD1H;
   logic CounterReloadXDH;

   // Create a history of Tap triggers in order to control the stepper
   // counter
   //
   `ip2211ringpll_ASYNC_RST_2MSFF_META(TapTriggerXD0H, dfx__SscModTrigNH, ClkModDfxXDH, DivEnXXL)
   `ip2211ringpll_ASYNC_RST_MSFF      (TapTriggerXD1H, TapTriggerXD0H,    ClkModDfxXDH, DivEnBXXL)

   assign ssc_mod_dfx__TriggerRegXDH = TapTriggerXD1H;

   // Reload the counter whenever the trigger changes (i.e. tap triggered
   // the stepper system)
   //
   always_comb begin : TAP_TRIGGER
      CounterReloadXDH = (TapTriggerXD0H ^ TapTriggerXD1H);
   end : TAP_TRIGGER

///=====================================================================================================================
/// Tap Controlled Stepper Counter
///=====================================================================================================================

   logic [5:0] CounterReloadValNH;

   // The counter counts a number of cycles set by a tap register before
   // stopping the SSC/Frac-N modulators so that the user can read the
   // value out on tap
   //
   //     SscModSteps  | Cycles To Count
   //   ---------------------------------
   //          00      |  1
   //          01      |  16
   //          10      |  32
   //          11      |  63
   //
   always_comb begin : COUNTER_RELOAD_VAL
      unique casez (dfx__SscModStepsNH)
         2'b00 : CounterReloadValNH = 6'd1;
         2'b01 : CounterReloadValNH = 6'd16;
         2'b10 : CounterReloadValNH = 6'd32;
         2'b11 : CounterReloadValNH = 6'd63;
         `ip2211ringpll_XDefault(CounterReloadValNH)
      endcase
   end : COUNTER_RELOAD_VAL

   logic DfxModEnXDH;
   logic [5:0] CountXDH;
   logic [5:0] CountNxtXDH;

   // The counter is enabled whenever the counter is not 0
   //
   always_comb begin : DFX_MODULE_EN
      DfxModEnXDH = !(CountXDH == 6'h0);
      ssc_mod_dfx__ModulatorEnNH = DfxModEnXDH;
   end : DFX_MODULE_EN

   // The counter always counts down to 0 and is reloaded whenever the tap
   // triggers a reload
   //
   always_comb begin : CNT_NXT_VAL
      CountNxtXDH = CounterReloadXDH ? CounterReloadValNH   :
                                       (CountXDH - 6'd1)    ;
   end : CNT_NXT_VAL
   
   // Counter Flops
   //
   `ip2211ringpll_EN_ASYNC_RST_MSFF(CountXDH, CountNxtXDH, ClkModDfxXDH, (CounterReloadXDH | DfxModEnXDH), DivEnBXXL)

///=====================================================================================================================
/// Clock Output Generation
///=====================================================================================================================
   
   logic DfxModEnXDL;
  
   // The DFX clock is enabled whenever the counter is not 0
   //
   // If the DFX module is disabled, the reference clock is passed directly
   //  to the output (by upstream muxing).  Otherwise, the Clock
   //   is a gated DFX clock generated by this module
   //
   `ip2211ringpll_LATCH_P(DfxModEnXDL, (DfxModEnXDH | ~dfx__SscDfxEnNH | ~LockXXnnnL), ClkModDfxXDH)
   `ip2211ringpll_CLKAND(ssc_mod_dfx__ClkModMXH, ClkModDfxXDH, DfxModEnXDL)

endmodule

`endif

`ifndef ip2211ringpll_SIGMA_DELTA_SV
`define ip2211ringpll_SIGMA_DELTA_SV

//`include "soc_macros.sv"

module ip2211ringpll_sigma_delta #(parameter SD_BITS = 16) (
   input  logic                 ClkModMXH,
   input  logic                 LockXXnnnL,
   input  logic                 reg_req_ack__MashStateResetMXH,
   input  logic [SD_BITS-1:0]   FractionMXH,
   output logic [SD_BITS-1:0]   ErrValMXH,
   output logic                 CarryMXH
);


   logic ResetXXL;
   
   always_comb begin : RESET_GEN
      ResetXXL = ~LockXXnnnL;
   end : RESET_GEN

   logic [SD_BITS-1:0] CarryErrValMXH;
   logic [SD_BITS:0] CarryErrValNxtMXH;

   always_comb begin : ACCUMULATOR_NXT
      CarryErrValNxtMXH = reg_req_ack__MashStateResetMXH ? '0                                       :
                                                           CarryErrValMXH[SD_BITS-1:0] + FractionMXH;
   end : ACCUMULATOR_NXT

   `ip2211ringpll_ASYNC_RST_MSFF(CarryErrValMXH, CarryErrValNxtMXH[SD_BITS-1:0], ClkModMXH, ResetXXL)

   always_comb begin : OUTPUT
      CarryMXH  = CarryErrValNxtMXH[SD_BITS];
      ErrValMXH = CarryErrValNxtMXH[SD_BITS-1:0];
   end : OUTPUT


endmodule

`endif

`ifndef ip2211ringpll_MASH_CARRY_SV
`define ip2211ringpll_MASH_CARRY_SV

//`include "soc_macros.sv"
//`include "ringpll_macros.sv"

module ip2211ringpll_mash_carry #(parameter CARRY_IN_BITS = 2, parameter bit NO_FLOPS=0) (
   input  logic                            ClkModMXH,
   input  logic                            LockXXnnnL,
   input  logic                            reg_req_ack__MashStateResetMXH,
   input  logic signed [CARRY_IN_BITS-1:0] CarryInMXH,
   input  logic signed [CARRY_IN_BITS-1:0] CarryInDelayMXH,
   input  logic                            SdStageCarryMXH,
   output logic signed [CARRY_IN_BITS:0]   CarryOutMXH,
   output logic signed [CARRY_IN_BITS:0]   CarryOutDelayMXH
);

///=====================================================================================================================
/// Reset Generation
///=====================================================================================================================
   logic ResetXXL;

   always_comb begin : RESET_GEN
      ResetXXL = ~LockXXnnnL;
   end : RESET_GEN


   // add 1 carry each stage
   //
   localparam CARRY_OUT_BITS = CARRY_IN_BITS+1;

   if (!NO_FLOPS) begin : DELAY_FLOPS
      // Generate a delayed version of the ip2211ringpll_mash_carry stage's carry out
      //
      `ip2211ringpll_ASYNC_RST_MSFF(CarryOutDelayMXH, reg_req_ack__MashStateResetMXH ? '0 : CarryOutMXH, ClkModMXH, ResetXXL)
   end : DELAY_FLOPS

   // Calculate the CarryOut
   //
   always_comb begin : CARRY_OUT
      CarryOutMXH = `ip2211ringpll_SX(CarryInMXH,      $bits(CarryOutMXH)) -
                    `ip2211ringpll_SX(CarryInDelayMXH, $bits(CarryOutMXH)) +
                    `ip2211ringpll_ZX(SdStageCarryMXH, $bits(CarryOutMXH)) ;
   end : CARRY_OUT


endmodule

`endif

`ifndef ip2211ringpll_MASH_MOD_SV
`define ip2211ringpll_MASH_MOD_SV

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "sigma_delta.sv"
//`include "mash_carry.sv"
//`include "ringpll_macros.sv"
`ifndef ip2211ringpll_SVA_OFF
//`include "intel_checkers.vs"
`endif

module ip2211ringpll_mash_mod 
//#(parameter FRAC_BITS = 24, parameter RATIO_BITS = 10, parameter ORDER=2) 
(
   input  logic                    ssc_mod_dfx__ClkModMXH,
   input  logic                    LockXXnnnL,
   input  logic                    reg_req_ack__MashStateResetMXH,
   input  logic                    dfx__mash_order_plus_one,
   input  logic [9:0]   ratio_async_mux__RatioMXH,
   input  logic [23:0]    ratio_async_mux__FractionMXH,
   output logic [9:0]   mash__RatioMXH,
   output logic                    mash__HalfIntMXH,
   output logic                    mash__PllModOnNH
);

 
   // Local parameter declaration to track sigma delta bits
   //
   //localparam SD_BITS = FRAC_BITS - 1;
   localparam SD_BITS = 23;

///=====================================================================================================================
/// Reset Generation
///=====================================================================================================================
   logic ResetXXL;

   always_comb begin : RESET_GEN
      ResetXXL = ~LockXXnnnL;
   end : RESET_GEN

///=====================================================================================================================
/// Static Modulator Enabled Signal
///=====================================================================================================================
   always_comb begin : MOD_ENABLED
      mash__PllModOnNH = |(ratio_async_mux__FractionMXH[22:0]);
   end : MOD_ENABLED

///=====================================================================================================================
/// Clock Rename
///=====================================================================================================================

   logic ClkModMXH;

   assign ClkModMXH = ssc_mod_dfx__ClkModMXH;

///========================================================================================================
/// Sigma Delta Modulators
///========================================================================================================
   
   genvar g_order;
   logic [2:0] [22:0] ErrValMXH;
   logic [2:0] CarryMXH;
   logic ClkLastOrderMXH;
   
   //=============================================================================
   // Sigma Delta
   //
   //  The sigma delta modulators are generated based on the requested
   //  ORDER parameter.  ORDER+1 sigma deltas are generated so that the
   //  user can select post-silicon if they want order or order+1.
   //
   //  The sigmal deltas are configured in a cascaded fashion so that the
   //  accumulator value of the previous sigma delta is fed to the desired
   //  input step of the next sigma delta.
   //
   //  Since the downstream dividers support half integer ratios, the
   //  sigma delta's internal accumulator will be width fractional bits - 1
   //
   //=============================================================================

   // Generate 1st order sigma delta
   //
   ip2211ringpll_sigma_delta #(.SD_BITS(23))  sigma_delta_ord_1 (
         .FractionMXH   ( ratio_async_mux__FractionMXH[22:0]   ),
         .ErrValMXH     ( ErrValMXH[0]                                ),
         .CarryMXH      ( CarryMXH[0]                                 ),
         .*
   );

   // Generate requested order of mash by duplicating the sigma deltas and
   // cascading
   //
   for (g_order=1; g_order<2; g_order++) begin : SIGMA_DELTA_BLOCKS
      ip2211ringpll_sigma_delta #(.SD_BITS(23)) ip2211ringpll_sigma_delta (
         .FractionMXH   ( ErrValMXH[g_order-1]   ),
         .ErrValMXH     ( ErrValMXH[g_order]     ),
         .CarryMXH      ( CarryMXH[g_order]      ),
         .*
      );
   end : SIGMA_DELTA_BLOCKS
 
   // Disable n+1 order sigma delta clock when 
   `ip2211ringpll_CLKAND(ClkLastOrderMXH, ClkModMXH, dfx__mash_order_plus_one)

   // Generate Last Order MASH+1
   //
   logic [22:0] FractionLastOrderMXH;

   always_comb begin : FRACTION_LAST_ORDER
      FractionLastOrderMXH = dfx__mash_order_plus_one ? ErrValMXH[1] : {23{1'b0}};
   end : FRACTION_LAST_ORDER

   // Generate n+1 order sigma delta
   //
   ip2211ringpll_sigma_delta #(.SD_BITS(23))  sigma_delta_ord_np1 (
         .ClkModMXH     ( ClkLastOrderMXH      ),
         .FractionMXH   ( FractionLastOrderMXH ),
         .ErrValMXH     ( ErrValMXH[2]     ),
         .CarryMXH      ( CarryMXH[2]      ),
         .*
   );

///========================================================================================================
/// Carry State Hold
///========================================================================================================

   // each stage adds 1 carry starting from 2 bits (value + sign)
   //   therefore, the governing equation for carry bits for any given
   //   stage is:
   //    x + 2
   //    x represents stage number (starting from the 0th stage)
  
   // accounting for order + 1 (example order = 2 means last stage is 3rd
   // order)
   //
   localparam MAX_CARRY_WIDTH = (2 + 1) + 1;

   logic signed [2:0] [MAX_CARRY_WIDTH-1:0] CarryDeltaMXH;
   logic signed [2:1] [MAX_CARRY_WIDTH-2:0] CarryDeltaDelayMXH;
   logic CarryDelayLastStageMXH;
   
   always_comb CarryDeltaMXH[2][1:0] = {1'b0,CarryMXH[2]};

   // Generate delayed carry for input to the last stage carry delta calculation
   //
   `ip2211ringpll_ASYNC_RST_MSFF(CarryDelayLastStageMXH, CarryDeltaMXH[2][0], ClkModMXH, ResetXXL)
   assign CarryDeltaDelayMXH[2][1:0] = {1'b0,CarryDelayLastStageMXH};

   for (g_order=1;g_order>=0; g_order--) begin : MASH_CARRY_BLOCKS
      localparam CARRY_IN_BITS = (1)-g_order + 2;
      if (g_order==0) begin : NO_FLOPS
         // Last stage does not have any flops for delay
         //
         ip2211ringpll_mash_carry #(.NO_FLOPS(1),.CARRY_IN_BITS(CARRY_IN_BITS)) mash_carry_stage_1 (
	    .ClkModMXH        (  ClkModMXH                                        ),
	    .LockXXnnnL       (  LockXXnnnL                                       ),
	    .reg_req_ack__MashStateResetMXH ( reg_req_ack__MashStateResetMXH      ),
            .CarryInMXH       (  CarryDeltaMXH     [g_order+1][CARRY_IN_BITS-1:0] ),
            .CarryInDelayMXH  (  CarryDeltaDelayMXH[g_order+1][CARRY_IN_BITS-1:0] ),
            .SdStageCarryMXH  (  CarryMXH          [g_order]                      ),
            .CarryOutMXH      (  CarryDeltaMXH     [g_order]  [CARRY_IN_BITS  :0] ),
            .CarryOutDelayMXH (                                                   )
         );
      end : NO_FLOPS
      else begin : FLOPS
         // 1st stage carry comes from last order sigma delta
         //
         ip2211ringpll_mash_carry #(.NO_FLOPS(0),.CARRY_IN_BITS(CARRY_IN_BITS)) mash_carry_stage   (
	    .ClkModMXH        (  ClkModMXH                                        ),
	    .LockXXnnnL       (  LockXXnnnL                                       ),
	    .reg_req_ack__MashStateResetMXH ( reg_req_ack__MashStateResetMXH      ),
            .CarryInMXH       (  CarryDeltaMXH     [g_order+1][CARRY_IN_BITS-1:0] ),
            .CarryInDelayMXH  (  CarryDeltaDelayMXH[g_order+1][CARRY_IN_BITS-1:0] ),
            .SdStageCarryMXH  (  CarryMXH          [g_order]                      ),
            .CarryOutMXH      (  CarryDeltaMXH     [g_order]  [CARRY_IN_BITS  :0] ),
            .CarryOutDelayMXH (  CarryDeltaDelayMXH[g_order]  [CARRY_IN_BITS  :0] )
         );
      end : FLOPS
   end : MASH_CARRY_BLOCKS

///========================================================================================================
/// Ratio Generation
///========================================================================================================
   
   logic [10:0] ConstNMXH;
   logic signed [10:0] DeltaNMXH;

   // Define the constant N portion to be the MSB of the fraction (half
   // integer) and the ratio
   //
   always_comb begin : RATIO_IN_N
      //ConstNMXH = {ratio_async_mux__RatioMXH, ratio_async_mux__FractionMXH[FRAC_BITS-1]};
      ConstNMXH = {ratio_async_mux__RatioMXH, ratio_async_mux__FractionMXH[23]};
      // Sign extend
      DeltaNMXH = `ip2211ringpll_SX(CarryDeltaMXH[0], $bits(DeltaNMXH));
   end : RATIO_IN_N

   // Derive the ratio and half integer switch by combining the constant
   // portion and the delta N from the sigma delta
   //
   always_comb begin : RATIO_GEN
      {mash__RatioMXH, mash__HalfIntMXH} = ConstNMXH + DeltaNMXH;
   end : RATIO_GEN

///========================================================================================================
/// Assertions
///========================================================================================================

   `ifndef ip2211ringpll_SVA_OFF
      `ip2211ringpll_ASSERTS_MUST(R_mash_mod_illegal_delta_order_plus_one,
                    (integer'(DeltaNMXH)<=int'(1 << 2)) && (integer'(DeltaNMXH)> (-1 * int'(1 << 2))),
                    posedge ClkModMXH,
                    ResetXXL | (dfx__mash_order_plus_one != 1'b1),
                  `ip2211ringpll_ERR_MSG("[LJPLL] mash modulator is not operating correctly due to invalid delta for order 3"));
      
      `ip2211ringpll_ASSERTS_MUST(R_mash_mod_illegal_delta_order_plus_zero,
                    (integer'(DeltaNMXH)<=int'(1 << (1))) && (integer'(DeltaNMXH)> (-1 * int'(1 << (1)))),
                    posedge ClkModMXH,
                    ResetXXL | (dfx__mash_order_plus_one != 1'b0),
                  `ip2211ringpll_ERR_MSG("[LJPLL] mash modulator is not operating correctly due to invalid delta for order 2"));
   `endif

endmodule

`endif

`ifndef ip2211ringpll_TLCTRL_SIP_SV 
`define ip2211ringpll_TLCTRL_SIP_SV 

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "ljpll_dfx.vh"
//`include "ringpll_macros.sv"
`ifndef ip2211ringpll_SVA_OFF
//`include "intel_checkers.vs"
`endif

typedef enum logic [2:0] {
   TLFSM_X          = 3'bxxx,
   TLFSM_OFF        = 3'b000,
   TLFSM_TL         = 3'b001,
   TLFSM_PLL        = 3'b111,
   TLFSM_LL         = 3'b010
} t_TlCtrlFsm;

module ip2211ringpll_tlctrl_sip
(
   input  logic                ClkRefXXH,
   input  logic                reset_sync__Reset_b_XXnnnL,
   input  logic  	       dfx__tllm_en, 
   input  logic                lock_detector__EarlyLockXXnnnH,
   output logic                tlctrl_sip__LockRstXXnnnH,
   output logic [1:0]          tlctrl_sip__StateXXnnnH,
   output logic                tlctrl_sip__TightLoopXXnnnH,
   output logic                tlctrl_sip__GateClkDistXXnnnL,
   output logic                EarlyLockXXnnnH,
   input logic                idfx_fscan_clkungate
);




  logic tllm_prchg_mode;
  assign tllm_prchg_mode = 1'b0;  // This feature is not supported in RingPll

  logic [1:0] tllm_sw_latency;
  assign tllm_sw_latency = 2'b00;  // This feature is not supported in RingPll

///========================================================================================================
/// Reset generation 
///========================================================================================================
   
   logic ResetXXnnnL;

   always_comb begin : RESET_GEN
      ResetXXnnnL = ~reset_sync__Reset_b_XXnnnL;
   end : RESET_GEN

///========================================================================================================
/// Gated clock generation 
///========================================================================================================
   t_TlCtrlFsm      StateXXnnnH;
   logic            ClkRefGateXXH;
   logic            ClockEnXXnnnH;
   logic            ClockEnXXnnnL;

   // Enable the clock under the following conditions:
   //   -- TLLM is enabled and we are not in the  LL state
   //   -- TLLM is disabled and we are not in the OFF state 
   //   -- TLLM is in an intermediate state
   //
   always_comb ClockEnXXnnnH = (~dfx__tllm_en & (StateXXnnnH != TLFSM_OFF)) |
                               ( dfx__tllm_en & (StateXXnnnH != TLFSM_LL) ) |
                               ( (StateXXnnnH != TLFSM_OFF) &
                                 (StateXXnnnH != TLFSM_LL)                       ) ;

   `ip2211ringpll_LATCH_P(ClockEnXXnnnL, ClockEnXXnnnH, ClkRefXXH)
   // Disable the clock whenever we are in reset since everything
   //   downstream on ClkRefGateXXH is async reset.  This reduces power
   //   consumption when the circuit is in reset.
   //
//idfx_fscan_clkungate change added for scan
   `ip2211ringpll_CLKAND(ClkRefGateXXH, ClkRefXXH, ((ClockEnXXnnnL & reset_sync__Reset_b_XXnnnL) || idfx_fscan_clkungate))

///========================================================================================================
/// PLL Tight Loop Mode State Control FSM
///
///  The PLL tight loop mode state control FSM sequences through the
///   following states to enable the PLL to lock first in tight loop
///   and then in long loop.
///
///  TLFSM_OFF         : PLL is off or tight loop lock mode is not enabled.
///                      The FSM will remain in this state until the PLL is
///                      enabled and tight loop lock mode is enabled.
///
///  TLFSM_TL          : PLL has been enabled. Force tightloop. Depending on configured precharge mode,
///                      either gate clock to distribution (tllm_prchg_mode 1) or 
///                      inject PLL clock into distribution (tllm_prchg_mode 0).
///                      This state terminates on early lock acquisition.
///
///  TLFSM_PLL         : Early lock has been acquired in tight loop. Switch
///                      the distribution clock to ungated PLL clock. This
///                      state terminates after counting a number of BCLKs.
///
///  TLFSM_LL          : The distrubution is in "steady state", switch from
///                      tight loop to long loop.
///
///  The following is a summary of the FSM outputs and what they do.
///
///  TightLoopXXnnnH     : Forces tight loop when output is 1 
///  GateClkDistXXnnnH   : Gates the clock to distribution
///  LockReadyXXnnnH     : Indicates that the lock signals can pass
///                        directly to its fanout
///  LockRstXXnnnH       : Hold lock counter reset 
///  WaitCntEnXXnnnH     : Enable the wait counter for switching latency
///                        of TLFSM_PLL -> TLFSM_LL 
///  
///========================================================================================================
   
   t_TlCtrlFsm  NxtStateXXnnnH;
   logic        LockReadyXXnnnH;
   logic        WaitDoneXXnnnH;
   logic        WaitCntEnXXnnnH;
   logic        GateClkDistXXnnnH;

   always_comb begin : TLCTRL_FSM

      unique casez (StateXXnnnH)

         TLFSM_OFF : begin
            NxtStateXXnnnH                      = TLFSM_TL;
            GateClkDistXXnnnH                   = 1'b0;
            LockReadyXXnnnH                     = 1'b1;
            WaitCntEnXXnnnH                     = 1'b0;
         end

         TLFSM_TL  : begin
            NxtStateXXnnnH                      = lock_detector__EarlyLockXXnnnH ? TLFSM_PLL : StateXXnnnH;
            GateClkDistXXnnnH                   = tllm_prchg_mode;
            LockReadyXXnnnH                     = 1'b0;
            WaitCntEnXXnnnH                     = 1'b0;
         end

         TLFSM_PLL : begin
            NxtStateXXnnnH                      = WaitDoneXXnnnH ? TLFSM_LL : StateXXnnnH;
            GateClkDistXXnnnH                   = 1'b0;
            LockReadyXXnnnH                     = 1'b0;
            // This should actually come from an ISO'd DistPwrGoodRL
            //   WaitCntEnXXnnnH = powergood (dig) & sync(DistPwrGoodRL)
            //     This would allow you to potentially boot the pll before
            //     distpwrgood = 1
            WaitCntEnXXnnnH                     = 1'b1;
         end

         TLFSM_LL  : begin
            NxtStateXXnnnH                      = TLFSM_OFF;
            GateClkDistXXnnnH                   = 1'b0;
            LockReadyXXnnnH                     = 1'b1;
            WaitCntEnXXnnnH                     = 1'b0;
         end

         default   : begin
            `ifndef ip2211ringpll_SVA_OFF
//               `ip2211ringpll_ASSERTC_FORBIDDEN(Illegal_Case_select, !($isunknown(StateXXnnnH)), `ip2211ringpll_ERR_MSG("Illegal case selector: 'StateXXnnnH' = %h", StateXXnnnH));
            `endif
         `ifndef ip2211ringpll_NO_VCSSIM
         if (^(StateXXnnnH) === 1'bX) begin
            //NxtStateXXnnnH                      = 'x;
            NxtStateXXnnnH                      = TLFSM_X;
            GateClkDistXXnnnH                   = 'x;
            LockReadyXXnnnH                     = 'x;
            WaitCntEnXXnnnH                     = 'x;
         end else begin
         `endif
            NxtStateXXnnnH                      = TLFSM_OFF;
            GateClkDistXXnnnH                   = 1'b0;
            LockReadyXXnnnH                     = 1'b1;
            WaitCntEnXXnnnH                     = 1'b0;
         `ifndef ip2211ringpll_NO_VCSSIM
         end
         `endif
         end
      endcase
      
      // Glitch protect with encoding
      //
      tlctrl_sip__TightLoopXXnnnH         = StateXXnnnH[0];
      tlctrl_sip__LockRstXXnnnH           = StateXXnnnH[2];

   end : TLCTRL_FSM

   `ip2211ringpll_ASYNC_RSTD_MSFF(StateXXnnnH, NxtStateXXnnnH, ClkRefGateXXH, ResetXXnnnL, TLFSM_OFF)
   assign tlctrl_sip__StateXXnnnH = StateXXnnnH[1:0];

///========================================================================================================
/// Early Lock Override 
///========================================================================================================

   always_comb begin : EARLY_LOCK_OVERRIDE

      // Gate Lock To Downstream Logic
      //
      EarlyLockXXnnnH = (LockReadyXXnnnH) ? lock_detector__EarlyLockXXnnnH : 1'b0;
   
   end : EARLY_LOCK_OVERRIDE

///========================================================================================================
/// Wait Counter - Control Transition From TL -> LL 
///========================================================================================================

   logic [3:0] WaitCntXXnnnH;

   `ip2211ringpll_EN_ASYNC_RST_MSFF(WaitCntXXnnnH, WaitCntXXnnnH + 4'b1, ClkRefGateXXH, WaitCntEnXXnnnH, ResetXXnnnL)

   always_comb begin : WAIT_CNT_DECODE

      unique casez (tllm_sw_latency[1:0])
         2'b00 :  WaitDoneXXnnnH = (WaitCntXXnnnH[0]   == 1'd1);  // Ref * 2
         2'b01 :  WaitDoneXXnnnH = (WaitCntXXnnnH[1:0] == 2'd3);  // Ref * 4
         2'b10 :  WaitDoneXXnnnH = (WaitCntXXnnnH[2:0] == 3'd7);  // Ref * 8
         2'b11 :  WaitDoneXXnnnH = (WaitCntXXnnnH[3:0] == 4'd15); // Ref * 16
         `ip2211ringpll_XDefault(WaitDoneXXnnnH)
      endcase
   
   end : WAIT_CNT_DECODE

///========================================================================================================
/// Convert GateClkDist to Low Phase ClkRef
///========================================================================================================

   logic ClkRefXXH_b;
   
   // Drive GateClkDist out on low phase in order to receive the ungate
   //   signal deterministically in the HIP
   //
   `ip2211ringpll_CLKINV(ClkRefXXH_b, ClkRefXXH)
   `ip2211ringpll_ASYNC_RST_LATCH(tlctrl_sip__GateClkDistXXnnnL, GateClkDistXXnnnH, ClkRefXXH_b, ResetXXnnnL)

///========================================================================================================
/// SV Assertions
///========================================================================================================

`ifndef ip2211ringpll_SVA_OFF
   // Check that EarlyLockQual does not glitch - this SVA is pretty useless
   //
   `ip2211ringpll_ASSERTS_GRAY_CODE(GLITCH_tlfsm_earlylockqual, {lock_detector__EarlyLockXXnnnH, StateXXnnnH[0]}, posedge ClkRefXXH, ~reset_sync__Reset_b_XXnnnL, `ip2211ringpll_ERR_MSG("EarlyLockQualXXnnnH has glitched - driver is in ip2211ringpll_tlctrl_sip"));

   // Check that the gate distribution signal asserts when precharge mode
   // is 1 and the FSM is in Tight Loop
   //
   `ip2211ringpll_ASSERTS_MUST(R_tlfsm_gate_dist_clk_when_prchg_1, (tlctrl_sip__GateClkDistXXnnnL | ~tllm_prchg_mode | StateXXnnnH!=TLFSM_TL), posedge ClkRefXXH, ~reset_sync__Reset_b_XXnnnL, `ip2211ringpll_ERR_MSG("Tight Loop Lock Mode FSM not gating the clock distribution when requested!"));
   
   // Check that the gate distribution signal is 0 when the FSM is not in
   // the TL state
   //
   `ip2211ringpll_ASSERTS_MUST(R_tlfsm_gate_dist_clk_outside_tight_loop, (~tlctrl_sip__GateClkDistXXnnnL | StateXXnnnH==TLFSM_TL), posedge ClkRefXXH, ~reset_sync__Reset_b_XXnnnL, `ip2211ringpll_ERR_MSG("Tight Loop Lock Mode FSM is gating the clock when the FSM is not in the tight loop mode!"));

`endif


endmodule // module ip2211ringpll_tlctrl_sip

`endif // ip2211ringpll_TLCTRL_SIP_SV 


`ifndef ip2211ringpll_GLOBAL_ALIGN_SV
`define ip2211ringpll_GLOBAL_ALIGN_SV

module ip2211ringpll_global_align (
   input  logic tlctrl_sip__GateClkDistXXnnnL,
   //input  logic dfx__GlobalAlignXXL,
   output logic global_align__GateClkDistXXnnnL
);


   always_comb begin : GLOBAL_ALIGN
       // Uncomment this OR gate when DFX GlobalAlign is used. - 03-02-2017
      //global_align__GateClkDistXXnnnL = dfx__GlobalAlignXXL | tlctrl_sip__GateClkDistXXnnnL;
      global_align__GateClkDistXXnnnL = tlctrl_sip__GateClkDistXXnnnL;
   end : GLOBAL_ALIGN


endmodule

`endif


//`celldefine
`ifndef ip2211ringpll_LJPLL_SIP_SV
`define ip2211ringpll_LJPLL_SIP_SV

`ifndef ip2211ringpll_SVA_OFF
//`include "intel_checkers.vs"
`endif
//`include "soc_macros.sv"
//`include "ljpll_dfx.vh"

//`include "reg_req_ack.sv"
//`include "sync_reset_clkgen.sv"
//`include "ratio_async_mux.sv"
//`include "lock_detector.sv"
//`include "unlock_counter.sv"
//`include "ljpll_reset_sync.sv"
//`include "ljpll_dfx.sv"
//`include "lock_timer.sv"
//`include "startup_gen.sv"
//`include "vctl_trim_fsm.sv"
//`include "idv_fublet.sv"
//`include "ljpll_idv.sv"
//`include "adc_ctl.sv"
//`include "ssc_mod_dfx.sv"
//`include "ssc_mod.sv"
//`include "mash_mod.sv"
//`include "tlctrl_sip.sv"
//`include "global_align.sv"
////`include "cp_ctrl_block.sv"
////`include "lpf_ctrl_block.sv"
////`include "iref_ctrl_block.sv"

module ip2211ringpll_ljpll_sip 
//#(                 parameter RATIO_BITS    = 10,
//                   parameter FRAC_BITS     = 24,
//                   parameter MASH_ORDER    = 2,
//                   parameter IDV_ADDR_BITS = 10,
//                   parameter IDV_CB_BITS   = 2,
//                   parameter IDV_PG_BITS   = 2,
//                   parameter FMOD_BITS     = 9,
//                   parameter bit SSC_EN    = 1,
//                   parameter bit TLLM_EN   = 1)
 (
   input  logic                         ClkRefXXH,
   input  logic                         Reset_b_NnnnH,
   input  logic                         PllDistPwrGoodNnnnH,
   input  logic                         BypassNnnnH,
   input  logic [9:0]    		RatioNnnnH,
   input  logic [23:0]    		FractionNnnnH,
   input  logic                         pll_fbgen__ClkFbMXH,
   input  logic                         pll_core__PfdLockRstNnnnH,
   input  logic [9:0]                   view_adc__dig_out,
   input  logic                         view_adc__done,
//   input  logic                         pllen,                  // new -nd

   output logic                         reset_sync__BypassXXnnnL,
   output logic                         reset_sync__Reset_b_XXnnnL,
   output logic                         reset_sync__BypassEnXXnnnL,
   output logic                         dfx__powergood,
   output logic				dfx__reset_b,

   output logic [1:0]                   dfx__ViewDigEnNnnnH,
   output logic [1:0]                   dfx__ViewAnaEnNnnnH,
   output logic [1:0] [4:0]             dfx__ViewSelNnnnH,
   input  logic [1:0]                   view_mux__ViewOutNnnnH,
   output logic                         ssc__DirectionMXH,
   output logic [9:0]    		mash__RatioMXH,
   output logic                         mash__HalfIntMXH,

   // IDV control bits
   //
   output logic                         idv_fub__IdvGateEnNH,
   output logic [3:0]                   idv__RdacCtlTH,
   output logic [3:0]                   idv__PgCtlTH,
   output logic [2:0]                   idv__CbCtlTH,

   output logic                         startup_gen__VctlRdacEnXXH,
   output logic                         startup_gen__PfdEnXXH,
   output logic                         vctl_trim_fsm__VctlRdacShortXXH,
   output logic                         EarlyLockXXnnnH,
   output logic                         LockXXnnnL,

   // TAP programming to SIP via RTDR-DFX modules.
   //
   //input  t_ljpll_dfx_in_ifc            dfx_in,
   //output t_ljpll_dfx_out_ifc           dfx_out,
   input  t_ljpll_tap_in_ifc            tap_in,
   output t_ljpll_tap_out_ifc           tap_out,

   input  logic                         ClkIdvIH,

   // View Signals to HIP
   //
   output logic                         lock_detector__RawLockXXnnnL,
   output logic                         ssc_mod_dfx__ClkModMXH,

   // Tap decode to HIP
   //
   output logic                         adc_ctl__StartXXH,
   output logic                         adc_ctl__Reset_bXXL,
   output logic [1:0]                   dfx__adc_clkdiv,
   output logic                         dfx__adc_freeze,
   output logic                         dfx__adc_chop_en,
   output logic                         dfx__adc_use_vref,
   output logic [2:0]                   dfx__adc_sel_in,

   // Fuse decode to HIP
   //
   output logic                         dfx__tight_loop,
   output logic [4:0]                   dfx__cp1_trim,
   output logic [4:0]                   dfx__cp2_trim,
   output logic [4:0]                   dfx__skadj_ctrl,
   output logic [3:0]                   dfx__lockthresh,
   output logic [5:0]                   dfx__dca_ctrl,
   output logic [1:0]                   dfx__dca_cb,

   // Tight loop lock mode
   //
   output logic                         tlctrl_sip__TightLoopXXnnnH,

//--------------------------------------------------------------------
   // Brought these in for over writing via TAP
   //
   input  logic                         fz_tight_loopb,         // Part of DFX_IN bus
   input  logic [4:0]                   fz_cp1trim,             // Part of DFX_IN bus
   input  logic [4:0]                   fz_cp2trim,             // Part of DFX_IN bus
   input  logic [1:0]                   fz_dca_cb,              // Part of DFX_IN bus
   input  logic [5:0]                   fz_dca_ctrl,            // Part of DFX_IN bus
   input  logic [2:0]                   fz_lockcnt,             // Part of DFX_IN bus
   input  logic                         fz_lockforce,           // Part of DFX_IN bus
   input  logic                         fz_lockstickyb,         // Part of DFX_IN bus
   input  logic [3:0]                   fz_lockthresh,          // Part of DFX_IN bus
   input  logic [4:0]                   fz_skadj,               // Part of DFX_IN bus
   input  logic [1:0]                   fz_cpnbias,        //NEW fuse: CP nbias tuning			// part of dfx_in
   input  logic [4:0]                   fz_irefgen,    //NEW fuse: Iref current			// part of dfx_in
   input  logic                         fz_nopfdpwrgate,   //NEW fuse: Disable ip2211ringpll_PFD power gating			// part of dfx_in
   input  logic                         fz_lpfclksel,      //NEW fuse: LPF clock selection			// part of dfx_in
   input  logic [1:0]                   fz_pfddly,         //NEW fuse: ip2211ringpll_PFD power gating delay section			// part of dfx_in
   input  logic [4:0]                   fz_spare,          //NEW fuse: spare bits			// part of dfx_in
   input  logic [5:0]                   fz_startup,    //NEW fuse: PLL startup circuit tuning			// part of dfx_in
   input  logic				fz_vcosel,
   input  logic [10:0]                  fz_vcotrim,        //NEW fuse: ip2211ringpll_VCO trim			// part of dfx_in
   input  logic [1:0]                   fz_ldo_vinvoltsel,      //new -nd			// part of dfx_in
   input  logic                         fz_ldo_bypass,          //new -nd			// part of dfx_in
   input  logic                         fz_ldo_extrefsel,       //new -nd			// part of dfx_in
   input  logic                         fz_ldo_faststart,       //new -nd			// part of dfx_in
   input  logic [3:0]                   fz_ldo_fbtrim,          //new -nd			// part of dfx_in
   input  logic [3:0]                   fz_ldo_reftrim,         //new -nd			// part of dfx_in
   input  logic [2:0]                   fz_pfd_pw,              // Part of DFX_IN bus

   input  logic                         mash_order_plus_one,    // Part of DFX_IN bus
   input  logic [8:0]                   ssc_cyc_to_peak_m1,         // Part of DFX_IN bus
   input  logic                         ssc_en,                 // Part of DFX_IN bus
   input  logic [23:0]                  ssc_frac_step,          // Part of DFX_IN bus

   input  logic                         ldo_enable,             //new -nd
   input  logic [5:0]                   mdiv_ratio,             //new -nd
   input  logic [1:0]                   vcodiv_ratio,           //new -nd
   input  logic [9:0]                   zdiv0_ratio,            //new -nd
   input  logic                         zdiv0_ratio_p5,         //new -nd
   input  logic [9:0]                   zdiv1_ratio,            //new -nd
   input  logic                         zdiv1_ratio_p5,         //new -nd
          // IDV interface
   input  logic                         idvdisable_bi,          // new -nd
   input  logic                         idvfreqai,              // new -nd
   input  logic                         idvfreqbi,              // new -nd
   input  logic                         idvpulsei,              // new -nd
   input  logic                         idvtclki,              // new -nd
   input  logic                         idvtctrli,             // new -nd
   input  logic                         idvtdi,                 // new -nd
   input  logic                         idvtresi,               // new -nd
//   input  logic                         clkidvih,               // new -nd

   output logic                         idvdisable_bo,  // part of dfx_out
   output logic                         idvfreqao,              // part of dfx_out
   output logic                         idvfreqbo,              // part of dfx_out
   output logic                         idvpulseo,              // part of dfx_out
   output logic                         idvtclko,               // part of dfx_out
   output logic                         idvtctrlo,              // part of dfx_out
   output logic                         idvtdo,         // part of dfx_out
   output logic                         idvtreso,               // part of dfx_out

   output logic                         dfx__ldo_enable_a,           // new -nd
   output logic                         dfx__ta_ldo_hiz_debug,       // new -nd
   output logic                         dfx__ta_ldo_idq_debug,       // new -nd
   output logic [4:0]                   dfx__ta_spare,               // new -nd
   output logic [1:0]                   dfx__fz_ldo_vinvoltsel_a,    // new -nd
   output logic                         dfx__fz_ldo_bypass_a,        // new -nd
   output logic                         dfx__fz_ldo_extrefsel_a,     // new -nd
   output logic                         dfx__fz_ldo_faststart_a,     // new -nd
   output logic [3:0]                   dfx__fz_ldo_fbtrim_a,        // new -nd
   output logic [3:0]                   dfx__fz_ldo_reftrim_a,       // new -nd
   output logic [5:0]                   dfx__mdiv_ratio_a,           // new -nd
   output logic [1:0]                   dfx__vcodiv_ratio_a,         // new -nd
   output logic [9:0]                   dfx__zdiv0_ratio_a,          //new -nd
   output logic                         dfx__zdiv0_ratio_p5_a,       //new -nd
   output logic [9:0]                   dfx__zdiv1_ratio_a,          //new -nd
   output logic                         dfx__zdiv1_ratio_p5_a,       //new -nd
   output logic [1:0]                   dfx__cpnbias,           //new -nd
   output logic [4:0]                   dfx__fz_irefgen_a,           //new -nd
   output  logic                        dfx__fz_lpfclksel_a,         //new -nd
   output  logic                        dfx__fz_nopfdpwrgate_a,      //new -nd
   output  logic [2:0]                  dfx__fz_pfd_pw_a,            //new -nd
   output  logic [1:0]                  dfx__fz_pfddly_a,            //new -nd
   output  logic [4:0]                  dfx__fz_spare_a,             //new -nd
   output  logic [5:0]                  dfx__fz_startup_a,           //new -nd
   output  logic                        dfx__fz_vcosel_a,            //new -nd
   output  logic [10:0]                 dfx__fz_vcotrim_a,           //new -nd

//--------------------------------------------------------------------
   // Global Alignment
   //
   output logic                         global_align__GateClkDistXXnnnL,
  //Scan interface
   input   logic [2:0]                   idfx_fscan_sdi,
   input   logic                         idfx_fscan_mode,
   input   logic                         idfx_fscan_shiften,
   input   logic                         idfx_fscan_rstbypen,
   input   logic                         idfx_fscan_byprstb,
   input   logic                         idfx_fscan_clkungate,
   output  logic [2:0]                   odfx_fscan_sdo

);

   //=============================================================================
   // Internal Wire Declaration
   //
   //    Declare wires for internal connectivity grouped by driver
   //=============================================================================

   // DFX
   //
   logic [14:0] 			     view_freq_count;
   t_ljpll_dfx_out_ifc           	     dfx_out;
   logic                                     dfx__bypass;
   logic [9:0] 				     dfx__RatioStepNH;
   logic [23:0]                              dfx__FracStepNH;
   logic                                     dfx__ssc_en;
   logic [1:0]                               dfx__ssc_mode;
   logic [8:0]                     	     dfx__ssc_cyc_to_peak_m1;
   logic                                     dfx__mash_order_plus_one;
   logic [9:0]                		     dfx__ratio;
   logic [23:0]                		     dfx__fraction;
//   logic [2:0]                               dfx__cp_mode;
//   logic [1:0]                               dfx__lpf_itrim;
//   logic [1:0]                               dfx__sr_lpf_mode;
   logic                                     dfx__GlobalAlignXXL;
   logic                                     dfx__openloop;
//   logic [3:0]                               dfx__startup_rdac;
   logic [3:0]                               dfx__vco_trim_pg;
   logic [2:0]                               dfx__vco_trim_cb;
//   logic [2:0]                               dfx__iref_mode;
//   logic [2:0]                               dfx__startcnt;
   logic                                     dfx__SscModTrigNH;
   logic  [1:0]                              dfx__SscModStepsNH;
   logic                                     dfx__SscDfxEnNH;
   logic  [1:0]                              dfx__SscModClkDivNH;
   logic                                     dfx__start_mode;
   logic                                     dfx__ratio_update_req;
   logic                                     dfx__ssc_prof_update_req;
   logic                                     dfx__disable_run_upd;
//   logic [10:0]                 	     dfx__fz_vcotrim_a;           //new -nd
   logic                                     dfx__tllm_en;		  //new -nd  fz_spare[3] is used.
   logic				     dfx__fz_lockforce_a;
   logic [2:0]				     dfx__fz_lockcnt_a;
   logic				     dfx__start_measurement;

   logic [3:0]				     dfx__ta_vctlrdac;
   logic				     dfx__ta_openloop2;

   // Startup Generator
   //
   logic                                     startup_gen__VctlTrimEnXXH;
   logic                                     startup_gen__ForcePullUpXXH;
   logic                         	     startup_gen__VctlRdacEnXXH_pre;
   logic                         	     startup_gen__PfdEnXXH_pre;

   // VCTL pump controller
   //
   logic                                     vctl_trim_fsm__TrimDoneXXH;
   //logic                                     vctl_trim_fsm__VctlRdacShortXXH;

   // IREF controller
   //
   logic                                    iref_ctrl__IrefDoneXXH;

   // Unlock Counter
   //
   logic [1:0]                               unlock_counter__UnlockCountXXnnnH;

   // Lock Timer
   //
   logic [11:0]                              lock_timer__LockTimeCntXXnnnH;

   // IDV Fublet
   //
   t_ljpll_idv_out_ifc                       idv_fub__idv_out;
   logic                                     idv_fub__IdvDisableTH;
   //logic [IDV_ADDR_BITS-1:0]                 idv_fub__IdvAddrTH;
   logic [9:0]                               idv_fub__IdvAddrTH;
   logic [3:0]                               idv__RdacCtlTH_pre;

   // Reg Req/Ack
   //
   logic                                     reg_req_ack__SscProfUpdReqMXH;
   logic                                     reg_req_ack__SscProfUpdAckMXH;
   logic                                     reg_req_ack__RatioUpdReqMXH;
   logic                                     reg_req_ack__RatioUpdAckMXH;
   logic                                     reg_req_ack__MashStateResetMXH;

   // Sync Reset Clkgen
   //
   logic                                     sync_reset_clkgen__ClkFbGateMXH;

   // SSC
   //
   logic [9:0]                               ssc__RatioMXH;
   logic [23:0]                              ssc__FractionMXH;
   logic                                     ssc__ProfUpdateMXH;
   logic                                     ssc__RatioUpdateMXH;

   // Ratio Async Mux
   //
   logic  [9:0]                              ratio_async_mux__RatioMXH;
   logic  [23:0]                             ratio_async_mux__FractionMXH;

   // MASH
   //
   logic                                     mash__PllModOnNH;

   // Lock Detector
   //
   logic                                     lock_detector__EarlyLockXXnnnH;

   // Tight loop lock mode
   logic                                     tlctrl_sip__LockRstXXnnnH_pre;
   logic                                     tlctrl_sip__TightLoopXXnnnH_pre;
   logic  [1:0]                              tlctrl_sip__StateXXnnnH_pre;
   logic                                     tlctrl_sip__GateClkDistXXnnnL_pre;

   logic                                     tlctrl_sip__LockRstXXnnnH;
   logic  [1:0]                              tlctrl_sip__StateXXnnnH;
   logic                                     tlctrl_sip__GateClkDistXXnnnL;

   logic                                     tlctrl_sip__EarlyLockXXnnnH;
   logic                                     reset_sync__Reset_b_XXnnnL_pre;

   // SSC DFX Module
   //
   logic                                     ssc_mod_dfx__TriggerRegXDH;
   logic                                     ssc_mod_dfx__ModulatorEnNH;

   logic 				     pll_core__CompOutNnnnH;
//   logic 				     cp_ctrl__cp_disable_fb_samp;
//   logic 				     cp_ctrl__cp_en_fb_amp;
//   logic 				     cp_ctrl__cp_sel_fb_amp;
//   logic 				     cp_ctrl__cp_iref_alt_mode;
   logic 				     lpf_ctrl__lpf_pg_en;
   logic [1:0] 				     lpf_ctrl__lpf_itrim;
   logic 				     vctl_trim_fsm__CmpEnXXH;
   logic 				     vctl_trim_fsm__PullUpNnnnH;
   logic 				     vctl_trim_fsm__PullDnNnnnH;

   logic 				     iref_ctrl__HighIModeNH;
   logic 				     iref_ctrl__RModeNH;
   logic 				     iref_ctrl__AmpDisableNH;
   logic 				     iref_ctrl__VcoClkSelNH;
   logic 				     iref_ctrl__VcoDiv16EnNH;
   logic 				     iref_ctrl__VcoDiv32EnNH;
//   logic 				     dfx__pfd_chop_en;
//   logic [2:0] 				     dfx__pfd_chop_val;
//   logic [1:0] 				     dfx__pvd_mode;
   logic [2:0] 				     dfx__pfd_residual_pw;
   logic 				     dfx__lockstickyb;
//   logic [2:0] 				     dfx__iref_ctune;
//   logic [3:0] 				     dfx__iref_ftune;
//   logic [3:0] 				     dfx__ro_freq_sel;
//   logic 				     dfx__lp_cp_en;


//ADC_CTL

   logic [1:0] 				     dfx__adc_start_cnt;
   logic 				     dfx__adc_start;

   logic                    vctl_trim_fsm__VctlRdacShortXXH_pre;
   // Tying LDO related tap signals
   //assign dfx__ta_ldo_hiz_debug = 1'b0;
   //assign dfx__ta_ldo_idq_debug = 1'b0;

   //=============================================================================
   // Submodule Declarations
   //
   //   Declare the top level SIP hierarchy of LJPLL
   //
   //   The top level hierarchy is as follows:
   //    -sip
   //    --ip2211ringpll_lock_detector
   //    --ip2211ringpll_lock_timer
   //    --dfx
   //    --reset_sync
   //    --startup_counter
   //    --tight loop lock control
   //=============================================================================

   // Lock Detector
   //   Detects the lock condition and generates a lock signal
   //
   ip2211ringpll_lock_detector ip2211ringpll_lock_detector
     (  
	.fz_lockforce                      (dfx__fz_lockforce_a),
	.fz_lockcnt                        (dfx__fz_lockcnt_a), 
	
	.ClkRefXXH                         (ClkRefXXH),
	.dfx__openloop                     (dfx__openloop),
	.dfx__GlobalAlignXXL               (dfx__GlobalAlignXXL),
	.pll_core__PfdLockRstNnnnH         (pll_core__PfdLockRstNnnnH),
	.reset_sync__Reset_b_XXnnnL        (reset_sync__Reset_b_XXnnnL),
	.reset_sync__BypassXXnnnL          (reset_sync__BypassXXnnnL),
	.reset_sync__BypassEnXXnnnL        (reset_sync__BypassEnXXnnnL),
	.startup_gen__PfdEnXXH             (dfx__reset_b),
	.tlctrl_sip__LockRstXXnnnH         (tlctrl_sip__LockRstXXnnnH),
	
	.lock_detector__RawLockXXnnnL      (lock_detector__RawLockXXnnnL),
	.lock_detector__EarlyLockXXnnnH    (lock_detector__EarlyLockXXnnnH),
	.LockXXnnnL                        (LockXXnnnL),
        .idfx_fscan_rstbypen               (idfx_fscan_rstbypen),
        .idfx_fscan_byprstb                (idfx_fscan_byprstb),
        .idfx_fscan_clkungate              (idfx_fscan_clkungate) 
     );

   // Lock Timer
   //   Starts when the PLL is enabled and counts the number of ref clocks that
   //   it takes before the lock condition is reached
   //
   ip2211ringpll_lock_timer ip2211ringpll_lock_timer
     (   
.* 
     );

   // Unlock Counter
   //    Counts up every time an unlock is detected - used for debug
   //
   ip2211ringpll_unlock_counter ip2211ringpll_unlock_counter  
     (   
.* 
     );

      // DFX Overrides
      //   Provides override muxes for various settings of the PLL
      //   for the purpose of DFX
      //
   ip2211ringpll_ljpll_dfx dfx  
	//	#(.RATIO_BITS(RATIO_BITS),
        //           .FRAC_BITS (FRAC_BITS),
        //           .FMOD_BITS(FMOD_BITS))         
 	//					dfx        ( .* );
     (  
//Inputs
//
	.tap_in                                (tap_in),
	.Reset_b_NnnnH                         (Reset_b_NnnnH),
	.PllDistPwrGoodNnnnH                   (PllDistPwrGoodNnnnH),
	.BypassNnnnH                           (BypassNnnnH),
	.RatioNnnnH                            (RatioNnnnH),
	.FractionNnnnH                         (FractionNnnnH),
	.unlock_counter__UnlockCountXXnnnH     (unlock_counter__UnlockCountXXnnnH),
	.lock_timer__LockTimeCntXXnnnH         (lock_timer__LockTimeCntXXnnnH),
	.lock_detector__RawLockXXnnnL          (lock_detector__RawLockXXnnnL),
	.tlctrl_sip__StateXXnnnH               (tlctrl_sip__StateXXnnnH),
	.view_adc__dig_out                     (view_adc__dig_out),
	.adc_ctl__StartXXH                     (adc_ctl__StartXXH),
	.view_adc__done                        (view_adc__done),
	.LockXXnnnL                            (LockXXnnnL),
	.mash__RatioMXH                        (mash__RatioMXH),
	.mash__HalfIntMXH                      (mash__HalfIntMXH),
	.ssc_mod_dfx__TriggerRegXDH            (ssc_mod_dfx__TriggerRegXDH),
	.ssc_mod_dfx__ModulatorEnNH            (ssc_mod_dfx__ModulatorEnNH),
	.iref_ctrl__IrefDoneXXH                (1'b0),
	.startup_gen__PfdEnXXH                 (startup_gen__PfdEnXXH),
        .view_freq_count                       (view_freq_count),
	.reset_sync__Reset_b_XXnnnL            (reset_sync__Reset_b_XXnnnL),
	.idv_fub__idv_out                      (8'b00000000),
	.reg_req_ack__RatioUpdAckMXH           (reg_req_ack__RatioUpdAckMXH),
	.reg_req_ack__SscProfUpdAckMXH         (reg_req_ack__SscProfUpdAckMXH),
	.view_mux__ViewOutNnnnH                (view_mux__ViewOutNnnnH),
	.fz_tight_loopb                        (fz_tight_loopb),
	.fz_cp1trim                            (fz_cp1trim),
	.fz_cp2trim                            (fz_cp2trim),
	.fz_dca_cb                             (fz_dca_cb),
	.fz_dca_ctrl                           (fz_dca_ctrl),
	.fz_lockcnt			       (fz_lockcnt),
	.fz_lockforce			       (fz_lockforce),
	.fz_lockstickyb                        (fz_lockstickyb),
	.fz_lockthresh                         (fz_lockthresh),
	.fz_skadj                              (fz_skadj),
	.fz_vcosel                             (fz_vcosel),
	.fz_cpnbias                            (fz_cpnbias),
	.fz_irefgen                            (fz_irefgen),
	.fz_nopfdpwrgate                       (fz_nopfdpwrgate),
	.fz_lpfclksel                          (fz_lpfclksel),
	.fz_pfddly                             (fz_pfddly),
	.fz_spare                              (fz_spare),
	.fz_startup                            (fz_startup),
	.fz_vcotrim                            (fz_vcotrim),
	.fz_ldo_vinvoltsel                     (fz_ldo_vinvoltsel),
	.fz_ldo_bypass                         (fz_ldo_bypass),
	.fz_ldo_extrefsel                      (fz_ldo_extrefsel),
	.fz_ldo_faststart                      (fz_ldo_faststart),
	.fz_ldo_fbtrim                         (fz_ldo_fbtrim),
	.fz_ldo_reftrim                        (fz_ldo_reftrim),
	.fz_pfd_pw                             (fz_pfd_pw),
	.mash_order_plus_one                   (mash_order_plus_one),
	.ssc_cyc_to_peak_m1                    (ssc_cyc_to_peak_m1),
	.ssc_en                                (ssc_en),
	.ssc_frac_step                         (ssc_frac_step),
	.ldo_enable                            (ldo_enable),
	.mdiv_ratio                            (mdiv_ratio),
	.vcodiv_ratio                          (vcodiv_ratio),
	.zdiv0_ratio                           (zdiv0_ratio),
	.zdiv0_ratio_p5                        (zdiv0_ratio_p5),
	.zdiv1_ratio                           (zdiv1_ratio),
	.zdiv1_ratio_p5                        (zdiv1_ratio_p5),
	
	// Outputs
	//
	.dfx_out                                (dfx_out),
	.tap_out                                (tap_out),
	.dfx__openloop                          (dfx__openloop),
	.dfx__ViewDigEnNnnnH                    (dfx__ViewDigEnNnnnH),
	.dfx__ViewAnaEnNnnnH                    (dfx__ViewAnaEnNnnnH),
	.dfx__ViewSelNnnnH                      (dfx__ViewSelNnnnH),
	.dfx__adc_clkdiv                        (dfx__adc_clkdiv),
	.dfx__adc_start                         (dfx__adc_start),
	.dfx__adc_start_cnt                     (dfx__adc_start_cnt),
	.dfx__adc_freeze                        (dfx__adc_freeze),
	.dfx__adc_chop_en                       (dfx__adc_chop_en),
	.dfx__adc_use_vref                      (dfx__adc_use_vref),
	.dfx__adc_sel_in                        (dfx__adc_sel_in),
	.dfx__GlobalAlignXXL                    (dfx__GlobalAlignXXL),
	.dfx__disable_run_upd                   (dfx__disable_run_upd),
	.dfx__mash_order_plus_one               (dfx__mash_order_plus_one),
	.dfx__ssc_en                            (dfx__ssc_en),
	//.dfx__ssc_mode                          (dfx__ssc_mode),
	//.dfx__cp_mode                           (dfx__cp_mode),
	//.dfx__lp_cp_en                          (dfx__lp_cp_en),
	//.dfx__lpf_itrim                         (dfx__lpf_itrim),
	//.dfx__sr_lpf_mode                       (dfx__sr_lpf_mode),
	//.dfx__startup_rdac                      (dfx__startup_rdac),
	//.dfx__iref_mode                         (dfx__iref_mode),
	//.dfx__startcnt                          (dfx__startcnt),
	.dfx__SscModTrigNH                      (dfx__SscModTrigNH),
	.dfx__SscModStepsNH                     (dfx__SscModStepsNH),
	.dfx__SscDfxEnNH                        (dfx__SscDfxEnNH),
	.dfx__SscModClkDivNH                    (dfx__SscModClkDivNH),
	//.dfx__start_mode                        (dfx__start_mode),
	.dfx__tight_loop                        (dfx__tight_loop),
	//.dfx__pfd_chop_en                       (dfx__pfd_chop_en),
	//.dfx__pfd_chop_val                      (dfx__pfd_chop_val),
	.dfx__pfd_residual_pw                   (dfx__pfd_residual_pw),
	.dfx__cp1_trim                          (dfx__cp1_trim),
	.dfx__cp2_trim                          (dfx__cp2_trim),
	.dfx__skadj_ctrl                        (dfx__skadj_ctrl),
	.dfx__fz_lockforce_a                    (dfx__fz_lockforce_a),
	.dfx__fz_lockcnt_a                      (dfx__fz_lockcnt_a),
	.dfx__lockthresh                        (dfx__lockthresh),
	.dfx__lockstickyb                       (dfx__lockstickyb),
	//.dfx__iref_ctune                        (dfx__iref_ctune),
	//.dfx__iref_ftune                        (dfx__iref_ftune),
	//.dfx__ro_freq_sel                       (dfx__ro_freq_sel),
	.dfx__dca_ctrl                          (dfx__dca_ctrl),
	.dfx__dca_cb                            (dfx__dca_cb),
	.dfx__tllm_en                           (dfx__tllm_en),
	//.dfx__RatioStepNH                       (dfx__RatioStepNH),
	.dfx__FracStepNH                        (dfx__FracStepNH),
	.dfx__ssc_cyc_to_peak_m1                (dfx__ssc_cyc_to_peak_m1),
	.dfx__ratio_update_req                  (dfx__ratio_update_req),
	.dfx__ssc_prof_update_req               (dfx__ssc_prof_update_req),
	.dfx__ldo_enable_a                      (dfx__ldo_enable_a),
        .dfx__ta_ldo_hiz_debug			(dfx__ta_ldo_hiz_debug),
        .dfx__ta_ldo_idq_debug			(dfx__ta_ldo_idq_debug),
        .dfx__ta_spare   			(dfx__ta_spare),
        .dfx__ta_vctlrdac			(dfx__ta_vctlrdac),
	.dfx__ta_openloop2			(dfx__ta_openloop2),
	.dfx__fz_ldo_vinvoltsel_a               (dfx__fz_ldo_vinvoltsel_a),
	.dfx__fz_ldo_bypass_a                   (dfx__fz_ldo_bypass_a),
	.dfx__fz_ldo_extrefsel_a                (dfx__fz_ldo_extrefsel_a),
	.dfx__fz_ldo_faststart_a                (dfx__fz_ldo_faststart_a),
	.dfx__fz_ldo_fbtrim_a                   (dfx__fz_ldo_fbtrim_a),
	.dfx__fz_ldo_reftrim_a                  (dfx__fz_ldo_reftrim_a),
	.dfx__mdiv_ratio_a                      (dfx__mdiv_ratio_a),
	.dfx__vcodiv_ratio_a                    (dfx__vcodiv_ratio_a),
	.dfx__zdiv0_ratio_a                     (dfx__zdiv0_ratio_a),
	.dfx__zdiv0_ratio_p5_a                  (dfx__zdiv0_ratio_p5_a),
	.dfx__zdiv1_ratio_a                     (dfx__zdiv1_ratio_a),
	.dfx__zdiv1_ratio_p5_a                  (dfx__zdiv1_ratio_p5_a),
	.dfx__cpnbias                           (dfx__cpnbias),
	.dfx__fz_irefgen_a                      (dfx__fz_irefgen_a),
	.dfx__fz_lpfclksel_a                    (dfx__fz_lpfclksel_a),
	.dfx__fz_nopfdpwrgate_a                 (dfx__fz_nopfdpwrgate_a),
	.dfx__fz_pfd_pw_a                       (dfx__fz_pfd_pw_a),
	.dfx__fz_pfddly_a                       (dfx__fz_pfddly_a),
	.dfx__fz_spare_a                        (dfx__fz_spare_a),
	.dfx__fz_startup_a                      (dfx__fz_startup_a),
	.dfx__fz_vcosel_a                       (dfx__fz_vcosel_a),
	.dfx__fz_vcotrim_a                      (dfx__fz_vcotrim_a),
	.dfx__start_measurement			(dfx__start_measurement),
	.dfx__reset_b                           (dfx__reset_b),
	.dfx__powergood                         (dfx__powergood),
	.dfx__bypass                            (dfx__bypass),
	.dfx__ratio                             (dfx__ratio),
	.dfx__fraction                          (dfx__fraction)
      );
   
      // Reset Syncronization
      //   Syncronization logic for the reset
      //
      //   This block allows the reset to drive asyncronously but will
      //   deassert reset syncronous to the reference clock
      //
      ip2211ringpll_ljpll_reset_sync reset_sync 
      (   
	  .ClkRefXXH			(ClkRefXXH),
	  .dfx__reset_b			(dfx__reset_b),
	  .dfx__bypass			(dfx__bypass),
	  .dfx__ldo_enable_a		(dfx__ldo_enable_a),
	  .ldo_timer			(dfx__fz_spare_a[1:0]),
	  .reset_sync__BypassXXnnnL	(reset_sync__BypassXXnnnL),
	  .reset_sync__Reset_b_XXnnnL	(reset_sync__Reset_b_XXnnnL_pre),
	  .reset_sync__BypassEnXXnnnL	(reset_sync__BypassEnXXnnnL),	
          .idfx_fscan_rstbypen               (idfx_fscan_rstbypen),
          .idfx_fscan_byprstb                (idfx_fscan_byprstb)
      );
   
      // Startup Counter
      //    Controls PLL startup by controlling the vctl rdac and charge pump
      //    enables. In addition, the IREF mode is also controlled from this
      //    unit.
      //
      ip2211ringpll_startup_gen ip2211ringpll_startup_gen
      (   
	  .ClkRefXXH			(ClkRefXXH),
	  .reset_sync__Reset_b_XXnnnL	(reset_sync__Reset_b_XXnnnL),
//	  .dfx__openloop			(dfx__openloop),
//	  .dfx__start_mode		(dfx__start_mode),
//	  .iref_ctrl__IrefDoneXXH		(iref_ctrl__IrefDoneXXH),
//	  .vctl_trim_fsm__TrimDoneXXH	(vctl_trim_fsm__TrimDoneXXH),
	
	  .startup_gen__ForcePullUpXXH	(startup_gen__ForcePullUpXXH),
	  .startup_gen__VctlTrimEnXXH	(startup_gen__VctlTrimEnXXH),
	  .startup_gen__VctlRdacEnXXH	(startup_gen__VctlRdacEnXXH_pre),
	  .startup_gen__PfdEnXXH	(startup_gen__PfdEnXXH_pre)
       );

      // If openloop2 TAP bit is set then drive values accordingly.
      // This gives a way to test ip2211ringpll_VCO openloop in regular TAP mode, in addition to the IDV openloop test.
      // The testchip won't have an IDV chain.
      //
	  assign startup_gen__VctlRdacEnXXH = dfx__ta_openloop2 ? 1'b1 : startup_gen__VctlRdacEnXXH_pre;
	  assign startup_gen__PfdEnXXH      = dfx__ta_openloop2 ? 1'b0 : startup_gen__PfdEnXXH_pre;


      // Charge Pump Controller
      //   This is a swappable block that can drive controls to the charge
      //   pump through the HIP interface.  All logic controlling the
      //   charge pump based on PLL state is inside this block.
      //
      //cp_ctrl_block                               cp_ctrl          ( .* );

      // IREF Controller
      //   This block controls the IREF startup counter and IREF mode. The
      //   IREF always starts on PLL enable
      //
      //iref_ctrl_block                             iref_ctrl        ( .* );

      // SR-LPF Controller
      //   This is a swappable block that can drive controls to the sample
      //   reset loop filter through the HIP interface.  All logic controlling the
      //   SR-LPF based on PLL state is inside this block.
      //
      //lpf_ctrl_block                              lpf_ctrl         ( .* );

      // IDV Fublet
      //    This block is the controller and address decode for IDV.  The IDV
      //    clock (from PLL PVD) feeds into this block to be distributed to
      //    the IDV chain.
      //
      //ip2211ringpll_idv_fublet  #(.IDV_ADDR_BITS(IDV_ADDR_BITS)) idv_fub         ( .dfx__idv_in ( dfx_in.idv ),
      ip2211ringpll_idv_fublet idv_fub
		//#(.IDV_ADDR_BITS(IDV_ADDR_BITS)) 
      (  
	 .* 
      );

      // LJPLL IDV
      //   This block decodes the IDV address for the LJPLL and sends the
      //   results to the AIP if IDV is enabled
      //
   assign dfx__vco_trim_pg = dfx__fz_vcotrim_a[9:6];
   assign dfx__vco_trim_cb = dfx__fz_vcotrim_a[2:0];

      ip2211ringpll_ljpll_idv                                   idv              ( 
			   	.dfx__openloop			(dfx__openloop),
   				//.dfx__startup_rdac		(dfx__startup_rdac),
   				.dfx__vco_trim_pg		(dfx__vco_trim_pg),
   				.dfx__vco_trim_cb		(dfx__vco_trim_cb),
   				.idv_fub__IdvAddrTH		(idv_fub__IdvAddrTH),
   				.idv_fub__IdvDisableTH		(idv_fub__IdvDisableTH),

   				//.idv__RdacCtlTH			(idv__RdacCtlTH),
   				.idv__RdacCtlTH			(idv__RdacCtlTH_pre),
   				.idv__CbCtlTH			(idv__CbCtlTH),
   				.idv__PgCtlTH			(idv__PgCtlTH)
				);

      // If openloop2 TAP bit is high then drive TAP vctlrdac[3:0] on output idv__RdacCtlTH bus. This
      // will override any settings from the IDV ip2211ringpll_VCO block.
      //
	assign idv__RdacCtlTH = dfx__ta_openloop2 ? dfx__ta_vctlrdac : idv__RdacCtlTH_pre;

//Mux added for scan
assign reset_sync__Reset_b_XXnnnL = idfx_fscan_rstbypen ? idfx_fscan_byprstb :  reset_sync__Reset_b_XXnnnL_pre;

      // LJPLL VCTL Trim FSM
      //   Controls the PLL startup sequence in any mode
      //
      ip2211ringpll_vctl_trim_fsm                               ip2211ringpll_vctl_trim_fsm    ( 
		.ClkRefXXH			(ClkRefXXH),
		.reset_sync__Reset_b_XXnnnL	(reset_sync__Reset_b_XXnnnL),
		.dfx__openloop			(dfx__openloop),
		.startup_gen__VctlTrimEnXXH	(startup_gen__VctlTrimEnXXH),
		.startup_gen__ForcePullUpXXH	(startup_gen__ForcePullUpXXH),
		.iref_ctrl__IrefDoneXXH		(1'b0),
		.pll_core__CompOutNnnnH		(1'b0),

		.vctl_trim_fsm__VctlRdacShortXXH (vctl_trim_fsm__VctlRdacShortXXH_pre),
		.vctl_trim_fsm__TrimDoneXXH	(vctl_trim_fsm__TrimDoneXXH),
		.vctl_trim_fsm__CmpEnXXH	(vctl_trim_fsm__CmpEnXXH),
		.vctl_trim_fsm__PullUpNnnnH	(vctl_trim_fsm__PullUpNnnnH),
		.vctl_trim_fsm__PullDnNnnnH	(vctl_trim_fsm__PullDnNnnnH),
                .idfx_fscan_byprstb             (idfx_fscan_byprstb),
                .idfx_fscan_rstbypen            (idfx_fscan_rstbypen) 
	 );

	// If openloop2 TAP bit is high then drive 1 on the following signal.
	//
      assign vctl_trim_fsm__VctlRdacShortXXH = dfx__ta_openloop2 ? 1'b1 : vctl_trim_fsm__VctlRdacShortXXH_pre;


      // ADC controller
      //   Controls the startup of the ADC inside the HIP
      //
      ip2211ringpll_adc_ctl ip2211ringpll_adc_ctl          
	( 
          .ClkRefXXH,

   	  .dfx__adc_start,
   	  .dfx__adc_start_cnt,

          .adc_ctl__StartXXH,
          .adc_ctl__Reset_bXXL,
          .idfx_fscan_rstbypen,
          .idfx_fscan_byprstb,
        .idfx_fscan_clkungate              (idfx_fscan_clkungate) 
	);

      // Reg Req/Ack Controller
      //   Controls the req/ack for register updates that occur when the PLL
      //   is enabled and locked.
      //
      ip2211ringpll_reg_req_ack ip2211ringpll_reg_req_ack      
	( 
	  .ssc_mod_dfx__ClkModMXH,
	  .LockXXnnnL,
	  .dfx__disable_run_upd,
	  .dfx__ratio_update_req,
	  .dfx__ssc_prof_update_req,
	  .ssc__ProfUpdateMXH,
	  .ssc__RatioUpdateMXH,
	  
	  .reg_req_ack__SscProfUpdReqMXH,
	  .reg_req_ack__SscProfUpdAckMXH,
	  .reg_req_ack__RatioUpdReqMXH,
	  .reg_req_ack__RatioUpdAckMXH,
	  .reg_req_ack__MashStateResetMXH
	);

      // Sync Reset Clkgen
      //   Used to generate a clock which can be used to reset syncronous
      //   flops that are clocked on the feedback clock in the SIP
      //
      ip2211ringpll_sync_reset_clkgen ip2211ringpll_sync_reset_clkgen
	( 
	  .ClkRefXXH,
	  .pll_fbgen__ClkFbMXH,
	  .reset_sync__BypassEnXXnnnL,
	  .EarlyLockXXnnnH,
	  .LockXXnnnL,	  
	  .sync_reset_clkgen__ClkFbGateMXH,
          .idfx_fscan_rstbypen,
          .idfx_fscan_byprstb,
        .idfx_fscan_clkungate              (idfx_fscan_clkungate) 
	);

      //if (SSC_EN) begin : SSC_MOD
      if (1'b1) begin : SSC_MOD
//         ip2211ringpll_ssc_mod 
//		//#(.RATIO_BITS(RATIO_BITS),
//                //   .FRAC_BITS(FRAC_BITS),
//                //   .FMOD_BITS(FMOD_BITS))         
//						ssc              ( .* );
         ip2211ringpll_ssc_mod ssc
	   (  
	      .ssc_mod_dfx__ClkModMXH		(ssc_mod_dfx__ClkModMXH),
	      .LockXXnnnL			(LockXXnnnL),
  
	      .dfx__RatioStepNH			(10'b0000000000),
	      .dfx__FracStepNH			(dfx__FracStepNH),
              .dfx__ssc_en			(dfx__ssc_en),
              .dfx__ssc_mode			(2'b00),
	      .dfx__ssc_cyc_to_peak_m1		(dfx__ssc_cyc_to_peak_m1),
              .reg_req_ack__SscProfUpdReqMXH	(reg_req_ack__SscProfUpdReqMXH),
              .reg_req_ack__SscProfUpdAckMXH	(reg_req_ack__SscProfUpdAckMXH),
              .reg_req_ack__RatioUpdReqMXH	(reg_req_ack__RatioUpdReqMXH),
              .reg_req_ack__RatioUpdAckMXH	(reg_req_ack__RatioUpdAckMXH),

	      .dfx__ratio			(dfx__ratio),
	      .dfx__fraction			(dfx__fraction),
	      .ssc__RatioMXH			(ssc__RatioMXH),
	      .ssc__FractionMXH			(ssc__FractionMXH),
              .ssc__DirectionMXH		(ssc__DirectionMXH),
	      .ssc__ProfUpdateMXH		(ssc__ProfUpdateMXH),
	      .ssc__RatioUpdateMXH		(ssc__RatioUpdateMXH)
	   );
      end : SSC_MOD
      else begin : NO_SSC


      ///=====================================================================================================================
      /// Ratio/Frac MUX
      ///=====================================================================================================================

        // Create a syncronizer for ratio/fb
        //
        `ip2211ringpll_EN_MSFF(ssc__RatioMXH, dfx__ratio, ssc_mod_dfx__ClkModMXH,       ssc__RatioUpdateMXH)
        `ip2211ringpll_EN_MSFF(ssc__FractionMXH, dfx__fraction, ssc_mod_dfx__ClkModMXH, ssc__RatioUpdateMXH)

         always_comb begin : SSC_PASS_THRU
            ssc__DirectionMXH    = 1'b0;
            ssc__ProfUpdateMXH   = 1'b0;
            ssc__RatioUpdateMXH  = ~LockXXnnnL | (reg_req_ack__RatioUpdReqMXH & ~reg_req_ack__RatioUpdAckMXH);
         end : SSC_PASS_THRU
      end : NO_SSC

      // Ratio Async Mux
      //   Allows dfx__ratio / dfx__fraction passthrough before lock so
      //   that syncronous flops on feedback clock can reset
      //
//      ip2211ringpll_ratio_async_mux  
//			//#(.RATIO_BITS(RATIO_BITS),
//                        //.FRAC_BITS(FRAC_BITS))   
//					ip2211ringpll_ratio_async_mux  ( .* );
      ip2211ringpll_ratio_async_mux  ip2211ringpll_ratio_async_mux  
	( 
          .reset_sync__BypassXXnnnL,
          .LockXXnnnL,
	  .dfx__ratio,
	  .ssc__RatioMXH,
	  .dfx__fraction,
	  .ssc__FractionMXH,
	  .ratio_async_mux__RatioMXH,
	  .ratio_async_mux__FractionMXH,
          .mdiv_ratio (dfx__mdiv_ratio_a)
	);

      //if ((FRAC_BITS>1) || SSC_EN) begin : MASH_MOD
      if ((24>1) || 1'b1) begin : MASH_MOD

      // SSC/FRAC-N DFX Module
      //   This IP provides DFX hooks for the frac-n/ssc modulators in
      //   order to debug this feature
      //
      ip2211ringpll_ssc_mod_dfx ip2211ringpll_ssc_mod_dfx
	( 
	  .sync_reset_clkgen__ClkFbGateMXH,
	  .LockXXnnnL,
	  .dfx__SscModTrigNH,
	  .dfx__SscModStepsNH,
	  .dfx__SscDfxEnNH,
	  .dfx__SscModClkDivNH,
	  .ssc_mod_dfx__TriggerRegXDH,
	  .ssc_mod_dfx__ModulatorEnNH,
	  .ssc_mod_dfx__ClkModMXH
	);

      // MASH modulator
      //   Adds FRAC-N capability to the PLL which is required for the SSC
      //   profiles requested in some SOC projects.  The SSC profile may
      //   have deltaR < 1
      //
//      ip2211ringpll_mash_mod 
//		//#(.FRAC_BITS(FRAC_BITS),
//                // .RATIO_BITS(RATIO_BITS),
//                // .ORDER(MASH_ORDER))              
//						mash             ( .* );

      ip2211ringpll_mash_mod mash 
	( 
	  .ssc_mod_dfx__ClkModMXH,
	  .LockXXnnnL,
	  .reg_req_ack__MashStateResetMXH,
	  .dfx__mash_order_plus_one,
	  .ratio_async_mux__RatioMXH,
	  .ratio_async_mux__FractionMXH,
	  .mash__RatioMXH,
	  .mash__HalfIntMXH,
	  .mash__PllModOnNH
	);

      end : MASH_MOD
      else begin : FRAC_ASSIGN

         assign ssc_mod_dfx__ClkModMXH = sync_reset_clkgen__ClkFbGateMXH;
         assign ssc_mod_dfx__TriggerRegXDH = 1'b0;
         assign ssc_mod_dfx__ModulatorEnNH = 1'b0;
         assign mash__RatioMXH   = ratio_async_mux__RatioMXH;
         assign mash__HalfIntMXH = ratio_async_mux__FractionMXH[23];
         assign mash__PllModOnNH = 1'b0;
      end : FRAC_ASSIGN


      //if (TLLM_EN) begin : TLLM_ENABLED
      // Tight loop lock mode control
      //   Tight loop lock mode FSM
      //
      ip2211ringpll_tlctrl_sip ip2211ringpll_tlctrl_sip
	( 
	  .ClkRefXXH(ClkRefXXH),
	  .reset_sync__Reset_b_XXnnnL(reset_sync__Reset_b_XXnnnL),
	  .dfx__tllm_en(dfx__tllm_en),
	  .lock_detector__EarlyLockXXnnnH(lock_detector__EarlyLockXXnnnH),
	  .tlctrl_sip__LockRstXXnnnH(tlctrl_sip__LockRstXXnnnH_pre),
	  .tlctrl_sip__StateXXnnnH(tlctrl_sip__StateXXnnnH_pre),
	  .tlctrl_sip__TightLoopXXnnnH(tlctrl_sip__TightLoopXXnnnH_pre),
	  .tlctrl_sip__GateClkDistXXnnnL(tlctrl_sip__GateClkDistXXnnnL_pre),
	  .EarlyLockXXnnnH(tlctrl_sip__EarlyLockXXnnnH),
        .idfx_fscan_clkungate              (idfx_fscan_clkungate) 
	  );
      //end : TLLM_ENABLED
      //else begin : TLLM_DISABLED
      //   assign tlctrl_sip__TightLoopXXnnnH       = 1'b0;
      //   assign tlctrl_sip__GateClkDistXXnnnL     = 1'b0;
      //   assign tlctrl_sip__LockRstXXnnnH         = 1'b0;
      //   assign tlctrl_sip__StateXXnnnH           = 2'b0;
      //   assign EarlyLockXXnnnH                   = lock_detector__EarlyLockXXnnnH;
      //end : TLLM_DISABLED

	// If TLLM is enabled then use the output of TLCTRL otherwise lock detector output.
	//
	// TLLM MUX
	//
	assign EarlyLockXXnnnH = (dfx__tllm_en) ? tlctrl_sip__EarlyLockXXnnnH : lock_detector__EarlyLockXXnnnH;
	assign tlctrl_sip__TightLoopXXnnnH = (dfx__tllm_en) ? tlctrl_sip__TightLoopXXnnnH_pre : 1'b0;
	assign tlctrl_sip__GateClkDistXXnnnL = (dfx__tllm_en) ? tlctrl_sip__GateClkDistXXnnnL_pre : 1'b0;
	assign tlctrl_sip__LockRstXXnnnH = (dfx__tllm_en) ? tlctrl_sip__LockRstXXnnnH_pre : 1'b0;
	assign tlctrl_sip__StateXXnnnH = (dfx__tllm_en) ? tlctrl_sip__StateXXnnnH_pre : 2'b00;



      // Global Alignment
      //   This IP ORs the external global alignment point with the gate
      //   signal from the Tight Loop Lock Mode SIP
      //
      ip2211ringpll_global_align ip2211ringpll_global_align
	( 
	  .tlctrl_sip__GateClkDistXXnnnL,
	  //.dfx__GlobalAlignXXL,
	  .global_align__GateClkDistXXnnnL
	);


   ///=========================================================================================
   // TAP measurement 
   // viewmux0 is being observed and count value is sent out on tap_out.
   // tap_out: logic [14:0]  view_freq_count
   // tap_in:  logic         start_measurement;   
   //
   
   logic        start_measurement_pre;
   logic 	start_measurement, measurement_refclk, measurement_viewclk;
   logic 	viewout0_clk;
   logic 	refclkcount_clk, viewclkcount_clk;
   logic 	refclkcountergate;
   logic 	refclk_cnt_rst, refclk_cnt_done, refclk_cnt_done_sticky;
   logic 	refclk_cnt_rst_pre;
   logic [7:0] 	refclk_cnt, refclk_cnt_next;
   logic [14:0] viewfreqcount;
   logic [14:0] viewout_cnt, viewout_cnt_next;
   logic 	localreset;
   logic 	localreset_pre;

   assign localreset_pre = dfx__reset_b;
 //Mux added for scan 
assign localreset = idfx_fscan_rstbypen ? idfx_fscan_byprstb : localreset_pre;
 
   assign viewout0_clk = view_mux__ViewOutNnnnH[0];
   
   // ip2211ringpll_MSFF to move from tck to refclk domain
   //
  
   assign start_measurement_pre = dfx__start_measurement & LockXXnnnL;
   `ip2211ringpll_ASYNC_RST_2MSFF_META(start_measurement, start_measurement_pre, ClkRefXXH, localreset)
   
   assign refclkcountergate = (start_measurement & ~refclk_cnt_done_sticky);
   //`ip2211ringpll_MAKE_CLK_GEN (refclkcount_clk, refclkcountergate, idfx_fscan_clkungate, ClkRefXXH)
 
 //idfx_fscan_clkungate control added for scan 
   `ip2211ringpll_MAKE_CLK_GEN (refclkcount_clk, refclkcountergate, idfx_fscan_clkungate , ClkRefXXH) 

   assign refclk_cnt_rst_pre = ~dfx__reset_b || ~start_measurement; 

   // Generate 128 refclk window to do measurements.
   //
   assign  refclk_cnt_next = refclk_cnt + 8'b00000001;
   `ip2211ringpll_ASYNC_RST_MSFF(refclk_cnt[7:0], refclk_cnt_next[7:0], refclkcount_clk, refclk_cnt_rst)
   assign refclk_cnt_done = (refclk_cnt == (8'd128 - 8'd1));//One less than 128
   `ip2211ringpll_ASYNC_RST_MSFF(refclk_cnt_done_sticky, (refclk_cnt_done_sticky | refclk_cnt_done), refclkcount_clk, refclk_cnt_rst)
  
 //Mux added for scan 
assign refclk_cnt_rst = idfx_fscan_rstbypen ? ~idfx_fscan_byprstb : refclk_cnt_rst_pre; 
 
   assign measurement_refclk = ~refclk_cnt_rst & ~refclk_cnt_done_sticky;
   
   // ip2211ringpll_MSFF to move from refclk to viewout[0] domain
   //
   `ip2211ringpll_ASYNC_RST_2MSFF_META(measurement_viewclk, measurement_refclk, viewout0_clk, localreset)

   // Count signal coming in on view bus bit 0 here.
   // Measure all rising edges that arrive while we are in 128 refcycle measurement window.
   //

   //`ip2211ringpll_MAKE_CLK_GEN (viewclkcount_clk, measurement_viewclk, idfx_fscan_clkungate, viewout0_clk)
 
 //idfx_fscan_clkungate control added for scan 
   `ip2211ringpll_MAKE_CLK_GEN (viewclkcount_clk, measurement_viewclk, idfx_fscan_clkungate , viewout0_clk) 

   assign  viewout_cnt_next = viewout_cnt + 15'b000000000000001;
   `ip2211ringpll_ASYNC_RST_MSFF(viewout_cnt[14:0], viewout_cnt_next[14:0], viewclkcount_clk, refclk_cnt_rst)

   // When refclk window is done then capture the viewout_cnt into a register on tck domain.
   //
   assign view_freq_count[14:0] = viewout_cnt[14:0]; 

///========================================================================================================
/// Assertions
///========================================================================================================
      `ifndef ip2211ringpll_SVA_OFF
      `ip2211ringpll_ASSERTS_MUST(R_ssc_mod_ratio_in_eq_ratio_out_at_en,
                        reset_sync__BypassXXnnnL | ({ssc__RatioMXH, ssc__FractionMXH} == {dfx__ratio, dfx__fraction}),
                        posedge (LockXXnnnL === 1'b1),
                        1'b0,
                     `ip2211ringpll_ERR_MSG("[LJPLL] SSC ratio out is not equal to ratio in at PLLEN when not in bypass mode"));
      `endif

endmodule

`endif
 

`ifndef ip2211ringpll_RINGPLL_SIP_SV
`define ip2211ringpll_RINGPLL_SIP_SV

`ifdef INTC_SYNTHESIS
`define ip2211ringpll_SVA_OFF 
`define ip2211ringpll_SVA_LIB_SVA2005 
`define ip2211ringpll_NO_VCSSIM
`define ip2211ringpll_INTC_NO_PWR_PINS
`endif

`ifndef ip2211ringpll_SVA_OFF
//`include "intel_checkers.vs"
`endif
//`include "soc_macros.sv"
//`include "ljpll_dfx.vh"

//`include "tcu_tpsb_stap_data_reg.sv"
//`include "ljpll_sip.sv"
////`include "ip22_ringpll_sip_defines.vh" // This is needed for Synthesis. 

module ip22_ringpll_sip 
//#(
//			parameter RATIO_BITS,
//                   	parameter FRAC_BITS,
//                   	parameter IDV_ADDR_BITS,
//                   	parameter FMOD_BITS,
//		   	parameter RTDR_WIDTH,
//			parameter SSC_EN,
//			parameter TLLM_EN,
//			parameter IDV_CB_BITS,
//                        parameter IDV_PG_BITS,
//		   	parameter TAP_OUT_WIDTH,
//		   	parameter TAP_IN_WIDTH)
 (
   `ifndef ip2211ringpll_INTC_NO_PWR_PINS
      input  wire                       vccdig,                 // Digital supply
      input  wire                       vss,                    // Ground
   `endif

   // LDO signals
   input  logic				ldo_enable,		//new -nd
   input  logic	[1:0]			fz_ldo_vinvoltsel,	//new -nd		// Part of DFX_IN bus
   input  logic				fz_ldo_bypass,		//new -nd		// Part of DFX_IN bus
   input  logic                         fz_ldo_extrefsel,	//new -nd		// Part of DFX_IN bus
   input  logic                         fz_ldo_faststart,	//new -nd		// Part of DFX_IN bus
   input  logic [3:0]                   fz_ldo_fbtrim,		//new -nd		// Part of DFX_IN bus
   input  logic [3:0]                   fz_ldo_reftrim,		//new -nd		// Part of DFX_IN bus

   input  logic [1:0]                   view_mux_viewoutnnnnh,

   input  logic                         pll_core_pfdlockrstnnnnh,
   input  logic                         pll_fbgen_clkfbmxh,
   input  logic                         clkrefxxh,
   input  logic                         bypassnnnnh,
   input  logic                         reset_b_nnnnh,

   input  logic                         plldistpwrgoodnnnnh,
   input  logic [9:0]    		rationnnnh,
   input  logic [23:0]    		fractionnnnnh,
   input  logic [5:0]    		mdiv_ratio,		//new -nd
   input  logic				mash_order_plus_one,    // Part of DFX_IN bus
   input  logic [8:0]			ssccyctopeakm1,     // Part of DFX_IN bus
   input  logic				ssc_en,    		// Part of DFX_IN bus
   input  logic [23:0] 			ssc_frac_step,		// Part of DFX_IN bus	

   input  logic [1:0]			vcodiv_ratio,		//new -nd
   input  logic [9:0]			zdiv0_ratio,		//new -nd
   input  logic 			zdiv0_ratio_p5,		//new -nd
   input  logic [9:0]			zdiv1_ratio,		//new -nd
   input  logic 			zdiv1_ratio_p5,		//new -nd
  
   input  logic [4:0]			fz_cp1trim,		// Part of DFX_IN bus
   input  logic [4:0]			fz_cp2trim,		// Part of DFX_IN bus
   input  logic [1:0]			fz_cpnbias,		// Part of DFX_IN bus
   input  logic [1:0]			fz_dca_cb,		// Part of DFX_IN bus
   input  logic [5:0]			fz_dca_ctrl,		// Part of DFX_IN bus
   input  logic [4:0]			fz_irefgen,		// Part of DFX_IN bus
   input  logic [2:0]			fz_lockcnt,		// Part of DFX_IN bus
   input  logic 			fz_lockforce,		// Part of DFX_IN bus
   input  logic 			fz_lockstickyb,		// Part of DFX_IN bus
   input  logic [3:0]			fz_lockthresh,		// Part of DFX_IN bus
   input  logic 			fz_lpfclksel,		// Part of DFX_IN bus
   input  logic 			fz_nopfdpwrgate,	// Part of DFX_IN bus
   input  logic [2:0]			fz_pfd_pw,		// Part of DFX_IN bus
   input  logic [1:0]			fz_pfddly,		// Part of DFX_IN bus
   input  logic [4:0]			fz_skadj,		// Part of DFX_IN bus

   input  logic [4:0]			fz_spare,		// Part of DFX_IN bus 
								//fz_spare[1:0] = LDO timer count
								//fz_spare[2] = disable_auto_bypass,
								//fz_spare[3] = TLLM Enable 
								//fz_spare[4] = free
								//
   input  logic [5:0]			fz_startup,		// Part of DFX_IN bus
   input  logic 			fz_tight_loopb,		// Part of DFX_IN bus
   input  logic 			fz_vcosel,		// Part of DFX_IN bus
   input  logic [10:0]			fz_vcotrim,		// Part of DFX_IN bus


  // IDV interface
   input  logic				idvdisable_bi,		// new -nd
   input  logic                         idvfreqai,		// new -nd
   input  logic                         idvfreqbi,		// new -nd
   input  logic                         idvpulsei,		// new -nd
   input  logic                         idvtclki,		// new -nd
   input  logic                         idvtctrli,		// new -nd
   input  logic                         idvtdi,			// new -nd
   input  logic                         idvtresi,		// new -nd

   output logic                         idvdisable_bo,	// part of dfx_out 
   output logic                         idvfreqao,		// part of dfx_out 
   output logic                         idvfreqbo,		// part of dfx_out 
   output logic                         idvpulseo,		// part of dfx_out 
   output logic                         idvtclko,		// part of dfx_out 
   output logic                         idvtctrlo,		// part of dfx_out 
   output logic                         idvtdo,		// part of dfx_out 
   output logic                         idvtreso,		// part of dfx_out 


   // RTDR interface
   //
   output logic                         tdo,
   input  logic                         tck,
   //input  logic                         sync_reset,
   input  logic                         tcapturedr, // stap_rtdr_capture tclkdr
   input  logic                         tdi,
   input  logic                         treg_en, // tap_rtdr_irdecoder_drselect
   input  logic                         trst_n, //stap_reset_b,
   input  logic                         tshiftdr,
   input  logic                         tupdatedr,


   input  logic [9:0]                   view_adc_dig_out,
   input  logic                         view_adc_done,
   input  logic				clkidvih,		// new -nd

   output logic				ldo_enable_a,		// new -nd
   output logic				ta_ldo_hiz_debug,	// new -nd
   output logic				ta_ldo_idq_debug,	// new -nd

   output logic [1:0]			fz_ldo_vinvoltsel_a,	// new -nd
   output logic				fz_ldo_bypass_a,	// new -nd
   output logic                         fz_ldo_extrefsel_a,     // new -nd
   output logic                         fz_ldo_faststart_a,     // new -nd
   output logic [3:0]                   fz_ldo_fbtrim_a,        // new -nd
   output logic [3:0]                   fz_ldo_reftrim_a,       // new -nd

   output logic                         dfx_powergood,

   output logic                         reset_sync_bypassxxnnnl,
   output logic                         reset_sync_bypassenxxnnnl,
   output logic                         reset_sync_reset_b_xxnnnl,

   output logic [9:0]    		mash_ratiomxh,
   output logic                         mash_halfintmxh,
   output logic [5:0]    		mdiv_ratio_a,		// new -nd

   output logic [1:0]    		vcodiv_ratio_a,		// new -nd
   output logic [9:0]			zdiv0_ratio_a,		//new -nd
   output logic 			zdiv0_ratio_p5_a,	//new -nd
   output logic [9:0]			zdiv1_ratio_a,		//new -nd
   output logic 			zdiv1_ratio_p5_a,	//new -nd

   output logic [4:0]			ta_spare,

   output logic                         idv_fub_idvgateennh,
   output logic [4:0]                   dfx_cp1_trim,
   output logic [4:0]                   dfx_cp2_trim,
   output logic [1:0]                   fz_cpnbias_a, 		//new -nd
   output logic [1:0]                   fz_dca_cb_a,
   output logic [5:0]                   dfx_dca_ctrl,
   output logic [4:0]			fz_irefgen_a,		//new -nd 



   output logic [3:0]                   dfx_lockthresh,
   output  logic 			fz_lpfclksel_a,		//new -nd	
   output  logic 			fz_nopfdpwrgate_a,	//new -nd
   output  logic [2:0]			fz_pfd_pw_a,		//new -nd
   output  logic [1:0]			fz_pfddly_a,		//new -nd
   output logic [4:0]                   dfx_skadj_ctrl,
   output  logic [4:0]			fz_spare_a,		//new -nd
   output  logic [5:0]			fz_startup_a,		//new -nd
   output logic                         dfx_tight_loop,
   output  logic 			fz_vcosel_a,		//new -nd
   output  logic [10:0]			fz_vcotrim_a,		//new -nd


   // Tight loop lock mode
   //
   output logic                         tlctrl_sip_tightloopxxnnnh,

   output logic                         adc_ctl_startxxh,
   output logic                         adc_ctl_reset_bxxl,
   output logic [1:0]                   dfx_adc_clkdiv,
   output logic                         dfx_adc_freeze,
   output logic                         dfx_adc_chop_en,
   output logic                         dfx_adc_use_vref,
   output logic [2:0]                   dfx_adc_sel_in,

   // LOCK signals
   //
   output logic                         lock_detector_rawlockxxnnnl,
   output logic                         lockxxnnnl,
   output logic                         earlylockxxnnnh,

   output logic [3:0]                   idv_rdacctlth,
   output logic                         startup_gen_vctlrdacenxxh,
   output logic                         startup_gen_pfdenxxh,

   output logic                         ssc_directionmxh,
   output logic                         ssc_mod_dfx_clkmodmxh,
   output logic                         vctl_trim_fsm_vctlrdacshortxxh,

   output logic [1:0]                   dfx_viewdigennnnnh,
   output logic [1:0]                   dfx_viewanaennnnnh,
   output logic [4:0]                   dfx_viewselnnnnh0,
   output logic [4:0]                   dfx_viewselnnnnh1,

   //Scan interface
   input   logic [2:0]                   idfx_fscan_sdi,
   input   logic                         idfx_fscan_mode,
   input   logic                         idfx_fscan_shiften,
   input   logic                         idfx_fscan_rstbypen,
   input   logic                         idfx_fscan_byprstb,
   input   logic                         idfx_fscan_clkungate,
   output  logic [2:0]                   odfx_fscan_sdo,

   // Global Alignment
   //
   output logic                         global_align_gateclkdistxxnnnl

);

   //=============================================================================
   // Internal Wire Declaration
   //
   //    Declare wires for internal connectivity grouped by driver
   //=============================================================================

//   logic                                     startup_gen__VctlTrimEnXXH;
   logic [3:0]                   idv__PgCtlTH;
   logic [2:0]                   idv__CbCtlTH;


   t_ljpll_tap_in_ifc            tap_in;
   t_ljpll_tap_out_ifc           tap_out;
       parameter RTDR_WIDTH = $bits(tap_in) + $bits(tap_out);
       parameter TAP_IN_WIDTH = $bits(tap_in);
       parameter TAP_OUT_WIDTH = $bits(tap_out);
   logic [RTDR_WIDTH - $bits(tap_out) - 1 : 0] data_out_dummy;
   logic [RTDR_WIDTH - $bits(tap_in) - 1 : 0] data_in_dummy;

   logic [10:0]                 fz_vcotrim_int;
//   logic 			pllen;

   // Delaying lock going to top level ringpll
   logic                         lock_int;
   logic                         lock_int1;
   logic                         lock_int2;
   logic                         lock_int3;
   logic                         lock_int4;
   logic			 dfx_reset_b;
   logic			 dfx_reset_b_pre;

   logic 			disable_auto_bypass;
   logic			reset_sync__BypassXXnnnL_int;

   //=============================================================================
   // Submodule Declarations
   //
   //   Declare the top level SIP hierarchy of LJPLL
   //
   //   The top level hierarchy is as follows:
   //    -ip22_ringpll_sip
   //    	--ip2211ringpll_ljpll_sip
   //    	--ip2211ringpll_tcu_tpsb_stap_data_reg
   //=============================================================================

// Name change, fuse mapping
//
assign fz_vcotrim_a[10]  = fz_vcotrim_int[10];  // Spare bit right now
assign fz_vcotrim_a[9:6] = idv__PgCtlTH;
assign fz_vcotrim_a[5:3] = fz_vcotrim_int[5:3]; 
assign fz_vcotrim_a[2:0] = idv__CbCtlTH; 
//assign pllen = reset_b_nnnnh;
//assign ta_spare = 5'b0;	// Assigning TAP spare bits to 0 for now.

//assign startup_gen__VctlTrimEnXXH = startup_gen_vctlrdacenxxh;

// AUTO BYPASS feature
// dfx_tight_loop=1 means full loop mode, disable auto bypass for full loop since
// we need the clock going out ungated in this case.
//
//assign disable_auto_bypass = fz_spare[2];
assign disable_auto_bypass = fz_spare[2] || dfx_tight_loop;


assign reset_sync_bypassxxnnnl = (reset_sync__BypassXXnnnL_int || (~(disable_auto_bypass || lock_int)));

wire [1:0][4:0] dfx__ViewSelNnnnH;
assign dfx_viewselnnnnh0[4:0] = dfx__ViewSelNnnnH[0][4:0]; 
assign dfx_viewselnnnnh1[4:0] = dfx__ViewSelNnnnH[1][4:0]; 

// Delay LOCK signal
// Lock is asserted with 1.5-cycle delay to allow smooth transition during auto-bypass
// from refclk to pllclk.
//
        `ip2211ringpll_ASYNC_RST_MSFF(lock_int1, lock_int, clkrefxxh, ~dfx_reset_b)
        `ip2211ringpll_ASYNC_RST_MSFF(lock_int2, lock_int1, clkrefxxh, ~dfx_reset_b)
        `ip2211ringpll_ASYNC_RST_MSFF(lock_int3, lock_int2, clkrefxxh, ~dfx_reset_b)
        `ip2211ringpll_ASYNC_RST_MSFF(lock_int4, lock_int3, clkrefxxh, ~dfx_reset_b)
        `ip2211ringpll_ASYNC_RST_MSFF(lockxxnnnl, lock_int4, clkrefxxh, ~dfx_reset_b)

assign dfx_reset_b = idfx_fscan_rstbypen ? idfx_fscan_byprstb : dfx_reset_b_pre;
	// SIP instantiation
	ip2211ringpll_ljpll_sip 
		   //#(.RATIO_BITS(RATIO_BITS),
                   //.FRAC_BITS (FRAC_BITS),
                   //.IDV_ADDR_BITS(10),
                   //.IDV_CB_BITS(2),
                   //.IDV_PG_BITS(2),
                   //.SSC_EN(SSC_EN),
                   //.FMOD_BITS(FMOD_BITS),
                   //.TLLM_EN(TLLM_EN)) 
	           // sip	(.*);

		sip (
                         .ClkRefXXH 			(clkrefxxh),
                         .Reset_b_NnnnH 		(reset_b_nnnnh),
                         .PllDistPwrGoodNnnnH		(plldistpwrgoodnnnnh),
                         .BypassNnnnH			(bypassnnnnh),
       			 .RatioNnnnH			(rationnnnh),
       			 .FractionNnnnH			(fractionnnnnh),
            		 //.ssc_cyc_to_peak_m1		(dfx__ssc_cyc_to_peak_m1),
                         .pll_fbgen__ClkFbMXH		(pll_fbgen_clkfbmxh),
                         .pll_core__PfdLockRstNnnnH	(pll_core_pfdlockrstnnnnh),
                       	 .view_adc__dig_out		(view_adc_dig_out),
                      	 .view_adc__done		(view_adc_done),
//                      	 .pllen				(reset_b_nnnnh),//pllen

                         //.reset_sync__BypassXXnnnL	(reset_sync__BypassXXnnnL),
                         .reset_sync__BypassXXnnnL	(reset_sync__BypassXXnnnL_int),
                         .reset_sync__Reset_b_XXnnnL	(reset_sync_reset_b_xxnnnl),
                      	 .reset_sync__BypassEnXXnnnL	(reset_sync_bypassenxxnnnl),
                         .dfx__powergood		(dfx_powergood),
			 .dfx__reset_b			(dfx_reset_b_pre),

                      	 .dfx__ViewDigEnNnnnH		(dfx_viewdigennnnnh),
                      	 .dfx__ViewAnaEnNnnnH		(dfx_viewanaennnnnh),
                 	 .dfx__ViewSelNnnnH		(dfx__ViewSelNnnnH),
                      	 .view_mux__ViewOutNnnnH	({view_mux_viewoutnnnnh[1],view_mux_viewoutnnnnh[0]}),
                      	 .ssc__DirectionMXH		(ssc_directionmxh),
       			 .mash__RatioMXH		(mash_ratiomxh),
                      	 .mash__HalfIntMXH		(mash_halfintmxh),

   			// IDV control bits
   			//
                      	 .idv_fub__IdvGateEnNH		(idv_fub_idvgateennh),
                      	 .idv__RdacCtlTH		(idv_rdacctlth),
                      	 .idv__PgCtlTH			(idv__PgCtlTH),
                      	 .idv__CbCtlTH			(idv__CbCtlTH),

                      	 .startup_gen__VctlRdacEnXXH	(startup_gen_vctlrdacenxxh),
                      	 .startup_gen__PfdEnXXH		(startup_gen_pfdenxxh),
                      	 .vctl_trim_fsm__VctlRdacShortXXH	(vctl_trim_fsm_vctlrdacshortxxh),
                      	 .EarlyLockXXnnnH		(earlylockxxnnnh),

                      	 //.LockXXnnnL			(LockXXnnnL),
                      	 .LockXXnnnL			(lock_int),

   			// TAP programming to SIP via RTDR-DFX modules.
   			//
               		 //.dfx_in			(dfx_in),
              	 	 //.dfx_out			(dfx_out),
          		 .tap_in			(tap_in),
          		 .tap_out			(tap_out),

                      	 .ClkIdvIH			(clkidvih),

   			// View Signals to HIP
   			//
                      	 .lock_detector__RawLockXXnnnL	(lock_detector_rawlockxxnnnl),
                      	 .ssc_mod_dfx__ClkModMXH	(ssc_mod_dfx_clkmodmxh),

   			// Tap decode to HIP
   			//
                      	 .adc_ctl__StartXXH		(adc_ctl_startxxh),
                      	 .adc_ctl__Reset_bXXL		(adc_ctl_reset_bxxl),
                      	 .dfx__adc_clkdiv		(dfx_adc_clkdiv),
                      	 .dfx__adc_freeze		(dfx_adc_freeze),
                      	 .dfx__adc_chop_en		(dfx_adc_chop_en),
                      	 .dfx__adc_use_vref		(dfx_adc_use_vref),
                      	 .dfx__adc_sel_in		(dfx_adc_sel_in),

                         .dfx__tight_loop		(dfx_tight_loop),
                      	 .dfx__cp1_trim			(dfx_cp1_trim),
                      	 .dfx__cp2_trim			(dfx_cp2_trim),
                      	 .dfx__skadj_ctrl		(dfx_skadj_ctrl),
                      	 .dfx__lockthresh		(dfx_lockthresh),
                         .dfx__dca_ctrl			(dfx_dca_ctrl),
                      	 .dfx__dca_cb			(fz_dca_cb_a),

   			// Tight loop lock mode
   			//
                      	 .tlctrl_sip__TightLoopXXnnnH	(tlctrl_sip_tightloopxxnnnh),
		     
 			//--------------------------------------------------------------------
   			// Brought these in for over writing via TAP
   			//
		     	.fz_tight_loopb			(fz_tight_loopb),	// Part of DFX_IN bus
			.fz_cp1trim			(fz_cp1trim),		// Part of DFX_IN bus
			.fz_cp2trim			(fz_cp2trim),		// Part of DFX_IN bus
			.fz_dca_cb			(fz_dca_cb),		// Part of DFX_IN bus
			.fz_dca_ctrl			(fz_dca_ctrl),		// Part of DFX_IN bus
			.fz_lockcnt			(fz_lockcnt),		// Part of DFX_IN bus
			.fz_lockforce			(fz_lockforce),		// Part of DFX_IN bus
			.fz_lockstickyb			(fz_lockstickyb),	// Part of DFX_IN bus
			.fz_lockthresh			(fz_lockthresh),	// Part of DFX_IN bus
			.fz_skadj			(fz_skadj),		// Part of DFX_IN bus

                     	.fz_cpnbias			(fz_cpnbias),        	//NEW fuse: CP nbias tuning // part of dfx_in
                     	.fz_irefgen			(fz_irefgen),    	//NEW fuse: Iref current    // part of dfx_in
                     	.fz_nopfdpwrgate		(fz_nopfdpwrgate),   	//NEW fuse: Disable ip2211ringpll_PFD power gating                  // part of dfx_in
                     	.fz_lpfclksel			(fz_lpfclksel),      	//NEW fuse: LPF clock selection                       // part of dfx_in
                     	.fz_pfddly			(fz_pfddly),         	//NEW fuse: ip2211ringpll_PFD power gating delay section                    // part of dfx_in
                     	.fz_spare			(fz_spare),          	//NEW fuse: spare bits                        // part of dfx_in
                     	.fz_startup			(fz_startup),    	//NEW fuse: PLL startup circuit tuning                    // part of dfx_in
                     	.fz_vcotrim			(fz_vcotrim),        	//NEW fuse: ip2211ringpll_VCO trim                  // part of dfx_in
			.fz_vcosel			(fz_vcosel),
                     	.fz_ldo_vinvoltsel		(fz_ldo_vinvoltsel),      //new -nd                       // part of dfx_in
                     	.fz_ldo_bypass			(fz_ldo_bypass),          //new -nd                       // part of dfx_in
                     	.fz_ldo_extrefsel		(fz_ldo_extrefsel),       //new -nd                       // part of dfx_in
                     	.fz_ldo_faststart		(fz_ldo_faststart),       //new -nd                       // part of dfx_in
                     	.fz_ldo_fbtrim			(fz_ldo_fbtrim),          //new -nd                       // part of dfx_in
                     	.fz_ldo_reftrim			(fz_ldo_reftrim),         //new -nd                       // part of dfx_in
   		     	.fz_pfd_pw         		(fz_pfd_pw),

                     	.mash_order_plus_one 		(mash_order_plus_one),
                     	.ssc_cyc_to_peak_m1		(ssccyctopeakm1),
               	     	.ssc_en				(ssc_en),
                     	.ssc_frac_step			(ssc_frac_step),

  			// Brought these in for over writing via TAP
   			//
                        .ldo_enable			(ldo_enable),             //new -nd
                      	.mdiv_ratio			(mdiv_ratio),             //new -nd
                      	.vcodiv_ratio			(vcodiv_ratio),           //new -nd
                      	.zdiv0_ratio			(zdiv0_ratio),            //new -nd
                      	.zdiv0_ratio_p5			(zdiv0_ratio_p5),         //new -nd
                      	.zdiv1_ratio			(zdiv1_ratio),            //new -nd
                        .zdiv1_ratio_p5			(zdiv1_ratio_p5),         //new -nd

          		// IDV interface
                        .idvdisable_bi			(idvdisable_bi),          // new -nd
                        .idvfreqai			(idvfreqai),              // new -nd
                        .idvfreqbi			(idvfreqbi),              // new -nd
                        .idvpulsei			(idvpulsei),              // new -nd
                        .idvtclki			(idvtclki),              // new -nd
                        .idvtctrli			(idvtctrli),             // new -nd
                        .idvtdi				(idvtdi),                 // new -nd
                        .idvtresi			(idvtresi),               // new -nd
//                        .clkidvih			(clkidvih),               // new -nd

                        .idvdisable_bo			(idvdisable_bo),  // part of dfx_out
                      	.idvfreqao			(idvfreqao),              // part of dfx_out
                      	.idvfreqbo			(idvfreqbo),              // part of dfx_out
                      	.idvpulseo			(idvpulseo),              // part of dfx_out
                      	.idvtclko			(idvtclko),               // part of dfx_out
                      	.idvtctrlo			(idvtctrlo),              // part of dfx_out
                      	.idvtdo				(idvtdo),         // part of dfx_out
                      	.idvtreso			(idvtreso),               // part of dfx_out

                        .dfx__ldo_enable_a		(ldo_enable_a),           // new -nd
                        .dfx__ta_ldo_hiz_debug		(ta_ldo_hiz_debug),       // new -nd
                        .dfx__ta_ldo_idq_debug		(ta_ldo_idq_debug),       // new -nd
                        .dfx__ta_spare			(ta_spare),		  // new -nd
                      	.dfx__fz_ldo_vinvoltsel_a	(fz_ldo_vinvoltsel_a),    // new -nd
                        .dfx__fz_ldo_bypass_a		(fz_ldo_bypass_a),        // new -nd
                        .dfx__fz_ldo_extrefsel_a	(fz_ldo_extrefsel_a),     // new -nd
                        .dfx__fz_ldo_faststart_a	(fz_ldo_faststart_a),     // new -nd
                      	.dfx__fz_ldo_fbtrim_a		(fz_ldo_fbtrim_a),        // new -nd
                      	.dfx__fz_ldo_reftrim_a		(fz_ldo_reftrim_a),       // new -nd
                     	.dfx__mdiv_ratio_a		(mdiv_ratio_a),           // new -nd
                     	.dfx__vcodiv_ratio_a		(vcodiv_ratio_a),         // new -nd
                      	.dfx__zdiv0_ratio_a		(zdiv0_ratio_a),          //new -nd
                        .dfx__zdiv0_ratio_p5_a		(zdiv0_ratio_p5_a),       //new -nd
                      	.dfx__zdiv1_ratio_a		(zdiv1_ratio_a),          //new -nd
                        .dfx__zdiv1_ratio_p5_a		(zdiv1_ratio_p5_a),       //new -nd
                      	.dfx__cpnbias			(fz_cpnbias_a),           //new -nd
                      	.dfx__fz_irefgen_a		(fz_irefgen_a),           //new -nd
                        .dfx__fz_lpfclksel_a		(fz_lpfclksel_a),         //new -nd
                        .dfx__fz_nopfdpwrgate_a		(fz_nopfdpwrgate_a),      //new -nd
                     	.dfx__fz_pfd_pw_a		(fz_pfd_pw_a),            //new -nd
                     	.dfx__fz_pfddly_a		(fz_pfddly_a),            //new -nd
                     	.dfx__fz_spare_a		(fz_spare_a),             //new -nd
                     	.dfx__fz_startup_a		(fz_startup_a),           //new -nd
                        .dfx__fz_vcosel_a		(fz_vcosel_a),            //new -nd
                    	.dfx__fz_vcotrim_a		(fz_vcotrim_int),           //new -nd

   			// Global Alignment
   			//
                      	.global_align__GateClkDistXXnnnL	(global_align_gateclkdistxxnnnl),
                        .idfx_fscan_sdi               (idfx_fscan_sdi       ), 
                        .idfx_fscan_mode              (idfx_fscan_mode      ),
                        .idfx_fscan_shiften           (idfx_fscan_shiften   ),
                        .idfx_fscan_rstbypen          (idfx_fscan_rstbypen  ),
                        .idfx_fscan_byprstb           (idfx_fscan_byprstb   ),
                        .idfx_fscan_clkungate         (idfx_fscan_clkungate ), 
                        .odfx_fscan_sdo               (odfx_fscan_sdo       )

		);

        assign data_out_dummy = '0;
   
      	// RTDR - TAP
     	ip2211ringpll_tcu_tpsb_stap_data_reg #(
                          .DATA_REG_STAP_SIZE_OF_EACH_TEST_DATA_REGISTER(RTDR_WIDTH),
                          .DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS(0)
                              )  ljpll_rtdr (

                        .sync_reset(1'b0),
                        .ftap_tck(tck),
                        .ftap_tdi(tdi),
                        .reset_b(trst_n),
                        .stap_irdecoder_drselect(treg_en),
                        .stap_fsm_capture_dr(tcapturedr),
                        .stap_fsm_shift_dr(tshiftdr),
                        .stap_fsm_update_dr(tupdatedr),
                        .tdr_data_in({tap_out, tap_in}),
                        .data_reg_tdo(tdo),
                        .tdr_data_out({data_in_dummy,tap_in})
                        //.tdr_data_out(rtdr_data_out)
                        //.tdr_data_out()       // Disconnected and driven for testing by TB dut.tap_in. Connect it later. -
                                              );


///=========================================================================================
/// Assertions
///=========================================================================================

endmodule

`endif	// `ifdef ip22_ringpll_sip

// collage-pragma translate_on

//`celldefine		// For ICF delivery only.

`ifndef ip2211ringpll_RINGPLL_SV
`define ip2211ringpll_RINGPLL_SV

//UNINCLUDED DUE TO INWAY REQUIREMENTS //`include "Timescale.v"
//`include "ljpll_dfx.vh"

//`include "soc_macros.sv"
//`include "soc_clock_macros.sv"
//`include "soc_power_macros.sv"
//`include "ringpll_macros.sv"

`ifndef ip2211ringpll_SVA_OFF
//`include "intel_checkers.vs"
`endif

//`include "ip2211ringpll_hip.sv"
//UNINCLUDED DUE TO INWAY REQUIREMENTS //`include "ip22_ringpll_sip.sv"
//UNINCLUDED DUE TO INWAY REQUIREMENTS //`include "ldopgd.sv"

module ringpll
//#(
   //parameter bit SYNC_GEN_EN = 1,
   //parameter bit [4:0] SYNC_GEN_PIPE_STAGE = 5'd7,
   //parameter bit SSC_EN  = 1,
   //parameter bit TLLM_EN = 1,
   //parameter     RATIO_BITS = 10, 
   //parameter     FMOD_BITS = 9
//)
(

   `ifndef ip2211ringpll_INTC_NO_PWR_PINS
      input  			vnnaon_nom,             // Always ON supply
      input  			vccdig_nom,                 // Digital supply
      input  			vccldo_hv,                 // LDO input supply (1.1V nominal)
      input  			vccdist_nom,                // Digital supply for output clocks and clkpostdist input
      input  			vss,                	// Ground 
   `endif
   // LDO
   input	  	powergood_vnn,		// Power good control signal
   input    		ldo_vref,               //NEW PIN: LDO reference voltage (0.6v) (Domain: analog)
   input 	  	ldo_enable,          	//NEW PIN: Enable LDO
   input [1:0]                  fz_ldo_vinvoltsel,      //  fz_ldo_1p24v  //NEW PIN: set to 1 if using 1.24v ldo input
   input 			fz_ldo_faststart,       //NEW PIN: Enables LDO fast startup mode
   input 			fz_ldo_bypass,          //NEW PIN: Enables LDO bypass
   input 			fz_ldo_extrefsel,       //NEW PIN: Selects external voltage ref (ldo_vref)
   input [3:0]                  fz_ldo_fbtrim,          //NEW PIN: Adjust LDO feedback divider
   input [3:0]                  fz_ldo_reftrim,         //NEW PIN: Adjust LDO internal voltage ref

   input  			clkref,                 //ClkRefXXH,
   input  			bypass,                 //BypassNnnnH,
   input  			pllen,                  //Reset_b_NnnnH,
   input  			pllfwen_b,		// NEW: PLL Firewall enable (0 = output inactive)

   input  [9:0]                 ratio,                  //RatioNnnnH,  // parameter     RATIO_BITS = 10
   input  [23:0]                fraction,               //FractionNnnnH,
   input  [5:0]                 mdiv_ratio,             // NEW: Refclk divider 
   input 			mash_order_plus_one,    // dfx_in
   input  [8:0]                 ssc_cyc_to_peak_m1,     // SscCycToPeakm1,   //parameter     FMOD_BITS = 9
   input  			ssc_en,                 // dfx_in
   input  [23:0]                ssc_frac_step,          // dfx_in Frac delta/step
   input  [1:0]                 vcodiv_ratio,           // NEW: Post ip2211ringpll_VCO divider (1,2,4,8)
   input  [9:0]                 zdiv0_ratio,            // NEW: post pll divider for clkpll0 (N.5 dividerl max = 1024.5) // parameter     RATIO_BITS = 10
   input 			zdiv0_ratio_p5,         // NEW: point five for clkpll0
   input  [9:0]                 zdiv1_ratio,            // NEW: post pll divider for clkpll1 (N.5 dividerl max = 1024.5) // parameter     RATIO_BITS = 10
   input 			zdiv1_ratio_p5,         // NEW: point five for clkpll0

   // FUSES: input  t_ljpll_dfx_in_ifc       dfx_in,
   input [4:0]                 	fz_cp1trim,             //dfx_in_fuse_cp1_trim,
   input [4:0]                 	fz_cp2trim,             //dfx_in_fuse_cp2_trim,
   input [1:0]                  fz_cpnbias,             //NEW fuse: CP nbias tuning
   input [1:0]                  fz_dca_cb,              //dfx_in_fuse_dca_cb,
   input [5:0]                  fz_dca_ctrl,            //dfx_in_fuse_dca_ctrl,

   input [4:0]                  fz_irefgen,             //NEW fuse: Iref current
   input [2:0]                  fz_lockcnt,             //dfx_in_fuse_lockcnt,
   input 			fz_lockforce,           //dfx_in_fuse_tie_lockrst_zero,
   input 			fz_lockstickyb,         //NEW fuse: Lock detect sticky enable bar Fusedefault value = 0
   input [3:0]                  fz_lockthresh,          //dfx_in_fuse_lockthresh,
   input 			fz_lpfclksel,           //NEW fuse: LPF clock selection
   input 			fz_nopfdpwrgate,        //NEW fuse: Disable ip2211ringpll_PFD power gating
   input [2:0]                  fz_pfd_pw,              //dfx_in_fuse_pfd_residual_pw,
   input [1:0]                  fz_pfddly,              //NEW fuse: ip2211ringpll_PFD power gating delay section
   input [4:0]                 	fz_skadj,               //dfx_in_fuse_skadj_ctrl,
   input [4:0]                  fz_spare,               //NEW fuse: spare bits
   input [5:0]                  fz_startup,             //NEW fuse: PLL startup circuit tuning
   input 			fz_tight_loopb,         //dfx_in_fuse_tight_loop,
   input 			fz_vcosel,              //NEW fuse: ip2211ringpll_VCO select (0=low freq., 1=high freq range)
   input [10:0]                 fz_vcotrim,             //NEW fuse: ip2211ringpll_VCO trim

   // IDV
   input 			idvdisable_bi,
   input 			idvfreqai,
   input 			idvfreqbi,
   input 			idvpulsei,
   input 			idvtclki,
   input 			idvtctrli,
   input 			idvtdi,
   input 			idvtresi,
   // IDV output
   output 			idvdisable_bo,          //dfx_out_idv_idvdisable_bo,
   output 			idvfreqao,              //dfx_out_idv_idvfreqao,
   output 			idvfreqbo,              //dfx_out_idv_idvfreqbo,
   output 			idvpulseo,              //dfx_out_idv_idvpulseo
   output 			idvtclko,               //dfx_out_idv_idvtclko,
   output 			idvtctrlo,              //dfx_out_idv_idvtctrlo,
   output 			idvtdo,                 //dfx_out_idv_idvtdo,
   output 			idvtreso,               //dfx_out_idv_idvtreso,

   // RTDR interface
   //
   output 			tdo,
   input  			tck,
   input  			tcapturedr, 		//tclkdr, //stap_rtdr_irdecoder_drselect,
   input  			tdi,
   input  			treg_en, 		//stap_rtdr_capture,
   input  			trst_n, 		//stap_reset_b,
   input  			tshiftdr,
   input  			tupdatedr,

 //Scan interface
  input   [2:0]                 idfx_fscan_sdi,
  input   			idfx_fscan_mode,
  input   			idfx_fscan_shiften,
  input   			idfx_fscan_rstbypen,
  input   			idfx_fscan_byprstb,
  input   			idfx_fscan_clkungate,
  output  [2:0]                 odfx_fscan_sdo,

   //input ta_ldo_hiz_debug,
   //input ta_ldo_idq_debug,
   // updated interface to include analog output pins
   //
   //output t_ljpll_dfx_out_ifc      dfx_out
   //output tri [1:0]                     viewanabus,             //ViewAnaBusNH,
   output [1:0]                 viewanabus,             //ViewAnaBusNH,
   input  			clkpostdist,            //ClkPostDistMH,
   output 			lock,                   //LockXXnnnL,
   output 			clkpll,
   output 			clkpll0,		// NEW: zdiv0 output
   output 			clkpll1,		// NEW: zdiv1 output
   output [1:0]                 view_dig_out            //dfx_out_view_view_dig_out

);

//`ifdef INTEL_EMULATION
//logic [2:0] count;
//logic lck;
//always_ff@(posedge clkpll or negedge pllen) begin
//  
//	if(~pllen) begin
//	count = 3'b000;
//	lck = 1'b0;
//	end
//
//	else if (count < 3'b101 ) begin
//	count = count + 1'b1;
//    	lck = 1'b0;
//    	end
//
//	else begin 
//	count = count;
//	lck = 1'b1;
//	end
//
//end
//
//assign lock = lck;
//
//bit [31:0] num1;
//bit [31:0] num2;
//bit [31:0] num3;
//
//assign num1 = 32'h77359400;
//
//assign num2 = 32'h1dcd6500;
//
////assign num3 
//assign num3 = 32'h1dcd6500;
//
//  emu_clk_osc emu_ip22_ringpll_1 (
//        .enable(pllen),
//        .numerator(num1), //Need to fill in this from the clk_ref, ratio and half_int
//        .denominator(1'b1), //Need to fill in this from the clk_ref, ratio and half_int
//        .clk_out(clkpll1));
//
//  emu_clk_osc emu_ip22_ringpll_2 (
//        .enable(pllen),
//        .numerator(num2), //Need to fill in this from the clk_ref, ratio and half_int
//        .denominator(1'b1), //Need to fill in this from the clk_ref, ratio and half_int
//        .clk_out(clkpll0));
//
//  emu_clk_osc emu_ip22_ringpll_3 (
//        .enable(pllen),
//        .numerator(num3), //Need to fill in this from the clk_ref, ratio and half_int
//        .denominator(1'b1), //Need to fill in this from the clk_ref, ratio and half_int
//        .clk_out(clkpll));
//
//
//`else

`ifndef INTC_COLLAGE

/// HSD 1805126747 The bmod needs to have timing paths defined so that the timing extracted from the .lib (i.e. the SDF) 
/// can be correctly annotated for timing aware gate level simulations.

specify
        (clkref => clkpll) = (0:0:0, 0:0:0);
        (clkref => clkpll0) = (0:0:0, 0:0:0);
        (clkref => clkpll1) = (0:0:0, 0:0:0);
        (clkref => idvdisable_bo) = (0:0:0, 0:0:0);
        (clkref => idvfreqao) = (0:0:0, 0:0:0);
        (clkref => idvfreqbo) = (0:0:0, 0:0:0);
        (clkref => idvpulseo) = (0:0:0, 0:0:0);
        (clkref => idvtclko) = (0:0:0, 0:0:0);
        (clkref => idvtctrlo) = (0:0:0, 0:0:0);
        (clkref => idvtdo) = (0:0:0, 0:0:0);
        (clkref => idvtreso) = (0:0:0, 0:0:0);
        (clkref => lock) = (0:0:0, 0:0:0);
        (clkref => tdo) = (0:0:0, 0:0:0);
        (clkref => viewanabus[0]) = (0:0:0, 0:0:0);
        (clkref => viewanabus[1]) = (0:0:0, 0:0:0);
        (clkref => view_dig_out[1]) = (0:0:0, 0:0:0);
        (clkref => view_dig_out[0]) = (0:0:0, 0:0:0);
endspecify

///========================================================================================================
/// Local parameters
///========================================================================================================


   //=============================================================================
   // Internal Wire Declaration
   //
   //    Declare wires for internal connectivity grouped by driver
   //=============================================================================
   
   t_ljpll_dfx_in_ifc       dfx_in;
   t_ljpll_dfx_out_ifc      dfx_out;
   t_ljpll_tap_in_ifc       tap_in;
   t_ljpll_tap_out_ifc      tap_out;
 
      parameter RTDR_WIDTH = $bits(tap_in) + $bits(tap_out);
      parameter TAP_IN_WIDTH = $bits(tap_in);
      parameter TAP_OUT_WIDTH = $bits(tap_out);
      parameter DFX_IN_WIDTH = $bits(dfx_in);
      parameter DFX_OUT_WIDTH = $bits(dfx_out);
 
   logic [RTDR_WIDTH - $bits(tap_out) - 1 : 0] data_out_dummy;
   logic [RTDR_WIDTH - $bits(tap_in) - 1 : 0] data_in_dummy;
   //logic [RTDR_WIDTH-1:0] rtdr_data_out;


   // PLL core
   //
   logic       pll_core__PfdLockRstNnnnH;
   logic       pll_core__CompOutNnnnH;
   logic       ClkIdvIH;

   // ODCS
   //
   //logic       odcs_dig__odcsrisetrig;
   //logic       odcs_dig__odcsfalltrig;
   //logic [4:0] odcs_dll__DlyLineSettingNH;

   // OPSP
   //
   //logic       odcs_opsp__RiseSampNH;
   //logic       odcs_opsp__FallSampNH;

   // STM
   //
   //logic       stm_ifdim__StmTrigStatusNH;

   // Charge Pump Controller
   //
   logic                 cp_ctrl__cp_disable_fb_samp;
   logic                 cp_ctrl__cp_en_fb_amp;
   logic                 cp_ctrl__cp_sel_fb_amp;
   logic                 cp_ctrl__cp_iref_alt_mode;
  
   // SR LPF controller
   //
   logic                         lpf_ctrl__lpf_pg_en;
   logic [1:0]                   lpf_ctrl__lpf_itrim;

   // IREF controller
   //
   logic                         iref_ctrl__HighIModeNH;
   logic                         iref_ctrl__RModeNH;
   logic                         iref_ctrl__AmpDisableNH;
   logic                         iref_ctrl__VcoClkSelNH;
   logic                         iref_ctrl__VcoDiv16EnNH;
   logic                         iref_ctrl__VcoDiv32EnNH;


   // IDV controller to AIP
   //
   logic [3:0]                   idv__RdacCtlTH;
   logic [3:0]                   idv__PgCtlTH;
   logic [1:0]                   idv__CbCtlTH;

   // Startup Generator
   //
   logic                 startup_gen__VctlRdacEnXXH;
   logic                 startup_gen__PfdEnXXH;
  
   // VCTL pullup/pulldn controller
   //
   logic                 vctl_trim_fsm__CmpEnXXH;
   logic                 vctl_trim_fsm__VctlRdacShortXXH;
   logic                 vctl_trim_fsm__PullUpNnnnH;
   logic                 vctl_trim_fsm__PullDnNnnnH;

   // PLL Feedback Divider
   //
   logic                 pll_fbgen__ClkFbMXH;

   // View Pins
   //
   logic [1:0] view_mux__ViewOutNnnnH;

   // View ADC
   //
   logic [9:0] view_adc__dig_out;
   logic       view_adc__done;

   // Reset sync
   //
   logic reset_sync__BypassXXnnnL;
   logic reset_sync__Reset_b_XXnnnL;
   logic reset_sync__BypassEnXXnnnL;
 
   // Lock Detector
   //
   logic lock_detector__RawLockXXnnnL;
   logic EarlyLockXXnnnH;

   // SSC Modulator Clock Out
   //
   logic ssc_mod_dfx__ClkModMXH;

   // ADC control
   //
   logic                      adc_ctl__StartXXH;
   logic                      adc_ctl__Reset_bXXL;
  
   // SSC profile generator
   //
   logic                           ssc__DirectionMXH;

   // MASH modulator
   //
   logic [9:0] mash__RatioMXH;
   logic                           mash__HalfIntMXH;

   // IDV controller
   //
   logic idv_fub__IdvGateEnNH;

   // DFX unit to pllljhip
   //
//   t_ljpll_dfx_in_ifc   dfx_in;
//   t_ljpll_dfx_out_ifc  dfx_out;
//   t_ljpll_tap_in_ifc       ljpll_tap_in_ifc;
//   t_ljpll_tap_out_ifc      ljpll_tap_out_ifc;


   logic                      dfx__powergood;
   logic                      dfx__tight_loop;
   logic                      dfx__pfd_chop_en; 
   logic [2:0]                dfx__pfd_chop_val; 
   logic [1:0]                dfx__pvd_mode; 
   logic [2:0]                dfx__pfd_residual_pw;
   logic [4:0]                dfx__cp1_trim;
   logic [4:0]                dfx__cp2_trim;
   logic [4:0]                dfx__skadj_ctrl;
   logic [3:0]                dfx__lockthresh;
   logic [1:0]                dfx__adc_clkdiv;
   logic                      dfx__adc_freeze;
   logic                      dfx__adc_chop_en;
   logic                      dfx__adc_use_vref;
   logic [2:0]                dfx__adc_sel_in;
   logic [2:0]                dfx__iref_ctune;
   logic [3:0]                dfx__iref_ftune;
   logic [1:0]                dfx__ViewAnaEnNnnnH;
   logic [1:0]                dfx__ViewDigEnNnnnH;
   //logic [1:0] [4:0]          dfx__ViewSelNnnnH;
   logic [1:0]                viewdigennh;
   logic [1:0]                viewanaennh;
   logic [4:0]                viewsel0;
   logic [4:0]                viewsel1;

//   t_opsp_config              dfx__opsp_config;
//   logic [1:0]                dfx__odcs_tuner_cb;
   logic [3:0]                dfx__ro_freq_sel;
   logic [5:0]                dfx__dca_ctrl;
//   logic [1:0]                dfx__dca_cb;
   logic [1:0]                fz_dca_cb_a;
   logic                      dfx__lp_cp_en;


   // Tight loop lock control
   //
   logic                         tlctrl_sip__TightLoopXXnnnH;

   logic [4:0]                   ta_spare;

   // Global Alignment
   //
   //logic                         global_align__GateClkDistXXnnnL;
    logic			 tllm_gate_clk_trunk;    //connected to SIP:global_align__gateclkdistxxnnnl
   

   // LDO
   logic                  ta_ldo_hiz_debug;       // new -nd
   logic                  ta_ldo_idq_debug;       // new -nd
//   logic                  ldo_enable;             //new -nd
//   logic [1:0]            fz_ldo_vinvoltsel;      //new -nd
//   logic                  fz_ldo_bypass;          //new -nd
//   logic                  fz_ldo_extrefsel;       //new -nd
//   logic                  fz_ldo_faststart;       //new -nd
//   logic [3:0]            fz_ldo_fbtrim;          //new -nd
//   logic [3:0]            fz_ldo_reftrim;         //new -nd

  // New - ip22_ringpll_sip related
//   logic [5:0]                   mdiv_ratio;             //new -nd
//   logic [1:0]                   vcodiv_ratio;           //new -nd
//   logic [9:0]                   zdiv0_ratio;            //new -nd
//   logic                         zdiv0_ratio_p5;         //new -nd
//   logic [9:0]                   zdiv1_ratio;            //new -nd
//   logic                         zdiv1_ratio_p5;         //new -nd

//   logic                         idvdisable_bi;          // new -nd
//   logic                         idvfreqai;              // new -nd
//   logic                         idvfreqbi;              // new -nd
//   logic                         idvpulsei;              // new -nd
//   logic                         idvtclki;              // new -nd
//   logic                         idvtctrli;             // new -nd
//   logic                         idvtdi;                 // new -nd
//   logic                         idvtresi;               // new -nd

   logic                         clkidvih;               // new -nd
//   logic                         pllen;                  // new -nd

   logic                         ldo_enable_a;           // new -nd
   logic [1:0]                   fz_ldo_vinvoltsel_a;    // new -nd
   logic                         fz_ldo_bypass_a;        // new -nd
   logic                         fz_ldo_extrefsel_a;     // new -nd
   logic                         fz_ldo_faststart_a;     // new -nd
   logic [3:0]                   fz_ldo_fbtrim_a;        // new -nd
   logic [3:0]                   fz_ldo_reftrim_a;       // new -nd
   logic [5:0]                   mdiv_ratio_a;           // new -nd
   logic [1:0]                   vcodiv_ratio_a;         // new -nd
   logic [9:0]                   zdiv0_ratio_a;          //new -nd
   logic                         zdiv0_ratio_p5_a;       //new -nd
   logic [9:0]                   zdiv1_ratio_a;          //new -nd
   logic                         zdiv1_ratio_p5_a;       //new -nd

 //  logic [1:0]                   dfx__cpnbias;           //new -nd
   logic [1:0]                   fz_cpnbias_a;           //new -nd
   logic [4:0]                   fz_irefgen_a;           //new -nd
    logic                        fz_lpfclksel_a;         //new -nd
    logic                        fz_nopfdpwrgate_a;      //new -nd
    logic [2:0]                  fz_pfd_pw_a;            //new -nd
    logic [1:0]                  fz_pfddly_a;            //new -nd
    logic [4:0]                  fz_spare_a;             //new -nd
    logic [5:0]                  fz_startup_a;           //new -nd
    logic                        fz_vcosel_a;            //new -nd
    logic [10:0]                 fz_vcotrim_a;           //new -nd


   // LDO analog dft pins
   logic                         anadft_ldo;
   logic                         anadft_ldovref;
   logic                         anadft_ldovfb;

   logic			 powergood_vccdig;

   //=============================================================================
   // Submodule Declarations
   //
   //   Declare the top level hierarchy of LJPLL
   //
   //   The top level hierarchy is as follows:
   //    -ljpll
   //    --sip
   //    --hip
   //=============================================================================
// Following will go via SIP to RTDR to TDO
//   output logic                    dfx_out_tap_pll_enable,
//   output logic                    dfx_out_dist_pwr_good,
//   output logic                    dfx_out_iref_done,
//   output logic                    dfx_out_pfd_en,
//   output logic [1:0]                   dfx_out_unlock_count,
//   output logic [11:0]                   dfx_out_lock_time,
//   output logic [7:0]                   dfx_out_pll_ratio,
//   output logic                    dfx_out_pll_half_int,
//   output logic                    dfx_out_lock,
//   output logic                    dfx_out_raw_lock,
//   output logic [9:0]                   dfx_out_adc_dig_out,
//   output logic                    dfx_out_adc_start,
//   output logic                    dfx_out_adc_done,
//   output logic                    dfx_out_ssc_mod_dfx_run,
//   output logic                    dfx_out_ssc_mod_dfx_trig,
//   output logic [1:0]                   dfx_out_tctrlfsmstate,
   //=============================================================================

 


//     ip2211ringpll_tcu_tpsb_stap_data_reg #(
//                          .DATA_REG_STAP_SIZE_OF_EACH_TEST_DATA_REGISTER(RTDR_WIDTH),
//                          .DATA_REG_STAP_RESET_VALUES_OF_TEST_DATA_REGISTERS(0)
//                              )  ljpll_rtdr (
//   
//                	.sync_reset(1'b0),
//                        .ftap_tck(tck),
//                        .ftap_tdi(tdi),
//                        .reset_b(trst_n),
//                        .stap_irdecoder_drselect(tclkdr),
//                        .stap_fsm_capture_dr(treg_en),
//                        .stap_fsm_shift_dr(tshiftdr),
//                        .stap_fsm_update_dr(tupdatedr),
//                        .tdr_data_in({tap_out, data_out_dummy}),
//                        .data_reg_tdo(tdo),
//                        .tdr_data_out({data_in_dummy,tap_in})
//                        //.tdr_data_out(rtdr_data_out)
//                        //.tdr_data_out()	// Disconnected and driven for testing by TB dut.tap_in. Connect it later. -
//                                              );

	//assign tap_in = rtdr_data_out[TAP_IN_WIDTH-1:0];
	//assign tap_in = 185'b0; 

	assign powergood_vccdig = powergood_vnn; // level shifted from AON to vccdig domain


	// LDO
	//ip2211ringpll_ldopgd			iip2211ringpll_ldopgd (
	ip2211ringpll_ldopgd			ipll_ldo (
					`ifndef ip2211ringpll_INTC_NO_PWR_PINS
						.vnnaon_nom	(vnnaon_nom),
						.vccdig		(vccdig_nom),
						.vccldo		(vccldo_hv),
						.vccpll		(vccpll),
      			.vssx 		(vss),
					`endif
            .powergood_vccdig (powergood_vccdig), 
						.powergood_vnn		(powergood_vnn),
						.ldo_vref	        (ldo_vref),
						.viewana		(anadft_ldo),
						.fz_ldo_vinvoltsel	(fz_ldo_vinvoltsel_a),
						.fz_ldo_faststart	(fz_ldo_faststart_a),
						.clkref			(clkref),
						.fz_ldo_bypass		(fz_ldo_bypass_a),
						.fz_ldo_extrefsel	(fz_ldo_extrefsel_a),
						.fz_ldo_fbtrim		(fz_ldo_fbtrim_a),
						.fz_ldo_reftrim		(fz_ldo_reftrim_a),
            .fz_spare_4_strong_ladder_en (fz_spare_a[4]), //Need fix ,  instatiation was wrong 
						.ldo_enable		(ldo_enable_a),
   							// LDO analog dft pins
                				.anadft_ldovref		(anadft_ldovref),
                				.anadft_ldovfb		(anadft_ldovfb),
						.ta_ldo_hiz_debug	(ta_ldo_hiz_debug),
						.ta_ldo_idq_debug	(ta_ldo_idq_debug)
					);


      // Soft IP
      //   Synthesizable support logic for the LJPLL
      //   Includes (SIP + RTDR)
      ip22_ringpll_sip  
		   //#(.RATIO_BITS($bits(ratio)),
                   //.FRAC_BITS ($bits(fraction)),
		   //.RTDR_WIDTH(RTDR_WIDTH),
		   //.TAP_OUT_WIDTH(TAP_OUT_WIDTH),
		   //.TAP_IN_WIDTH(TAP_IN_WIDTH),
                   //.IDV_ADDR_BITS(10),
                   //.IDV_CB_BITS(2),
                   //.IDV_PG_BITS(2),
                   //.SSC_EN(1),
                   //.FMOD_BITS(9),
                   //.TLLM_EN(1))                 
				iip2211ringpll_sip       ( 
   					`ifndef ip2211ringpll_INTC_NO_PWR_PINS
      					.vccdig 					(vccdig_nom), 
      					.vss 						(vss),
   					`endif
					.ldo_enable				(ldo_enable),
					.fz_ldo_vinvoltsel			(fz_ldo_vinvoltsel),    // part of dfx_in
					.fz_ldo_bypass				(fz_ldo_bypass),    // part of dfx_in
					.fz_ldo_extrefsel			(fz_ldo_extrefsel),    // part of dfx_in
					.fz_ldo_faststart			(fz_ldo_faststart),    // part of dfx_in
					.fz_ldo_fbtrim				(fz_ldo_fbtrim),    // part of dfx_in
					.fz_ldo_reftrim				(fz_ldo_reftrim),    // part of dfx_in

					.view_mux_viewoutnnnnh 		(view_mux__ViewOutNnnnH),
					.pll_core_pfdlockrstnnnnh 		(pll_core__PfdLockRstNnnnH),
					.pll_fbgen_clkfbmxh 			(pll_fbgen__ClkFbMXH),
					.clkrefxxh 				(clkref),
					.bypassnnnnh 				(bypass),
					.reset_b_nnnnh 				(pllen),
					//.plldistpwrgoodnnnnh 			(pllen),
					.plldistpwrgoodnnnnh 			(powergood_vccdig),
					.rationnnnh 				(ratio),
					.fractionnnnnh 				(fraction),

					.mdiv_ratio				(mdiv_ratio),
					.mash_order_plus_one			(mash_order_plus_one),
					.ssccyctopeakm1				(ssc_cyc_to_peak_m1),
					.ssc_en					(ssc_en),
					.ssc_frac_step				(ssc_frac_step),

					.vcodiv_ratio				(vcodiv_ratio),
					.zdiv0_ratio				(zdiv0_ratio),
					.zdiv0_ratio_p5				(zdiv0_ratio_p5),
					.zdiv1_ratio				(zdiv1_ratio),
					.zdiv1_ratio_p5				(zdiv1_ratio_p5),


					.fz_cp1trim				(fz_cp1trim),
					.fz_cp2trim				(fz_cp2trim),
					.fz_cpnbias				(fz_cpnbias),
					.fz_dca_cb				(fz_dca_cb),
					.fz_dca_ctrl				(fz_dca_ctrl),
					.fz_irefgen				(fz_irefgen),
					.fz_lockcnt				(fz_lockcnt),
					.fz_lockforce				(fz_lockforce),
					.fz_lockstickyb				(fz_lockstickyb),
					.fz_lockthresh				(fz_lockthresh),
					.fz_lpfclksel				(fz_lpfclksel),
					.fz_nopfdpwrgate			(fz_nopfdpwrgate),
					.fz_pfd_pw				(fz_pfd_pw),
					.fz_pfddly				(fz_pfddly),
					.fz_skadj				(fz_skadj),	
					.fz_spare				(fz_spare),
					.fz_startup				(fz_startup),
					.fz_tight_loopb				(fz_tight_loopb),
					.fz_vcosel				(fz_vcosel),
					.fz_vcotrim				(fz_vcotrim),

					.idvdisable_bi				(idvdisable_bi),
					.idvfreqai				(idvfreqai),
					.idvfreqbi				(idvfreqbi),
					.idvpulsei				(idvpulsei),
					.idvtclki				(idvtclki),
					.idvtctrli				(idvtctrli),
					.idvtdi					(idvtdi),
					.idvtresi				(idvtresi),

                       			.idvdisable_bo                  	(idvdisable_bo),  // part of dfx_out
                        		.idvfreqao                      	(idvfreqao),      // part of dfx_out
                        		.idvfreqbo                      	(idvfreqbo),      // part of dfx_out
                        		.idvpulseo                      	(idvpulseo),      // part of dfx_out
                        		.idvtclko                       	(idvtclko),       // part of dfx_out
                        		.idvtctrlo                      	(idvtctrlo),      // part of dfx_out
                        		.idvtdo                         	(idvtdo),         // part of dfx_out
                        		.idvtreso                       	(idvtreso),       // part of dfx_out

					// RTDR interface
   					//
					.tdo					(tdo),
					.tck					(tck),
					//.sync_reset				(sync_reset),
					//.sync_reset				(1'b0),
					.tcapturedr				(tcapturedr),
					.tdi					(tdi),
					.treg_en				(treg_en),
					.trst_n					(trst_n),
					.tshiftdr				(tshiftdr),
					.tupdatedr				(tupdatedr),

					.view_adc_dig_out 			(view_adc__dig_out),
					.view_adc_done 			(view_adc__done),
					.clkidvih 				(ClkIdvIH),
						
					.ldo_enable_a				(ldo_enable_a),
					.ta_ldo_hiz_debug			(ta_ldo_hiz_debug),
					.ta_ldo_idq_debug			(ta_ldo_idq_debug),
					.fz_ldo_vinvoltsel_a			(fz_ldo_vinvoltsel_a),
					.fz_ldo_bypass_a			(fz_ldo_bypass_a),
					.fz_ldo_extrefsel_a			(fz_ldo_extrefsel_a),
					.fz_ldo_faststart_a			(fz_ldo_faststart_a),
					.fz_ldo_fbtrim_a			(fz_ldo_fbtrim_a),
					.fz_ldo_reftrim_a			(fz_ldo_reftrim_a),
					.dfx_powergood 			(dfx__powergood),


					.reset_sync_bypassxxnnnl 		(reset_sync__BypassXXnnnL),
					.reset_sync_bypassenxxnnnl 		(reset_sync__BypassEnXXnnnL),
					.reset_sync_reset_b_xxnnnl 		(reset_sync__Reset_b_XXnnnL),
					.mash_ratiomxh 			(mash__RatioMXH),
					.mash_halfintmxh 			(mash__HalfIntMXH),
					.mdiv_ratio_a				(mdiv_ratio_a),

					.vcodiv_ratio_a				(vcodiv_ratio_a),
					.zdiv0_ratio_a				(zdiv0_ratio_a),
					.zdiv0_ratio_p5_a			(zdiv0_ratio_p5_a),
					.zdiv1_ratio_a				(zdiv1_ratio_a),
					.zdiv1_ratio_p5_a			(zdiv1_ratio_p5_a),
					.ta_spare				(ta_spare),

					.idv_fub_idvgateennh 			(idv_fub__IdvGateEnNH),
					.dfx_cp1_trim 				(dfx__cp1_trim),
					.dfx_cp2_trim 				(dfx__cp2_trim),
					.fz_cpnbias_a				(fz_cpnbias_a),
					.fz_dca_cb_a				(fz_dca_cb_a),
					.dfx_dca_ctrl				(dfx__dca_ctrl),
					.fz_irefgen_a				(fz_irefgen_a),

					.dfx_lockthresh 			(dfx__lockthresh),
					.fz_lpfclksel_a				(fz_lpfclksel_a),
					.fz_nopfdpwrgate_a			(fz_nopfdpwrgate_a),
					.fz_pfd_pw_a				(fz_pfd_pw_a),
					.fz_pfddly_a				(fz_pfddly_a),
					.dfx_skadj_ctrl 			(dfx__skadj_ctrl),
					.fz_spare_a				(fz_spare_a),
					.fz_startup_a				(fz_startup_a),
					.dfx_tight_loop			(dfx__tight_loop),
					.fz_vcosel_a				(fz_vcosel_a),
					.fz_vcotrim_a				(fz_vcotrim_a),

					.tlctrl_sip_tightloopxxnnnh 		(tlctrl_sip__TightLoopXXnnnH),
					.adc_ctl_startxxh 			(adc_ctl__StartXXH),
					.adc_ctl_reset_bxxl 			(adc_ctl__Reset_bXXL),
					.dfx_adc_clkdiv 			(dfx__adc_clkdiv),
					.dfx_adc_freeze 			(dfx__adc_freeze),
					.dfx_adc_chop_en 			(dfx__adc_chop_en),
					.dfx_adc_use_vref 			(dfx__adc_use_vref),
					.dfx_adc_sel_in 			(dfx__adc_sel_in),
					.lock_detector_rawlockxxnnnl 		(lock_detector__RawLockXXnnnL),
					.lockxxnnnl 				(lock),
					.earlylockxxnnnh 			(EarlyLockXXnnnH),

					.idv_rdacctlth 			(idv__RdacCtlTH),
					.startup_gen_vctlrdacenxxh 		(startup_gen__VctlRdacEnXXH),
					.startup_gen_pfdenxxh 			(startup_gen__PfdEnXXH),


					.ssc_directionmxh 			(ssc__DirectionMXH),
					.ssc_mod_dfx_clkmodmxh 		(ssc_mod_dfx__ClkModMXH),
					.vctl_trim_fsm_vctlrdacshortxxh 	(vctl_trim_fsm__VctlRdacShortXXH),

					.dfx_viewdigennnnnh 			(dfx__ViewDigEnNnnnH),
					.dfx_viewanaennnnnh 			(dfx__ViewAnaEnNnnnH),
					//.dfx__ViewSelNnnnH 			(dfx__ViewSelNnnnH),
					.dfx_viewselnnnnh0			(viewsel0),
					.dfx_viewselnnnnh1			(viewsel1),

                                         //Scan interface
                                         .idfx_fscan_sdi,
                                         .idfx_fscan_mode,
                                         .idfx_fscan_shiften,
                                         .idfx_fscan_rstbypen,
                                         .idfx_fscan_byprstb,
                                         .idfx_fscan_clkungate,
                                         .odfx_fscan_sdo,

					.global_align_gateclkdistxxnnnl 	(tllm_gate_clk_trunk)			
				);

        // Output driver. This is being driven into SIP as well.
        assign view_dig_out = view_mux__ViewOutNnnnH;
logic hip_sync_rst;
//synchronizing powergood signal
     `ip2211ringpll_ASYNC_RST_2MSFF_META(hip_sync_rst, dfx__powergood,clkref, reset_sync__Reset_b_XXnnnL)


  
      
      // PLL Hard IP
      //   This block instantiates the PLL hard IP block that is delivered
      //   from the analog HIP team
      //
      //cpfljfulla                                    pll_hip         (
      ip2211ringpll_hip     iip2211ringpll_hip         (
  					`ifndef ip2211ringpll_INTC_NO_PWR_PINS
               	.vccdig			(vccdig_nom),
               	.vccpll			(vccpll),
               	.vccdist		(vccdist_nom),
               	.vccvdd2	        (vccldo_hv),
		.vss			(vss),
   					`endif
               	.vccref			(ldo_vref),
               .clkrefxxh               (   clkref                                            ),
               .clkpostdistmh           (   clkpostdist                                       ),
               //.reset_b_xxl           (   reset_sync__Reset_b_XXnnnL                        ),
               .reset_b_xxl             (   (hip_sync_rst)   ),//********8
               .bypassxxl               (   reset_sync__BypassXXnnnL                          ),
               .bypassenxxl             (   reset_sync__BypassEnXXnnnL                        ),
               .powergood               (   dfx__powergood                                    ),
               .ratio                   (   mash__RatioMXH                                    ),
	       .ratio_halfint           (   mash__HalfIntMXH                                  ),

	       .ratiozdiv0		(   zdiv0_ratio_a                                     ),
	       .zdiv0ratiop5            (   zdiv0_ratio_p5_a                                  ),
	       .ratiozdiv1		(   zdiv1_ratio_a                                     ),
	       .zdiv1ratiop5            (   zdiv1_ratio_p5_a                                  ),

               .adc_startxxh            (   adc_ctl__StartXXH                                 ),
               .adc_reset_bxxl          (   adc_ctl__Reset_bXXL                               ),
               .adc_clkdiv              (   dfx__adc_clkdiv                                   ),
               .adc_freeze              (   dfx__adc_freeze                                   ),
               .adc_chop_en             (   dfx__adc_chop_en                                  ),
               .adc_use_vref            (   dfx__adc_use_vref                                 ),
               .adc_sel_in              (   dfx__adc_sel_in                                   ),

               .clkfbmxh                (   pll_fbgen__ClkFbMXH                               ),
               .rawlockxxl              (   lock_detector__RawLockXXnnnL                      ),
               .lockxxl                 (   lock                                              ),
               .earlylockxxh            (   EarlyLockXXnnnH                                   ),


		// New pins
		.fz_lpfclksel		 (    fz_lpfclksel_a                                    ),
		.fz_nopfdpwrgate	 (    fz_nopfdpwrgate_a                                 ),
		.fz_tight_loopb		 (    dfx__tight_loop                                   ),
		.fz_vcosel		 (    fz_vcosel_a                                       ),
		.fz_cp1trim		 (    dfx__cp1_trim                                     ),
		.fz_cp2trim		 (    dfx__cp2_trim                                     ),
		.fz_cpnbias		 (    fz_cpnbias_a                                      ),
		.fz_dca_cb		 (    fz_dca_cb_a                                       ),
		.fz_dca_ctrl		 (    dfx__dca_ctrl                                     ),
		.fz_irefgen		 (    fz_irefgen_a                                      ),
		.fz_lockthresh		 (    dfx__lockthresh                                   ),
		.fz_pfd_pw		 (    fz_pfd_pw_a                                       ),
		.fz_pfddly		 (    fz_pfddly_a                                       ),
		.fz_skadj		 (    dfx__skadj_ctrl                                   ),
		.fz_spare		 (    fz_spare_a                                        ),
		.fz_startup		 (    fz_startup_a                                      ),
		.fz_vcotrim		 (    fz_vcotrim_a                                      ),

   		// LDO analog dft pins
                .anadft_ldovref		 (    anadft_ldovref					),
                .anadft_ldo		 (    anadft_ldo					),
                .anadft_ldovfb		 (    anadft_ldovfb					),

                .ssc_reload              (    ssc__DirectionMXH                                 ),
                .mod_clk_to_view         (     ssc_mod_dfx__ClkModMXH                            ),
                .vctlrdacctlnh           (     idv__RdacCtlTH                                    ),
                .vctlrdacennl            (     startup_gen__VctlRdacEnXXH                        ),
                .rdactovctlennh          (     vctl_trim_fsm__VctlRdacShortXXH                   ),
                .pfdennh                 (     startup_gen__PfdEnXXH                             ),

                .viewdigennh             (     dfx__ViewDigEnNnnnH                               ),
                .viewanaennh             (     dfx__ViewAnaEnNnnnH                               ),
                .viewsel0                (     viewsel0                                          ),
                .viewsel1                (     viewsel1                                          ),
                .viewoutnh               (    view_mux__ViewOutNnnnH                            ),
                .viewanabusnh            (     viewanabus                                        ),


                .tllm_force_tight_loop   (   tlctrl_sip__TightLoopXXnnnH                       ),
                .tllm_gate_clk_trunk     (   tllm_gate_clk_trunk                               ),

                .idv_gate_en             (     idv_fub__IdvGateEnNH                              ),
                .clkidvih                (     ClkIdvIH                                          ),

		.ta_spare		(     ta_spare                                         ),
	        .vcodiv_ratio		(   vcodiv_ratio_a                                    ),
	        .mdiv_ratio		(   mdiv_ratio_a                                      ),

                .adc_dig_out             (     view_adc__dig_out                                 ),
                .adc_done                (     view_adc__done                                    ),


                .pfdlockrstnh            (     pll_core__PfdLockRstNnnnH                         ),
	        .clkplldiv0              (   clkpll0                                           ),
	        .clkplldiv1              (   clkpll1                                           ),
                .clkpllmh                (     clkpll                                            )
          
              );

`endif // ifndef INTC_COLLAGE

 
   ///============================================================================
   /// SV Assertions
   ///============================================================================
   `ifndef ip2211ringpll_SVA_OFF
     
      //localparam FUSE_STRUCT_WIDTH = $bits(dfx_in.fuse);
      localparam FUSE_STRUCT_WIDTH = $bits(dfx_in.fuse);

      logic sva_output_en;
      logic sva_bypass_mode;
      logic sva_bypass_mode_pre;
      logic sva_reset;

      //assign sva_output_en = reset_sync__Reset_b_XXnnnL | (reset_sync__BypassXXnnnL & reset_sync__BypassEnXXnnnL);
      assign sva_output_en = reset_sync__Reset_b_XXnnnL | (bypass & reset_sync__BypassEnXXnnnL);
      //assign sva_bypass_mode = (reset_sync__BypassXXnnnL & reset_sync__BypassEnXXnnnL) & lock;
      assign sva_bypass_mode_pre = (reset_sync__BypassXXnnnL & reset_sync__BypassEnXXnnnL) & lock;
      //`ip2211ringpll_MSFF(sva_bypass_mode, sva_bypass_mode_pre, clkref)

      assign sva_reset     = ~sva_output_en;

      always @ (posedge clkref or posedge sva_reset) begin
	if (sva_reset) 
		sva_bypass_mode <= 1'b0;
	else
		sva_bypass_mode <= sva_bypass_mode_pre;
      end

      // LJPLL should not have X inputs when enabled
      //
      `ip2211ringpll_ASSERTS_KNOWN_DRIVEN(R_ljpll_X_inputs,
         //{clkref, pllen, PllDistPwrGoodNnnnH, 
         {clkref, pllen, pllen, 
         //BypassNnnnH, RatioNnnnH, FractionNnnnH, dfx_in.fuse, dfx_in.tap, dfx_in.register, dfx_in.odcs, dfx_in.ip2211ringpll_global_align},
         //bypass, ratio, fraction, dfx_in.fuse, tap_in,dfx_in.register, 1'b0, 1'b0},
         //bypass, ratio, fraction, 1'b0, tap_in,1'b0, 1'b0, 1'b0},
         bypass, ratio, fraction, 1'b0, 1'b0,1'b0, 1'b0, 1'b0},
         clkref, sva_reset,
      `ip2211ringpll_ERR_MSG("[LJPLL] X inputs to ljpll after powerup"));
 
      // LJPLL should not have X outputs after lock
      //
      `ip2211ringpll_ASSERTS_KNOWN_DRIVEN(R_ljpll_X_after_lock1,
         {EarlyLockXXnnnH, lock, clkpll,
         //dfx_out.tap, dfx_out.view.view_dig_out},
         //tap_in, view_dig_out},
         1'b0, view_dig_out},
         clkref, ~lock,
      `ip2211ringpll_ERR_MSG("[LJPLL] undriven outputs after lock"));
      
      // LJPLL should not have X outputs after lock
      //
      //`ip2211ringpll_ASSERTS_KNOWN_DRIVEN(R_ljpll_X_after_lock_sync,
      //   {ClkSyncMXH, SyncOutMnnnH},
      //   clkref, (~lock | ~SYNC_GEN_EN),
      //`ip2211ringpll_ERR_MSG("[LJPLL] undriven outputs after lock"));
     
      // IDV specific known drivens
      //
      //`ip2211ringpll_ASSERTS_KNOWN_DRIVEN(R_ljpll_X_inputs_idv,
      //{dfx_in.idv},
      //   clkref, sva_reset,
      //`ip2211ringpll_ERR_MSG("[LJPLL] IDV has X inputs to ljpll after powerup"));
      `ip2211ringpll_ASSERTS_KNOWN_DRIVEN(R_ljpll_X_inputs_idv,
         {idvtclki,idvtdi,idvtresi,idvtctrli,idvdisable_bi,idvfreqai,idvfreqbi,idvpulsei},
         clkref, sva_reset,
      `ip2211ringpll_ERR_MSG("[LJPLL] IDV has X inputs to ljpll after powerup"));
      
      //`ip2211ringpll_ASSERTS_KNOWN_DRIVEN(R_ljpll_X_after_lock_idv,
      //{dfx_out.idv},
      //  clkref, ~lock,
      //`ip2211ringpll_ERR_MSG("[LJPLL] undriven IDV outputs after lock"));
      `ip2211ringpll_ASSERTS_KNOWN_DRIVEN(R_ljpll_X_after_lock_idv,
         {idvtclko,idvtdo,idvtreso,idvtctrlo,idvdisable_bo,idvfreqao,idvfreqbo,idvpulseo},
         clkref, ~lock,
      `ip2211ringpll_ERR_MSG("[LJPLL] undriven IDV outputs after lock"));
      
      // Ratio may not change after pll is enabled (dynamic ratio
      //   change is not supported)
      //
      `ip2211ringpll_ASSERTS_STABLE(R_ljpll_dynamic_ratio,
                      {ratio,fraction},
                      $rose(reset_sync__Reset_b_XXnnnL),
                      lock,
                      posedge clkref,
                      sva_reset,
      `ip2211ringpll_ERR_MSG("[LJPLL] Ratio change after pllen but before lock is not supported"));

      // Fuse values may not change after pll is enabled
      //
      `ip2211ringpll_ASSERTS_STABLE(R_ljpll_fuse_stable,
                      dfx_in.fuse[FUSE_STRUCT_WIDTH-1:6], // ignore dca_ctrl
                      $rose(reset_sync__Reset_b_XXnnnL),
                      1'b0,
                      posedge clkref,
                      sva_reset,
      `ip2211ringpll_ERR_MSG("[LJPLL] Fuse bus changed when the PLL was enabled"));

      // Ratio must be >= 2 for proper PLL functionality
      //
      `ip2211ringpll_ASSERTS_FORBIDDEN(R_ljpll_illegal_ratio,
                         ratio < { {$bits(ratio)-2{1'b0}} , 2'h2 },
                         posedge reset_sync__Reset_b_XXnnnL,
                         1'b0,
      `ip2211ringpll_ERR_MSG("[LJPLL] PLL ratio must be >=2"));
      
      // PLL output clock must be clkref in bypass mode
      //
      `ip2211ringpll_ASSERTC_SAME(R_ljpll_bypass_clkout,
                    clkref,
                    clkpll,
                    ~sva_bypass_mode,
      `ip2211ringpll_ERR_MSG("[LJPLL] PLL output clock is expected to be reference clock in bypass mode but it is not"));

      // Earlylock must be asserted any time lock is asserted
      //
      `ip2211ringpll_ASSERTC_MUST(R_ljpll_earlylock_error,
                    (EarlyLockXXnnnH===1'b1),
                    ~lock,
      `ip2211ringpll_ERR_MSG("[LJPLL] PLL early lock is not asserted at time of lock"));

      // The PLL must lock within 104 reference clock cycles in normal
      //   operation (spec)
      //
      `ip2211ringpll_ASSERTS_TRIGGER(R_pllen2lock_sequence,
                       $rose(sva_output_en),
                       ##[8:190] $rose(lock),
                       posedge clkref,
                       //dfx_in.tap.openloop | sva_reset | reset_sync__BypassXXnnnL | dfx_in.ip2211ringpll_global_align ,
                       //tap_in.openloop | sva_reset | reset_sync__BypassXXnnnL ,
                       tap_in.openloop | sva_reset | sva_bypass_mode ,
      `ip2211ringpll_ERR_MSG("[LJPLL] The PLL is expected to lock within 190 reference clock cycles"));
      
      // The PLL must lock within 5 reference clock cycles in bypass mode
      //
      `ip2211ringpll_ASSERTS_TRIGGER(R_pllbypen2lock_sequence,
                       $rose(sva_output_en),
                       ##[0:5] $rose(lock),
                       posedge clkref,
                       //dfx_in.tap.openloop | sva_reset | ~reset_sync__BypassXXnnnL,
                       //tap_in.openloop | sva_reset | ~reset_sync__BypassXXnnnL,
                       tap_in.openloop | sva_reset | ~sva_bypass_mode,
      `ip2211ringpll_ERR_MSG("[LJPLL] The PLL is expected to lock within 104 reference clock cycles"));

      // The sync generator must be disabled when we are operating in
      //   FRAC-N or SSC mode
      //
//      `ip2211ringpll_ASSERTC_MUST(R_syncgen_disabled_ssc_frac_mode, 
                    //~(SYNC_GEN_EN & ((dfx_in.register.ssc_en & SSC_EN)  | (|fraction))),
//                    ~(((ssc_en)  | (|fraction))),
//                    ~reset_sync__Reset_b_XXnnnL,
//      `ip2211ringpll_ERR_MSG("[LJPLL] The SYNC_GEN_EN parameter should be tied OFF when the LJPLL is expected to use Frac-N or SSC. This enables power savings and prevents mistakes."));

      // Global align is not supported when the sync generator is enabled
      //
      //`ip2211ringpll_ASSERTC_MUST(R_syncgen_disabled_global_align, 
      //              ~(SYNC_GEN_EN & (dfx_in.ip2211ringpll_global_align)),
      //              ~reset_sync__Reset_b_XXnnnL,
      //`ip2211ringpll_ERR_MSG("[LJPLL] The SYNC_GEN_EN parameter should be tied OFF when the LJPLL is expected to use the global align feature"));

   `endif

///========================================================================================================
/// Module End
///========================================================================================================
//`endif
endmodule

`endif

//`endcelldefine


