VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO Noise_injection_block_modified_v13
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN Noise_injection_block_modified_v13 0 0 ;
  SIZE 18.576 BY 189.7985 ;
  SYMMETRY X Y R90 ;
  PIN Random
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m2 ;
        RECT 0 189.7345 0.3215 189.7785 ;
    END
  END Random
  PIN Iout
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER m3 ;
        RECT 1.5995 189.7545 1.6435 189.7985 ;
    END
  END Iout
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER m3 ;
        RECT 0.4455 0.2035 0.4895 189.3885 ;
    END
    PORT
      LAYER m3 ;
        RECT 18.0865 0.4945 18.1305 189.3885 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER m3 ;
        RECT 0.811 0.225 0.855 189.5685 ;
    END
    PORT
      LAYER m3 ;
        RECT 17.721 0.5445 17.765 189.5685 ;
    END
  END vss
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 2.4125 0.044 2.4565 ;
    END
  END S[0]
  PIN S[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 129.8525 0.044 129.8965 ;
    END
  END S[10]
  PIN S[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 18.532 129.8525 18.576 129.8965 ;
    END
  END S[11]
  PIN S[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 144.9725 0.044 145.0165 ;
    END
  END S[12]
  PIN S[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 159.0125 0.044 159.0565 ;
    END
  END S[13]
  PIN S[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 177.3725 0.044 177.4165 ;
    END
  END S[14]
  PIN S[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 18.532 177.3725 18.576 177.4165 ;
    END
  END S[15]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 16.4525 0.044 16.4965 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 34.8125 0.044 34.8565 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 18.532 34.8125 18.576 34.8565 ;
    END
  END S[3]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 49.9325 0.044 49.9765 ;
    END
  END S[4]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 63.9725 0.044 64.0165 ;
    END
  END S[5]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 82.3325 0.044 82.3765 ;
    END
  END S[6]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 18.532 82.3325 18.576 82.3765 ;
    END
  END S[7]
  PIN S[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 97.4525 0.044 97.4965 ;
    END
  END S[8]
  PIN S[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER m6 ;
        RECT 0 111.4925 0.044 111.5365 ;
    END
  END S[9]
  PIN VB[0]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m6 ;
        RECT 0 0.0055 0.448 0.0955 ;
    END
  END VB[0]
  PIN VB[1]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m6 ;
        RECT 0 47.5255 0.25 47.6155 ;
    END
  END VB[1]
  PIN VB[2]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m6 ;
        RECT 0 95.0455 0.25 95.1355 ;
    END
  END VB[2]
  PIN VB[3]
    DIRECTION INPUT ;
    USE ANALOG ;
    PORT
      LAYER m6 ;
        RECT 0 142.5655 0.358 142.6555 ;
    END
  END VB[3]
  OBS
    LAYER m1 SPACING 0.04 ;
      RECT 0 0 18.576 189.7985 ;
    LAYER m5 SPACING 0.046 ;
      RECT 0 0 18.576 189.7985 ;
    LAYER m2 ;
      RECT 0.3815 189.7345 8.4375 189.7785 ;
    LAYER m2 SPACING 0.046 ;
      RECT 0.4015 0 18.576 189.7985 ;
      RECT 0 0 18.576 189.6545 ;
    LAYER m3 ;
      RECT 1.5995 37.0345 1.6435 189.6545 ;
      RECT 0.4455 189.4945 0.4895 189.5945 ;
    LAYER m3 SPACING 0.046 ;
      RECT 1.7235 189.6485 18.576 189.7985 ;
      RECT 18.2105 0 18.576 189.7985 ;
      RECT 0.4175 189.6485 1.5195 189.7985 ;
      RECT 0.935 0 17.641 189.6745 ;
      RECT 17.845 189.4685 18.576 189.7985 ;
      RECT 0.4175 189.4685 0.731 189.7985 ;
      RECT 0.5695 0 0.731 189.7985 ;
      RECT 0 189.4685 0.731 189.6385 ;
      RECT 17.845 0 18.0065 189.7985 ;
      RECT 0 0 0.3655 189.6385 ;
      RECT 0 177.3145 0.397 177.4745 ;
      RECT 0 49.8745 0.3975 50.0345 ;
      RECT 0.935 0 18.0065 0.4645 ;
      RECT 0.935 0 18.576 0.4145 ;
      RECT 0.5695 0 18.576 0.145 ;
      RECT 0 0 18.576 0.1235 ;
    LAYER m4 SPACING 0.046 ;
      RECT 1.7395 189.6645 18.576 189.7985 ;
      RECT 18.2265 0 18.576 189.7985 ;
      RECT 0 189.6645 1.5035 189.7985 ;
      RECT 0.951 0 1.5035 189.7985 ;
      RECT 17.861 189.4845 18.576 189.7985 ;
      RECT 1.7395 0 17.625 189.7985 ;
      RECT 0 189.4845 0.715 189.7985 ;
      RECT 0.5855 0 0.715 189.7985 ;
      RECT 0.951 0 17.625 189.6585 ;
      RECT 17.861 0 17.9905 189.7985 ;
      RECT 0 0 0.3495 189.7985 ;
      RECT 18.1575 177.3725 18.576 177.4165 ;
      RECT 0 177.3725 0.455 177.4165 ;
      RECT 0 159.0125 0.378 159.0565 ;
      RECT 0 144.9725 0.374 145.0165 ;
      RECT 18.1685 129.8525 18.576 129.8965 ;
      RECT 0 129.8525 0.3565 129.8965 ;
      RECT 0 111.4925 0.3755 111.5365 ;
      RECT 18.1605 82.3325 18.576 82.3765 ;
      RECT 0 82.3325 0.373 82.3765 ;
      RECT 0 63.9725 0.3815 64.0165 ;
      RECT 0 49.9325 0.4555 49.9765 ;
      RECT 18.188 34.8125 18.576 34.8565 ;
      RECT 0 34.8125 0.3525 34.8565 ;
      RECT 0 16.4525 0.3755 16.4965 ;
      RECT 0 2.4125 0.3775 2.4565 ;
      RECT 0.951 0 17.9905 0.4485 ;
      RECT 0.951 0 18.576 0.3985 ;
      RECT 0.5855 0 18.576 0.129 ;
      RECT 0 0 18.576 0.1075 ;
    LAYER m8 SPACING 0.18 ;
      RECT 0 0 18.576 189.7985 ;
    LAYER m6 ;
      RECT 7.0425 0.005 7.1325 0.38 ;
      RECT 11.4435 0.005 11.5335 0.322 ;
      RECT 0.548 0.0055 7.1325 0.0955 ;
      RECT 7.0425 0.005 11.5335 0.095 ;
      RECT 17.787 34.8125 18.432 34.8565 ;
      RECT 17.825 82.3325 18.432 82.3765 ;
      RECT 17.825 129.8525 18.432 129.8965 ;
      RECT 17.8185 177.3725 18.432 177.4165 ;
      RECT 0.35 47.5255 7.0425 47.6155 ;
      RECT 0.35 95.0455 7.0425 95.1355 ;
      RECT 0.458 142.5655 7.0425 142.6555 ;
      RECT 0.144 49.9325 0.4255 49.9765 ;
      RECT 0.144 177.3725 0.425 177.4165 ;
      RECT 0.144 63.9725 0.3515 64.0165 ;
      RECT 0.144 159.0125 0.348 159.0565 ;
      RECT 0.144 2.4125 0.3475 2.4565 ;
      RECT 0.144 16.4525 0.3455 16.4965 ;
      RECT 0.144 111.4925 0.3455 111.5365 ;
      RECT 0.144 144.9725 0.344 145.0165 ;
      RECT 0.144 82.3325 0.343 82.3765 ;
      RECT 0.144 129.8525 0.3265 129.8965 ;
      RECT 0.144 34.8125 0.3225 34.8565 ;
      RECT 0.144 97.4525 0.3165 97.4965 ;
    LAYER m6 SPACING 0.046 ;
      RECT 0 177.6225 18.576 189.7985 ;
      RECT 0.25 142.8615 18.326 189.7985 ;
      RECT 0 159.2625 18.576 177.1665 ;
      RECT 0.564 130.1025 18.576 177.1665 ;
      RECT 0 145.2225 18.576 158.8065 ;
      RECT 0 142.8615 18.576 144.7665 ;
      RECT 0 130.1025 18.576 142.3595 ;
      RECT 0.25 95.3415 18.326 142.3595 ;
      RECT 0 111.7425 18.576 129.6465 ;
      RECT 0.456 82.5825 18.576 129.6465 ;
      RECT 0 97.7025 18.576 111.2865 ;
      RECT 0 95.3415 18.576 97.2465 ;
      RECT 0 82.5825 18.576 94.8395 ;
      RECT 0.25 47.8215 18.326 94.8395 ;
      RECT 0 64.2225 18.576 82.1265 ;
      RECT 0.456 35.0625 18.576 82.1265 ;
      RECT 0 50.1825 18.576 63.7665 ;
      RECT 0 47.8215 18.576 49.7265 ;
      RECT 0 35.0625 18.576 47.3195 ;
      RECT 0.25 0.3015 18.326 47.3195 ;
      RECT 0 16.7025 18.576 34.6065 ;
      RECT 0.654 0 18.576 34.6065 ;
      RECT 0 2.6625 18.576 16.2465 ;
      RECT 0 0.3015 18.576 2.2065 ;
    LAYER m7 SPACING 0.18 ;
      RECT 0 177.7565 18.576 189.7985 ;
      RECT 0.384 142.9955 18.192 189.7985 ;
      RECT 0 159.3965 18.576 177.0325 ;
      RECT 0.698 130.2365 18.576 177.0325 ;
      RECT 0 145.3565 18.576 158.6725 ;
      RECT 0 142.9955 18.576 144.6325 ;
      RECT 0 130.2365 18.576 142.2255 ;
      RECT 0.384 95.4755 18.192 142.2255 ;
      RECT 0 111.8765 18.576 129.5125 ;
      RECT 0.59 82.7165 18.576 129.5125 ;
      RECT 0 97.8365 18.576 111.1525 ;
      RECT 0 95.4755 18.576 97.1125 ;
      RECT 0 82.7165 18.576 94.7055 ;
      RECT 0.384 47.9555 18.192 94.7055 ;
      RECT 0 64.3565 18.576 81.9925 ;
      RECT 0.59 35.1965 18.576 81.9925 ;
      RECT 0 50.3165 18.576 63.6325 ;
      RECT 0 47.9555 18.576 49.5925 ;
      RECT 0 35.1965 18.576 47.1855 ;
      RECT 0.384 0.4355 18.192 47.1855 ;
      RECT 0 16.8365 18.576 34.4725 ;
      RECT 0.788 0 18.576 34.4725 ;
      RECT 0 2.7965 18.576 16.1125 ;
      RECT 0 0.4355 18.576 2.0725 ;
    LAYER gm0 SPACING 0.54 ;
      RECT 0 0 18.576 189.7985 ;
    LAYER gmz SPACING 0.54 ;
      RECT 0 0 18.576 189.7985 ;
    LAYER gmb SPACING 1 ;
      RECT 0 0 18.576 189.7985 ;
  END
END Noise_injection_block_modified_v13

END LIBRARY
